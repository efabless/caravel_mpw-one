magic
tech sky130A
magscale 1 2
timestamp 1625004094
<< nwell >>
rect 231772 997737 243593 998041
rect 283172 997737 294993 998041
rect 341772 997737 353593 998041
rect 577972 997737 589793 998041
rect 677737 944807 678041 956628
rect 39559 873172 39863 884993
rect 678733 862378 679465 863083
rect 688918 862857 693847 863143
rect 695297 863024 696080 863083
rect 681431 850034 682216 862084
rect 688918 858297 689204 862857
rect 689636 862238 690068 862857
rect 689636 860908 689804 862238
rect 689754 860293 689804 860908
rect 693561 858037 693847 862857
rect 694716 862441 696080 863024
rect 694716 862094 695964 862441
rect 694932 861805 695964 862094
rect 694932 861316 695256 861805
rect 694932 861301 695148 861316
rect 684453 851345 684811 853217
rect 684082 850034 684811 851345
rect 681431 846910 682669 850034
rect 683557 846910 684811 850034
rect 692119 850470 692253 853612
rect 687724 847175 688010 848933
rect 690639 847175 690809 848933
rect 692119 847175 692355 850470
rect 687724 847152 692355 847175
rect 694233 847152 694469 853612
rect 696449 850470 696633 853612
rect 696347 847152 696633 850470
rect 687724 846866 696633 847152
rect 703733 853792 705676 863083
rect 703733 846912 705677 853792
rect 706576 861723 713395 863083
rect 706576 847274 706938 861723
rect 711303 861497 713395 861723
rect 711303 849606 711695 861497
rect 712309 849606 713395 861497
rect 711303 847274 713395 849606
rect 706576 846913 713395 847274
rect 706576 846912 711646 846913
rect 39559 830772 39863 842593
rect 677737 804607 678041 816428
rect 5954 801287 11024 801288
rect 4205 800926 11024 801287
rect 4205 798594 6297 800926
rect 4205 786703 5291 798594
rect 5905 786703 6297 798594
rect 4205 786477 6297 786703
rect 10662 786477 11024 800926
rect 4205 785117 11024 786477
rect 11923 794408 13867 801288
rect 11924 785117 13867 794408
rect 20967 801048 29876 801334
rect 20967 797730 21253 801048
rect 20967 794588 21151 797730
rect 23131 794588 23367 801048
rect 25245 801025 29876 801048
rect 25245 797730 25481 801025
rect 26791 799267 26961 801025
rect 29590 799267 29876 801025
rect 25347 794588 25481 797730
rect 32789 798166 34043 801290
rect 34931 798166 36169 801290
rect 32789 796855 33518 798166
rect 32789 794983 33147 796855
rect 22452 786884 22668 786899
rect 22344 786395 22668 786884
rect 21636 786106 22668 786395
rect 21636 785759 22884 786106
rect 21520 785176 22884 785759
rect 23753 785343 24039 790163
rect 27796 787292 27846 787907
rect 27796 785962 27964 787292
rect 27532 785343 27964 785962
rect 28396 785343 28682 789903
rect 35384 786116 36169 798166
rect 21520 785117 22303 785176
rect 23753 785057 28682 785343
rect 38135 785117 38867 785822
rect 678733 774978 679465 775683
rect 688918 775457 693847 775743
rect 695297 775624 696080 775683
rect 681431 762634 682216 774684
rect 688918 770897 689204 775457
rect 689636 774838 690068 775457
rect 689636 773508 689804 774838
rect 689754 772893 689804 773508
rect 693561 770637 693847 775457
rect 694716 775041 696080 775624
rect 694716 774694 695964 775041
rect 694932 774405 695964 774694
rect 694932 773916 695256 774405
rect 694932 773901 695148 773916
rect 684453 763945 684811 765817
rect 684082 762634 684811 763945
rect 681431 759510 682669 762634
rect 683557 759510 684811 762634
rect 692119 763070 692253 766212
rect 687724 759775 688010 761533
rect 690639 759775 690809 761533
rect 692119 759775 692355 763070
rect 687724 759752 692355 759775
rect 694233 759752 694469 766212
rect 696449 763070 696633 766212
rect 696347 759752 696633 763070
rect 687724 759466 696633 759752
rect 703733 766392 705676 775683
rect 703733 759512 705677 766392
rect 706576 774323 713395 775683
rect 706576 759874 706938 774323
rect 711303 774097 713395 774323
rect 711303 762206 711695 774097
rect 712309 762206 713395 774097
rect 711303 759874 713395 762206
rect 706576 759513 713395 759874
rect 706576 759512 711646 759513
rect 5954 758087 11024 758088
rect 4205 757726 11024 758087
rect 4205 755394 6297 757726
rect 4205 743503 5291 755394
rect 5905 743503 6297 755394
rect 4205 743277 6297 743503
rect 10662 743277 11024 757726
rect 4205 741917 11024 743277
rect 11923 751208 13867 758088
rect 11924 741917 13867 751208
rect 20967 757848 29876 758134
rect 20967 754530 21253 757848
rect 20967 751388 21151 754530
rect 23131 751388 23367 757848
rect 25245 757825 29876 757848
rect 25245 754530 25481 757825
rect 26791 756067 26961 757825
rect 29590 756067 29876 757825
rect 25347 751388 25481 754530
rect 32789 754966 34043 758090
rect 34931 754966 36169 758090
rect 32789 753655 33518 754966
rect 32789 751783 33147 753655
rect 22452 743684 22668 743699
rect 22344 743195 22668 743684
rect 21636 742906 22668 743195
rect 21636 742559 22884 742906
rect 21520 741976 22884 742559
rect 23753 742143 24039 746963
rect 27796 744092 27846 744707
rect 27796 742762 27964 744092
rect 27532 742143 27964 742762
rect 28396 742143 28682 746703
rect 35384 742916 36169 754966
rect 21520 741917 22303 741976
rect 23753 741857 28682 742143
rect 38135 741917 38867 742622
rect 678733 730578 679465 731283
rect 688918 731057 693847 731343
rect 695297 731224 696080 731283
rect 681431 718234 682216 730284
rect 688918 726497 689204 731057
rect 689636 730438 690068 731057
rect 689636 729108 689804 730438
rect 689754 728493 689804 729108
rect 693561 726237 693847 731057
rect 694716 730641 696080 731224
rect 694716 730294 695964 730641
rect 694932 730005 695964 730294
rect 694932 729516 695256 730005
rect 694932 729501 695148 729516
rect 684453 719545 684811 721417
rect 684082 718234 684811 719545
rect 681431 715110 682669 718234
rect 683557 715110 684811 718234
rect 692119 718670 692253 721812
rect 687724 715375 688010 717133
rect 690639 715375 690809 717133
rect 692119 715375 692355 718670
rect 687724 715352 692355 715375
rect 694233 715352 694469 721812
rect 696449 718670 696633 721812
rect 696347 715352 696633 718670
rect 687724 715066 696633 715352
rect 703733 721992 705676 731283
rect 703733 715112 705677 721992
rect 706576 729923 713395 731283
rect 706576 715474 706938 729923
rect 711303 729697 713395 729923
rect 711303 717806 711695 729697
rect 712309 717806 713395 729697
rect 711303 715474 713395 717806
rect 706576 715113 713395 715474
rect 706576 715112 711646 715113
rect 5954 714887 11024 714888
rect 4205 714526 11024 714887
rect 4205 712194 6297 714526
rect 4205 700303 5291 712194
rect 5905 700303 6297 712194
rect 4205 700077 6297 700303
rect 10662 700077 11024 714526
rect 4205 698717 11024 700077
rect 11923 708008 13867 714888
rect 11924 698717 13867 708008
rect 20967 714648 29876 714934
rect 20967 711330 21253 714648
rect 20967 708188 21151 711330
rect 23131 708188 23367 714648
rect 25245 714625 29876 714648
rect 25245 711330 25481 714625
rect 26791 712867 26961 714625
rect 29590 712867 29876 714625
rect 25347 708188 25481 711330
rect 32789 711766 34043 714890
rect 34931 711766 36169 714890
rect 32789 710455 33518 711766
rect 32789 708583 33147 710455
rect 22452 700484 22668 700499
rect 22344 699995 22668 700484
rect 21636 699706 22668 699995
rect 21636 699359 22884 699706
rect 21520 698776 22884 699359
rect 23753 698943 24039 703763
rect 27796 700892 27846 701507
rect 27796 699562 27964 700892
rect 27532 698943 27964 699562
rect 28396 698943 28682 703503
rect 35384 699716 36169 711766
rect 21520 698717 22303 698776
rect 23753 698657 28682 698943
rect 38135 698717 38867 699422
rect 678733 686378 679465 687083
rect 688918 686857 693847 687143
rect 695297 687024 696080 687083
rect 681431 674034 682216 686084
rect 688918 682297 689204 686857
rect 689636 686238 690068 686857
rect 689636 684908 689804 686238
rect 689754 684293 689804 684908
rect 693561 682037 693847 686857
rect 694716 686441 696080 687024
rect 694716 686094 695964 686441
rect 694932 685805 695964 686094
rect 694932 685316 695256 685805
rect 694932 685301 695148 685316
rect 684453 675345 684811 677217
rect 684082 674034 684811 675345
rect 5954 671487 11024 671488
rect 4205 671126 11024 671487
rect 4205 668794 6297 671126
rect 4205 656903 5291 668794
rect 5905 656903 6297 668794
rect 4205 656677 6297 656903
rect 10662 656677 11024 671126
rect 4205 655317 11024 656677
rect 11923 664608 13867 671488
rect 11924 655317 13867 664608
rect 20967 671248 29876 671534
rect 20967 667930 21253 671248
rect 20967 664788 21151 667930
rect 23131 664788 23367 671248
rect 25245 671225 29876 671248
rect 25245 667930 25481 671225
rect 26791 669467 26961 671225
rect 29590 669467 29876 671225
rect 25347 664788 25481 667930
rect 32789 668366 34043 671490
rect 34931 668366 36169 671490
rect 681431 670910 682669 674034
rect 683557 670910 684811 674034
rect 692119 674470 692253 677612
rect 687724 671175 688010 672933
rect 690639 671175 690809 672933
rect 692119 671175 692355 674470
rect 687724 671152 692355 671175
rect 694233 671152 694469 677612
rect 696449 674470 696633 677612
rect 696347 671152 696633 674470
rect 687724 670866 696633 671152
rect 703733 677792 705676 687083
rect 703733 670912 705677 677792
rect 706576 685723 713395 687083
rect 706576 671274 706938 685723
rect 711303 685497 713395 685723
rect 711303 673606 711695 685497
rect 712309 673606 713395 685497
rect 711303 671274 713395 673606
rect 706576 670913 713395 671274
rect 706576 670912 711646 670913
rect 32789 667055 33518 668366
rect 32789 665183 33147 667055
rect 22452 657084 22668 657099
rect 22344 656595 22668 657084
rect 21636 656306 22668 656595
rect 21636 655959 22884 656306
rect 21520 655376 22884 655959
rect 23753 655543 24039 660363
rect 27796 657492 27846 658107
rect 27796 656162 27964 657492
rect 27532 655543 27964 656162
rect 28396 655543 28682 660103
rect 35384 656316 36169 668366
rect 21520 655317 22303 655376
rect 23753 655257 28682 655543
rect 38135 655317 38867 656022
rect 678733 642178 679465 642883
rect 688918 642657 693847 642943
rect 695297 642824 696080 642883
rect 681431 629834 682216 641884
rect 688918 638097 689204 642657
rect 689636 642038 690068 642657
rect 689636 640708 689804 642038
rect 689754 640093 689804 640708
rect 693561 637837 693847 642657
rect 694716 642241 696080 642824
rect 694716 641894 695964 642241
rect 694932 641605 695964 641894
rect 694932 641116 695256 641605
rect 694932 641101 695148 641116
rect 684453 631145 684811 633017
rect 684082 629834 684811 631145
rect 5954 628287 11024 628288
rect 4205 627926 11024 628287
rect 4205 625594 6297 627926
rect 4205 613703 5291 625594
rect 5905 613703 6297 625594
rect 4205 613477 6297 613703
rect 10662 613477 11024 627926
rect 4205 612117 11024 613477
rect 11923 621408 13867 628288
rect 11924 612117 13867 621408
rect 20967 628048 29876 628334
rect 20967 624730 21253 628048
rect 20967 621588 21151 624730
rect 23131 621588 23367 628048
rect 25245 628025 29876 628048
rect 25245 624730 25481 628025
rect 26791 626267 26961 628025
rect 29590 626267 29876 628025
rect 25347 621588 25481 624730
rect 32789 625166 34043 628290
rect 34931 625166 36169 628290
rect 681431 626710 682669 629834
rect 683557 626710 684811 629834
rect 692119 630270 692253 633412
rect 687724 626975 688010 628733
rect 690639 626975 690809 628733
rect 692119 626975 692355 630270
rect 687724 626952 692355 626975
rect 694233 626952 694469 633412
rect 696449 630270 696633 633412
rect 696347 626952 696633 630270
rect 687724 626666 696633 626952
rect 703733 633592 705676 642883
rect 703733 626712 705677 633592
rect 706576 641523 713395 642883
rect 706576 627074 706938 641523
rect 711303 641297 713395 641523
rect 711303 629406 711695 641297
rect 712309 629406 713395 641297
rect 711303 627074 713395 629406
rect 706576 626713 713395 627074
rect 706576 626712 711646 626713
rect 32789 623855 33518 625166
rect 32789 621983 33147 623855
rect 22452 613884 22668 613899
rect 22344 613395 22668 613884
rect 21636 613106 22668 613395
rect 21636 612759 22884 613106
rect 21520 612176 22884 612759
rect 23753 612343 24039 617163
rect 27796 614292 27846 614907
rect 27796 612962 27964 614292
rect 27532 612343 27964 612962
rect 28396 612343 28682 616903
rect 35384 613116 36169 625166
rect 21520 612117 22303 612176
rect 23753 612057 28682 612343
rect 38135 612117 38867 612822
rect 678733 597778 679465 598483
rect 688918 598257 693847 598543
rect 695297 598424 696080 598483
rect 681431 585434 682216 597484
rect 688918 593697 689204 598257
rect 689636 597638 690068 598257
rect 689636 596308 689804 597638
rect 689754 595693 689804 596308
rect 693561 593437 693847 598257
rect 694716 597841 696080 598424
rect 694716 597494 695964 597841
rect 694932 597205 695964 597494
rect 694932 596716 695256 597205
rect 694932 596701 695148 596716
rect 684453 586745 684811 588617
rect 684082 585434 684811 586745
rect 5954 585087 11024 585088
rect 4205 584726 11024 585087
rect 4205 582394 6297 584726
rect 4205 570503 5291 582394
rect 5905 570503 6297 582394
rect 4205 570277 6297 570503
rect 10662 570277 11024 584726
rect 4205 568917 11024 570277
rect 11923 578208 13867 585088
rect 11924 568917 13867 578208
rect 20967 584848 29876 585134
rect 20967 581530 21253 584848
rect 20967 578388 21151 581530
rect 23131 578388 23367 584848
rect 25245 584825 29876 584848
rect 25245 581530 25481 584825
rect 26791 583067 26961 584825
rect 29590 583067 29876 584825
rect 25347 578388 25481 581530
rect 32789 581966 34043 585090
rect 34931 581966 36169 585090
rect 681431 582310 682669 585434
rect 683557 582310 684811 585434
rect 692119 585870 692253 589012
rect 687724 582575 688010 584333
rect 690639 582575 690809 584333
rect 692119 582575 692355 585870
rect 687724 582552 692355 582575
rect 694233 582552 694469 589012
rect 696449 585870 696633 589012
rect 696347 582552 696633 585870
rect 687724 582266 696633 582552
rect 703733 589192 705676 598483
rect 703733 582312 705677 589192
rect 706576 597123 713395 598483
rect 706576 582674 706938 597123
rect 711303 596897 713395 597123
rect 711303 585006 711695 596897
rect 712309 585006 713395 596897
rect 711303 582674 713395 585006
rect 706576 582313 713395 582674
rect 706576 582312 711646 582313
rect 32789 580655 33518 581966
rect 32789 578783 33147 580655
rect 22452 570684 22668 570699
rect 22344 570195 22668 570684
rect 21636 569906 22668 570195
rect 21636 569559 22884 569906
rect 21520 568976 22884 569559
rect 23753 569143 24039 573963
rect 27796 571092 27846 571707
rect 27796 569762 27964 571092
rect 27532 569143 27964 569762
rect 28396 569143 28682 573703
rect 35384 569916 36169 581966
rect 21520 568917 22303 568976
rect 23753 568857 28682 569143
rect 38135 568917 38867 569622
rect 678733 553578 679465 554283
rect 688918 554057 693847 554343
rect 695297 554224 696080 554283
rect 5954 541887 11024 541888
rect 4205 541526 11024 541887
rect 4205 539194 6297 541526
rect 4205 527303 5291 539194
rect 5905 527303 6297 539194
rect 4205 527077 6297 527303
rect 10662 527077 11024 541526
rect 4205 525717 11024 527077
rect 11923 535008 13867 541888
rect 11924 525717 13867 535008
rect 20967 541648 29876 541934
rect 20967 538330 21253 541648
rect 20967 535188 21151 538330
rect 23131 535188 23367 541648
rect 25245 541625 29876 541648
rect 25245 538330 25481 541625
rect 26791 539867 26961 541625
rect 29590 539867 29876 541625
rect 25347 535188 25481 538330
rect 32789 538766 34043 541890
rect 34931 538766 36169 541890
rect 32789 537455 33518 538766
rect 32789 535583 33147 537455
rect 22452 527484 22668 527499
rect 22344 526995 22668 527484
rect 21636 526706 22668 526995
rect 21636 526359 22884 526706
rect 21520 525776 22884 526359
rect 23753 525943 24039 530763
rect 27796 527892 27846 528507
rect 27796 526562 27964 527892
rect 27532 525943 27964 526562
rect 28396 525943 28682 530503
rect 35384 526716 36169 538766
rect 681431 541234 682216 553284
rect 688918 549497 689204 554057
rect 689636 553438 690068 554057
rect 689636 552108 689804 553438
rect 689754 551493 689804 552108
rect 693561 549237 693847 554057
rect 694716 553641 696080 554224
rect 694716 553294 695964 553641
rect 694932 553005 695964 553294
rect 694932 552516 695256 553005
rect 694932 552501 695148 552516
rect 684453 542545 684811 544417
rect 684082 541234 684811 542545
rect 681431 538110 682669 541234
rect 683557 538110 684811 541234
rect 692119 541670 692253 544812
rect 687724 538375 688010 540133
rect 690639 538375 690809 540133
rect 692119 538375 692355 541670
rect 687724 538352 692355 538375
rect 694233 538352 694469 544812
rect 696449 541670 696633 544812
rect 696347 538352 696633 541670
rect 687724 538066 696633 538352
rect 703733 544992 705676 554283
rect 703733 538112 705677 544992
rect 706576 552923 713395 554283
rect 706576 538474 706938 552923
rect 711303 552697 713395 552923
rect 711303 540806 711695 552697
rect 712309 540806 713395 552697
rect 711303 538474 713395 540806
rect 706576 538113 713395 538474
rect 706576 538112 711646 538113
rect 21520 525717 22303 525776
rect 23753 525657 28682 525943
rect 38135 525717 38867 526422
rect 39559 485772 39863 497593
rect 677737 495807 678041 507628
rect 5954 414087 11024 414088
rect 4205 413726 11024 414087
rect 4205 411394 6297 413726
rect 4205 399503 5291 411394
rect 5905 399503 6297 411394
rect 4205 399277 6297 399503
rect 10662 399277 11024 413726
rect 4205 397917 11024 399277
rect 11923 407208 13867 414088
rect 11924 397917 13867 407208
rect 20967 413848 29876 414134
rect 20967 410530 21253 413848
rect 20967 407388 21151 410530
rect 23131 407388 23367 413848
rect 25245 413825 29876 413848
rect 25245 410530 25481 413825
rect 26791 412067 26961 413825
rect 29590 412067 29876 413825
rect 25347 407388 25481 410530
rect 32789 410966 34043 414090
rect 34931 410966 36169 414090
rect 32789 409655 33518 410966
rect 32789 407783 33147 409655
rect 22452 399684 22668 399699
rect 22344 399195 22668 399684
rect 21636 398906 22668 399195
rect 21636 398559 22884 398906
rect 21520 397976 22884 398559
rect 23753 398143 24039 402963
rect 27796 400092 27846 400707
rect 27796 398762 27964 400092
rect 27532 398143 27964 398762
rect 28396 398143 28682 402703
rect 35384 398916 36169 410966
rect 677737 409207 678041 421028
rect 21520 397917 22303 397976
rect 23753 397857 28682 398143
rect 38135 397917 38867 398622
rect 678733 379378 679465 380083
rect 688918 379857 693847 380143
rect 695297 380024 696080 380083
rect 5954 370887 11024 370888
rect 4205 370526 11024 370887
rect 4205 368194 6297 370526
rect 4205 356303 5291 368194
rect 5905 356303 6297 368194
rect 4205 356077 6297 356303
rect 10662 356077 11024 370526
rect 4205 354717 11024 356077
rect 11923 364008 13867 370888
rect 11924 354717 13867 364008
rect 20967 370648 29876 370934
rect 20967 367330 21253 370648
rect 20967 364188 21151 367330
rect 23131 364188 23367 370648
rect 25245 370625 29876 370648
rect 25245 367330 25481 370625
rect 26791 368867 26961 370625
rect 29590 368867 29876 370625
rect 25347 364188 25481 367330
rect 32789 367766 34043 370890
rect 34931 367766 36169 370890
rect 32789 366455 33518 367766
rect 32789 364583 33147 366455
rect 22452 356484 22668 356499
rect 22344 355995 22668 356484
rect 21636 355706 22668 355995
rect 21636 355359 22884 355706
rect 21520 354776 22884 355359
rect 23753 354943 24039 359763
rect 27796 356892 27846 357507
rect 27796 355562 27964 356892
rect 27532 354943 27964 355562
rect 28396 354943 28682 359503
rect 35384 355716 36169 367766
rect 681431 367034 682216 379084
rect 688918 375297 689204 379857
rect 689636 379238 690068 379857
rect 689636 377908 689804 379238
rect 689754 377293 689804 377908
rect 693561 375037 693847 379857
rect 694716 379441 696080 380024
rect 694716 379094 695964 379441
rect 694932 378805 695964 379094
rect 694932 378316 695256 378805
rect 694932 378301 695148 378316
rect 684453 368345 684811 370217
rect 684082 367034 684811 368345
rect 681431 363910 682669 367034
rect 683557 363910 684811 367034
rect 692119 367470 692253 370612
rect 687724 364175 688010 365933
rect 690639 364175 690809 365933
rect 692119 364175 692355 367470
rect 687724 364152 692355 364175
rect 694233 364152 694469 370612
rect 696449 367470 696633 370612
rect 696347 364152 696633 367470
rect 687724 363866 696633 364152
rect 703733 370792 705676 380083
rect 703733 363912 705677 370792
rect 706576 378723 713395 380083
rect 706576 364274 706938 378723
rect 711303 378497 713395 378723
rect 711303 366606 711695 378497
rect 712309 366606 713395 378497
rect 711303 364274 713395 366606
rect 706576 363913 713395 364274
rect 706576 363912 711646 363913
rect 21520 354717 22303 354776
rect 23753 354657 28682 354943
rect 38135 354717 38867 355422
rect 678733 335178 679465 335883
rect 688918 335657 693847 335943
rect 695297 335824 696080 335883
rect 5954 327487 11024 327488
rect 4205 327126 11024 327487
rect 4205 324794 6297 327126
rect 4205 312903 5291 324794
rect 5905 312903 6297 324794
rect 4205 312677 6297 312903
rect 10662 312677 11024 327126
rect 4205 311317 11024 312677
rect 11923 320608 13867 327488
rect 11924 311317 13867 320608
rect 20967 327248 29876 327534
rect 20967 323930 21253 327248
rect 20967 320788 21151 323930
rect 23131 320788 23367 327248
rect 25245 327225 29876 327248
rect 25245 323930 25481 327225
rect 26791 325467 26961 327225
rect 29590 325467 29876 327225
rect 25347 320788 25481 323930
rect 32789 324366 34043 327490
rect 34931 324366 36169 327490
rect 32789 323055 33518 324366
rect 32789 321183 33147 323055
rect 22452 313084 22668 313099
rect 22344 312595 22668 313084
rect 21636 312306 22668 312595
rect 21636 311959 22884 312306
rect 21520 311376 22884 311959
rect 23753 311543 24039 316363
rect 27796 313492 27846 314107
rect 27796 312162 27964 313492
rect 27532 311543 27964 312162
rect 28396 311543 28682 316103
rect 35384 312316 36169 324366
rect 681431 322834 682216 334884
rect 688918 331097 689204 335657
rect 689636 335038 690068 335657
rect 689636 333708 689804 335038
rect 689754 333093 689804 333708
rect 693561 330837 693847 335657
rect 694716 335241 696080 335824
rect 694716 334894 695964 335241
rect 694932 334605 695964 334894
rect 694932 334116 695256 334605
rect 694932 334101 695148 334116
rect 684453 324145 684811 326017
rect 684082 322834 684811 324145
rect 681431 319710 682669 322834
rect 683557 319710 684811 322834
rect 692119 323270 692253 326412
rect 687724 319975 688010 321733
rect 690639 319975 690809 321733
rect 692119 319975 692355 323270
rect 687724 319952 692355 319975
rect 694233 319952 694469 326412
rect 696449 323270 696633 326412
rect 696347 319952 696633 323270
rect 687724 319666 696633 319952
rect 703733 326592 705676 335883
rect 703733 319712 705677 326592
rect 706576 334523 713395 335883
rect 706576 320074 706938 334523
rect 711303 334297 713395 334523
rect 711303 322406 711695 334297
rect 712309 322406 713395 334297
rect 711303 320074 713395 322406
rect 706576 319713 713395 320074
rect 706576 319712 711646 319713
rect 21520 311317 22303 311376
rect 23753 311257 28682 311543
rect 38135 311317 38867 312022
rect 678733 290978 679465 291683
rect 688918 291457 693847 291743
rect 695297 291624 696080 291683
rect 5954 284287 11024 284288
rect 4205 283926 11024 284287
rect 4205 281594 6297 283926
rect 4205 269703 5291 281594
rect 5905 269703 6297 281594
rect 4205 269477 6297 269703
rect 10662 269477 11024 283926
rect 4205 268117 11024 269477
rect 11923 277408 13867 284288
rect 11924 268117 13867 277408
rect 20967 284048 29876 284334
rect 20967 280730 21253 284048
rect 20967 277588 21151 280730
rect 23131 277588 23367 284048
rect 25245 284025 29876 284048
rect 25245 280730 25481 284025
rect 26791 282267 26961 284025
rect 29590 282267 29876 284025
rect 25347 277588 25481 280730
rect 32789 281166 34043 284290
rect 34931 281166 36169 284290
rect 32789 279855 33518 281166
rect 32789 277983 33147 279855
rect 22452 269884 22668 269899
rect 22344 269395 22668 269884
rect 21636 269106 22668 269395
rect 21636 268759 22884 269106
rect 21520 268176 22884 268759
rect 23753 268343 24039 273163
rect 27796 270292 27846 270907
rect 27796 268962 27964 270292
rect 27532 268343 27964 268962
rect 28396 268343 28682 272903
rect 35384 269116 36169 281166
rect 681431 278634 682216 290684
rect 688918 286897 689204 291457
rect 689636 290838 690068 291457
rect 689636 289508 689804 290838
rect 689754 288893 689804 289508
rect 693561 286637 693847 291457
rect 694716 291041 696080 291624
rect 694716 290694 695964 291041
rect 694932 290405 695964 290694
rect 694932 289916 695256 290405
rect 694932 289901 695148 289916
rect 684453 279945 684811 281817
rect 684082 278634 684811 279945
rect 681431 275510 682669 278634
rect 683557 275510 684811 278634
rect 692119 279070 692253 282212
rect 687724 275775 688010 277533
rect 690639 275775 690809 277533
rect 692119 275775 692355 279070
rect 687724 275752 692355 275775
rect 694233 275752 694469 282212
rect 696449 279070 696633 282212
rect 696347 275752 696633 279070
rect 687724 275466 696633 275752
rect 703733 282392 705676 291683
rect 703733 275512 705677 282392
rect 706576 290323 713395 291683
rect 706576 275874 706938 290323
rect 711303 290097 713395 290323
rect 711303 278206 711695 290097
rect 712309 278206 713395 290097
rect 711303 275874 713395 278206
rect 706576 275513 713395 275874
rect 706576 275512 711646 275513
rect 21520 268117 22303 268176
rect 23753 268057 28682 268343
rect 38135 268117 38867 268822
rect 678733 246578 679465 247283
rect 688918 247057 693847 247343
rect 695297 247224 696080 247283
rect 5954 241087 11024 241088
rect 4205 240726 11024 241087
rect 4205 238394 6297 240726
rect 4205 226503 5291 238394
rect 5905 226503 6297 238394
rect 4205 226277 6297 226503
rect 10662 226277 11024 240726
rect 4205 224917 11024 226277
rect 11923 234208 13867 241088
rect 11924 224917 13867 234208
rect 20967 240848 29876 241134
rect 20967 237530 21253 240848
rect 20967 234388 21151 237530
rect 23131 234388 23367 240848
rect 25245 240825 29876 240848
rect 25245 237530 25481 240825
rect 26791 239067 26961 240825
rect 29590 239067 29876 240825
rect 25347 234388 25481 237530
rect 32789 237966 34043 241090
rect 34931 237966 36169 241090
rect 32789 236655 33518 237966
rect 32789 234783 33147 236655
rect 22452 226684 22668 226699
rect 22344 226195 22668 226684
rect 21636 225906 22668 226195
rect 21636 225559 22884 225906
rect 21520 224976 22884 225559
rect 23753 225143 24039 229963
rect 27796 227092 27846 227707
rect 27796 225762 27964 227092
rect 27532 225143 27964 225762
rect 28396 225143 28682 229703
rect 35384 225916 36169 237966
rect 681431 234234 682216 246284
rect 688918 242497 689204 247057
rect 689636 246438 690068 247057
rect 689636 245108 689804 246438
rect 689754 244493 689804 245108
rect 693561 242237 693847 247057
rect 694716 246641 696080 247224
rect 694716 246294 695964 246641
rect 694932 246005 695964 246294
rect 694932 245516 695256 246005
rect 694932 245501 695148 245516
rect 684453 235545 684811 237417
rect 684082 234234 684811 235545
rect 681431 231110 682669 234234
rect 683557 231110 684811 234234
rect 692119 234670 692253 237812
rect 687724 231375 688010 233133
rect 690639 231375 690809 233133
rect 692119 231375 692355 234670
rect 687724 231352 692355 231375
rect 694233 231352 694469 237812
rect 696449 234670 696633 237812
rect 696347 231352 696633 234670
rect 687724 231066 696633 231352
rect 703733 237992 705676 247283
rect 703733 231112 705677 237992
rect 706576 245923 713395 247283
rect 706576 231474 706938 245923
rect 711303 245697 713395 245923
rect 711303 233806 711695 245697
rect 712309 233806 713395 245697
rect 711303 231474 713395 233806
rect 706576 231113 713395 231474
rect 706576 231112 711646 231113
rect 21520 224917 22303 224976
rect 23753 224857 28682 225143
rect 38135 224917 38867 225622
rect 678733 202378 679465 203083
rect 688918 202857 693847 203143
rect 695297 203024 696080 203083
rect 5954 197887 11024 197888
rect 4205 197526 11024 197887
rect 4205 195194 6297 197526
rect 4205 183303 5291 195194
rect 5905 183303 6297 195194
rect 4205 183077 6297 183303
rect 10662 183077 11024 197526
rect 4205 181717 11024 183077
rect 11923 191008 13867 197888
rect 11924 181717 13867 191008
rect 20967 197648 29876 197934
rect 20967 194330 21253 197648
rect 20967 191188 21151 194330
rect 23131 191188 23367 197648
rect 25245 197625 29876 197648
rect 25245 194330 25481 197625
rect 26791 195867 26961 197625
rect 29590 195867 29876 197625
rect 25347 191188 25481 194330
rect 32789 194766 34043 197890
rect 34931 194766 36169 197890
rect 32789 193455 33518 194766
rect 32789 191583 33147 193455
rect 22452 183484 22668 183499
rect 22344 182995 22668 183484
rect 21636 182706 22668 182995
rect 21636 182359 22884 182706
rect 21520 181776 22884 182359
rect 23753 181943 24039 186763
rect 27796 183892 27846 184507
rect 27796 182562 27964 183892
rect 27532 181943 27964 182562
rect 28396 181943 28682 186503
rect 35384 182716 36169 194766
rect 681431 190034 682216 202084
rect 688918 198297 689204 202857
rect 689636 202238 690068 202857
rect 689636 200908 689804 202238
rect 689754 200293 689804 200908
rect 693561 198037 693847 202857
rect 694716 202441 696080 203024
rect 694716 202094 695964 202441
rect 694932 201805 695964 202094
rect 694932 201316 695256 201805
rect 694932 201301 695148 201316
rect 684453 191345 684811 193217
rect 684082 190034 684811 191345
rect 681431 186910 682669 190034
rect 683557 186910 684811 190034
rect 692119 190470 692253 193612
rect 687724 187175 688010 188933
rect 690639 187175 690809 188933
rect 692119 187175 692355 190470
rect 687724 187152 692355 187175
rect 694233 187152 694469 193612
rect 696449 190470 696633 193612
rect 696347 187152 696633 190470
rect 687724 186866 696633 187152
rect 703733 193792 705676 203083
rect 703733 186912 705677 193792
rect 706576 201723 713395 203083
rect 706576 187274 706938 201723
rect 711303 201497 713395 201723
rect 711303 189606 711695 201497
rect 712309 189606 713395 201497
rect 711303 187274 713395 189606
rect 706576 186913 713395 187274
rect 706576 186912 711646 186913
rect 21520 181717 22303 181776
rect 23753 181657 28682 181943
rect 38135 181717 38867 182422
rect 678733 158178 679465 158883
rect 688918 158657 693847 158943
rect 695297 158824 696080 158883
rect 681431 145834 682216 157884
rect 688918 154097 689204 158657
rect 689636 158038 690068 158657
rect 689636 156708 689804 158038
rect 689754 156093 689804 156708
rect 693561 153837 693847 158657
rect 694716 158241 696080 158824
rect 694716 157894 695964 158241
rect 694932 157605 695964 157894
rect 694932 157116 695256 157605
rect 694932 157101 695148 157116
rect 684453 147145 684811 149017
rect 684082 145834 684811 147145
rect 681431 142710 682669 145834
rect 683557 142710 684811 145834
rect 692119 146270 692253 149412
rect 687724 142975 688010 144733
rect 690639 142975 690809 144733
rect 692119 142975 692355 146270
rect 687724 142952 692355 142975
rect 694233 142952 694469 149412
rect 696449 146270 696633 149412
rect 696347 142952 696633 146270
rect 687724 142666 696633 142952
rect 703733 149592 705676 158883
rect 703733 142712 705677 149592
rect 706576 157523 713395 158883
rect 706576 143074 706938 157523
rect 711303 157297 713395 157523
rect 711303 145406 711695 157297
rect 712309 145406 713395 157297
rect 711303 143074 713395 145406
rect 706576 142713 713395 143074
rect 706576 142712 711646 142713
rect 39559 112572 39863 124393
rect 678733 113778 679465 114483
rect 688918 114257 693847 114543
rect 695297 114424 696080 114483
rect 681431 101434 682216 113484
rect 688918 109697 689204 114257
rect 689636 113638 690068 114257
rect 689636 112308 689804 113638
rect 689754 111693 689804 112308
rect 693561 109437 693847 114257
rect 694716 113841 696080 114424
rect 694716 113494 695964 113841
rect 694932 113205 695964 113494
rect 694932 112716 695256 113205
rect 694932 112701 695148 112716
rect 684453 102745 684811 104617
rect 684082 101434 684811 102745
rect 681431 98310 682669 101434
rect 683557 98310 684811 101434
rect 692119 101870 692253 105012
rect 687724 98575 688010 100333
rect 690639 98575 690809 100333
rect 692119 98575 692355 101870
rect 687724 98552 692355 98575
rect 694233 98552 694469 105012
rect 696449 101870 696633 105012
rect 696347 98552 696633 101870
rect 687724 98266 696633 98552
rect 703733 105192 705676 114483
rect 703733 98312 705677 105192
rect 706576 113123 713395 114483
rect 706576 98674 706938 113123
rect 711303 112897 713395 113123
rect 711303 101006 711695 112897
rect 712309 101006 713395 112897
rect 711303 98674 713395 101006
rect 706576 98313 713395 98674
rect 706576 98312 711646 98313
rect 79607 39559 91428 39863
rect 569807 39559 581628 39863
rect 623607 39559 635428 39863
rect 201778 38135 202483 38867
rect 310378 38135 311083 38867
rect 365178 38135 365883 38867
rect 419978 38135 420683 38867
rect 474778 38135 475483 38867
rect 529578 38135 530283 38867
rect 186310 35384 201484 36169
rect 294910 35384 310084 36169
rect 349710 35384 364884 36169
rect 404510 35384 419684 36169
rect 459310 35384 474484 36169
rect 514110 35384 529284 36169
rect 186310 34931 189434 35384
rect 294910 34931 298034 35384
rect 349710 34931 352834 35384
rect 404510 34931 407634 35384
rect 459310 34931 462434 35384
rect 514110 34931 517234 35384
rect 186310 33518 189434 34043
rect 294910 33518 298034 34043
rect 349710 33518 352834 34043
rect 404510 33518 407634 34043
rect 459310 33518 462434 34043
rect 514110 33518 517234 34043
rect 186310 33147 190745 33518
rect 294910 33147 299345 33518
rect 349710 33147 354145 33518
rect 404510 33147 408945 33518
rect 459310 33147 463745 33518
rect 514110 33147 518545 33518
rect 186310 32789 192617 33147
rect 294910 32789 301217 33147
rect 349710 32789 356017 33147
rect 404510 32789 410817 33147
rect 459310 32789 465617 33147
rect 514110 32789 520417 33147
rect 186266 29590 188333 29876
rect 294866 29590 296933 29876
rect 349666 29590 351733 29876
rect 404466 29590 406533 29876
rect 459266 29590 461333 29876
rect 514066 29590 516133 29876
rect 186266 26961 186575 29590
rect 197697 28396 202543 28682
rect 202257 27964 202543 28396
rect 200308 27846 202543 27964
rect 199693 27796 202543 27846
rect 201638 27532 202543 27796
rect 186266 26791 188333 26961
rect 186266 25481 186575 26791
rect 186266 25347 193012 25481
rect 186266 25245 189870 25347
rect 186266 23367 186552 25245
rect 202257 24039 202543 27532
rect 197437 23753 202543 24039
rect 294866 26961 295175 29590
rect 306297 28396 311143 28682
rect 310857 27964 311143 28396
rect 308908 27846 311143 27964
rect 308293 27796 311143 27846
rect 310238 27532 311143 27796
rect 294866 26791 296933 26961
rect 294866 25481 295175 26791
rect 294866 25347 301612 25481
rect 294866 25245 298470 25347
rect 294866 23367 295152 25245
rect 310857 24039 311143 27532
rect 306037 23753 311143 24039
rect 349666 26961 349975 29590
rect 361097 28396 365943 28682
rect 365657 27964 365943 28396
rect 363708 27846 365943 27964
rect 363093 27796 365943 27846
rect 365038 27532 365943 27796
rect 349666 26791 351733 26961
rect 349666 25481 349975 26791
rect 349666 25347 356412 25481
rect 349666 25245 353270 25347
rect 349666 23367 349952 25245
rect 365657 24039 365943 27532
rect 360837 23753 365943 24039
rect 404466 26961 404775 29590
rect 415897 28396 420743 28682
rect 420457 27964 420743 28396
rect 418508 27846 420743 27964
rect 417893 27796 420743 27846
rect 419838 27532 420743 27796
rect 404466 26791 406533 26961
rect 404466 25481 404775 26791
rect 404466 25347 411212 25481
rect 404466 25245 408070 25347
rect 404466 23367 404752 25245
rect 420457 24039 420743 27532
rect 415637 23753 420743 24039
rect 459266 26961 459575 29590
rect 470697 28396 475543 28682
rect 475257 27964 475543 28396
rect 473308 27846 475543 27964
rect 472693 27796 475543 27846
rect 474638 27532 475543 27796
rect 459266 26791 461333 26961
rect 459266 25481 459575 26791
rect 459266 25347 466012 25481
rect 459266 25245 462870 25347
rect 459266 23367 459552 25245
rect 475257 24039 475543 27532
rect 470437 23753 475543 24039
rect 514066 26961 514375 29590
rect 525497 28396 530343 28682
rect 530057 27964 530343 28396
rect 528108 27846 530343 27964
rect 527493 27796 530343 27846
rect 529438 27532 530343 27796
rect 514066 26791 516133 26961
rect 514066 25481 514375 26791
rect 514066 25347 520812 25481
rect 514066 25245 517670 25347
rect 514066 23367 514352 25245
rect 530057 24039 530343 27532
rect 525237 23753 530343 24039
rect 186266 23131 193012 23367
rect 294866 23131 301612 23367
rect 349666 23131 356412 23367
rect 404466 23131 411212 23367
rect 459266 23131 466012 23367
rect 514066 23131 520812 23367
rect 186266 21253 186552 23131
rect 201494 22668 202424 22884
rect 200701 22452 202424 22668
rect 200716 22344 202424 22452
rect 201205 22303 202424 22344
rect 201205 21636 202483 22303
rect 201841 21520 202483 21636
rect 186266 21151 189870 21253
rect 186266 20967 193012 21151
rect 294866 21253 295152 23131
rect 310094 22668 311024 22884
rect 309301 22452 311024 22668
rect 309316 22344 311024 22452
rect 309805 22303 311024 22344
rect 309805 21636 311083 22303
rect 310441 21520 311083 21636
rect 294866 21151 298470 21253
rect 294866 20967 301612 21151
rect 349666 21253 349952 23131
rect 364894 22668 365824 22884
rect 364101 22452 365824 22668
rect 364116 22344 365824 22452
rect 364605 22303 365824 22344
rect 364605 21636 365883 22303
rect 365241 21520 365883 21636
rect 349666 21151 353270 21253
rect 349666 20967 356412 21151
rect 404466 21253 404752 23131
rect 419694 22668 420624 22884
rect 418901 22452 420624 22668
rect 418916 22344 420624 22452
rect 419405 22303 420624 22344
rect 419405 21636 420683 22303
rect 420041 21520 420683 21636
rect 404466 21151 408070 21253
rect 404466 20967 411212 21151
rect 459266 21253 459552 23131
rect 474494 22668 475424 22884
rect 473701 22452 475424 22668
rect 473716 22344 475424 22452
rect 474205 22303 475424 22344
rect 474205 21636 475483 22303
rect 474841 21520 475483 21636
rect 459266 21151 462870 21253
rect 459266 20967 466012 21151
rect 514066 21253 514352 23131
rect 529294 22668 530224 22884
rect 528501 22452 530224 22668
rect 528516 22344 530224 22452
rect 529005 22303 530224 22344
rect 529005 21636 530283 22303
rect 529641 21520 530283 21636
rect 514066 21151 517670 21253
rect 514066 20967 520812 21151
rect 132534 11924 147666 13867
rect 186312 11924 202483 13867
rect 294912 11924 311083 13867
rect 349712 11924 365883 13867
rect 404512 11924 420683 13867
rect 459312 11924 475483 13867
rect 514112 11924 530283 13867
rect 186312 11923 193192 11924
rect 294912 11923 301792 11924
rect 349712 11923 356592 11924
rect 404512 11923 411392 11924
rect 459312 11923 466192 11924
rect 514112 11923 520992 11924
rect 132476 10662 147703 11024
rect 132476 6297 132981 10662
rect 147265 6297 147703 10662
rect 132476 5958 147703 6297
rect 186312 10662 202483 11024
rect 186312 6297 186674 10662
rect 201123 6297 202483 10662
rect 186312 5954 202483 6297
rect 294912 10662 311083 11024
rect 294912 6297 295274 10662
rect 309723 6297 311083 10662
rect 294912 5954 311083 6297
rect 349712 10662 365883 11024
rect 349712 6297 350074 10662
rect 364523 6297 365883 10662
rect 349712 5954 365883 6297
rect 404512 10662 420683 11024
rect 404512 6297 404874 10662
rect 419323 6297 420683 10662
rect 404512 5954 420683 6297
rect 459312 10662 475483 11024
rect 459312 6297 459674 10662
rect 474123 6297 475483 10662
rect 459312 5954 475483 6297
rect 514112 10662 530283 11024
rect 514112 6297 514474 10662
rect 528923 6297 530283 10662
rect 514112 5954 530283 6297
rect 186313 5905 202483 5954
rect 186313 5291 189006 5905
rect 200897 5291 202483 5905
rect 186313 4205 202483 5291
rect 294913 5905 311083 5954
rect 294913 5291 297606 5905
rect 309497 5291 311083 5905
rect 294913 4205 311083 5291
rect 349713 5905 365883 5954
rect 349713 5291 352406 5905
rect 364297 5291 365883 5905
rect 349713 4205 365883 5291
rect 404513 5905 420683 5954
rect 404513 5291 407206 5905
rect 419097 5291 420683 5905
rect 404513 4205 420683 5291
rect 459313 5905 475483 5954
rect 459313 5291 462006 5905
rect 473897 5291 475483 5905
rect 459313 4205 475483 5291
rect 514113 5905 530283 5954
rect 514113 5291 516806 5905
rect 528697 5291 530283 5905
rect 514113 4205 530283 5291
<< pwell >>
rect 230099 997787 231657 1002358
rect 281499 997787 283057 1002358
rect 677787 956743 682358 958301
rect 35242 871499 39813 873057
rect 696187 861957 703671 863043
rect 696187 861140 696851 861957
rect 696591 855123 696851 861140
rect 697993 861853 703671 861957
rect 697993 855123 698310 861853
rect 696591 853832 697197 855123
rect 696591 853682 696652 853832
rect 696795 847646 697197 853832
rect 697764 852424 698310 855123
rect 697504 847646 698310 852424
rect 696795 847427 698310 847646
rect 702627 854951 703671 861853
rect 702627 849618 703463 854951
rect 702627 847427 703671 849618
rect 696795 846942 703671 847427
rect 705737 846942 706513 863058
rect 677787 816543 682358 818101
rect 11087 785142 11863 801258
rect 13929 800773 20805 801258
rect 13929 798582 14973 800773
rect 14137 793249 14973 798582
rect 13929 786347 14973 793249
rect 19290 800554 20805 800773
rect 19290 795776 20096 800554
rect 19290 793077 19836 795776
rect 20403 794368 20805 800554
rect 20948 794368 21009 794518
rect 20403 793077 21009 794368
rect 19290 786347 19607 793077
rect 13929 786243 19607 786347
rect 20749 787060 21009 793077
rect 20749 786243 21413 787060
rect 13929 785157 21413 786243
rect 696187 774557 703671 775643
rect 696187 773740 696851 774557
rect 696591 767723 696851 773740
rect 697993 774453 703671 774557
rect 697993 767723 698310 774453
rect 696591 766432 697197 767723
rect 696591 766282 696652 766432
rect 696795 760246 697197 766432
rect 697764 765024 698310 767723
rect 697504 760246 698310 765024
rect 696795 760027 698310 760246
rect 702627 767551 703671 774453
rect 702627 762218 703463 767551
rect 702627 760027 703671 762218
rect 696795 759542 703671 760027
rect 705737 759542 706513 775658
rect 11087 741942 11863 758058
rect 13929 757573 20805 758058
rect 13929 755382 14973 757573
rect 14137 750049 14973 755382
rect 13929 743147 14973 750049
rect 19290 757354 20805 757573
rect 19290 752576 20096 757354
rect 19290 749877 19836 752576
rect 20403 751168 20805 757354
rect 20948 751168 21009 751318
rect 20403 749877 21009 751168
rect 19290 743147 19607 749877
rect 13929 743043 19607 743147
rect 20749 743860 21009 749877
rect 20749 743043 21413 743860
rect 13929 741957 21413 743043
rect 696187 730157 703671 731243
rect 696187 729340 696851 730157
rect 696591 723323 696851 729340
rect 697993 730053 703671 730157
rect 697993 723323 698310 730053
rect 696591 722032 697197 723323
rect 696591 721882 696652 722032
rect 696795 715846 697197 722032
rect 697764 720624 698310 723323
rect 697504 715846 698310 720624
rect 696795 715627 698310 715846
rect 702627 723151 703671 730053
rect 702627 717818 703463 723151
rect 702627 715627 703671 717818
rect 696795 715142 703671 715627
rect 705737 715142 706513 731258
rect 11087 698742 11863 714858
rect 13929 714373 20805 714858
rect 13929 712182 14973 714373
rect 14137 706849 14973 712182
rect 13929 699947 14973 706849
rect 19290 714154 20805 714373
rect 19290 709376 20096 714154
rect 19290 706677 19836 709376
rect 20403 707968 20805 714154
rect 20948 707968 21009 708118
rect 20403 706677 21009 707968
rect 19290 699947 19607 706677
rect 13929 699843 19607 699947
rect 20749 700660 21009 706677
rect 20749 699843 21413 700660
rect 13929 698757 21413 699843
rect 696187 685957 703671 687043
rect 696187 685140 696851 685957
rect 696591 679123 696851 685140
rect 697993 685853 703671 685957
rect 697993 679123 698310 685853
rect 696591 677832 697197 679123
rect 696591 677682 696652 677832
rect 11087 655342 11863 671458
rect 13929 670973 20805 671458
rect 13929 668782 14973 670973
rect 14137 663449 14973 668782
rect 13929 656547 14973 663449
rect 19290 670754 20805 670973
rect 19290 665976 20096 670754
rect 19290 663277 19836 665976
rect 20403 664568 20805 670754
rect 696795 671646 697197 677832
rect 697764 676424 698310 679123
rect 697504 671646 698310 676424
rect 696795 671427 698310 671646
rect 702627 678951 703671 685853
rect 702627 673618 703463 678951
rect 702627 671427 703671 673618
rect 696795 670942 703671 671427
rect 705737 670942 706513 687058
rect 20948 664568 21009 664718
rect 20403 663277 21009 664568
rect 19290 656547 19607 663277
rect 13929 656443 19607 656547
rect 20749 657260 21009 663277
rect 20749 656443 21413 657260
rect 13929 655357 21413 656443
rect 696187 641757 703671 642843
rect 696187 640940 696851 641757
rect 696591 634923 696851 640940
rect 697993 641653 703671 641757
rect 697993 634923 698310 641653
rect 696591 633632 697197 634923
rect 696591 633482 696652 633632
rect 11087 612142 11863 628258
rect 13929 627773 20805 628258
rect 13929 625582 14973 627773
rect 14137 620249 14973 625582
rect 13929 613347 14973 620249
rect 19290 627554 20805 627773
rect 19290 622776 20096 627554
rect 19290 620077 19836 622776
rect 20403 621368 20805 627554
rect 696795 627446 697197 633632
rect 697764 632224 698310 634923
rect 697504 627446 698310 632224
rect 696795 627227 698310 627446
rect 702627 634751 703671 641653
rect 702627 629418 703463 634751
rect 702627 627227 703671 629418
rect 696795 626742 703671 627227
rect 705737 626742 706513 642858
rect 20948 621368 21009 621518
rect 20403 620077 21009 621368
rect 19290 613347 19607 620077
rect 13929 613243 19607 613347
rect 20749 614060 21009 620077
rect 20749 613243 21413 614060
rect 13929 612157 21413 613243
rect 696187 597357 703671 598443
rect 696187 596540 696851 597357
rect 696591 590523 696851 596540
rect 697993 597253 703671 597357
rect 697993 590523 698310 597253
rect 696591 589232 697197 590523
rect 696591 589082 696652 589232
rect 11087 568942 11863 585058
rect 13929 584573 20805 585058
rect 13929 582382 14973 584573
rect 14137 577049 14973 582382
rect 13929 570147 14973 577049
rect 19290 584354 20805 584573
rect 19290 579576 20096 584354
rect 19290 576877 19836 579576
rect 20403 578168 20805 584354
rect 696795 583046 697197 589232
rect 697764 587824 698310 590523
rect 697504 583046 698310 587824
rect 696795 582827 698310 583046
rect 702627 590351 703671 597253
rect 702627 585018 703463 590351
rect 702627 582827 703671 585018
rect 696795 582342 703671 582827
rect 705737 582342 706513 598458
rect 20948 578168 21009 578318
rect 20403 576877 21009 578168
rect 19290 570147 19607 576877
rect 13929 570043 19607 570147
rect 20749 570860 21009 576877
rect 20749 570043 21413 570860
rect 13929 568957 21413 570043
rect 11087 525742 11863 541858
rect 13929 541373 20805 541858
rect 13929 539182 14973 541373
rect 14137 533849 14973 539182
rect 13929 526947 14973 533849
rect 19290 541154 20805 541373
rect 19290 536376 20096 541154
rect 19290 533677 19836 536376
rect 20403 534968 20805 541154
rect 20948 534968 21009 535118
rect 20403 533677 21009 534968
rect 19290 526947 19607 533677
rect 13929 526843 19607 526947
rect 20749 527660 21009 533677
rect 20749 526843 21413 527660
rect 13929 525757 21413 526843
rect 696187 553157 703671 554243
rect 696187 552340 696851 553157
rect 696591 546323 696851 552340
rect 697993 553053 703671 553157
rect 697993 546323 698310 553053
rect 696591 545032 697197 546323
rect 696591 544882 696652 545032
rect 696795 538846 697197 545032
rect 697764 543624 698310 546323
rect 697504 538846 698310 543624
rect 696795 538627 698310 538846
rect 702627 546151 703671 553053
rect 702627 540818 703463 546151
rect 702627 538627 703671 540818
rect 696795 538142 703671 538627
rect 705737 538142 706513 554258
rect 677787 507743 682358 509301
rect 35242 484099 39813 485657
rect 11087 397942 11863 414058
rect 13929 413573 20805 414058
rect 13929 411382 14973 413573
rect 14137 406049 14973 411382
rect 13929 399147 14973 406049
rect 19290 413354 20805 413573
rect 19290 408576 20096 413354
rect 19290 405877 19836 408576
rect 20403 407168 20805 413354
rect 20948 407168 21009 407318
rect 20403 405877 21009 407168
rect 19290 399147 19607 405877
rect 13929 399043 19607 399147
rect 20749 399860 21009 405877
rect 20749 399043 21413 399860
rect 13929 397957 21413 399043
rect 11087 354742 11863 370858
rect 13929 370373 20805 370858
rect 13929 368182 14973 370373
rect 14137 362849 14973 368182
rect 13929 355947 14973 362849
rect 19290 370154 20805 370373
rect 19290 365376 20096 370154
rect 19290 362677 19836 365376
rect 20403 363968 20805 370154
rect 20948 363968 21009 364118
rect 20403 362677 21009 363968
rect 19290 355947 19607 362677
rect 13929 355843 19607 355947
rect 20749 356660 21009 362677
rect 20749 355843 21413 356660
rect 13929 354757 21413 355843
rect 696187 378957 703671 380043
rect 696187 378140 696851 378957
rect 696591 372123 696851 378140
rect 697993 378853 703671 378957
rect 697993 372123 698310 378853
rect 696591 370832 697197 372123
rect 696591 370682 696652 370832
rect 696795 364646 697197 370832
rect 697764 369424 698310 372123
rect 697504 364646 698310 369424
rect 696795 364427 698310 364646
rect 702627 371951 703671 378853
rect 702627 366618 703463 371951
rect 702627 364427 703671 366618
rect 696795 363942 703671 364427
rect 705737 363942 706513 380058
rect 11087 311342 11863 327458
rect 13929 326973 20805 327458
rect 13929 324782 14973 326973
rect 14137 319449 14973 324782
rect 13929 312547 14973 319449
rect 19290 326754 20805 326973
rect 19290 321976 20096 326754
rect 19290 319277 19836 321976
rect 20403 320568 20805 326754
rect 20948 320568 21009 320718
rect 20403 319277 21009 320568
rect 19290 312547 19607 319277
rect 13929 312443 19607 312547
rect 20749 313260 21009 319277
rect 20749 312443 21413 313260
rect 13929 311357 21413 312443
rect 696187 334757 703671 335843
rect 696187 333940 696851 334757
rect 696591 327923 696851 333940
rect 697993 334653 703671 334757
rect 697993 327923 698310 334653
rect 696591 326632 697197 327923
rect 696591 326482 696652 326632
rect 696795 320446 697197 326632
rect 697764 325224 698310 327923
rect 697504 320446 698310 325224
rect 696795 320227 698310 320446
rect 702627 327751 703671 334653
rect 702627 322418 703463 327751
rect 702627 320227 703671 322418
rect 696795 319742 703671 320227
rect 705737 319742 706513 335858
rect 11087 268142 11863 284258
rect 13929 283773 20805 284258
rect 13929 281582 14973 283773
rect 14137 276249 14973 281582
rect 13929 269347 14973 276249
rect 19290 283554 20805 283773
rect 19290 278776 20096 283554
rect 19290 276077 19836 278776
rect 20403 277368 20805 283554
rect 20948 277368 21009 277518
rect 20403 276077 21009 277368
rect 19290 269347 19607 276077
rect 13929 269243 19607 269347
rect 20749 270060 21009 276077
rect 20749 269243 21413 270060
rect 13929 268157 21413 269243
rect 696187 290557 703671 291643
rect 696187 289740 696851 290557
rect 696591 283723 696851 289740
rect 697993 290453 703671 290557
rect 697993 283723 698310 290453
rect 696591 282432 697197 283723
rect 696591 282282 696652 282432
rect 696795 276246 697197 282432
rect 697764 281024 698310 283723
rect 697504 276246 698310 281024
rect 696795 276027 698310 276246
rect 702627 283551 703671 290453
rect 702627 278218 703463 283551
rect 702627 276027 703671 278218
rect 696795 275542 703671 276027
rect 705737 275542 706513 291658
rect 11087 224942 11863 241058
rect 13929 240573 20805 241058
rect 13929 238382 14973 240573
rect 14137 233049 14973 238382
rect 13929 226147 14973 233049
rect 19290 240354 20805 240573
rect 19290 235576 20096 240354
rect 19290 232877 19836 235576
rect 20403 234168 20805 240354
rect 20948 234168 21009 234318
rect 20403 232877 21009 234168
rect 19290 226147 19607 232877
rect 13929 226043 19607 226147
rect 20749 226860 21009 232877
rect 20749 226043 21413 226860
rect 13929 224957 21413 226043
rect 696187 246157 703671 247243
rect 696187 245340 696851 246157
rect 696591 239323 696851 245340
rect 697993 246053 703671 246157
rect 697993 239323 698310 246053
rect 696591 238032 697197 239323
rect 696591 237882 696652 238032
rect 696795 231846 697197 238032
rect 697764 236624 698310 239323
rect 697504 231846 698310 236624
rect 696795 231627 698310 231846
rect 702627 239151 703671 246053
rect 702627 233818 703463 239151
rect 702627 231627 703671 233818
rect 696795 231142 703671 231627
rect 705737 231142 706513 247258
rect 11087 181742 11863 197858
rect 13929 197373 20805 197858
rect 13929 195182 14973 197373
rect 14137 189849 14973 195182
rect 13929 182947 14973 189849
rect 19290 197154 20805 197373
rect 19290 192376 20096 197154
rect 19290 189677 19836 192376
rect 20403 190968 20805 197154
rect 20948 190968 21009 191118
rect 20403 189677 21009 190968
rect 19290 182947 19607 189677
rect 13929 182843 19607 182947
rect 20749 183660 21009 189677
rect 20749 182843 21413 183660
rect 13929 181757 21413 182843
rect 696187 201957 703671 203043
rect 696187 201140 696851 201957
rect 696591 195123 696851 201140
rect 697993 201853 703671 201957
rect 697993 195123 698310 201853
rect 696591 193832 697197 195123
rect 696591 193682 696652 193832
rect 696795 187646 697197 193832
rect 697764 192424 698310 195123
rect 697504 187646 698310 192424
rect 696795 187427 698310 187646
rect 702627 194951 703671 201853
rect 702627 189618 703463 194951
rect 702627 187427 703671 189618
rect 696795 186942 703671 187427
rect 705737 186942 706513 203058
rect 696187 157757 703671 158843
rect 696187 156940 696851 157757
rect 696591 150923 696851 156940
rect 697993 157653 703671 157757
rect 697993 150923 698310 157653
rect 696591 149632 697197 150923
rect 696591 149482 696652 149632
rect 696795 143446 697197 149632
rect 697764 148224 698310 150923
rect 697504 143446 698310 148224
rect 696795 143227 698310 143446
rect 702627 150751 703671 157653
rect 702627 145418 703463 150751
rect 702627 143227 703671 145418
rect 696795 142742 703671 143227
rect 705737 142742 706513 158858
rect 35242 110899 39813 112457
rect 696187 113357 703671 114443
rect 696187 112540 696851 113357
rect 696591 106523 696851 112540
rect 697993 113253 703671 113357
rect 697993 106523 698310 113253
rect 696591 105232 697197 106523
rect 696591 105082 696652 105232
rect 696795 99046 697197 105232
rect 697764 103824 698310 106523
rect 697504 99046 698310 103824
rect 696795 98827 698310 99046
rect 702627 106351 703671 113253
rect 702627 101018 703463 106351
rect 702627 98827 703671 101018
rect 696795 98342 703671 98827
rect 705737 98342 706513 114458
rect 635543 35242 637101 39813
rect 200540 21009 202443 21413
rect 193082 20948 202443 21009
rect 309140 21009 311043 21413
rect 301682 20948 311043 21009
rect 363940 21009 365843 21413
rect 356482 20948 365843 21009
rect 418740 21009 420643 21413
rect 411282 20948 420643 21009
rect 473540 21009 475443 21413
rect 466082 20948 475443 21009
rect 528340 21009 530243 21413
rect 520882 20948 530243 21009
rect 193232 20805 202443 20948
rect 301832 20805 311043 20948
rect 356632 20805 365843 20948
rect 411432 20805 420643 20948
rect 466232 20805 475443 20948
rect 521032 20805 530243 20948
rect 186342 20749 202443 20805
rect 135906 20653 147626 20654
rect 132574 20401 147626 20653
rect 132574 20154 133214 20401
rect 135906 20154 147626 20401
rect 132574 19495 147626 20154
rect 132574 15173 132888 19495
rect 147313 15173 147626 19495
rect 132574 14137 147626 15173
rect 132574 13929 135218 14137
rect 139250 13929 147626 14137
rect 186342 20403 194523 20749
rect 186342 20096 187046 20403
rect 186342 19836 191824 20096
rect 186342 19607 194523 19836
rect 201357 19607 202443 20749
rect 186342 19290 202443 19607
rect 186342 14973 186827 19290
rect 201253 14973 202443 19290
rect 186342 14137 202443 14973
rect 186342 13929 189018 14137
rect 194351 13929 202443 14137
rect 294942 20749 311043 20805
rect 294942 20403 303123 20749
rect 294942 20096 295646 20403
rect 294942 19836 300424 20096
rect 294942 19607 303123 19836
rect 309957 19607 311043 20749
rect 294942 19290 311043 19607
rect 294942 14973 295427 19290
rect 309853 14973 311043 19290
rect 294942 14137 311043 14973
rect 294942 13929 297618 14137
rect 302951 13929 311043 14137
rect 349742 20749 365843 20805
rect 349742 20403 357923 20749
rect 349742 20096 350446 20403
rect 349742 19836 355224 20096
rect 349742 19607 357923 19836
rect 364757 19607 365843 20749
rect 349742 19290 365843 19607
rect 349742 14973 350227 19290
rect 364653 14973 365843 19290
rect 349742 14137 365843 14973
rect 349742 13929 352418 14137
rect 357751 13929 365843 14137
rect 404542 20749 420643 20805
rect 404542 20403 412723 20749
rect 404542 20096 405246 20403
rect 404542 19836 410024 20096
rect 404542 19607 412723 19836
rect 419557 19607 420643 20749
rect 404542 19290 420643 19607
rect 404542 14973 405027 19290
rect 419453 14973 420643 19290
rect 404542 14137 420643 14973
rect 404542 13929 407218 14137
rect 412551 13929 420643 14137
rect 459342 20749 475443 20805
rect 459342 20403 467523 20749
rect 459342 20096 460046 20403
rect 459342 19836 464824 20096
rect 459342 19607 467523 19836
rect 474357 19607 475443 20749
rect 459342 19290 475443 19607
rect 459342 14973 459827 19290
rect 474253 14973 475443 19290
rect 459342 14137 475443 14973
rect 459342 13929 462018 14137
rect 467351 13929 475443 14137
rect 514142 20749 530243 20805
rect 514142 20403 522323 20749
rect 514142 20096 514846 20403
rect 514142 19836 519624 20096
rect 514142 19607 522323 19836
rect 529157 19607 530243 20749
rect 514142 19290 530243 19607
rect 514142 14973 514627 19290
rect 529053 14973 530243 19290
rect 514142 14137 530243 14973
rect 514142 13929 516818 14137
rect 522151 13929 530243 14137
rect 132542 11087 147658 11863
rect 186342 11087 202458 11863
rect 294942 11087 311058 11863
rect 349742 11087 365858 11863
rect 404542 11087 420658 11863
rect 459342 11087 475458 11863
rect 514142 11087 530258 11863
<< obsli1 >>
rect 75581 1007253 89409 1033820
rect 123581 1007253 137409 1033820
rect 171581 1007253 185409 1033820
rect 229522 998007 243971 1037539
rect 280922 998007 295371 1037539
rect 339614 998007 353955 1037539
rect 425381 1007253 439209 1033820
rect 474781 1007253 488609 1033820
rect 526381 1007253 540209 1033820
rect 575814 998007 590155 1037539
rect 627581 1007253 641409 1033820
rect 229522 997813 231631 998007
rect 231807 997984 232009 998007
rect 243346 997984 243536 998007
rect 231807 997794 243536 997984
rect 280922 997813 283031 998007
rect 283207 997984 283409 998007
rect 294746 997984 294936 998007
rect 283207 997794 294936 997984
rect 341813 997978 342009 998007
rect 353352 997978 353530 998007
rect 341813 997800 353530 997978
rect 578013 997978 578209 998007
rect 589552 997978 589730 998007
rect 578013 997800 589730 997978
rect 3780 955781 30347 969609
rect 677813 956769 717539 958878
rect 678007 956593 717539 956769
rect 677794 956391 717539 956593
rect 677794 945054 677984 956391
rect 678007 945054 717539 956391
rect 677794 944864 717539 945054
rect 678007 944429 717539 944864
rect 44 913048 39396 927951
rect 678204 891449 717556 906352
rect 61 884936 39593 885371
rect 61 884746 39806 884936
rect 61 873409 39593 884746
rect 39616 873409 39806 884746
rect 61 873207 39806 873409
rect 61 873031 39593 873207
rect 61 870922 39787 873031
rect 696779 863017 703644 863023
rect 703855 863017 705630 863023
rect 678799 863000 679399 863017
rect 689044 863000 693721 863017
rect 695363 863000 696014 863017
rect 696213 863000 703645 863017
rect 703799 863000 705630 863017
rect 705763 863000 706487 863032
rect 706631 863017 711618 863023
rect 706631 863000 713329 863017
rect 677646 847000 717541 863000
rect 681497 846976 682603 847000
rect 683623 846976 684745 847000
rect 687850 846983 696516 847000
rect 696821 846968 703645 847000
rect 703799 846983 705611 847000
rect 705763 846968 706487 847000
rect 706643 846979 713329 847000
rect 61 842530 39593 842955
rect 61 842352 39800 842530
rect 61 831009 39593 842352
rect 39622 831009 39800 842352
rect 61 830813 39800 831009
rect 61 828614 39593 830813
rect 677813 816569 717539 818678
rect 678007 816393 717539 816569
rect 677794 816191 717539 816393
rect 677794 804854 677984 816191
rect 678007 804854 717539 816191
rect 677794 804664 717539 804854
rect 678007 804229 717539 804664
rect 4271 801200 10957 801221
rect 11113 801200 11837 801232
rect 11989 801200 13801 801217
rect 13955 801200 20779 801232
rect 21084 801200 29750 801217
rect 32855 801200 33977 801224
rect 34997 801200 36103 801224
rect 59 785200 39954 801200
rect 4271 785183 10969 785200
rect 5982 785177 10969 785183
rect 11113 785168 11837 785200
rect 11970 785183 13801 785200
rect 13955 785183 21387 785200
rect 21586 785183 22237 785200
rect 23879 785183 28556 785200
rect 38201 785183 38801 785200
rect 11970 785177 13745 785183
rect 13956 785177 20821 785183
rect 696779 775617 703644 775623
rect 703855 775617 705630 775623
rect 678799 775600 679399 775617
rect 689044 775600 693721 775617
rect 695363 775600 696014 775617
rect 696213 775600 703645 775617
rect 703799 775600 705630 775617
rect 705763 775600 706487 775632
rect 706631 775617 711618 775623
rect 706631 775600 713329 775617
rect 677646 759600 717541 775600
rect 681497 759576 682603 759600
rect 683623 759576 684745 759600
rect 687850 759583 696516 759600
rect 696821 759568 703645 759600
rect 703799 759583 705611 759600
rect 705763 759568 706487 759600
rect 706643 759579 713329 759600
rect 4271 758000 10957 758021
rect 11113 758000 11837 758032
rect 11989 758000 13801 758017
rect 13955 758000 20779 758032
rect 21084 758000 29750 758017
rect 32855 758000 33977 758024
rect 34997 758000 36103 758024
rect 59 742000 39954 758000
rect 4271 741983 10969 742000
rect 5982 741977 10969 741983
rect 11113 741968 11837 742000
rect 11970 741983 13801 742000
rect 13955 741983 21387 742000
rect 21586 741983 22237 742000
rect 23879 741983 28556 742000
rect 38201 741983 38801 742000
rect 11970 741977 13745 741983
rect 13956 741977 20821 741983
rect 696779 731217 703644 731223
rect 703855 731217 705630 731223
rect 678799 731200 679399 731217
rect 689044 731200 693721 731217
rect 695363 731200 696014 731217
rect 696213 731200 703645 731217
rect 703799 731200 705630 731217
rect 705763 731200 706487 731232
rect 706631 731217 711618 731223
rect 706631 731200 713329 731217
rect 677646 715200 717541 731200
rect 681497 715176 682603 715200
rect 683623 715176 684745 715200
rect 687850 715183 696516 715200
rect 696821 715168 703645 715200
rect 703799 715183 705611 715200
rect 705763 715168 706487 715200
rect 706643 715179 713329 715200
rect 4271 714800 10957 714821
rect 11113 714800 11837 714832
rect 11989 714800 13801 714817
rect 13955 714800 20779 714832
rect 21084 714800 29750 714817
rect 32855 714800 33977 714824
rect 34997 714800 36103 714824
rect 59 698800 39954 714800
rect 4271 698783 10969 698800
rect 5982 698777 10969 698783
rect 11113 698768 11837 698800
rect 11970 698783 13801 698800
rect 13955 698783 21387 698800
rect 21586 698783 22237 698800
rect 23879 698783 28556 698800
rect 38201 698783 38801 698800
rect 11970 698777 13745 698783
rect 13956 698777 20821 698783
rect 696779 687017 703644 687023
rect 703855 687017 705630 687023
rect 678799 687000 679399 687017
rect 689044 687000 693721 687017
rect 695363 687000 696014 687017
rect 696213 687000 703645 687017
rect 703799 687000 705630 687017
rect 705763 687000 706487 687032
rect 706631 687017 711618 687023
rect 706631 687000 713329 687017
rect 4271 671400 10957 671421
rect 11113 671400 11837 671432
rect 11989 671400 13801 671417
rect 13955 671400 20779 671432
rect 21084 671400 29750 671417
rect 32855 671400 33977 671424
rect 34997 671400 36103 671424
rect 59 655400 39954 671400
rect 677646 671000 717541 687000
rect 681497 670976 682603 671000
rect 683623 670976 684745 671000
rect 687850 670983 696516 671000
rect 696821 670968 703645 671000
rect 703799 670983 705611 671000
rect 705763 670968 706487 671000
rect 706643 670979 713329 671000
rect 4271 655383 10969 655400
rect 5982 655377 10969 655383
rect 11113 655368 11837 655400
rect 11970 655383 13801 655400
rect 13955 655383 21387 655400
rect 21586 655383 22237 655400
rect 23879 655383 28556 655400
rect 38201 655383 38801 655400
rect 11970 655377 13745 655383
rect 13956 655377 20821 655383
rect 696779 642817 703644 642823
rect 703855 642817 705630 642823
rect 678799 642800 679399 642817
rect 689044 642800 693721 642817
rect 695363 642800 696014 642817
rect 696213 642800 703645 642817
rect 703799 642800 705630 642817
rect 705763 642800 706487 642832
rect 706631 642817 711618 642823
rect 706631 642800 713329 642817
rect 4271 628200 10957 628221
rect 11113 628200 11837 628232
rect 11989 628200 13801 628217
rect 13955 628200 20779 628232
rect 21084 628200 29750 628217
rect 32855 628200 33977 628224
rect 34997 628200 36103 628224
rect 59 612200 39954 628200
rect 677646 626800 717541 642800
rect 681497 626776 682603 626800
rect 683623 626776 684745 626800
rect 687850 626783 696516 626800
rect 696821 626768 703645 626800
rect 703799 626783 705611 626800
rect 705763 626768 706487 626800
rect 706643 626779 713329 626800
rect 4271 612183 10969 612200
rect 5982 612177 10969 612183
rect 11113 612168 11837 612200
rect 11970 612183 13801 612200
rect 13955 612183 21387 612200
rect 21586 612183 22237 612200
rect 23879 612183 28556 612200
rect 38201 612183 38801 612200
rect 11970 612177 13745 612183
rect 13956 612177 20821 612183
rect 696779 598417 703644 598423
rect 703855 598417 705630 598423
rect 678799 598400 679399 598417
rect 689044 598400 693721 598417
rect 695363 598400 696014 598417
rect 696213 598400 703645 598417
rect 703799 598400 705630 598417
rect 705763 598400 706487 598432
rect 706631 598417 711618 598423
rect 706631 598400 713329 598417
rect 4271 585000 10957 585021
rect 11113 585000 11837 585032
rect 11989 585000 13801 585017
rect 13955 585000 20779 585032
rect 21084 585000 29750 585017
rect 32855 585000 33977 585024
rect 34997 585000 36103 585024
rect 59 569000 39954 585000
rect 677646 582400 717541 598400
rect 681497 582376 682603 582400
rect 683623 582376 684745 582400
rect 687850 582383 696516 582400
rect 696821 582368 703645 582400
rect 703799 582383 705611 582400
rect 705763 582368 706487 582400
rect 706643 582379 713329 582400
rect 4271 568983 10969 569000
rect 5982 568977 10969 568983
rect 11113 568968 11837 569000
rect 11970 568983 13801 569000
rect 13955 568983 21387 569000
rect 21586 568983 22237 569000
rect 23879 568983 28556 569000
rect 38201 568983 38801 569000
rect 11970 568977 13745 568983
rect 13956 568977 20821 568983
rect 696779 554217 703644 554223
rect 703855 554217 705630 554223
rect 678799 554200 679399 554217
rect 689044 554200 693721 554217
rect 695363 554200 696014 554217
rect 696213 554200 703645 554217
rect 703799 554200 705630 554217
rect 705763 554200 706487 554232
rect 706631 554217 711618 554223
rect 706631 554200 713329 554217
rect 4271 541800 10957 541821
rect 11113 541800 11837 541832
rect 11989 541800 13801 541817
rect 13955 541800 20779 541832
rect 21084 541800 29750 541817
rect 32855 541800 33977 541824
rect 34997 541800 36103 541824
rect 59 525800 39954 541800
rect 677646 538200 717541 554200
rect 681497 538176 682603 538200
rect 683623 538176 684745 538200
rect 687850 538183 696516 538200
rect 696821 538168 703645 538200
rect 703799 538183 705611 538200
rect 705763 538168 706487 538200
rect 706643 538179 713329 538200
rect 4271 525783 10969 525800
rect 5982 525777 10969 525783
rect 11113 525768 11837 525800
rect 11970 525783 13801 525800
rect 13955 525783 21387 525800
rect 21586 525783 22237 525800
rect 23879 525783 28556 525800
rect 38201 525783 38801 525800
rect 11970 525777 13745 525783
rect 13956 525777 20821 525783
rect 677813 507769 717539 509878
rect 678007 507593 717539 507769
rect 677794 507391 717539 507593
rect 61 497536 39593 497971
rect 61 497346 39806 497536
rect 61 486009 39593 497346
rect 39616 486009 39806 497346
rect 677794 496054 677984 507391
rect 678007 496054 717539 507391
rect 677794 495864 717539 496054
rect 678007 495429 717539 495864
rect 61 485807 39806 486009
rect 61 485631 39593 485807
rect 61 483522 39787 485631
rect 44 441248 39396 456151
rect 678204 451649 717556 466552
rect 678007 420987 717539 423186
rect 677800 420791 717539 420987
rect 4271 414000 10957 414021
rect 11113 414000 11837 414032
rect 11989 414000 13801 414017
rect 13955 414000 20779 414032
rect 21084 414000 29750 414017
rect 32855 414000 33977 414024
rect 34997 414000 36103 414024
rect 59 398000 39954 414000
rect 677800 409448 677978 420791
rect 678007 409448 717539 420791
rect 677800 409270 717539 409448
rect 678007 408845 717539 409270
rect 4271 397983 10969 398000
rect 5982 397977 10969 397983
rect 11113 397968 11837 398000
rect 11970 397983 13801 398000
rect 13955 397983 21387 398000
rect 21586 397983 22237 398000
rect 23879 397983 28556 398000
rect 38201 397983 38801 398000
rect 11970 397977 13745 397983
rect 13956 397977 20821 397983
rect 696779 380017 703644 380023
rect 703855 380017 705630 380023
rect 678799 380000 679399 380017
rect 689044 380000 693721 380017
rect 695363 380000 696014 380017
rect 696213 380000 703645 380017
rect 703799 380000 705630 380017
rect 705763 380000 706487 380032
rect 706631 380017 711618 380023
rect 706631 380000 713329 380017
rect 4271 370800 10957 370821
rect 11113 370800 11837 370832
rect 11989 370800 13801 370817
rect 13955 370800 20779 370832
rect 21084 370800 29750 370817
rect 32855 370800 33977 370824
rect 34997 370800 36103 370824
rect 59 354800 39954 370800
rect 677646 364000 717541 380000
rect 681497 363976 682603 364000
rect 683623 363976 684745 364000
rect 687850 363983 696516 364000
rect 696821 363968 703645 364000
rect 703799 363983 705611 364000
rect 705763 363968 706487 364000
rect 706643 363979 713329 364000
rect 4271 354783 10969 354800
rect 5982 354777 10969 354783
rect 11113 354768 11837 354800
rect 11970 354783 13801 354800
rect 13955 354783 21387 354800
rect 21586 354783 22237 354800
rect 23879 354783 28556 354800
rect 38201 354783 38801 354800
rect 11970 354777 13745 354783
rect 13956 354777 20821 354783
rect 696779 335817 703644 335823
rect 703855 335817 705630 335823
rect 678799 335800 679399 335817
rect 689044 335800 693721 335817
rect 695363 335800 696014 335817
rect 696213 335800 703645 335817
rect 703799 335800 705630 335817
rect 705763 335800 706487 335832
rect 706631 335817 711618 335823
rect 706631 335800 713329 335817
rect 4271 327400 10957 327421
rect 11113 327400 11837 327432
rect 11989 327400 13801 327417
rect 13955 327400 20779 327432
rect 21084 327400 29750 327417
rect 32855 327400 33977 327424
rect 34997 327400 36103 327424
rect 59 311400 39954 327400
rect 677646 319800 717541 335800
rect 681497 319776 682603 319800
rect 683623 319776 684745 319800
rect 687850 319783 696516 319800
rect 696821 319768 703645 319800
rect 703799 319783 705611 319800
rect 705763 319768 706487 319800
rect 706643 319779 713329 319800
rect 4271 311383 10969 311400
rect 5982 311377 10969 311383
rect 11113 311368 11837 311400
rect 11970 311383 13801 311400
rect 13955 311383 21387 311400
rect 21586 311383 22237 311400
rect 23879 311383 28556 311400
rect 38201 311383 38801 311400
rect 11970 311377 13745 311383
rect 13956 311377 20821 311383
rect 696779 291617 703644 291623
rect 703855 291617 705630 291623
rect 678799 291600 679399 291617
rect 689044 291600 693721 291617
rect 695363 291600 696014 291617
rect 696213 291600 703645 291617
rect 703799 291600 705630 291617
rect 705763 291600 706487 291632
rect 706631 291617 711618 291623
rect 706631 291600 713329 291617
rect 4271 284200 10957 284221
rect 11113 284200 11837 284232
rect 11989 284200 13801 284217
rect 13955 284200 20779 284232
rect 21084 284200 29750 284217
rect 32855 284200 33977 284224
rect 34997 284200 36103 284224
rect 59 268200 39954 284200
rect 677646 275600 717541 291600
rect 681497 275576 682603 275600
rect 683623 275576 684745 275600
rect 687850 275583 696516 275600
rect 696821 275568 703645 275600
rect 703799 275583 705611 275600
rect 705763 275568 706487 275600
rect 706643 275579 713329 275600
rect 4271 268183 10969 268200
rect 5982 268177 10969 268183
rect 11113 268168 11837 268200
rect 11970 268183 13801 268200
rect 13955 268183 21387 268200
rect 21586 268183 22237 268200
rect 23879 268183 28556 268200
rect 38201 268183 38801 268200
rect 11970 268177 13745 268183
rect 13956 268177 20821 268183
rect 696779 247217 703644 247223
rect 703855 247217 705630 247223
rect 678799 247200 679399 247217
rect 689044 247200 693721 247217
rect 695363 247200 696014 247217
rect 696213 247200 703645 247217
rect 703799 247200 705630 247217
rect 705763 247200 706487 247232
rect 706631 247217 711618 247223
rect 706631 247200 713329 247217
rect 4271 241000 10957 241021
rect 11113 241000 11837 241032
rect 11989 241000 13801 241017
rect 13955 241000 20779 241032
rect 21084 241000 29750 241017
rect 32855 241000 33977 241024
rect 34997 241000 36103 241024
rect 59 225000 39954 241000
rect 677646 231200 717541 247200
rect 681497 231176 682603 231200
rect 683623 231176 684745 231200
rect 687850 231183 696516 231200
rect 696821 231168 703645 231200
rect 703799 231183 705611 231200
rect 705763 231168 706487 231200
rect 706643 231179 713329 231200
rect 4271 224983 10969 225000
rect 5982 224977 10969 224983
rect 11113 224968 11837 225000
rect 11970 224983 13801 225000
rect 13955 224983 21387 225000
rect 21586 224983 22237 225000
rect 23879 224983 28556 225000
rect 38201 224983 38801 225000
rect 11970 224977 13745 224983
rect 13956 224977 20821 224983
rect 696779 203017 703644 203023
rect 703855 203017 705630 203023
rect 678799 203000 679399 203017
rect 689044 203000 693721 203017
rect 695363 203000 696014 203017
rect 696213 203000 703645 203017
rect 703799 203000 705630 203017
rect 705763 203000 706487 203032
rect 706631 203017 711618 203023
rect 706631 203000 713329 203017
rect 4271 197800 10957 197821
rect 11113 197800 11837 197832
rect 11989 197800 13801 197817
rect 13955 197800 20779 197832
rect 21084 197800 29750 197817
rect 32855 197800 33977 197824
rect 34997 197800 36103 197824
rect 59 181800 39954 197800
rect 677646 187000 717541 203000
rect 681497 186976 682603 187000
rect 683623 186976 684745 187000
rect 687850 186983 696516 187000
rect 696821 186968 703645 187000
rect 703799 186983 705611 187000
rect 705763 186968 706487 187000
rect 706643 186979 713329 187000
rect 4271 181783 10969 181800
rect 5982 181777 10969 181783
rect 11113 181768 11837 181800
rect 11970 181783 13801 181800
rect 13955 181783 21387 181800
rect 21586 181783 22237 181800
rect 23879 181783 28556 181800
rect 38201 181783 38801 181800
rect 11970 181777 13745 181783
rect 13956 181777 20821 181783
rect 696779 158817 703644 158823
rect 703855 158817 705630 158823
rect 678799 158800 679399 158817
rect 689044 158800 693721 158817
rect 695363 158800 696014 158817
rect 696213 158800 703645 158817
rect 703799 158800 705630 158817
rect 705763 158800 706487 158832
rect 706631 158817 711618 158823
rect 706631 158800 713329 158817
rect 677646 142800 717541 158800
rect 681497 142776 682603 142800
rect 683623 142776 684745 142800
rect 687850 142783 696516 142800
rect 696821 142768 703645 142800
rect 703799 142783 705611 142800
rect 705763 142768 706487 142800
rect 706643 142779 713329 142800
rect 61 124336 39593 124771
rect 61 124146 39806 124336
rect 61 112809 39593 124146
rect 39616 112809 39806 124146
rect 696779 114417 703644 114423
rect 703855 114417 705630 114423
rect 678799 114400 679399 114417
rect 689044 114400 693721 114417
rect 695363 114400 696014 114417
rect 696213 114400 703645 114417
rect 703799 114400 705630 114417
rect 705763 114400 706487 114432
rect 706631 114417 711618 114423
rect 706631 114400 713329 114417
rect 61 112607 39806 112809
rect 61 112431 39593 112607
rect 61 110322 39787 112431
rect 677646 98400 717541 114400
rect 681497 98376 682603 98400
rect 683623 98376 684745 98400
rect 687850 98383 696516 98400
rect 696821 98368 703645 98400
rect 703799 98383 705611 98400
rect 705763 98368 706487 98400
rect 706643 98379 713329 98400
rect 44 68048 39396 82951
rect 79670 39622 91387 39800
rect 79670 39593 79848 39622
rect 91191 39593 91387 39622
rect 79245 61 93586 39593
rect 132600 19721 147600 39963
rect 186400 38801 202400 39954
rect 186400 38201 202417 38801
rect 186400 36103 202400 38201
rect 186376 34997 202400 36103
rect 186400 33977 202400 34997
rect 186376 32855 202400 33977
rect 186400 29750 202400 32855
rect 186383 28556 202400 29750
rect 186383 23879 202417 28556
rect 186383 22237 202400 23879
rect 186383 21586 202417 22237
rect 186383 21387 202400 21586
rect 186383 21084 202417 21387
rect 186400 20821 202417 21084
rect 186400 20779 202423 20821
rect 132600 13955 147653 19721
rect 186368 13956 202423 20779
rect 186368 13955 202417 13956
rect 132600 11837 147600 13955
rect 186400 13801 202400 13955
rect 186383 13745 202417 13801
rect 186383 11989 202423 13745
rect 186400 11970 202423 11989
rect 186400 11837 202400 11970
rect 132568 11113 147632 11837
rect 186368 11113 202432 11837
rect 132600 156 147600 11113
rect 186400 10969 202400 11113
rect 186400 10957 202423 10969
rect 186379 5982 202423 10957
rect 186379 4271 202417 5982
rect 186400 59 202400 4271
rect 241249 44 256152 39396
rect 295000 38801 311000 39954
rect 349800 38801 365800 39954
rect 404600 38801 420600 39954
rect 459400 38801 475400 39954
rect 514200 38801 530200 39954
rect 569870 39622 581587 39800
rect 569870 39593 570048 39622
rect 581391 39593 581587 39622
rect 623664 39616 635393 39806
rect 623664 39593 623854 39616
rect 635191 39593 635393 39616
rect 635569 39593 637678 39787
rect 295000 38201 311017 38801
rect 349800 38201 365817 38801
rect 404600 38201 420617 38801
rect 459400 38201 475417 38801
rect 514200 38201 530217 38801
rect 295000 36103 311000 38201
rect 349800 36103 365800 38201
rect 404600 36103 420600 38201
rect 459400 36103 475400 38201
rect 514200 36103 530200 38201
rect 294976 34997 311000 36103
rect 349776 34997 365800 36103
rect 404576 34997 420600 36103
rect 459376 34997 475400 36103
rect 514176 34997 530200 36103
rect 295000 33977 311000 34997
rect 349800 33977 365800 34997
rect 404600 33977 420600 34997
rect 459400 33977 475400 34997
rect 514200 33977 530200 34997
rect 294976 32855 311000 33977
rect 349776 32855 365800 33977
rect 404576 32855 420600 33977
rect 459376 32855 475400 33977
rect 514176 32855 530200 33977
rect 295000 29750 311000 32855
rect 349800 29750 365800 32855
rect 404600 29750 420600 32855
rect 459400 29750 475400 32855
rect 514200 29750 530200 32855
rect 294983 28556 311000 29750
rect 349783 28556 365800 29750
rect 404583 28556 420600 29750
rect 459383 28556 475400 29750
rect 514183 28556 530200 29750
rect 294983 23879 311017 28556
rect 349783 23879 365817 28556
rect 404583 23879 420617 28556
rect 459383 23879 475417 28556
rect 514183 23879 530217 28556
rect 294983 22237 311000 23879
rect 349783 22237 365800 23879
rect 404583 22237 420600 23879
rect 459383 22237 475400 23879
rect 514183 22237 530200 23879
rect 294983 21586 311017 22237
rect 349783 21586 365817 22237
rect 404583 21586 420617 22237
rect 459383 21586 475417 22237
rect 514183 21586 530217 22237
rect 294983 21387 311000 21586
rect 349783 21387 365800 21586
rect 404583 21387 420600 21586
rect 459383 21387 475400 21586
rect 514183 21387 530200 21586
rect 294983 21084 311017 21387
rect 349783 21084 365817 21387
rect 404583 21084 420617 21387
rect 459383 21084 475417 21387
rect 514183 21084 530217 21387
rect 295000 20821 311017 21084
rect 349800 20821 365817 21084
rect 404600 20821 420617 21084
rect 459400 20821 475417 21084
rect 514200 20821 530217 21084
rect 295000 20779 311023 20821
rect 349800 20779 365823 20821
rect 404600 20779 420623 20821
rect 459400 20779 475423 20821
rect 514200 20779 530223 20821
rect 294968 13956 311023 20779
rect 349768 13956 365823 20779
rect 404568 13956 420623 20779
rect 459368 13956 475423 20779
rect 514168 13956 530223 20779
rect 294968 13955 311017 13956
rect 349768 13955 365817 13956
rect 404568 13955 420617 13956
rect 459368 13955 475417 13956
rect 514168 13955 530217 13956
rect 295000 13801 311000 13955
rect 349800 13801 365800 13955
rect 404600 13801 420600 13955
rect 459400 13801 475400 13955
rect 514200 13801 530200 13955
rect 294983 13745 311017 13801
rect 349783 13745 365817 13801
rect 404583 13745 420617 13801
rect 459383 13745 475417 13801
rect 514183 13745 530217 13801
rect 294983 11989 311023 13745
rect 349783 11989 365823 13745
rect 404583 11989 420623 13745
rect 459383 11989 475423 13745
rect 514183 11989 530223 13745
rect 295000 11970 311023 11989
rect 349800 11970 365823 11989
rect 404600 11970 420623 11989
rect 459400 11970 475423 11989
rect 514200 11970 530223 11989
rect 295000 11837 311000 11970
rect 349800 11837 365800 11970
rect 404600 11837 420600 11970
rect 459400 11837 475400 11970
rect 514200 11837 530200 11970
rect 294968 11113 311032 11837
rect 349768 11113 365832 11837
rect 404568 11113 420632 11837
rect 459368 11113 475432 11837
rect 514168 11113 530232 11837
rect 295000 10969 311000 11113
rect 349800 10969 365800 11113
rect 404600 10969 420600 11113
rect 459400 10969 475400 11113
rect 514200 10969 530200 11113
rect 295000 10957 311023 10969
rect 349800 10957 365823 10969
rect 404600 10957 420623 10969
rect 459400 10957 475423 10969
rect 514200 10957 530223 10969
rect 294979 5982 311023 10957
rect 349779 5982 365823 10957
rect 404579 5982 420623 10957
rect 459379 5982 475423 10957
rect 514179 5982 530223 10957
rect 294979 4271 311017 5982
rect 349779 4271 365817 5982
rect 404579 4271 420617 5982
rect 459379 4271 475417 5982
rect 514179 4271 530217 5982
rect 295000 59 311000 4271
rect 349800 59 365800 4271
rect 404600 59 420600 4271
rect 459400 59 475400 4271
rect 514200 59 530200 4271
rect 569445 61 583786 39593
rect 623229 61 637678 39593
<< metal1 >>
rect 673730 855380 673736 855432
rect 673788 855420 673794 855432
rect 675386 855420 675392 855432
rect 673788 855392 675392 855420
rect 673788 855380 673794 855392
rect 675386 855380 675392 855392
rect 675444 855380 675450 855432
rect 42242 787992 42248 788044
rect 42300 788032 42306 788044
rect 42426 788032 42432 788044
rect 42300 788004 42432 788032
rect 42300 787992 42306 788004
rect 42426 787992 42432 788004
rect 42484 787992 42490 788044
rect 673730 773304 673736 773356
rect 673788 773344 673794 773356
rect 675202 773344 675208 773356
rect 673788 773316 675208 773344
rect 673788 773304 673794 773316
rect 675202 773304 675208 773316
rect 675260 773344 675266 773356
rect 675386 773344 675392 773356
rect 675260 773316 675392 773344
rect 675260 773304 675266 773316
rect 675386 773304 675392 773316
rect 675444 773304 675450 773356
rect 673730 769088 673736 769140
rect 673788 769128 673794 769140
rect 675202 769128 675208 769140
rect 673788 769100 675208 769128
rect 673788 769088 673794 769100
rect 675202 769088 675208 769100
rect 675260 769128 675266 769140
rect 675386 769128 675392 769140
rect 675260 769100 675392 769128
rect 675260 769088 675266 769100
rect 675386 769088 675392 769100
rect 675444 769088 675450 769140
rect 673730 728560 673736 728612
rect 673788 728600 673794 728612
rect 675386 728600 675392 728612
rect 673788 728572 675392 728600
rect 673788 728560 673794 728572
rect 675386 728560 675392 728572
rect 675444 728560 675450 728612
rect 673454 724004 673460 724056
rect 673512 724044 673518 724056
rect 675386 724044 675392 724056
rect 673512 724016 675392 724044
rect 673512 724004 673518 724016
rect 675386 724004 675392 724016
rect 675444 724004 675450 724056
rect 673454 684292 673460 684344
rect 673512 684332 673518 684344
rect 675294 684332 675300 684344
rect 673512 684304 675300 684332
rect 673512 684292 673518 684304
rect 675294 684292 675300 684304
rect 675352 684292 675358 684344
rect 673822 680076 673828 680128
rect 673880 680116 673886 680128
rect 675386 680116 675392 680128
rect 673880 680088 675392 680116
rect 673880 680076 673886 680088
rect 675386 680076 675392 680088
rect 675444 680076 675450 680128
rect 673822 640092 673828 640144
rect 673880 640132 673886 640144
rect 675294 640132 675300 640144
rect 673880 640104 675300 640132
rect 673880 640092 673886 640104
rect 675294 640092 675300 640104
rect 675352 640092 675358 640144
rect 673730 635740 673736 635792
rect 673788 635780 673794 635792
rect 675294 635780 675300 635792
rect 673788 635752 675300 635780
rect 673788 635740 673794 635752
rect 675294 635740 675300 635752
rect 675352 635740 675358 635792
rect 673730 596096 673736 596148
rect 673788 596136 673794 596148
rect 675202 596136 675208 596148
rect 673788 596108 675208 596136
rect 673788 596096 673794 596108
rect 675202 596096 675208 596108
rect 675260 596136 675266 596148
rect 675386 596136 675392 596148
rect 675260 596108 675392 596136
rect 675260 596096 675266 596108
rect 675386 596096 675392 596108
rect 675444 596096 675450 596148
rect 673730 590792 673736 590844
rect 673788 590832 673794 590844
rect 675202 590832 675208 590844
rect 673788 590804 675208 590832
rect 673788 590792 673794 590804
rect 675202 590792 675208 590804
rect 675260 590832 675266 590844
rect 675386 590832 675392 590844
rect 675260 590804 675392 590832
rect 675260 590792 675266 590804
rect 675386 590792 675392 590804
rect 675444 590792 675450 590844
rect 41782 576512 41788 576564
rect 41840 576552 41846 576564
rect 42242 576552 42248 576564
rect 41840 576524 42248 576552
rect 41840 576512 41846 576524
rect 42242 576512 42248 576524
rect 42300 576552 42306 576564
rect 42426 576552 42432 576564
rect 42300 576524 42432 576552
rect 42300 576512 42306 576524
rect 42426 576512 42432 576524
rect 42484 576512 42490 576564
rect 673730 551488 673736 551540
rect 673788 551528 673794 551540
rect 675202 551528 675208 551540
rect 673788 551500 675208 551528
rect 673788 551488 673794 551500
rect 675202 551488 675208 551500
rect 675260 551488 675266 551540
rect 673454 547000 673460 547052
rect 673512 547040 673518 547052
rect 675202 547040 675208 547052
rect 673512 547012 675208 547040
rect 673512 547000 673518 547012
rect 675202 547000 675208 547012
rect 675260 547040 675266 547052
rect 675386 547040 675392 547052
rect 675260 547012 675392 547040
rect 675260 547000 675266 547012
rect 675386 547000 675392 547012
rect 675444 547000 675450 547052
rect 673546 372784 673552 372836
rect 673604 372824 673610 372836
rect 675386 372824 675392 372836
rect 673604 372796 675392 372824
rect 673604 372784 673610 372796
rect 675386 372784 675392 372796
rect 675444 372784 675450 372836
rect 673546 333072 673552 333124
rect 673604 333112 673610 333124
rect 675294 333112 675300 333124
rect 673604 333084 675300 333112
rect 673604 333072 673610 333084
rect 675294 333072 675300 333084
rect 675352 333072 675358 333124
rect 673730 328244 673736 328296
rect 673788 328284 673794 328296
rect 675386 328284 675392 328296
rect 673788 328256 675392 328284
rect 673788 328244 673794 328256
rect 675386 328244 675392 328256
rect 675444 328244 675450 328296
rect 42242 313080 42248 313132
rect 42300 313120 42306 313132
rect 42300 313092 42380 313120
rect 42300 313080 42306 313092
rect 42352 312928 42380 313092
rect 42334 312876 42340 312928
rect 42392 312876 42398 312928
rect 673730 289280 673736 289332
rect 673788 289320 673794 289332
rect 675386 289320 675392 289332
rect 673788 289292 675392 289320
rect 673788 289280 673794 289292
rect 675386 289280 675392 289292
rect 675444 289280 675450 289332
rect 42334 284112 42340 284164
rect 42392 284112 42398 284164
rect 42352 283960 42380 284112
rect 673730 284044 673736 284096
rect 673788 284084 673794 284096
rect 675386 284084 675392 284096
rect 673788 284056 675392 284084
rect 673788 284044 673794 284056
rect 675386 284044 675392 284056
rect 675444 284044 675450 284096
rect 42334 283908 42340 283960
rect 42392 283908 42398 283960
rect 673730 244604 673736 244656
rect 673788 244644 673794 244656
rect 675386 244644 675392 244656
rect 673788 244616 675392 244644
rect 673788 244604 673794 244616
rect 675386 244604 675392 244616
rect 675444 244604 675450 244656
rect 673730 239640 673736 239692
rect 673788 239680 673794 239692
rect 675386 239680 675392 239692
rect 673788 239652 675392 239680
rect 673788 239640 673794 239652
rect 675386 239640 675392 239652
rect 675444 239640 675450 239692
rect 673730 200404 673736 200456
rect 673788 200444 673794 200456
rect 675386 200444 675392 200456
rect 673788 200416 675392 200444
rect 673788 200404 673794 200416
rect 675386 200404 675392 200416
rect 675444 200404 675450 200456
rect 673730 195780 673736 195832
rect 673788 195820 673794 195832
rect 675386 195820 675392 195832
rect 673788 195792 675392 195820
rect 673788 195780 673794 195792
rect 675386 195780 675392 195792
rect 675444 195780 675450 195832
rect 673730 156272 673736 156324
rect 673788 156312 673794 156324
rect 675386 156312 675392 156324
rect 673788 156284 675392 156312
rect 673788 156272 673794 156284
rect 675386 156272 675392 156284
rect 675444 156272 675450 156324
rect 673822 151716 673828 151768
rect 673880 151756 673886 151768
rect 675294 151756 675300 151768
rect 673880 151728 675300 151756
rect 673880 151716 673886 151728
rect 675294 151716 675300 151728
rect 675352 151716 675358 151768
rect 673822 111800 673828 111852
rect 673880 111840 673886 111852
rect 675386 111840 675392 111852
rect 673880 111812 675392 111840
rect 673880 111800 673886 111812
rect 675386 111800 675392 111812
rect 675444 111800 675450 111852
rect 673638 107312 673644 107364
rect 673696 107352 673702 107364
rect 675294 107352 675300 107364
rect 673696 107324 675300 107352
rect 673696 107312 673702 107324
rect 675294 107312 675300 107324
rect 675352 107312 675358 107364
rect 673638 46968 673644 46980
rect 527468 46940 673644 46968
rect 527468 46912 527496 46940
rect 673638 46928 673644 46940
rect 673696 46928 673702 46980
rect 527450 46860 527456 46912
rect 527508 46860 527514 46912
rect 42334 45568 42340 45620
rect 42392 45608 42398 45620
rect 143626 45608 143632 45620
rect 42392 45580 143632 45608
rect 42392 45568 42398 45580
rect 143626 45568 143632 45580
rect 143684 45568 143690 45620
rect 143626 44140 143632 44192
rect 143684 44180 143690 44192
rect 145098 44180 145104 44192
rect 143684 44152 145104 44180
rect 143684 44140 143690 44152
rect 145098 44140 145104 44152
rect 145156 44180 145162 44192
rect 195330 44180 195336 44192
rect 145156 44152 195336 44180
rect 145156 44140 145162 44152
rect 195330 44140 195336 44152
rect 195388 44180 195394 44192
rect 199654 44180 199660 44192
rect 195388 44152 199660 44180
rect 195388 44140 195394 44152
rect 199654 44140 199660 44152
rect 199712 44140 199718 44192
rect 363046 44316 363052 44328
rect 303586 44288 303936 44316
rect 199838 44208 199844 44260
rect 199896 44248 199902 44260
rect 303586 44248 303614 44288
rect 303908 44260 303936 44288
rect 361546 44288 363052 44316
rect 199896 44220 303614 44248
rect 199896 44208 199902 44220
rect 303890 44208 303896 44260
rect 303948 44248 303954 44260
rect 308214 44248 308220 44260
rect 303948 44220 308220 44248
rect 303948 44208 303954 44220
rect 308214 44208 308220 44220
rect 308272 44248 308278 44260
rect 358722 44248 358728 44260
rect 308272 44220 358728 44248
rect 308272 44208 308278 44220
rect 358722 44208 358728 44220
rect 358780 44248 358786 44260
rect 361546 44248 361574 44288
rect 363046 44276 363052 44288
rect 363104 44316 363110 44328
rect 413554 44316 413560 44328
rect 363104 44288 413560 44316
rect 363104 44276 363110 44288
rect 413554 44276 413560 44288
rect 413612 44316 413618 44328
rect 417878 44316 417884 44328
rect 413612 44288 417884 44316
rect 413612 44276 413618 44288
rect 417878 44276 417884 44288
rect 417936 44316 417942 44328
rect 468294 44316 468300 44328
rect 417936 44288 468300 44316
rect 417936 44276 417942 44288
rect 468294 44276 468300 44288
rect 468352 44316 468358 44328
rect 472618 44316 472624 44328
rect 468352 44288 472624 44316
rect 468352 44276 468358 44288
rect 472618 44276 472624 44288
rect 472676 44316 472682 44328
rect 472676 44288 523172 44316
rect 472676 44276 472682 44288
rect 358780 44220 361574 44248
rect 358780 44208 358786 44220
rect 523144 44192 523172 44288
rect 523126 44140 523132 44192
rect 523184 44180 523190 44192
rect 527450 44180 527456 44192
rect 523184 44152 527456 44180
rect 523184 44140 523190 44152
rect 527450 44140 527456 44152
rect 527508 44140 527514 44192
rect 409322 41760 409328 41812
rect 409380 41800 409386 41812
rect 412358 41800 412364 41812
rect 409380 41772 412364 41800
rect 409380 41760 409386 41772
rect 412358 41760 412364 41772
rect 412416 41800 412422 41812
rect 415210 41800 415216 41812
rect 412416 41772 415216 41800
rect 412416 41760 412422 41772
rect 415210 41760 415216 41772
rect 415268 41760 415274 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
<< via1 >>
rect 673736 855380 673788 855432
rect 675392 855380 675444 855432
rect 42248 787992 42300 788044
rect 42432 787992 42484 788044
rect 673736 773304 673788 773356
rect 675208 773304 675260 773356
rect 675392 773304 675444 773356
rect 673736 769088 673788 769140
rect 675208 769088 675260 769140
rect 675392 769088 675444 769140
rect 673736 728560 673788 728612
rect 675392 728560 675444 728612
rect 673460 724004 673512 724056
rect 675392 724004 675444 724056
rect 673460 684292 673512 684344
rect 675300 684292 675352 684344
rect 673828 680076 673880 680128
rect 675392 680076 675444 680128
rect 673828 640092 673880 640144
rect 675300 640092 675352 640144
rect 673736 635740 673788 635792
rect 675300 635740 675352 635792
rect 673736 596096 673788 596148
rect 675208 596096 675260 596148
rect 675392 596096 675444 596148
rect 673736 590792 673788 590844
rect 675208 590792 675260 590844
rect 675392 590792 675444 590844
rect 41788 576512 41840 576564
rect 42248 576512 42300 576564
rect 42432 576512 42484 576564
rect 673736 551488 673788 551540
rect 675208 551488 675260 551540
rect 673460 547000 673512 547052
rect 675208 547000 675260 547052
rect 675392 547000 675444 547052
rect 673552 372784 673604 372836
rect 675392 372784 675444 372836
rect 673552 333072 673604 333124
rect 675300 333072 675352 333124
rect 673736 328244 673788 328296
rect 675392 328244 675444 328296
rect 42248 313080 42300 313132
rect 42340 312876 42392 312928
rect 673736 289280 673788 289332
rect 675392 289280 675444 289332
rect 42340 284112 42392 284164
rect 673736 284044 673788 284096
rect 675392 284044 675444 284096
rect 42340 283908 42392 283960
rect 673736 244604 673788 244656
rect 675392 244604 675444 244656
rect 673736 239640 673788 239692
rect 675392 239640 675444 239692
rect 673736 200404 673788 200456
rect 675392 200404 675444 200456
rect 673736 195780 673788 195832
rect 675392 195780 675444 195832
rect 673736 156272 673788 156324
rect 675392 156272 675444 156324
rect 673828 151716 673880 151768
rect 675300 151716 675352 151768
rect 673828 111800 673880 111852
rect 675392 111800 675444 111852
rect 673644 107312 673696 107364
rect 675300 107312 675352 107364
rect 673644 46928 673696 46980
rect 527456 46860 527508 46912
rect 42340 45568 42392 45620
rect 143632 45568 143684 45620
rect 143632 44140 143684 44192
rect 145104 44140 145156 44192
rect 195336 44140 195388 44192
rect 199660 44140 199712 44192
rect 199844 44208 199896 44260
rect 303896 44208 303948 44260
rect 308220 44208 308272 44260
rect 358728 44208 358780 44260
rect 363052 44276 363104 44328
rect 413560 44276 413612 44328
rect 417884 44276 417936 44328
rect 468300 44276 468352 44328
rect 472624 44276 472676 44328
rect 523132 44140 523184 44192
rect 527456 44140 527508 44192
rect 409328 41760 409380 41812
rect 412364 41760 412416 41812
rect 415216 41760 415268 41812
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
<< obsm1 >>
rect 75850 1006851 89088 1007371
rect 123850 1006851 137088 1007371
rect 171850 1006851 185088 1007371
rect 229437 998007 243983 1037545
rect 280837 998007 295383 1037545
rect 339437 998007 354124 1037545
rect 425650 1006851 438888 1007371
rect 475050 1006851 488288 1007371
rect 526650 1006851 539888 1007371
rect 575637 998007 590324 1037545
rect 627850 1006851 641088 1007371
rect 230125 997826 231171 998007
rect 231807 997984 232070 998007
tri 232070 997984 232093 998007 sw
tri 243285 997984 243308 998007 se
rect 243308 997984 243536 998007
rect 231807 997794 243536 997984
rect 281525 997826 282571 998007
rect 283207 997984 283470 998007
tri 283470 997984 283493 998007 sw
tri 294685 997984 294708 998007 se
rect 294708 997984 294936 998007
rect 283207 997794 294936 997984
rect 341807 997984 342070 998007
tri 342070 997984 342093 998007 sw
tri 353285 997984 353308 998007 se
rect 353308 997984 353536 998007
rect 341807 997794 353536 997984
rect 578007 997984 578270 998007
tri 578270 997984 578293 998007 sw
tri 589485 997984 589508 998007 se
rect 589508 997984 589736 998007
rect 578007 997794 589736 997984
rect 585778 996452 585842 996464
rect 674742 996452 674806 996464
rect 585778 996424 674806 996452
rect 585778 996412 585842 996424
rect 674742 996412 674806 996424
rect 42242 996384 42306 996396
rect 339494 996384 339558 996396
rect 673546 996384 673610 996396
rect 42242 996356 673610 996384
rect 42242 996344 42306 996356
rect 339494 996344 339558 996356
rect 673546 996344 673610 996356
rect 44910 990128 44974 990140
rect 673638 990128 673702 990140
rect 44910 990100 673702 990128
rect 44910 990088 44974 990100
rect 673638 990088 673702 990100
rect 42334 990060 42398 990072
rect 673454 990060 673518 990072
rect 42334 990032 673518 990060
rect 42334 990020 42398 990032
rect 673454 990020 673518 990032
rect 30229 956050 30749 969288
rect 678007 958275 717545 958963
rect 677826 957229 717545 958275
rect 678007 956593 717545 957229
rect 677794 956330 717545 956593
rect 677794 945092 677984 956330
tri 677984 956307 678007 956330 nw
tri 677984 945092 678007 945115 sw
rect 678007 945092 717545 956330
rect 677794 944864 717545 945092
rect 678007 944417 717545 944864
rect 24523 929387 40977 930187
tri 40977 929387 41777 930187 sw
rect 24523 928240 41777 929387
rect 32 924313 39593 928000
rect 39756 924313 41777 928240
rect 32 917185 41777 924313
rect 32 916331 39600 917185
rect 32 913024 39593 916331
rect 678007 903069 717568 906376
rect 678000 902215 717568 903069
rect 675823 895087 717568 902215
rect 675823 891160 677844 895087
rect 678007 891400 717568 895087
rect 675823 890013 693077 891160
tri 675823 889213 676623 890013 ne
rect 676623 889213 693077 890013
rect 55 884936 39593 885383
rect 55 884708 39806 884936
rect 55 873470 39593 884708
tri 39593 884685 39616 884708 ne
tri 39593 873470 39616 873493 se
rect 39616 873470 39806 884708
rect 55 873207 39806 873470
rect 55 872571 39593 873207
rect 55 871525 39774 872571
rect 55 870837 39593 871525
rect 689038 863000 693727 863023
rect 695550 863000 695896 863029
rect 696779 863000 703644 863023
rect 703855 863000 711618 863023
rect 42426 861200 42490 861212
rect 44174 861200 44238 861212
rect 42426 861172 44238 861200
rect 42426 861160 42490 861172
rect 44174 861160 44238 861172
rect 673546 859160 673610 859172
rect 675386 859160 675450 859172
rect 673546 859132 675450 859160
rect 673546 859120 673610 859132
rect 675386 859120 675450 859132
rect 673638 856100 673702 856112
rect 675386 856100 675450 856112
rect 673638 856072 675450 856100
rect 673638 856060 673702 856072
rect 675386 856060 675450 856072
rect 673454 849708 673518 849720
rect 675386 849708 675450 849720
rect 673454 849680 675450 849708
rect 673454 849668 673518 849680
rect 675386 849668 675450 849680
rect 676231 847000 717600 863000
rect 681497 846977 682603 847000
rect 683624 846977 684745 847000
rect 687844 846988 696516 847000
rect 687844 846977 692186 846988
tri 692186 846977 692197 846988 nw
rect 696779 846971 703644 847000
rect 703855 846971 711618 847000
rect 713380 846996 713795 847000
rect 55 842536 39593 843124
rect 55 842308 39806 842536
rect 55 831070 39593 842308
tri 39593 842285 39616 842308 ne
tri 39593 831070 39616 831093 se
rect 39616 831070 39806 842308
rect 55 830807 39806 831070
rect 55 828437 39593 830807
rect 678007 818075 717545 818763
rect 677826 817029 717545 818075
rect 678007 816393 717545 817029
rect 677794 816130 717545 816393
rect 677794 804892 677984 816130
tri 677984 816107 678007 816130 nw
tri 677984 804892 678007 804915 sw
rect 678007 804892 717545 816130
rect 677794 804664 717545 804892
rect 678007 804217 717545 804664
rect 675294 803808 675358 803820
rect 677594 803808 677658 803820
rect 675294 803780 677658 803808
rect 675294 803768 675358 803780
rect 677594 803768 677658 803780
rect 3805 801200 4220 801204
rect 5982 801200 13745 801229
rect 13956 801200 20821 801229
tri 25403 801212 25414 801223 se
rect 25414 801212 29756 801223
rect 21084 801200 29756 801212
rect 32855 801200 33976 801223
rect 34997 801200 36103 801223
rect 0 785200 41369 801200
rect 42242 801020 42306 801032
rect 42610 801020 42674 801032
rect 42242 800992 42674 801020
rect 42242 800980 42306 800992
rect 42610 800980 42674 800992
rect 41782 798572 41846 798584
rect 42334 798572 42398 798584
rect 41782 798544 42398 798572
rect 41782 798532 41846 798544
rect 42334 798532 42398 798544
rect 41782 792112 41846 792124
rect 42426 792112 42490 792124
rect 41782 792084 42490 792112
rect 41782 792072 41846 792084
rect 42426 792072 42490 792084
rect 41782 789120 41846 789132
rect 42610 789120 42674 789132
rect 41782 789092 42674 789120
rect 41782 789080 41846 789092
rect 42610 789080 42674 789092
rect 5982 785177 13745 785200
rect 13956 785177 20821 785200
rect 21704 785171 22050 785200
rect 23873 785177 28562 785200
rect 689038 775600 693727 775623
rect 695550 775600 695896 775629
rect 696779 775600 703644 775623
rect 703855 775600 711618 775623
rect 673546 772800 673610 772812
rect 675386 772800 675450 772812
rect 673546 772772 675450 772800
rect 673546 772760 673610 772772
rect 675386 772760 675450 772772
rect 673638 769672 673702 769684
rect 673914 769672 673978 769684
rect 675386 769672 675450 769684
rect 673638 769644 675450 769672
rect 673638 769632 673702 769644
rect 673914 769632 673978 769644
rect 675386 769632 675450 769644
rect 675202 767632 675266 767644
rect 675386 767632 675450 767644
rect 675202 767604 675450 767632
rect 675202 767592 675266 767604
rect 675386 767592 675450 767604
rect 673454 761308 673518 761320
rect 674006 761308 674070 761320
rect 675386 761308 675450 761320
rect 673454 761280 675450 761308
rect 673454 761268 673518 761280
rect 674006 761268 674070 761280
rect 675386 761268 675450 761280
rect 675202 760220 675266 760232
rect 675386 760220 675450 760232
rect 675202 760192 675450 760220
rect 675202 760180 675266 760192
rect 675386 760180 675450 760192
rect 676231 759600 717600 775600
rect 681497 759577 682603 759600
rect 683624 759577 684745 759600
rect 687844 759588 696516 759600
rect 687844 759577 692186 759588
tri 692186 759577 692197 759588 nw
rect 696779 759571 703644 759600
rect 703855 759571 711618 759600
rect 713380 759596 713795 759600
rect 3805 758000 4220 758004
rect 5982 758000 13745 758029
rect 13956 758000 20821 758029
tri 25403 758012 25414 758023 se
rect 25414 758012 29756 758023
rect 21084 758000 29756 758012
rect 32855 758000 33976 758023
rect 34997 758000 36103 758023
rect 0 742000 41369 758000
rect 41782 756276 41846 756288
rect 42334 756276 42398 756288
rect 42610 756276 42674 756288
rect 41782 756248 42674 756276
rect 41782 756236 41846 756248
rect 42334 756236 42398 756248
rect 42610 756236 42674 756248
rect 41782 748320 41846 748332
rect 42518 748320 42582 748332
rect 41782 748292 42582 748320
rect 41782 748280 41846 748292
rect 42518 748280 42582 748292
rect 41782 744852 41846 744864
rect 42426 744852 42490 744864
rect 42702 744852 42766 744864
rect 41782 744824 42766 744852
rect 41782 744812 41846 744824
rect 42426 744812 42490 744824
rect 42702 744812 42766 744824
rect 5982 741977 13745 742000
rect 13956 741977 20821 742000
rect 21704 741971 22050 742000
rect 23873 741977 28562 742000
rect 689038 731200 693727 731223
rect 695550 731200 695896 731229
rect 696779 731200 703644 731223
rect 703855 731200 711618 731223
rect 673546 728396 673610 728408
rect 675386 728396 675450 728408
rect 673546 728368 675450 728396
rect 673546 728356 673610 728368
rect 675386 728356 675450 728368
rect 673914 725268 673978 725280
rect 675386 725268 675450 725280
rect 673914 725240 675450 725268
rect 673914 725228 673978 725240
rect 675386 725228 675450 725240
rect 673638 717856 673702 717868
rect 674006 717856 674070 717868
rect 675386 717856 675450 717868
rect 673638 717828 675450 717856
rect 673638 717816 673702 717828
rect 674006 717816 674070 717828
rect 675386 717816 675450 717828
rect 676231 715200 717600 731200
rect 681497 715177 682603 715200
rect 683624 715177 684745 715200
rect 687844 715188 696516 715200
rect 687844 715177 692186 715188
tri 692186 715177 692197 715188 nw
rect 696779 715171 703644 715200
rect 703855 715171 711618 715200
rect 713380 715196 713795 715200
rect 3805 714800 4220 714804
rect 5982 714800 13745 714829
rect 13956 714800 20821 714829
tri 25403 714812 25414 714823 se
rect 25414 714812 29756 714823
rect 21084 714800 29756 714812
rect 32855 714800 33976 714823
rect 34997 714800 36103 714823
rect 0 698800 41369 714800
rect 41782 713096 41846 713108
rect 42610 713096 42674 713108
rect 41782 713068 42674 713096
rect 41782 713056 41846 713068
rect 42610 713056 42674 713068
rect 41782 704800 41846 704812
rect 42518 704800 42582 704812
rect 41782 704772 42582 704800
rect 41782 704760 41846 704772
rect 42518 704760 42582 704772
rect 41782 701672 41846 701684
rect 42426 701672 42490 701684
rect 41782 701644 42490 701672
rect 41782 701632 41846 701644
rect 42426 701632 42490 701644
rect 5982 698777 13745 698800
rect 13956 698777 20821 698800
rect 21704 698771 22050 698800
rect 23873 698777 28562 698800
rect 689038 687000 693727 687023
rect 695550 687000 695896 687029
rect 696779 687000 703644 687023
rect 703855 687000 711618 687023
rect 673546 683108 673610 683120
rect 673730 683108 673794 683120
rect 675386 683108 675450 683120
rect 673546 683080 675450 683108
rect 673546 683068 673610 683080
rect 673730 683068 673794 683080
rect 675386 683068 675450 683080
rect 673546 680456 673610 680468
rect 673914 680456 673978 680468
rect 675386 680456 675450 680468
rect 673546 680428 675450 680456
rect 673546 680416 673610 680428
rect 673914 680416 673978 680428
rect 675386 680416 675450 680428
rect 675202 678824 675266 678836
rect 675386 678824 675450 678836
rect 675202 678796 675450 678824
rect 675202 678784 675266 678796
rect 675386 678784 675450 678796
rect 673638 673656 673702 673668
rect 674006 673656 674070 673668
rect 675386 673656 675450 673668
rect 673638 673628 675450 673656
rect 673638 673616 673702 673628
rect 674006 673616 674070 673628
rect 675386 673616 675450 673628
rect 3805 671400 4220 671404
rect 5982 671400 13745 671429
rect 13956 671400 20821 671429
tri 25403 671412 25414 671423 se
rect 25414 671412 29756 671423
rect 21084 671400 29756 671412
rect 32855 671400 33976 671423
rect 34997 671400 36103 671423
rect 0 655400 41369 671400
rect 676231 671000 717600 687000
rect 681497 670977 682603 671000
rect 683624 670977 684745 671000
rect 687844 670988 696516 671000
rect 687844 670977 692186 670988
tri 692186 670977 692197 670988 nw
rect 696779 670971 703644 671000
rect 703855 670971 711618 671000
rect 713380 670996 713795 671000
rect 41782 668760 41846 668772
rect 42610 668760 42674 668772
rect 41782 668732 42674 668760
rect 41782 668720 41846 668732
rect 42610 668720 42674 668732
rect 41782 661348 41846 661360
rect 42518 661348 42582 661360
rect 41782 661320 42582 661348
rect 41782 661308 41846 661320
rect 42518 661308 42582 661320
rect 41782 659308 41846 659320
rect 42426 659308 42490 659320
rect 42702 659308 42766 659320
rect 41782 659280 42766 659308
rect 41782 659268 41846 659280
rect 42426 659268 42490 659280
rect 42702 659268 42766 659280
rect 5982 655377 13745 655400
rect 13956 655377 20821 655400
rect 21704 655371 22050 655400
rect 23873 655377 28562 655400
rect 689038 642800 693727 642823
rect 695550 642800 695896 642829
rect 696779 642800 703644 642823
rect 703855 642800 711618 642823
rect 673638 638908 673702 638920
rect 675386 638908 675450 638920
rect 673638 638880 675450 638908
rect 673638 638868 673702 638880
rect 675386 638868 675450 638880
rect 673546 636324 673610 636336
rect 675386 636324 675450 636336
rect 673546 636296 675450 636324
rect 673546 636284 673610 636296
rect 675386 636284 675450 636296
rect 675202 634624 675266 634636
rect 675386 634624 675450 634636
rect 675202 634596 675450 634624
rect 675202 634584 675266 634596
rect 675386 634584 675450 634596
rect 673454 629456 673518 629468
rect 674006 629456 674070 629468
rect 675386 629456 675450 629468
rect 673454 629428 675450 629456
rect 673454 629416 673518 629428
rect 674006 629416 674070 629428
rect 675386 629416 675450 629428
rect 3805 628200 4220 628204
rect 5982 628200 13745 628229
rect 13956 628200 20821 628229
tri 25403 628212 25414 628223 se
rect 25414 628212 29756 628223
rect 21084 628200 29756 628212
rect 32855 628200 33976 628223
rect 34997 628200 36103 628223
rect 0 612200 41369 628200
rect 676231 626800 717600 642800
rect 681497 626777 682603 626800
rect 683624 626777 684745 626800
rect 687844 626788 696516 626800
rect 687844 626777 692186 626788
tri 692186 626777 692197 626788 nw
rect 696779 626771 703644 626800
rect 703855 626771 711618 626800
rect 713380 626796 713795 626800
rect 41782 625512 41846 625524
rect 42610 625512 42674 625524
rect 41782 625484 42674 625512
rect 41782 625472 41846 625484
rect 42610 625472 42674 625484
rect 41782 618168 41846 618180
rect 42518 618168 42582 618180
rect 41782 618140 42582 618168
rect 41782 618128 41846 618140
rect 42518 618128 42582 618140
rect 41782 615040 41846 615052
rect 42702 615040 42766 615052
rect 41782 615012 42766 615040
rect 41782 615000 41846 615012
rect 42260 614712 42288 615012
rect 42702 615000 42766 615012
rect 42242 614660 42306 614712
rect 5982 612177 13745 612200
rect 13956 612177 20821 612200
rect 21704 612171 22050 612200
rect 23873 612177 28562 612200
rect 689038 598400 693727 598423
rect 695550 598400 695896 598429
rect 696779 598400 703644 598423
rect 703855 598400 711618 598423
rect 673638 595184 673702 595196
rect 675386 595184 675450 595196
rect 673638 595156 675450 595184
rect 673638 595144 673702 595156
rect 675386 595144 675450 595156
rect 673546 591920 673610 591932
rect 675386 591920 675450 591932
rect 673546 591892 675450 591920
rect 673546 591880 673610 591892
rect 675386 591880 675450 591892
rect 3805 585000 4220 585004
rect 5982 585000 13745 585029
rect 13956 585000 20821 585029
tri 25403 585012 25414 585023 se
rect 25414 585012 29756 585023
rect 21084 585000 29756 585012
rect 32855 585000 33976 585023
rect 34997 585000 36103 585023
rect 0 569000 41369 585000
rect 673454 584168 673518 584180
rect 673914 584168 673978 584180
rect 675386 584168 675450 584180
rect 673454 584140 675450 584168
rect 673454 584128 673518 584140
rect 673914 584128 673978 584140
rect 675386 584128 675450 584140
rect 41782 583284 41846 583296
rect 42610 583284 42674 583296
rect 41782 583256 42674 583284
rect 41782 583244 41846 583256
rect 42610 583244 42674 583256
rect 676231 582400 717600 598400
rect 681497 582377 682603 582400
rect 683624 582377 684745 582400
rect 687844 582388 696516 582400
rect 687844 582377 692186 582388
tri 692186 582377 692197 582388 nw
rect 696779 582371 703644 582400
rect 703855 582371 711618 582400
rect 713380 582396 713795 582400
rect 41782 575940 41846 575952
rect 42518 575940 42582 575952
rect 41782 575912 42582 575940
rect 41782 575900 41846 575912
rect 42518 575900 42582 575912
rect 41782 571860 41846 571872
rect 42426 571860 42490 571872
rect 41782 571832 42490 571860
rect 41782 571820 41846 571832
rect 42426 571820 42490 571832
rect 5982 568977 13745 569000
rect 13956 568977 20821 569000
rect 21704 568971 22050 569000
rect 23873 568977 28562 569000
rect 689038 554200 693727 554223
rect 695550 554200 695896 554229
rect 696779 554200 703644 554223
rect 703855 554200 711618 554223
rect 673638 551392 673702 551404
rect 675386 551392 675450 551404
rect 673638 551364 675450 551392
rect 673638 551352 673702 551364
rect 675386 551352 675450 551364
rect 673546 548264 673610 548276
rect 675386 548264 675450 548276
rect 673546 548236 675450 548264
rect 673546 548224 673610 548236
rect 675386 548224 675450 548236
rect 3805 541800 4220 541804
rect 5982 541800 13745 541829
rect 13956 541800 20821 541829
tri 25403 541812 25414 541823 se
rect 25414 541812 29756 541823
rect 21084 541800 29756 541812
rect 32855 541800 33976 541823
rect 34997 541800 36103 541823
rect 0 525800 41369 541800
rect 673914 540920 673978 540932
rect 675386 540920 675450 540932
rect 673914 540892 675450 540920
rect 673914 540880 673978 540892
rect 675386 540880 675450 540892
rect 41782 540104 41846 540116
rect 42610 540104 42674 540116
rect 41782 540076 42674 540104
rect 41782 540064 41846 540076
rect 42610 540064 42674 540076
rect 676231 538200 717600 554200
rect 681497 538177 682603 538200
rect 683624 538177 684745 538200
rect 687844 538188 696516 538200
rect 687844 538177 692186 538188
tri 692186 538177 692197 538188 nw
rect 696779 538171 703644 538200
rect 703855 538171 711618 538200
rect 713380 538196 713795 538200
rect 41782 531808 41846 531820
rect 42518 531808 42582 531820
rect 42702 531808 42766 531820
rect 41782 531780 42766 531808
rect 41782 531768 41846 531780
rect 42518 531768 42582 531780
rect 42702 531768 42766 531780
rect 41782 528680 41846 528692
rect 42426 528680 42490 528692
rect 41782 528652 42490 528680
rect 41782 528640 41846 528652
rect 42426 528640 42490 528652
rect 5982 525777 13745 525800
rect 13956 525777 20821 525800
rect 21704 525771 22050 525800
rect 23873 525777 28562 525800
rect 678007 509275 717545 509963
rect 677826 508229 717545 509275
rect 678007 507593 717545 508229
rect 677794 507330 717545 507593
rect 675294 499508 675358 499520
rect 676122 499508 676186 499520
rect 675294 499480 676186 499508
rect 675294 499468 675358 499480
rect 676122 499468 676186 499480
rect 55 497536 39593 497983
rect 55 497308 39806 497536
rect 55 486070 39593 497308
tri 39593 497285 39616 497308 ne
tri 39593 486070 39616 486093 se
rect 39616 486070 39806 497308
rect 677794 496092 677984 507330
tri 677984 507307 678007 507330 nw
tri 677984 496092 678007 496115 sw
rect 678007 496092 717545 507330
rect 677794 495864 717545 496092
rect 678007 495417 717545 495864
rect 676122 494884 676186 494896
rect 677962 494884 678026 494896
rect 676122 494856 678026 494884
rect 676122 494844 676186 494856
rect 677962 494844 678026 494856
rect 55 485807 39806 486070
rect 55 485171 39593 485807
rect 55 484125 39774 485171
rect 55 483437 39593 484125
rect 678007 463269 717568 466576
rect 678000 462415 717568 463269
rect 24523 457587 40977 458387
tri 40977 457587 41777 458387 sw
rect 24523 456440 41777 457587
rect 32 452513 39593 456200
rect 39756 452513 41777 456440
rect 32 445385 41777 452513
rect 675823 455287 717568 462415
rect 675823 451360 677844 455287
rect 678007 451600 717568 455287
rect 675823 450213 693077 451360
tri 675823 449413 676623 450213 ne
rect 676623 449413 693077 450213
rect 32 444531 39600 445385
rect 32 441224 39593 444531
rect 674006 422260 674070 422272
rect 674742 422260 674806 422272
rect 674006 422232 674806 422260
rect 674006 422220 674070 422232
rect 674742 422220 674806 422232
rect 678007 420993 717545 423363
rect 677794 420730 717545 420993
rect 674006 419200 674070 419212
rect 677502 419200 677566 419212
rect 674006 419172 677566 419200
rect 674006 419160 674070 419172
rect 677502 419160 677566 419172
rect 3805 414000 4220 414004
rect 5982 414000 13745 414029
rect 13956 414000 20821 414029
tri 25403 414012 25414 414023 se
rect 25414 414012 29756 414023
rect 21084 414000 29756 414012
rect 32855 414000 33976 414023
rect 34997 414000 36103 414023
rect 0 398000 41369 414000
rect 41782 411312 41846 411324
rect 42518 411312 42582 411324
rect 41782 411284 42582 411312
rect 41782 411272 41846 411284
rect 42518 411272 42582 411284
rect 677794 409492 677984 420730
tri 677984 420707 678007 420730 nw
tri 677984 409492 678007 409515 sw
rect 678007 409492 717545 420730
rect 677794 409264 717545 409492
rect 678007 408676 717545 409264
rect 41782 404920 41846 404932
rect 42702 404920 42766 404932
rect 41782 404892 42766 404920
rect 41782 404880 41846 404892
rect 42702 404880 42766 404892
rect 41782 401928 41846 401940
rect 42426 401928 42490 401940
rect 41782 401900 42490 401928
rect 41782 401888 41846 401900
rect 42426 401888 42490 401900
rect 5982 397977 13745 398000
rect 13956 397977 20821 398000
rect 21704 397971 22050 398000
rect 23873 397977 28562 398000
rect 689038 380000 693727 380023
rect 695550 380000 695896 380029
rect 696779 380000 703644 380023
rect 703855 380000 711618 380023
rect 673914 376156 673978 376168
rect 675386 376156 675450 376168
rect 673914 376128 675450 376156
rect 673914 376116 673978 376128
rect 675386 376116 675450 376128
rect 673730 373096 673794 373108
rect 675386 373096 675450 373108
rect 673730 373068 675450 373096
rect 673730 373056 673794 373068
rect 675386 373056 675450 373068
rect 3805 370800 4220 370804
rect 5982 370800 13745 370829
rect 13956 370800 20821 370829
tri 25403 370812 25414 370823 se
rect 25414 370812 29756 370823
rect 21084 370800 29756 370812
rect 32855 370800 33976 370823
rect 34997 370800 36103 370823
rect 0 354800 41369 370800
rect 41782 369084 41846 369096
rect 42518 369084 42582 369096
rect 41782 369056 42582 369084
rect 41782 369044 41846 369056
rect 42518 369044 42582 369056
rect 674006 365752 674070 365764
rect 675386 365752 675450 365764
rect 674006 365724 675450 365752
rect 674006 365712 674070 365724
rect 675386 365712 675450 365724
rect 676231 364000 717600 380000
rect 681497 363977 682603 364000
rect 683624 363977 684745 364000
rect 687844 363988 696516 364000
rect 687844 363977 692186 363988
tri 692186 363977 692197 363988 nw
rect 696779 363971 703644 364000
rect 703855 363971 711618 364000
rect 713380 363996 713795 364000
rect 41782 361332 41846 361344
rect 42610 361332 42674 361344
rect 41782 361304 42674 361332
rect 41782 361292 41846 361304
rect 42610 361292 42674 361304
rect 41782 357660 41846 357672
rect 42426 357660 42490 357672
rect 42702 357660 42766 357672
rect 41782 357632 42766 357660
rect 41782 357620 41846 357632
rect 42426 357620 42490 357632
rect 42702 357620 42766 357632
rect 5982 354777 13745 354800
rect 13956 354777 20821 354800
rect 21704 354771 22050 354800
rect 23873 354777 28562 354800
rect 689038 335800 693727 335823
rect 695550 335800 695896 335829
rect 696779 335800 703644 335823
rect 703855 335800 711618 335823
rect 673730 333996 673794 334008
rect 675202 333996 675266 334008
rect 673730 333968 675266 333996
rect 673730 333956 673794 333968
rect 675202 333956 675266 333968
rect 673454 331956 673518 331968
rect 673914 331956 673978 331968
rect 675386 331956 675450 331968
rect 673454 331928 675450 331956
rect 673454 331916 673518 331928
rect 673914 331916 673978 331928
rect 675386 331916 675450 331928
rect 673546 328896 673610 328908
rect 675202 328896 675266 328908
rect 675386 328896 675450 328908
rect 673546 328868 675450 328896
rect 673546 328856 673610 328868
rect 675202 328856 675266 328868
rect 675386 328856 675450 328868
rect 3805 327400 4220 327404
rect 5982 327400 13745 327429
rect 13956 327400 20821 327429
tri 25403 327412 25414 327423 se
rect 25414 327412 29756 327423
rect 21084 327400 29756 327412
rect 32855 327400 33976 327423
rect 34997 327400 36103 327423
rect 0 311400 41369 327400
rect 41782 325700 41846 325712
rect 42518 325700 42582 325712
rect 41782 325672 42582 325700
rect 41782 325660 41846 325672
rect 42518 325660 42582 325672
rect 673638 322504 673702 322516
rect 674006 322504 674070 322516
rect 675386 322504 675450 322516
rect 673638 322476 675450 322504
rect 673638 322464 673702 322476
rect 674006 322464 674070 322476
rect 675386 322464 675450 322476
rect 676231 319800 717600 335800
rect 681497 319777 682603 319800
rect 683624 319777 684745 319800
rect 687844 319788 696516 319800
rect 687844 319777 692186 319788
tri 692186 319777 692197 319788 nw
rect 696779 319771 703644 319800
rect 703855 319771 711618 319800
rect 713380 319796 713795 319800
rect 41782 317404 41846 317416
rect 42610 317404 42674 317416
rect 41782 317376 42674 317404
rect 41782 317364 41846 317376
rect 42610 317364 42674 317376
rect 41782 314276 41846 314288
rect 42518 314276 42582 314288
rect 42702 314276 42766 314288
rect 41782 314248 42766 314276
rect 41782 314236 41846 314248
rect 42518 314236 42582 314248
rect 42702 314236 42766 314248
rect 5982 311377 13745 311400
rect 13956 311377 20821 311400
rect 21704 311371 22050 311400
rect 23873 311377 28562 311400
rect 689038 291600 693727 291623
rect 695550 291600 695896 291629
rect 696779 291600 703644 291623
rect 703855 291600 711618 291623
rect 673454 288776 673518 288788
rect 675386 288776 675450 288788
rect 673454 288748 675450 288776
rect 673454 288736 673518 288748
rect 675386 288736 675450 288748
rect 673546 285308 673610 285320
rect 675386 285308 675450 285320
rect 673546 285280 675450 285308
rect 673546 285268 673610 285280
rect 675386 285268 675450 285280
rect 3805 284200 4220 284204
rect 5982 284200 13745 284229
rect 13956 284200 20821 284229
tri 25403 284212 25414 284223 se
rect 25414 284212 29756 284223
rect 21084 284200 29756 284212
rect 32855 284200 33976 284223
rect 34997 284200 36103 284223
rect 0 268200 41369 284200
rect 41782 281568 41846 281580
rect 42426 281568 42490 281580
rect 42702 281568 42766 281580
rect 41782 281540 42766 281568
rect 41782 281528 41846 281540
rect 42426 281528 42490 281540
rect 42702 281528 42766 281540
rect 673638 277352 673702 277364
rect 675386 277352 675450 277364
rect 673638 277324 675450 277352
rect 673638 277312 673702 277324
rect 675386 277312 675450 277324
rect 676231 275600 717600 291600
rect 681497 275577 682603 275600
rect 683624 275577 684745 275600
rect 687844 275588 696516 275600
rect 687844 275577 692186 275588
tri 692186 275577 692197 275588 nw
rect 696779 275571 703644 275600
rect 703855 275571 711618 275600
rect 713380 275596 713795 275600
rect 41782 274700 41846 274712
rect 42610 274700 42674 274712
rect 41782 274672 42674 274700
rect 41782 274660 41846 274672
rect 42610 274660 42674 274672
rect 41782 272116 41846 272128
rect 42518 272116 42582 272128
rect 41782 272088 42582 272116
rect 41782 272076 41846 272088
rect 42518 272076 42582 272088
rect 5982 268177 13745 268200
rect 13956 268177 20821 268200
rect 21704 268171 22050 268200
rect 23873 268177 28562 268200
rect 689038 247200 693727 247223
rect 695550 247200 695896 247229
rect 696779 247200 703644 247223
rect 703855 247200 711618 247223
rect 673454 243760 673518 243772
rect 675386 243760 675450 243772
rect 673454 243732 675450 243760
rect 673454 243720 673518 243732
rect 675386 243720 675450 243732
rect 3805 241000 4220 241004
rect 5982 241000 13745 241029
rect 13956 241000 20821 241029
tri 25403 241012 25414 241023 se
rect 25414 241012 29756 241023
rect 21084 241000 29756 241012
rect 32855 241000 33976 241023
rect 34997 241000 36103 241023
rect 0 225000 41369 241000
rect 673546 240292 673610 240304
rect 675386 240292 675450 240304
rect 673546 240264 675450 240292
rect 673546 240252 673610 240264
rect 675386 240252 675450 240264
rect 41782 238320 41846 238332
rect 42426 238320 42490 238332
rect 42702 238320 42766 238332
rect 41782 238292 42766 238320
rect 41782 238280 41846 238292
rect 42426 238280 42490 238292
rect 42702 238280 42766 238292
rect 673638 233900 673702 233912
rect 675386 233900 675450 233912
rect 673638 233872 675450 233900
rect 673638 233860 673702 233872
rect 675386 233860 675450 233872
rect 41782 231928 41846 231940
rect 42610 231928 42674 231940
rect 41782 231900 42674 231928
rect 41782 231888 41846 231900
rect 42610 231888 42674 231900
rect 676231 231200 717600 247200
rect 681497 231177 682603 231200
rect 683624 231177 684745 231200
rect 687844 231188 696516 231200
rect 687844 231177 692186 231188
tri 692186 231177 692197 231188 nw
rect 696779 231171 703644 231200
rect 703855 231171 711618 231200
rect 713380 231196 713795 231200
rect 41782 228868 41846 228880
rect 42518 228868 42582 228880
rect 41782 228840 42582 228868
rect 41782 228828 41846 228840
rect 42518 228828 42582 228840
rect 5982 224977 13745 225000
rect 13956 224977 20821 225000
rect 21704 224971 22050 225000
rect 23873 224977 28562 225000
rect 689038 203000 693727 203023
rect 695550 203000 695896 203029
rect 696779 203000 703644 203023
rect 703855 203000 711618 203023
rect 673454 199152 673518 199164
rect 675386 199152 675450 199164
rect 673454 199124 675450 199152
rect 673454 199112 673518 199124
rect 675386 199112 675450 199124
rect 3805 197800 4220 197804
rect 5982 197800 13745 197829
rect 13956 197800 20821 197829
tri 25403 197812 25414 197823 se
rect 25414 197812 29756 197823
rect 21084 197800 29756 197812
rect 32855 197800 33976 197823
rect 34997 197800 36103 197823
rect 0 181800 41369 197800
rect 673546 197044 673610 197056
rect 675386 197044 675450 197056
rect 673546 197016 675450 197044
rect 673546 197004 673610 197016
rect 675386 197004 675450 197016
rect 41782 195140 41846 195152
rect 42426 195140 42490 195152
rect 41782 195112 42490 195140
rect 41782 195100 41846 195112
rect 42426 195100 42490 195112
rect 673638 189292 673702 189304
rect 675386 189292 675450 189304
rect 673638 189264 675450 189292
rect 673638 189252 673702 189264
rect 675386 189252 675450 189264
rect 41782 188748 41846 188760
rect 42518 188748 42582 188760
rect 42794 188748 42858 188760
rect 41782 188720 42858 188748
rect 41782 188708 41846 188720
rect 42518 188708 42582 188720
rect 42794 188708 42858 188720
rect 676231 187000 717600 203000
rect 681497 186977 682603 187000
rect 683624 186977 684745 187000
rect 687844 186988 696516 187000
rect 687844 186977 692186 186988
tri 692186 186977 692197 186988 nw
rect 696779 186971 703644 187000
rect 703855 186971 711618 187000
rect 713380 186996 713795 187000
rect 41782 185688 41846 185700
rect 42702 185688 42766 185700
rect 41782 185660 42766 185688
rect 41782 185648 41846 185660
rect 42702 185648 42766 185660
rect 42242 184396 42306 184408
rect 42702 184396 42766 184408
rect 42242 184368 42766 184396
rect 42242 184356 42306 184368
rect 42702 184356 42766 184368
rect 5982 181777 13745 181800
rect 13956 181777 20821 181800
rect 21704 181771 22050 181800
rect 23873 181777 28562 181800
rect 689038 158800 693727 158823
rect 695550 158800 695896 158829
rect 696779 158800 703644 158823
rect 703855 158800 711618 158823
rect 673454 155972 673518 155984
rect 673914 155972 673978 155984
rect 675386 155972 675450 155984
rect 673454 155944 675450 155972
rect 673454 155932 673518 155944
rect 673914 155932 673978 155944
rect 675386 155932 675450 155944
rect 673546 152844 673610 152856
rect 675386 152844 675450 152856
rect 673546 152816 675450 152844
rect 673546 152804 673610 152816
rect 675386 152804 675450 152816
rect 673730 144548 673794 144560
rect 675386 144548 675450 144560
rect 673730 144520 675450 144548
rect 673730 144508 673794 144520
rect 675386 144508 675450 144520
rect 676231 142800 717600 158800
rect 681497 142777 682603 142800
rect 683624 142777 684745 142800
rect 687844 142788 696516 142800
rect 687844 142777 692186 142788
tri 692186 142777 692197 142788 nw
rect 696779 142771 703644 142800
rect 703855 142771 711618 142800
rect 713380 142796 713795 142800
rect 55 124336 39593 124783
rect 55 124108 39806 124336
rect 55 112870 39593 124108
tri 39593 124085 39616 124108 ne
tri 39593 112870 39616 112893 se
rect 39616 112870 39806 124108
rect 42518 121496 42582 121508
rect 44174 121496 44238 121508
rect 42518 121468 44238 121496
rect 42518 121456 42582 121468
rect 44174 121456 44238 121468
rect 689038 114400 693727 114423
rect 695550 114400 695896 114429
rect 696779 114400 703644 114423
rect 703855 114400 711618 114423
rect 55 112607 39806 112870
rect 55 111971 39593 112607
rect 55 110925 39774 111971
rect 673454 111568 673518 111580
rect 673914 111568 673978 111580
rect 675386 111568 675450 111580
rect 673454 111540 675450 111568
rect 673454 111528 673518 111540
rect 673914 111528 673978 111540
rect 675386 111528 675450 111540
rect 55 110237 39593 110925
rect 673546 108440 673610 108452
rect 675386 108440 675450 108452
rect 673546 108412 675450 108440
rect 673546 108400 673610 108412
rect 675386 108400 675450 108412
rect 42426 106060 42490 106072
rect 44174 106060 44238 106072
rect 42426 106032 44238 106060
rect 42426 106020 42490 106032
rect 44174 106020 44238 106032
rect 676231 98400 717600 114400
rect 681497 98377 682603 98400
rect 683624 98377 684745 98400
rect 687844 98388 696516 98400
rect 687844 98377 692186 98388
tri 692186 98377 692197 98388 nw
rect 696779 98371 703644 98400
rect 703855 98371 711618 98400
rect 713380 98396 713795 98400
rect 31928 85187 32702 85239
rect 31928 84387 40900 85187
tri 40900 84387 41700 85187 sw
rect 31928 83240 41700 84387
rect 31928 83049 32702 83240
rect 32 79313 39593 83000
rect 39756 79313 41700 83240
rect 32 72099 41700 79313
rect 32 71331 39600 72099
rect 39796 71731 41700 72099
tri 39796 71331 40196 71731 ne
rect 40196 71331 41300 71731
tri 41300 71331 41700 71731 nw
rect 32 68024 39593 71331
rect 44818 46928 44882 46980
rect 200868 46940 297772 46968
rect 44836 46900 44864 46928
rect 200868 46912 200896 46940
rect 143534 46900 143598 46912
rect 44836 46872 143598 46900
rect 143534 46860 143598 46872
rect 200850 46860 200914 46912
rect 240888 46900 240916 46940
rect 297744 46912 297772 46940
rect 309428 46940 352604 46968
rect 309428 46912 309456 46940
rect 352576 46912 352604 46940
rect 364260 46940 407436 46968
rect 364260 46912 364288 46940
rect 407408 46912 407436 46940
rect 419092 46940 462176 46968
rect 419092 46912 419120 46940
rect 462148 46912 462176 46940
rect 473832 46940 517008 46968
rect 473832 46912 473860 46940
rect 516980 46912 517008 46940
rect 256234 46900 256298 46912
rect 240888 46872 256298 46900
rect 256234 46860 256298 46872
rect 297726 46860 297790 46912
rect 309410 46860 309474 46912
rect 352558 46860 352622 46912
rect 364242 46860 364306 46912
rect 407390 46860 407454 46912
rect 419074 46860 419138 46912
rect 462130 46860 462194 46912
rect 473814 46860 473878 46912
rect 516962 46860 517026 46912
rect 42242 45676 42306 45688
rect 140958 45676 141022 45688
rect 42242 45648 141022 45676
rect 42242 45636 42306 45648
rect 140958 45636 141022 45648
rect 186682 45608 186746 45620
rect 194686 45608 194750 45620
rect 186682 45580 194750 45608
rect 186682 45568 186746 45580
rect 194686 45568 194750 45580
rect 523770 45608 523834 45620
rect 673546 45608 673610 45620
rect 523770 45580 673610 45608
rect 523770 45568 523834 45580
rect 673546 45568 673610 45580
rect 44910 45540 44974 45552
rect 195974 45540 196038 45552
rect 44910 45512 196038 45540
rect 44910 45500 44974 45512
rect 195974 45500 196038 45512
rect 518710 45540 518774 45552
rect 673730 45540 673794 45552
rect 518710 45512 673794 45540
rect 518710 45500 518774 45512
rect 673730 45500 673794 45512
rect 349982 44452 350046 44464
rect 359366 44452 359430 44464
rect 414198 44452 414262 44464
rect 349982 44424 414262 44452
rect 349982 44412 350046 44424
rect 359366 44412 359430 44424
rect 414198 44412 414262 44424
rect 188522 44384 188586 44396
rect 192846 44384 192910 44396
rect 297082 44384 297146 44396
rect 299566 44384 299630 44396
rect 305730 44384 305794 44396
rect 468938 44384 469002 44396
rect 523770 44384 523834 44396
rect 188522 44356 201540 44384
rect 188522 44344 188586 44356
rect 192846 44344 192910 44356
rect 201512 44328 201540 44356
rect 284266 44356 322934 44384
rect 195974 44316 196038 44328
rect 201494 44316 201558 44328
rect 284266 44316 284294 44356
rect 297082 44344 297146 44356
rect 299566 44344 299630 44356
rect 305730 44344 305794 44356
rect 195974 44288 199792 44316
rect 195974 44276 196038 44288
rect 199764 44180 199792 44288
rect 201494 44288 284294 44316
rect 295242 44316 295306 44328
rect 303246 44316 303310 44328
rect 322906 44316 322934 44356
rect 468938 44356 523834 44384
rect 468938 44344 469002 44356
rect 523770 44344 523834 44356
rect 351914 44316 351978 44328
rect 354398 44316 354462 44328
rect 360562 44316 360626 44328
rect 295242 44288 303310 44316
rect 201494 44276 201558 44288
rect 295242 44276 295306 44288
rect 303246 44276 303310 44288
rect 322906 44288 360626 44316
rect 351914 44276 351978 44288
rect 354398 44276 354462 44288
rect 360562 44276 360626 44288
rect 406746 44248 406810 44260
rect 461486 44248 461550 44260
rect 516318 44248 516382 44260
rect 518710 44248 518774 44260
rect 380866 44220 518774 44248
rect 304534 44180 304598 44192
rect 349982 44180 350046 44192
rect 199764 44152 350046 44180
rect 304534 44140 304598 44152
rect 349982 44140 350046 44152
rect 350074 44180 350138 44192
rect 358078 44180 358142 44192
rect 350074 44152 358142 44180
rect 350074 44140 350138 44152
rect 358078 44140 358142 44152
rect 360562 44180 360626 44192
rect 380866 44180 380894 44220
rect 406746 44208 406810 44220
rect 461486 44208 461550 44220
rect 516318 44208 516382 44220
rect 518710 44208 518774 44220
rect 360562 44152 380894 44180
rect 414198 44180 414262 44192
rect 468938 44180 469002 44192
rect 414198 44152 469002 44180
rect 360562 44140 360626 44152
rect 414198 44140 414262 44152
rect 468938 44140 469002 44152
rect 579890 42752 579954 42764
rect 673454 42752 673518 42764
rect 579890 42724 673518 42752
rect 579890 42712 579954 42724
rect 673454 42712 673518 42724
rect 189258 41936 189322 41948
rect 191098 41936 191162 41948
rect 192294 41936 192358 41948
rect 193582 41936 193646 41948
rect 196434 41936 196498 41948
rect 189258 41908 196498 41936
rect 189258 41896 189322 41908
rect 191098 41896 191162 41908
rect 192294 41896 192358 41908
rect 193582 41896 193646 41908
rect 196434 41896 196498 41908
rect 198458 41936 198522 41948
rect 200114 41936 200178 41948
rect 198458 41908 200178 41936
rect 198458 41896 198522 41908
rect 200114 41896 200178 41908
rect 297910 41936 297974 41948
rect 300670 41936 300734 41948
rect 297910 41908 300734 41936
rect 297910 41896 297974 41908
rect 300670 41896 300734 41908
rect 302234 41936 302298 41948
rect 305270 41936 305334 41948
rect 306558 41936 306622 41948
rect 308674 41936 308738 41948
rect 302234 41908 308738 41936
rect 302234 41896 302298 41908
rect 305270 41896 305334 41908
rect 306558 41896 306622 41908
rect 308674 41896 308738 41908
rect 352650 41936 352714 41948
rect 355502 41936 355566 41948
rect 352650 41908 355566 41936
rect 352650 41896 352714 41908
rect 355502 41896 355566 41908
rect 356974 41936 357038 41948
rect 359826 41936 359890 41948
rect 361114 41936 361178 41948
rect 363506 41936 363570 41948
rect 356974 41908 363570 41936
rect 356974 41896 357038 41908
rect 359826 41896 359890 41908
rect 361114 41896 361178 41908
rect 363506 41896 363570 41908
rect 407482 41936 407546 41948
rect 410242 41936 410306 41948
rect 411530 41936 411594 41948
rect 414566 41936 414630 41948
rect 415854 41936 415918 41948
rect 418246 41936 418310 41948
rect 407482 41908 418310 41936
rect 407482 41896 407546 41908
rect 410242 41896 410306 41908
rect 411530 41896 411594 41908
rect 414566 41896 414630 41908
rect 415854 41896 415918 41908
rect 418246 41896 418310 41908
rect 462314 41936 462378 41948
rect 465074 41936 465138 41948
rect 466362 41936 466426 41948
rect 469398 41936 469462 41948
rect 470686 41936 470750 41948
rect 473078 41936 473142 41948
rect 462314 41908 473142 41936
rect 462314 41896 462378 41908
rect 465074 41896 465138 41908
rect 466362 41896 466426 41908
rect 469398 41896 469462 41908
rect 470686 41896 470750 41908
rect 473078 41896 473142 41908
rect 517054 41936 517118 41948
rect 519906 41936 519970 41948
rect 521194 41936 521258 41948
rect 524230 41936 524294 41948
rect 525518 41936 525582 41948
rect 527910 41936 527974 41948
rect 517054 41908 527974 41936
rect 517054 41896 517118 41908
rect 519906 41896 519970 41908
rect 521194 41896 521258 41908
rect 524230 41896 524294 41908
rect 525518 41896 525582 41908
rect 527910 41896 527974 41908
rect 146294 41868 146358 41880
rect 568850 41868 568914 41880
rect 579890 41868 579954 41880
rect 146294 41840 579954 41868
rect 146294 41828 146358 41840
rect 568850 41828 568914 41840
rect 579890 41828 579954 41840
rect 198918 41800 198982 41812
rect 307754 41800 307818 41812
rect 362494 41800 362558 41812
rect 168346 41772 380894 41800
rect 93762 41528 93826 41540
rect 168346 41528 168374 41772
rect 198918 41760 198982 41772
rect 307754 41760 307818 41772
rect 362494 41760 362558 41772
rect 93762 41500 168374 41528
rect 93762 41488 93826 41500
tri 239482 41369 239813 41700 se
rect 239813 41369 252469 41700
rect 135162 40236 135226 40248
rect 143534 40236 143598 40248
rect 135162 40208 143598 40236
rect 135162 40196 135226 40208
rect 143534 40196 143598 40208
rect 140990 40100 141054 40112
rect 143066 40100 143130 40112
rect 144546 40100 144610 40112
rect 146294 40100 146358 40112
rect 140990 40072 146358 40100
rect 140990 40060 141054 40072
rect 142586 40000 142614 40072
rect 143066 40060 143130 40072
rect 144546 40060 144610 40072
rect 146294 40060 146358 40072
rect 132600 39878 140940 39963
rect 140996 39934 141048 40000
rect 141104 39878 141313 39963
rect 141369 39934 141499 40000
rect 141555 39878 141898 39963
rect 141954 39934 142084 40000
rect 142140 39878 142517 39963
rect 79664 39616 91393 39806
rect 79664 39593 79892 39616
tri 79892 39593 79915 39616 nw
tri 91107 39593 91130 39616 ne
rect 91130 39593 91393 39616
rect 79076 55 93763 39593
rect 132600 37949 142517 39878
rect 142573 38005 142619 40000
rect 142675 39878 143012 39963
rect 143068 39934 143128 40000
rect 143184 39878 144517 39963
rect 144573 39934 144689 40000
rect 144745 39878 145035 39963
rect 145091 39934 145143 40000
rect 145199 39878 147600 39963
rect 142675 37949 147600 39878
rect 132600 20821 147600 37949
rect 186400 36103 202400 41369
rect 186377 34997 202400 36103
rect 186400 33976 202400 34997
rect 186377 32855 202400 33976
rect 186400 29756 202400 32855
tri 239013 40900 239482 41369 se
rect 239482 41300 252469 41369
tri 252469 41300 252869 41700 sw
rect 380866 41528 380894 41772
rect 417326 41800 417390 41812
rect 417252 41772 417390 41800
rect 417252 41528 417280 41772
rect 417326 41760 417390 41772
rect 472158 41800 472222 41812
rect 526714 41800 526778 41812
rect 472084 41772 472222 41800
rect 472084 41528 472112 41772
rect 472158 41760 472222 41772
rect 516106 41772 526778 41800
rect 516106 41528 516134 41772
rect 526714 41760 526778 41772
rect 380866 41500 516134 41528
rect 239482 40900 252869 41300
rect 239013 40196 252869 40900
rect 239013 39796 252469 40196
tri 252469 39796 252869 40196 nw
rect 239013 39756 252101 39796
rect 239013 32702 240960 39756
rect 244887 39600 252101 39756
rect 244887 39593 252869 39600
rect 238961 31928 241151 32702
rect 186377 28562 202400 29756
rect 186377 25414 202423 28562
tri 186377 25403 186388 25414 ne
rect 186388 23873 202423 25414
rect 186388 22050 202400 23873
rect 186388 21704 202429 22050
rect 186388 21084 202400 21704
rect 186400 20821 202400 21084
rect 132571 13956 147629 20821
rect 186371 13956 202423 20821
rect 132600 13745 147600 13956
rect 186400 13745 202400 13956
rect 132571 5982 147629 13745
rect 186371 5982 202423 13745
rect 132600 158 147600 5982
rect 186400 4220 202400 5982
rect 186396 3805 202400 4220
rect 186400 0 202400 3805
rect 241200 32 256176 39593
rect 295000 36103 311000 41369
rect 349800 36103 365800 41369
rect 404600 36103 420600 41369
rect 459400 36103 475400 41369
rect 514200 36103 530200 41369
rect 569864 39616 581593 39806
rect 569864 39593 570092 39616
tri 570092 39593 570115 39616 nw
tri 581307 39593 581330 39616 ne
rect 581330 39593 581593 39616
rect 623664 39616 635393 39806
rect 623664 39593 623892 39616
tri 623892 39593 623915 39616 nw
tri 635107 39593 635130 39616 ne
rect 635130 39593 635393 39616
rect 636029 39593 637075 39774
rect 294977 34997 311000 36103
rect 349777 34997 365800 36103
rect 404577 34997 420600 36103
rect 459377 34997 475400 36103
rect 514177 34997 530200 36103
rect 295000 33976 311000 34997
rect 349800 33976 365800 34997
rect 404600 33976 420600 34997
rect 459400 33976 475400 34997
rect 514200 33976 530200 34997
rect 294977 32855 311000 33976
rect 349777 32855 365800 33976
rect 404577 32855 420600 33976
rect 459377 32855 475400 33976
rect 514177 32855 530200 33976
rect 295000 29756 311000 32855
rect 349800 29756 365800 32855
rect 404600 29756 420600 32855
rect 459400 29756 475400 32855
rect 514200 29756 530200 32855
rect 294977 28562 311000 29756
rect 349777 28562 365800 29756
rect 404577 28562 420600 29756
rect 459377 28562 475400 29756
rect 514177 28562 530200 29756
rect 294977 25414 311023 28562
tri 294977 25403 294988 25414 ne
rect 294988 23873 311023 25414
rect 349777 25414 365823 28562
tri 349777 25403 349788 25414 ne
rect 349788 23873 365823 25414
rect 404577 25414 420623 28562
tri 404577 25403 404588 25414 ne
rect 404588 23873 420623 25414
rect 459377 25414 475423 28562
tri 459377 25403 459388 25414 ne
rect 459388 23873 475423 25414
rect 514177 25414 530223 28562
tri 514177 25403 514188 25414 ne
rect 514188 23873 530223 25414
rect 294988 22050 311000 23873
rect 349788 22050 365800 23873
rect 404588 22050 420600 23873
rect 459388 22050 475400 23873
rect 514188 22050 530200 23873
rect 294988 21704 311029 22050
rect 349788 21704 365829 22050
rect 404588 21704 420629 22050
rect 459388 21704 475429 22050
rect 514188 21704 530229 22050
rect 294988 21084 311000 21704
rect 349788 21084 365800 21704
rect 404588 21084 420600 21704
rect 459388 21084 475400 21704
rect 514188 21084 530200 21704
rect 295000 20821 311000 21084
rect 349800 20821 365800 21084
rect 404600 20821 420600 21084
rect 459400 20821 475400 21084
rect 514200 20821 530200 21084
rect 294971 13956 311023 20821
rect 349771 13956 365823 20821
rect 404571 13956 420623 20821
rect 459371 13956 475423 20821
rect 514171 13956 530223 20821
rect 295000 13745 311000 13956
rect 349800 13745 365800 13956
rect 404600 13745 420600 13956
rect 459400 13745 475400 13956
rect 514200 13745 530200 13956
rect 294971 5982 311023 13745
rect 349771 5982 365823 13745
rect 404571 5982 420623 13745
rect 459371 5982 475423 13745
rect 514171 5982 530223 13745
rect 295000 4220 311000 5982
rect 349800 4220 365800 5982
rect 404600 4220 420600 5982
rect 459400 4220 475400 5982
rect 514200 4220 530200 5982
rect 294996 3805 311000 4220
rect 349796 3805 365800 4220
rect 404596 3805 420600 4220
rect 459396 3805 475400 4220
rect 514196 3805 530200 4220
rect 295000 0 311000 3805
rect 349800 0 365800 3805
rect 404600 0 420600 3805
rect 459400 0 475400 3805
rect 514200 0 530200 3805
rect 569276 55 583963 39593
rect 623217 55 637763 39593
<< metal2 >>
rect 229499 997600 234279 998011
rect 239478 997600 244258 1002732
rect 280899 997600 285679 998011
rect 290878 997600 295658 1002732
rect 41713 800217 42193 800273
rect 41713 798377 42193 798433
rect 41713 797733 42193 797789
rect 41713 796537 42193 796593
rect 41713 795893 42193 795949
rect 41713 795341 42193 795397
rect 41713 794697 42193 794753
rect 41713 794053 42193 794109
rect 41713 793501 42193 793557
rect 41722 792269 42288 792282
rect 41713 792254 42288 792269
rect 41713 792213 42193 792254
rect 41713 791017 42193 791073
rect 41713 790373 42193 790429
rect 41713 789729 42193 789785
rect 41713 789177 42193 789233
rect 42260 788066 42288 792254
rect 41892 788050 42288 788066
rect 41892 788044 42300 788050
rect 41892 788038 42248 788044
rect 41892 787945 41920 788038
rect 42248 787986 42300 787992
rect 42260 787955 42288 787986
rect 41713 787889 42193 787945
rect 41713 787337 42193 787393
rect 41713 786693 42193 786749
rect 41713 786049 42193 786105
rect 41713 785497 42193 785553
rect 41713 757017 42193 757073
rect 41713 755177 42193 755233
rect 41713 754533 42193 754589
rect 41713 753337 42193 753393
rect 41713 752693 42193 752749
rect 41713 752141 42193 752197
rect 41713 751497 42193 751553
rect 41713 750853 42193 750909
rect 41713 750301 42193 750357
rect 42432 788044 42484 788050
rect 42432 787986 42484 787992
rect 42444 749578 42472 787986
rect 41800 749550 42472 749578
rect 41800 749069 41828 749550
rect 41713 749013 42193 749069
rect 41722 749006 41828 749013
rect 41713 747817 42193 747873
rect 41713 747173 42193 747229
rect 41713 746529 42193 746585
rect 41713 745977 42193 746033
rect 41713 744731 42193 744745
rect 42260 744731 42288 749550
rect 41713 744703 42288 744731
rect 41713 744689 42193 744703
rect 41713 744137 42193 744193
rect 41713 743493 42193 743549
rect 41713 742849 42193 742905
rect 41713 742297 42193 742353
rect 42260 728654 42288 744703
rect 42260 728626 42380 728654
rect 41713 713817 42193 713873
rect 41713 711977 42193 712033
rect 41713 711333 42193 711389
rect 41713 710137 42193 710193
rect 41713 709493 42193 709549
rect 41713 708941 42193 708997
rect 41713 708297 42193 708353
rect 41713 707653 42193 707709
rect 41713 707101 42193 707157
rect 41713 705855 42193 705869
rect 42352 705855 42380 728626
rect 41713 705827 42380 705855
rect 41713 705813 42193 705827
rect 41713 704617 42193 704673
rect 41713 703973 42193 704029
rect 41713 703329 42193 703385
rect 41713 702777 42193 702833
rect 41713 701489 42193 701545
rect 41892 701434 41920 701489
rect 42260 701434 42288 705827
rect 673736 855432 673788 855438
rect 673736 855374 673788 855380
rect 673748 773362 673776 855374
rect 673736 773356 673788 773362
rect 673736 773298 673788 773304
rect 673736 769140 673788 769146
rect 673736 769082 673788 769088
rect 673748 728618 673776 769082
rect 673736 728612 673788 728618
rect 673736 728554 673788 728560
rect 673460 724056 673512 724062
rect 673460 723998 673512 724004
rect 41892 701406 42288 701434
rect 41713 700937 42193 700993
rect 41713 700293 42193 700349
rect 41713 699649 42193 699705
rect 41713 699097 42193 699153
rect 42260 690014 42288 701406
rect 42260 689986 42380 690014
rect 41713 670417 42193 670473
rect 41713 668577 42193 668633
rect 41713 667933 42193 667989
rect 41713 666737 42193 666793
rect 41713 666093 42193 666149
rect 41713 665541 42193 665597
rect 41713 664897 42193 664953
rect 41713 664253 42193 664309
rect 41713 663701 42193 663757
rect 42352 662538 42380 689986
rect 41892 662510 42380 662538
rect 41892 662469 41920 662510
rect 41713 662413 42193 662469
rect 41713 661217 42193 661273
rect 41713 660573 42193 660629
rect 41713 659929 42193 659985
rect 41713 659377 42193 659433
rect 41713 658131 42193 658145
rect 42260 658131 42288 662510
rect 673472 684350 673500 723998
rect 673460 684344 673512 684350
rect 673460 684286 673512 684292
rect 41713 658103 42288 658131
rect 41713 658089 42193 658103
rect 41713 657537 42193 657593
rect 41713 656893 42193 656949
rect 41713 656249 42193 656305
rect 41713 655697 42193 655753
rect 42260 651374 42288 658103
rect 42260 651346 42380 651374
rect 41713 627217 42193 627273
rect 41713 625377 42193 625433
rect 41713 624733 42193 624789
rect 41713 623537 42193 623593
rect 41713 622893 42193 622949
rect 41713 622341 42193 622397
rect 41713 621697 42193 621753
rect 41713 621053 42193 621109
rect 41713 620501 42193 620557
rect 41713 619213 42193 619269
rect 41892 619154 41920 619213
rect 42352 619154 42380 651346
rect 41892 619126 42380 619154
rect 41713 618017 42193 618073
rect 41713 617373 42193 617429
rect 41713 616729 42193 616785
rect 41713 616177 42193 616233
rect 41713 614889 42193 614945
rect 41800 614802 41828 614889
rect 42260 614802 42288 619126
rect 41800 614774 42380 614802
rect 41713 614337 42193 614393
rect 41713 613693 42193 613749
rect 41713 613049 42193 613105
rect 41713 612497 42193 612553
rect 42352 604454 42380 614774
rect 42352 604426 42472 604454
rect 41713 584017 42193 584073
rect 41713 582177 42193 582233
rect 41713 581533 42193 581589
rect 41713 580337 42193 580393
rect 41713 579693 42193 579749
rect 41713 579141 42193 579197
rect 41713 578497 42193 578553
rect 41713 577853 42193 577909
rect 41713 577301 42193 577357
rect 41788 576564 41840 576570
rect 41788 576506 41840 576512
rect 42248 576564 42300 576570
rect 42248 576506 42300 576512
rect 41800 576069 41828 576506
rect 41713 576013 42193 576069
rect 41713 574817 42193 574873
rect 41713 574173 42193 574229
rect 41713 573529 42193 573585
rect 41713 572977 42193 573033
rect 41713 571731 42193 571745
rect 42260 571731 42288 576506
rect 42444 576570 42472 604426
rect 42432 576564 42484 576570
rect 42432 576506 42484 576512
rect 673828 680128 673880 680134
rect 673828 680070 673880 680076
rect 673840 640150 673868 680070
rect 673828 640144 673880 640150
rect 673828 640086 673880 640092
rect 673736 635792 673788 635798
rect 673736 635734 673788 635740
rect 673748 596154 673776 635734
rect 673736 596148 673788 596154
rect 673736 596090 673788 596096
rect 41713 571703 42380 571731
rect 41713 571689 42193 571703
rect 41713 571137 42193 571193
rect 41713 570493 42193 570549
rect 41713 569849 42193 569905
rect 41713 569297 42193 569353
rect 41713 540817 42193 540873
rect 41713 538977 42193 539033
rect 41713 538333 42193 538389
rect 41713 537137 42193 537193
rect 41713 536493 42193 536549
rect 41713 535941 42193 535997
rect 41713 535297 42193 535353
rect 41713 534653 42193 534709
rect 41713 534101 42193 534157
rect 41713 532855 42193 532869
rect 42352 532855 42380 571703
rect 41713 532827 42380 532855
rect 41713 532813 42193 532827
rect 41713 531617 42193 531673
rect 41713 530973 42193 531029
rect 41713 530329 42193 530385
rect 41713 529777 42193 529833
rect 41713 528489 42193 528545
rect 41892 528442 41920 528489
rect 42260 528442 42288 532827
rect 673736 590844 673788 590850
rect 673736 590786 673788 590792
rect 673748 551546 673776 590786
rect 673736 551540 673788 551546
rect 673736 551482 673788 551488
rect 673460 547052 673512 547058
rect 673460 546994 673512 547000
rect 41892 528414 42288 528442
rect 41713 527937 42193 527993
rect 41713 527293 42193 527349
rect 41713 526649 42193 526705
rect 41713 526097 42193 526153
rect 42260 419534 42288 528414
rect 42260 419506 42380 419534
rect 41713 413017 42193 413073
rect 41713 411177 42193 411233
rect 41713 410533 42193 410589
rect 41713 409337 42193 409393
rect 41713 408693 42193 408749
rect 41713 408141 42193 408197
rect 41713 407497 42193 407553
rect 41713 406853 42193 406909
rect 41713 406301 42193 406357
rect 42352 405498 42380 419506
rect 41800 405470 42380 405498
rect 41800 405069 41828 405470
rect 41713 405013 42193 405069
rect 41713 403817 42193 403873
rect 41713 403173 42193 403229
rect 41713 402529 42193 402585
rect 41713 401977 42193 402033
rect 41713 400738 42193 400745
rect 42260 400738 42288 405470
rect 41713 400710 42288 400738
rect 41713 400689 42193 400710
rect 41713 400137 42193 400193
rect 41713 399493 42193 399549
rect 41713 398849 42193 398905
rect 41713 398297 42193 398353
rect 42260 380894 42288 400710
rect 42260 380866 42380 380894
rect 41713 369817 42193 369873
rect 41713 367977 42193 368033
rect 41713 367333 42193 367389
rect 41713 366137 42193 366193
rect 41713 365493 42193 365549
rect 41713 364941 42193 364997
rect 41713 364297 42193 364353
rect 41713 363653 42193 363709
rect 41713 363101 42193 363157
rect 41713 361813 42193 361869
rect 41800 361574 41828 361813
rect 42352 361574 42380 380866
rect 41800 361546 42380 361574
rect 41713 360617 42193 360673
rect 41713 359973 42193 360029
rect 41713 359329 42193 359385
rect 41713 358777 42193 358833
rect 41713 357531 42193 357545
rect 42260 357531 42288 361546
rect 41713 357503 42380 357531
rect 41713 357489 42193 357503
rect 41713 356937 42193 356993
rect 41713 356293 42193 356349
rect 41713 355649 42193 355705
rect 41713 355097 42193 355153
rect 41713 326417 42193 326473
rect 41713 324577 42193 324633
rect 41713 323933 42193 323989
rect 41713 322737 42193 322793
rect 41713 322093 42193 322149
rect 41713 321541 42193 321597
rect 41713 320897 42193 320953
rect 41713 320253 42193 320309
rect 41713 319701 42193 319757
rect 41713 318413 42193 318469
rect 41892 318322 41920 318413
rect 42352 318322 42380 357503
rect 673472 380894 673500 546994
rect 677600 954121 678011 958901
rect 677600 944142 682732 948922
rect 675407 862647 675887 862703
rect 675407 862095 675887 862151
rect 675407 861451 675887 861507
rect 675407 860807 675887 860863
rect 675407 860282 675887 860311
rect 675312 860255 675887 860282
rect 675312 860254 675418 860255
rect 675312 855973 675340 860254
rect 675407 858967 675887 859023
rect 675407 858415 675887 858471
rect 675407 857771 675887 857827
rect 675407 857127 675887 857183
rect 675407 855973 675887 855987
rect 675312 855945 675887 855973
rect 675404 855931 675887 855945
rect 675404 855438 675432 855931
rect 675392 855432 675444 855438
rect 675392 855374 675444 855380
rect 675407 854643 675887 854699
rect 675407 854091 675887 854147
rect 675407 853447 675887 853503
rect 675407 852803 675887 852859
rect 675407 852251 675887 852307
rect 675407 851607 675887 851663
rect 675407 850411 675887 850467
rect 675407 849767 675887 849823
rect 675407 847927 675887 847983
rect 675208 773356 675260 773362
rect 675208 773298 675260 773304
rect 675220 769146 675248 773298
rect 675208 769140 675260 769146
rect 675208 769082 675260 769088
rect 675407 775247 675887 775303
rect 675407 774695 675887 774751
rect 675407 774051 675887 774107
rect 675407 773407 675887 773463
rect 675392 773356 675444 773362
rect 675392 773298 675444 773304
rect 675404 772911 675432 773298
rect 675404 772883 675887 772911
rect 675407 772855 675887 772883
rect 675407 771567 675887 771623
rect 675407 771015 675887 771071
rect 675407 770371 675887 770427
rect 675407 769727 675887 769783
rect 675392 769140 675444 769146
rect 675392 769082 675444 769088
rect 675404 768587 675432 769082
rect 675404 768559 675887 768587
rect 675407 768531 675887 768559
rect 675407 767243 675887 767299
rect 675407 766691 675887 766747
rect 675407 766047 675887 766103
rect 675407 765403 675887 765459
rect 675407 764851 675887 764907
rect 675407 764207 675887 764263
rect 675407 763011 675887 763067
rect 675407 762367 675887 762423
rect 675407 760527 675887 760583
rect 675407 730847 675887 730903
rect 675407 730295 675887 730351
rect 675407 729651 675887 729707
rect 675407 729007 675887 729063
rect 675392 728612 675444 728618
rect 675392 728554 675444 728560
rect 675404 728511 675432 728554
rect 675404 728498 675887 728511
rect 675312 728470 675887 728498
rect 675312 724690 675340 728470
rect 675407 728455 675887 728470
rect 675407 727167 675887 727223
rect 675407 726615 675887 726671
rect 675407 725971 675887 726027
rect 675407 725327 675887 725383
rect 675312 724662 675432 724690
rect 675404 724187 675432 724662
rect 675404 724131 675887 724187
rect 675404 724062 675432 724131
rect 675392 724056 675444 724062
rect 675392 723998 675444 724004
rect 675407 722843 675887 722899
rect 675407 722291 675887 722347
rect 675407 721647 675887 721703
rect 675407 721003 675887 721059
rect 675407 720451 675887 720507
rect 675407 719807 675887 719863
rect 675407 718611 675887 718667
rect 675407 717967 675887 718023
rect 675407 716127 675887 716183
rect 675407 686647 675887 686703
rect 675407 686095 675887 686151
rect 675407 685451 675887 685507
rect 675407 684807 675887 684863
rect 675312 684350 675340 684381
rect 675300 684344 675352 684350
rect 675407 684298 675887 684311
rect 675352 684292 675887 684298
rect 675300 684286 675887 684292
rect 675312 684270 675887 684286
rect 675312 680354 675340 684270
rect 675407 684255 675887 684270
rect 675407 682967 675887 683023
rect 675407 682415 675887 682471
rect 675407 681771 675887 681827
rect 675407 681127 675887 681183
rect 675312 680326 675432 680354
rect 675404 680134 675432 680326
rect 675392 680128 675444 680134
rect 675392 680070 675444 680076
rect 675404 679987 675432 680070
rect 675404 679932 675887 679987
rect 675407 679931 675887 679932
rect 675407 678643 675887 678699
rect 675407 678091 675887 678147
rect 675407 677447 675887 677503
rect 675407 676803 675887 676859
rect 675407 676251 675887 676307
rect 675407 675607 675887 675663
rect 675407 674411 675887 674467
rect 675407 673767 675887 673823
rect 675407 671927 675887 671983
rect 675407 642447 675887 642503
rect 675407 641895 675887 641951
rect 675407 641251 675887 641307
rect 675407 640607 675887 640663
rect 675312 640150 675340 640181
rect 675300 640144 675352 640150
rect 675407 640098 675887 640111
rect 675352 640092 675887 640098
rect 675300 640086 675887 640092
rect 675312 640070 675887 640086
rect 675312 635882 675340 640070
rect 675407 640055 675887 640070
rect 675407 638767 675887 638823
rect 675407 638215 675887 638271
rect 675407 637571 675887 637627
rect 675407 636927 675887 636983
rect 675312 635854 675432 635882
rect 675312 635798 675340 635854
rect 675300 635792 675352 635798
rect 675300 635734 675352 635740
rect 675404 635787 675432 635854
rect 675404 635732 675887 635787
rect 675407 635731 675887 635732
rect 675407 634443 675887 634499
rect 675407 633891 675887 633947
rect 675407 633247 675887 633303
rect 675407 632603 675887 632659
rect 675407 632051 675887 632107
rect 675407 631407 675887 631463
rect 675407 630211 675887 630267
rect 675407 629567 675887 629623
rect 675407 627727 675887 627783
rect 675208 596148 675260 596154
rect 675208 596090 675260 596096
rect 675220 590850 675248 596090
rect 675208 590844 675260 590850
rect 675208 590786 675260 590792
rect 675407 598047 675887 598103
rect 675407 597495 675887 597551
rect 675407 596851 675887 596907
rect 675407 596207 675887 596263
rect 675392 596148 675444 596154
rect 675392 596090 675444 596096
rect 675404 595711 675432 596090
rect 675404 595683 675887 595711
rect 675407 595655 675887 595683
rect 675407 594367 675887 594423
rect 675407 593815 675887 593871
rect 675407 593171 675887 593227
rect 675407 592527 675887 592583
rect 675407 591359 675887 591387
rect 675404 591331 675887 591359
rect 675404 590850 675432 591331
rect 675392 590844 675444 590850
rect 675392 590786 675444 590792
rect 675407 590043 675887 590099
rect 675407 589491 675887 589547
rect 675407 588847 675887 588903
rect 675407 588203 675887 588259
rect 675407 587651 675887 587707
rect 675407 587007 675887 587063
rect 675407 585811 675887 585867
rect 675407 585167 675887 585223
rect 675407 583327 675887 583383
rect 675407 553847 675887 553903
rect 675407 553295 675887 553351
rect 675407 552651 675887 552707
rect 675407 552007 675887 552063
rect 675220 551546 675248 551580
rect 675208 551540 675260 551546
rect 675407 551497 675887 551511
rect 675260 551488 675887 551497
rect 675208 551482 675887 551488
rect 675220 551469 675887 551482
rect 675220 547058 675248 551469
rect 675407 551455 675887 551469
rect 675407 550167 675887 550223
rect 675407 549615 675887 549671
rect 675407 548971 675887 549027
rect 675407 548327 675887 548383
rect 675407 547159 675887 547187
rect 675404 547131 675887 547159
rect 675404 547058 675432 547131
rect 675208 547052 675260 547058
rect 675208 546994 675260 547000
rect 675392 547052 675444 547058
rect 675392 546994 675444 547000
rect 675407 545843 675887 545899
rect 675407 545291 675887 545347
rect 675407 544647 675887 544703
rect 675407 544003 675887 544059
rect 675407 543451 675887 543507
rect 675407 542807 675887 542863
rect 675407 541611 675887 541667
rect 675407 540967 675887 541023
rect 675407 539127 675887 539183
rect 673472 380866 673592 380894
rect 673564 372842 673592 380866
rect 675407 379647 675887 379703
rect 675407 379095 675887 379151
rect 675407 378451 675887 378507
rect 675407 377807 675887 377863
rect 675407 377297 675887 377311
rect 675312 377269 675887 377297
rect 673552 372836 673604 372842
rect 673552 372778 673604 372784
rect 41892 318294 42380 318322
rect 41713 317217 42193 317273
rect 41713 316573 42193 316629
rect 41713 315929 42193 315985
rect 41713 315377 42193 315433
rect 41713 314089 42193 314145
rect 41722 314078 41920 314089
rect 41892 313970 41920 314078
rect 42260 313970 42288 318294
rect 41892 313942 42288 313970
rect 41713 313537 42193 313593
rect 42260 313138 42288 313942
rect 42248 313132 42300 313138
rect 42248 313074 42300 313080
rect 41713 312893 42193 312949
rect 41713 312249 42193 312305
rect 41713 311697 42193 311753
rect 42340 312928 42392 312934
rect 42340 312870 42392 312876
rect 42352 284170 42380 312870
rect 42340 284164 42392 284170
rect 42340 284106 42392 284112
rect 42340 283960 42392 283966
rect 42340 283902 42392 283908
rect 41713 283217 42193 283273
rect 41713 281377 42193 281433
rect 41713 280733 42193 280789
rect 41713 279537 42193 279593
rect 41713 278893 42193 278949
rect 41713 278341 42193 278397
rect 41713 277697 42193 277753
rect 41713 277053 42193 277109
rect 41713 276501 42193 276557
rect 42352 275346 42380 283902
rect 41800 275318 42380 275346
rect 41800 275269 41828 275318
rect 41713 275213 42193 275269
rect 41713 274017 42193 274073
rect 41713 273373 42193 273429
rect 41713 272729 42193 272785
rect 41713 272177 42193 272233
rect 41713 270931 42193 270945
rect 42260 270931 42288 275318
rect 673564 333130 673592 372778
rect 673552 333124 673604 333130
rect 673552 333066 673604 333072
rect 675312 372858 675340 377269
rect 675407 377255 675887 377269
rect 675407 375967 675887 376023
rect 675407 375415 675887 375471
rect 675407 374771 675887 374827
rect 675407 374127 675887 374183
rect 675407 372980 675887 372987
rect 675404 372931 675887 372980
rect 675404 372858 675432 372931
rect 675312 372842 675432 372858
rect 675312 372836 675444 372842
rect 675312 372830 675392 372836
rect 675392 372778 675444 372784
rect 41713 270903 42288 270931
rect 41713 270889 42193 270903
rect 41713 270337 42193 270393
rect 41713 269693 42193 269749
rect 41713 269049 42193 269105
rect 41713 268497 42193 268553
rect 42260 264974 42288 270903
rect 42260 264946 42380 264974
rect 41713 240017 42193 240073
rect 41713 238177 42193 238233
rect 41713 236337 42193 236393
rect 41713 235141 42193 235197
rect 41713 234497 42193 234553
rect 41713 233853 42193 233909
rect 41713 233301 42193 233357
rect 42352 232506 42380 264946
rect 41800 232478 42380 232506
rect 41800 232069 41828 232478
rect 41713 232013 42193 232069
rect 41713 230817 42193 230873
rect 41713 230173 42193 230229
rect 41713 229529 42193 229585
rect 41713 228977 42193 229033
rect 42260 227882 42288 232478
rect 41800 227854 42288 227882
rect 41800 227746 41828 227854
rect 41722 227745 41828 227746
rect 41713 227689 42193 227745
rect 41713 227137 42193 227193
rect 41713 226493 42193 226549
rect 42260 226334 42288 227854
rect 42260 226306 42380 226334
rect 41713 225849 42193 225905
rect 41713 225297 42193 225353
rect 41713 196817 42193 196873
rect 41713 194977 42193 195033
rect 41713 193137 42193 193193
rect 41713 191941 42193 191997
rect 41713 191297 42193 191353
rect 41713 190653 42193 190709
rect 41713 190101 42193 190157
rect 42352 188986 42380 226306
rect 673736 328296 673788 328302
rect 673736 328238 673788 328244
rect 41892 188958 42380 188986
rect 41892 188869 41920 188958
rect 41713 188813 42193 188869
rect 41713 187617 42193 187673
rect 41713 186973 42193 187029
rect 41713 186329 42193 186385
rect 41713 185777 42193 185833
rect 41713 184531 42193 184545
rect 42260 184531 42288 188958
rect 41713 184503 42380 184531
rect 41713 184489 42193 184503
rect 41713 183937 42193 183993
rect 41713 183293 42193 183349
rect 41713 182649 42193 182705
rect 41713 182097 42193 182153
rect 42352 45626 42380 184503
rect 673748 289338 673776 328238
rect 675407 371643 675887 371699
rect 675407 371091 675887 371147
rect 675407 370447 675887 370503
rect 675407 369803 675887 369859
rect 675407 368607 675887 368663
rect 675407 366767 675887 366823
rect 675407 364927 675887 364983
rect 675407 335447 675887 335503
rect 675407 334895 675887 334951
rect 675407 334251 675887 334307
rect 675407 333607 675887 333663
rect 675312 333130 675340 333180
rect 675300 333124 675352 333130
rect 675407 333097 675887 333111
rect 675352 333072 675887 333097
rect 675300 333069 675887 333072
rect 675300 333066 675352 333069
rect 675312 328658 675340 333066
rect 675407 333055 675887 333069
rect 675407 331767 675887 331823
rect 675407 331215 675887 331271
rect 675407 330571 675887 330627
rect 675407 329927 675887 329983
rect 675407 328780 675887 328787
rect 675404 328731 675887 328780
rect 675404 328658 675432 328731
rect 675312 328630 675432 328658
rect 675404 328302 675432 328630
rect 675392 328296 675444 328302
rect 675392 328238 675444 328244
rect 675407 327443 675887 327499
rect 675407 326891 675887 326947
rect 675407 326247 675887 326303
rect 675407 325603 675887 325659
rect 675407 324407 675887 324463
rect 675407 322567 675887 322623
rect 675407 320727 675887 320783
rect 675407 291247 675887 291303
rect 675407 290695 675887 290751
rect 675407 290051 675887 290107
rect 675407 289407 675887 289463
rect 673736 289332 673788 289338
rect 673736 289274 673788 289280
rect 675392 289332 675444 289338
rect 675392 289274 675444 289280
rect 675404 288911 675432 289274
rect 675404 288897 675887 288911
rect 675312 288869 675887 288897
rect 675312 285138 675340 288869
rect 675407 288855 675887 288869
rect 675407 287567 675887 287623
rect 675407 287015 675887 287071
rect 675407 286371 675887 286427
rect 675407 285727 675887 285783
rect 675312 285110 675432 285138
rect 675404 284587 675432 285110
rect 675404 284531 675887 284587
rect 675404 284102 675432 284531
rect 673736 284096 673788 284102
rect 673736 284038 673788 284044
rect 675392 284096 675444 284102
rect 675392 284038 675444 284044
rect 673748 244662 673776 284038
rect 675407 283243 675887 283299
rect 675407 282691 675887 282747
rect 675407 282047 675887 282103
rect 675407 281403 675887 281459
rect 675407 280207 675887 280263
rect 675407 278367 675887 278423
rect 675407 276527 675887 276583
rect 675407 246847 675887 246903
rect 675407 246295 675887 246351
rect 675407 245651 675887 245707
rect 675407 245007 675887 245063
rect 673736 244656 673788 244662
rect 673736 244598 673788 244604
rect 675392 244656 675444 244662
rect 675392 244598 675444 244604
rect 675404 244511 675432 244598
rect 675404 244455 675887 244511
rect 675404 243930 675432 244455
rect 675312 243902 675432 243930
rect 675312 240173 675340 243902
rect 675407 243167 675887 243223
rect 675407 242615 675887 242671
rect 675407 241971 675887 242027
rect 675407 241327 675887 241383
rect 675407 240173 675887 240187
rect 675312 240145 675887 240173
rect 675404 240131 675887 240145
rect 675404 239698 675432 240131
rect 673736 239692 673788 239698
rect 673736 239634 673788 239640
rect 675392 239692 675444 239698
rect 675392 239634 675444 239640
rect 673748 200462 673776 239634
rect 675407 238843 675887 238899
rect 675407 238291 675887 238347
rect 675407 237647 675887 237703
rect 675407 237003 675887 237059
rect 675407 235807 675887 235863
rect 675407 233967 675887 234023
rect 675407 232127 675887 232183
rect 675407 202647 675887 202703
rect 675407 202095 675887 202151
rect 675407 201451 675887 201507
rect 675407 200807 675887 200863
rect 673736 200456 673788 200462
rect 673736 200398 673788 200404
rect 675392 200456 675444 200462
rect 675392 200398 675444 200404
rect 675404 200311 675432 200398
rect 675404 200255 675887 200311
rect 675404 199730 675432 200255
rect 675312 199702 675432 199730
rect 675312 195973 675340 199702
rect 675407 198967 675887 199023
rect 675407 198415 675887 198471
rect 675407 197771 675887 197827
rect 675407 197127 675887 197183
rect 675407 195973 675887 195987
rect 675312 195945 675887 195973
rect 675404 195931 675887 195945
rect 675404 195838 675432 195931
rect 673736 195832 673788 195838
rect 673736 195774 673788 195780
rect 675392 195832 675444 195838
rect 675392 195774 675444 195780
rect 42340 45620 42392 45626
rect 42340 45562 42392 45568
rect 527456 46912 527508 46918
rect 527456 46854 527508 46860
rect 143632 45620 143684 45626
rect 143632 45562 143684 45568
rect 143644 44198 143672 45562
rect 143632 44192 143684 44198
rect 143632 44134 143684 44140
rect 145104 44192 145156 44198
rect 145104 44134 145156 44140
rect 145116 40202 145144 44134
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 195336 44192 195388 44198
rect 195336 44134 195388 44140
rect 195348 42193 195376 44134
rect 199844 44260 199896 44266
rect 199844 44202 199896 44208
rect 199660 44192 199712 44198
rect 199856 44146 199884 44202
rect 199712 44140 199884 44146
rect 199660 44134 199884 44140
rect 199672 44118 199884 44134
rect 199672 42193 199700 44118
rect 187327 41713 187383 42193
rect 194043 41713 194099 42193
rect 195331 41713 195387 42193
rect 199655 41713 199711 42193
rect 145091 39706 145143 40000
rect 303896 44260 303948 44266
rect 303896 44202 303948 44208
rect 303908 42193 303936 44202
rect 308220 44260 308272 44266
rect 308220 44202 308272 44208
rect 308232 42193 308260 44202
rect 358728 44260 358780 44266
rect 358728 44202 358780 44208
rect 358740 42193 358768 44202
rect 363052 44328 363104 44334
rect 363052 44270 363104 44276
rect 363064 42193 363092 44270
rect 411074 44432 411130 44441
rect 411074 44367 411130 44376
rect 411088 42193 411116 44367
rect 413560 44328 413612 44334
rect 413560 44270 413612 44276
rect 413572 42193 413600 44270
rect 417884 44328 417936 44334
rect 417884 44270 417936 44276
rect 417896 42193 417924 44270
rect 419722 44296 419778 44305
rect 419722 44231 419778 44240
rect 419736 42193 419764 44231
rect 465814 44432 465870 44441
rect 465814 44367 465870 44376
rect 465828 42193 465856 44367
rect 468300 44328 468352 44334
rect 468300 44270 468352 44276
rect 468312 42193 468340 44270
rect 472624 44328 472676 44334
rect 472624 44270 472676 44276
rect 472636 42193 472664 44270
rect 474462 44432 474518 44441
rect 474462 44367 474518 44376
rect 474476 42193 474504 44367
rect 518806 44296 518862 44305
rect 518806 44231 518862 44240
rect 518820 42193 518848 44231
rect 523132 44192 523184 44198
rect 523132 44134 523184 44140
rect 523144 42193 523172 44134
rect 524970 44296 525026 44305
rect 524970 44231 525026 44240
rect 524984 42193 525012 44231
rect 527468 44198 527496 46854
rect 527456 44192 527508 44198
rect 527456 44134 527508 44140
rect 527468 42193 527496 44134
rect 673748 156330 673776 195774
rect 675407 194643 675887 194699
rect 675407 194091 675887 194147
rect 675407 193447 675887 193503
rect 675407 192803 675887 192859
rect 675407 191607 675887 191663
rect 675407 189767 675887 189823
rect 675407 187927 675887 187983
rect 675407 158447 675887 158503
rect 675407 157895 675887 157951
rect 675407 157251 675887 157307
rect 675407 156607 675887 156663
rect 673736 156324 673788 156330
rect 673736 156266 673788 156272
rect 675392 156324 675444 156330
rect 675392 156266 675444 156272
rect 675404 156210 675432 156266
rect 675312 156182 675432 156210
rect 673828 151768 673880 151774
rect 673828 151710 673880 151716
rect 673644 107364 673696 107370
rect 673644 107306 673696 107312
rect 673656 46986 673684 107306
rect 673840 111858 673868 151710
rect 673828 111852 673880 111858
rect 673828 111794 673880 111800
rect 675312 151774 675340 156182
rect 675404 156111 675432 156182
rect 675404 156060 675887 156111
rect 675407 156055 675887 156060
rect 675407 154767 675887 154823
rect 675407 154215 675887 154271
rect 675407 153571 675887 153627
rect 675407 152927 675887 152983
rect 675300 151773 675352 151774
rect 675407 151773 675887 151787
rect 675300 151768 675887 151773
rect 675352 151745 675887 151768
rect 675407 151731 675887 151745
rect 675300 151710 675352 151716
rect 675312 151662 675340 151710
rect 675407 150443 675887 150499
rect 675407 149891 675887 149947
rect 675407 149247 675887 149303
rect 675407 148603 675887 148659
rect 675407 147407 675887 147463
rect 675407 145567 675887 145623
rect 675407 143727 675887 143783
rect 675407 114047 675887 114103
rect 675407 113495 675887 113551
rect 675407 112851 675887 112907
rect 675407 112207 675887 112263
rect 675392 111852 675444 111858
rect 675392 111794 675444 111800
rect 675404 111711 675432 111794
rect 675404 111697 675887 111711
rect 675312 111669 675887 111697
rect 675312 107386 675340 111669
rect 675407 111655 675887 111669
rect 675407 110367 675887 110423
rect 675407 109815 675887 109871
rect 675407 109171 675887 109227
rect 675407 108527 675887 108583
rect 675407 107386 675887 107387
rect 675312 107370 675887 107386
rect 675300 107364 675887 107370
rect 675352 107358 675887 107364
rect 675407 107331 675887 107358
rect 675300 107306 675352 107312
rect 675312 107275 675340 107306
rect 673644 46980 673696 46986
rect 673644 46922 673696 46928
rect 675407 106043 675887 106099
rect 675407 105491 675887 105547
rect 675407 104847 675887 104903
rect 675407 104203 675887 104259
rect 675407 103007 675887 103063
rect 675407 101167 675887 101223
rect 675407 99327 675887 99383
rect 302643 41713 302699 42193
rect 303908 41806 303987 42193
rect 303931 41713 303987 41806
rect 306967 41713 307023 42193
rect 308232 41806 308311 42193
rect 308255 41713 308311 41806
rect 310095 41713 310151 42193
rect 357443 41713 357499 42193
rect 358731 41713 358787 42193
rect 361767 41713 361823 42193
rect 363055 41713 363111 42193
rect 364895 41713 364951 42193
rect 405527 41713 405583 42193
rect 409207 41834 409263 42193
rect 409207 41818 409368 41834
rect 409207 41812 409380 41818
rect 409207 41806 409328 41812
rect 409207 41713 409263 41806
rect 409328 41754 409380 41760
rect 411047 41820 411116 42193
rect 411047 41713 411103 41820
rect 412243 41834 412299 42193
rect 412243 41818 412404 41834
rect 413531 41820 413600 42193
rect 415371 41834 415427 42193
rect 412243 41812 412416 41818
rect 412243 41806 412364 41812
rect 412243 41713 412299 41806
rect 412364 41754 412416 41760
rect 413531 41713 413587 41820
rect 415228 41818 415427 41834
rect 415216 41812 415427 41818
rect 415268 41806 415427 41812
rect 415216 41754 415268 41760
rect 415371 41713 415427 41806
rect 416567 41713 416623 42193
rect 417855 41820 417924 42193
rect 419695 41820 419764 42193
rect 417855 41713 417911 41820
rect 419695 41713 419751 41820
rect 460327 41713 460383 42193
rect 464007 41834 464063 42193
rect 464007 41818 464200 41834
rect 464007 41812 464212 41818
rect 464007 41806 464160 41812
rect 464007 41713 464063 41806
rect 464160 41754 464212 41760
rect 465828 41806 465903 42193
rect 465847 41713 465903 41806
rect 467043 41834 467099 42193
rect 467043 41818 467236 41834
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 467043 41713 467099 41806
rect 468312 41806 468387 42193
rect 470171 41834 470227 42193
rect 470060 41818 470227 41834
rect 467196 41754 467248 41760
rect 468331 41713 468387 41806
rect 470048 41812 470227 41818
rect 470100 41806 470227 41812
rect 470048 41754 470100 41760
rect 470171 41713 470227 41806
rect 471367 41713 471423 42193
rect 472636 41806 472711 42193
rect 474476 41806 474551 42193
rect 472655 41713 472711 41806
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 518807 41713 518863 42193
rect 520647 41713 520703 42193
rect 521843 41713 521899 42193
rect 523131 41713 523187 42193
rect 524971 41713 525027 42193
rect 526167 41713 526223 42193
rect 527455 41713 527511 42193
rect 529295 41713 529351 42193
<< via2 >>
rect 411074 44376 411130 44432
rect 419722 44240 419778 44296
rect 465814 44376 465870 44432
rect 474462 44376 474518 44432
rect 518806 44240 518862 44296
rect 524970 44240 525026 44296
<< obsm2 >>
rect 75850 1006851 89088 1007371
rect 123850 1006851 137088 1007371
rect 171850 1006851 185088 1007371
rect 229453 1002788 244258 1036615
rect 280853 1002788 295658 1036615
rect 229453 998067 239422 1002788
rect 234335 998007 239422 998067
rect 234579 997600 234979 997984
rect 280853 998067 290822 1002788
rect 285735 998007 290822 998067
rect 285979 997600 286379 997984
rect 339453 998007 354258 1036615
rect 425650 1006851 438888 1007371
rect 475050 1006851 488288 1007371
rect 526650 1006851 539888 1007371
rect 575653 998007 590458 1036615
rect 627850 1006851 641088 1007371
rect 339499 997600 344279 998007
rect 344579 997600 344979 997984
rect 349478 997600 354258 998007
rect 575699 997600 580479 998007
rect 580779 997600 581179 997984
rect 585678 997600 590458 998007
rect 585782 997455 585838 997529
rect 339498 997047 339554 997121
rect 339512 996402 339540 997047
rect 585796 996470 585824 997455
rect 585784 996406 585836 996470
rect 674748 996406 674800 996470
rect 42248 996338 42300 996402
rect 339500 996338 339552 996402
rect 673552 996338 673604 996402
rect 30229 956050 30749 969288
rect 7 928240 30281 930187
rect 30753 928000 31683 930228
rect 32033 928240 34915 930187
rect 7 927940 39593 928000
rect 7 923819 39600 927940
rect 7 923707 39593 923819
rect 7 917185 39600 923707
rect 7 917099 39593 917185
rect 7 913100 39600 917099
rect 7 913000 39593 913100
rect 30760 910805 31690 913000
rect 985 880878 40000 885658
rect 985 875679 39593 880878
rect 39616 875979 40000 876379
rect 985 870899 40000 875679
rect 985 870853 39593 870899
rect 985 838478 40000 843258
rect 985 833279 39593 838478
rect 39616 833579 40000 833979
rect 985 828499 40000 833279
rect 985 828453 39593 828499
rect 0 800973 41713 801183
rect 42260 801038 42288 996338
rect 44916 990082 44968 990146
rect 42340 990014 42392 990078
rect 42248 800974 42300 801038
rect 0 800805 41657 800973
rect 41713 800903 42193 800917
rect 41713 800875 42288 800903
rect 41713 800861 42193 800875
rect 0 800329 41713 800805
rect 0 800161 41657 800329
rect 0 799685 41713 800161
rect 0 799517 41657 799685
rect 41713 799573 42193 799629
rect 0 799133 41713 799517
rect 0 798965 41657 799133
rect 41722 799077 41828 799082
rect 41713 799021 42193 799077
rect 0 798489 41713 798965
rect 41800 798590 41828 799021
rect 41788 798526 41840 798590
rect 0 798321 41657 798489
rect 0 797845 41713 798321
rect 0 797677 41657 797845
rect 0 797293 41713 797677
rect 0 797125 41657 797293
rect 41713 797181 42193 797237
rect 0 796649 41713 797125
rect 0 796481 41657 796649
rect 0 796005 41713 796481
rect 0 795837 41657 796005
rect 0 795453 41713 795837
rect 0 795285 41657 795453
rect 0 794809 41713 795285
rect 0 794641 41657 794809
rect 0 794165 41713 794641
rect 0 793997 41657 794165
rect 0 793613 41713 793997
rect 0 793445 41657 793613
rect 0 792969 41713 793445
rect 42260 793098 42288 800875
rect 42352 798590 42380 990014
rect 44928 902534 44956 990082
rect 673460 990014 673512 990078
rect 44836 902506 44956 902534
rect 44836 885873 44864 902506
rect 44178 885799 44234 885873
rect 44822 885799 44878 885873
rect 44192 871049 44220 885799
rect 44178 870975 44234 871049
rect 44192 861218 44220 870975
rect 42432 861154 42484 861218
rect 44180 861154 44232 861218
rect 42340 798526 42392 798590
rect 41800 793070 42288 793098
rect 0 792801 41657 792969
rect 41800 792913 41828 793070
rect 41713 792857 42193 792913
rect 0 792325 41713 792801
rect 0 792157 41657 792325
rect 0 791681 41713 792157
rect 41788 792066 41840 792130
rect 0 791513 41657 791681
rect 41800 791625 41828 792066
rect 41713 791569 42193 791625
rect 0 791129 41713 791513
rect 0 790961 41657 791129
rect 0 790485 41713 790961
rect 0 790317 41657 790485
rect 0 789841 41713 790317
rect 0 789673 41657 789841
rect 0 789289 41713 789673
rect 0 789121 41657 789289
rect 0 788645 41713 789121
rect 41788 789074 41840 789138
rect 0 788477 41657 788645
rect 41800 788589 41828 789074
rect 41713 788533 42193 788589
rect 0 788001 41713 788477
rect 0 787833 41657 788001
rect 0 787449 41713 787833
rect 0 787281 41657 787449
rect 0 786805 41713 787281
rect 0 786637 41657 786805
rect 0 786161 41713 786637
rect 0 785993 41657 786161
rect 0 785609 41713 785993
rect 0 785441 41657 785609
rect 0 785242 41713 785441
rect 0 757773 41713 757983
rect 0 757605 41657 757773
rect 41713 757703 42193 757717
rect 41713 757675 42288 757703
rect 41713 757661 42193 757675
rect 0 757129 41713 757605
rect 0 756961 41657 757129
rect 0 756485 41713 756961
rect 0 756317 41657 756485
rect 41713 756373 42193 756429
rect 0 755933 41713 756317
rect 41788 756230 41840 756294
rect 0 755765 41657 755933
rect 41800 755877 41828 756230
rect 41713 755821 42193 755877
rect 0 755289 41713 755765
rect 0 755121 41657 755289
rect 0 754645 41713 755121
rect 0 754477 41657 754645
rect 0 754093 41713 754477
rect 0 753925 41657 754093
rect 41713 753981 42193 754037
rect 0 753449 41713 753925
rect 0 753281 41657 753449
rect 0 752805 41713 753281
rect 0 752637 41657 752805
rect 0 752253 41713 752637
rect 0 752085 41657 752253
rect 0 751609 41713 752085
rect 0 751441 41657 751609
rect 0 750965 41713 751441
rect 0 750797 41657 750965
rect 0 750413 41713 750797
rect 0 750245 41657 750413
rect 0 749769 41713 750245
rect 42260 749850 42288 757675
rect 42352 756294 42380 798526
rect 42444 792130 42472 861154
rect 673472 849726 673500 990014
rect 673564 859178 673592 996338
rect 673644 990082 673696 990146
rect 673552 859114 673604 859178
rect 673460 849662 673512 849726
rect 42616 800974 42668 801038
rect 42432 792066 42484 792130
rect 42444 792010 42472 792066
rect 42444 791982 42564 792010
rect 42340 756230 42392 756294
rect 41800 749822 42288 749850
rect 0 749601 41657 749769
rect 41800 749714 41828 749822
rect 41722 749713 41828 749714
rect 41713 749657 42193 749713
rect 0 749125 41713 749601
rect 0 748957 41657 749125
rect 0 748481 41713 748957
rect 0 748313 41657 748481
rect 41713 748369 42193 748425
rect 41800 748338 41828 748369
rect 0 747929 41713 748313
rect 41788 748274 41840 748338
rect 0 747761 41657 747929
rect 0 747285 41713 747761
rect 0 747117 41657 747285
rect 0 746641 41713 747117
rect 0 746473 41657 746641
rect 0 746089 41713 746473
rect 0 745921 41657 746089
rect 0 745445 41713 745921
rect 0 745277 41657 745445
rect 41713 745333 42193 745389
rect 0 744801 41713 745277
rect 41800 744870 41828 745333
rect 41788 744806 41840 744870
rect 0 744633 41657 744801
rect 42536 748338 42564 791982
rect 42628 789138 42656 800974
rect 42616 789074 42668 789138
rect 42628 786614 42656 789074
rect 42628 786586 42748 786614
rect 42616 756230 42668 756294
rect 42524 748274 42576 748338
rect 42432 744806 42484 744870
rect 0 744249 41713 744633
rect 0 744081 41657 744249
rect 0 743605 41713 744081
rect 0 743437 41657 743605
rect 0 742961 41713 743437
rect 0 742793 41657 742961
rect 0 742409 41713 742793
rect 0 742241 41657 742409
rect 0 742042 41713 742241
rect 0 714573 41713 714783
rect 0 714405 41657 714573
rect 41713 714461 42193 714517
rect 0 713929 41713 714405
rect 41892 714218 41920 714461
rect 41892 714190 42288 714218
rect 0 713761 41657 713929
rect 0 713285 41713 713761
rect 0 713117 41657 713285
rect 41713 713173 42193 713229
rect 0 712733 41713 713117
rect 41788 713050 41840 713114
rect 0 712565 41657 712733
rect 41800 712677 41828 713050
rect 41713 712621 42193 712677
rect 0 712089 41713 712565
rect 0 711921 41657 712089
rect 0 711445 41713 711921
rect 0 711277 41657 711445
rect 0 710893 41713 711277
rect 0 710725 41657 710893
rect 41713 710781 42193 710837
rect 0 710249 41713 710725
rect 0 710081 41657 710249
rect 0 709605 41713 710081
rect 0 709437 41657 709605
rect 0 709053 41713 709437
rect 0 708885 41657 709053
rect 0 708409 41713 708885
rect 0 708241 41657 708409
rect 0 707765 41713 708241
rect 0 707597 41657 707765
rect 0 707213 41713 707597
rect 0 707045 41657 707213
rect 0 706569 41713 707045
rect 0 706401 41657 706569
rect 41713 706499 42193 706513
rect 42260 706499 42288 714190
rect 41713 706471 42288 706499
rect 41713 706457 42193 706471
rect 0 705925 41713 706401
rect 0 705757 41657 705925
rect 0 705281 41713 705757
rect 0 705113 41657 705281
rect 41713 705169 42193 705225
rect 0 704729 41713 705113
rect 41800 704818 41828 705169
rect 41788 704754 41840 704818
rect 0 704561 41657 704729
rect 0 704085 41713 704561
rect 0 703917 41657 704085
rect 0 703441 41713 703917
rect 0 703273 41657 703441
rect 0 702889 41713 703273
rect 0 702721 41657 702889
rect 0 702245 41713 702721
rect 0 702077 41657 702245
rect 41713 702133 42193 702189
rect 0 701601 41713 702077
rect 41800 701690 41828 702133
rect 41788 701626 41840 701690
rect 0 701433 41657 701601
rect 42444 701690 42472 744806
rect 42536 704818 42564 748274
rect 42628 713114 42656 756230
rect 42720 744870 42748 786586
rect 673472 761326 673500 849662
rect 673564 772818 673592 859114
rect 673656 856118 673684 990082
rect 673644 856054 673696 856118
rect 673552 772754 673604 772818
rect 673460 761262 673512 761326
rect 42708 744806 42760 744870
rect 673564 728414 673592 772754
rect 673656 769690 673684 856054
rect 673644 769626 673696 769690
rect 673920 769626 673972 769690
rect 673552 728350 673604 728414
rect 42616 713050 42668 713114
rect 42524 704754 42576 704818
rect 42432 701626 42484 701690
rect 0 701049 41713 701433
rect 0 700881 41657 701049
rect 0 700405 41713 700881
rect 0 700237 41657 700405
rect 0 699761 41713 700237
rect 0 699593 41657 699761
rect 0 699209 41713 699593
rect 0 699041 41657 699209
rect 0 698842 41713 699041
rect 0 671173 41713 671383
rect 0 671005 41657 671173
rect 41713 671061 42193 671117
rect 0 670529 41713 671005
rect 41800 670694 41828 671061
rect 41800 670666 42288 670694
rect 0 670361 41657 670529
rect 0 669885 41713 670361
rect 0 669717 41657 669885
rect 41713 669773 42193 669829
rect 0 669333 41713 669717
rect 0 669165 41657 669333
rect 41713 669221 42193 669277
rect 0 668689 41713 669165
rect 41800 668778 41828 669221
rect 41788 668714 41840 668778
rect 0 668521 41657 668689
rect 0 668045 41713 668521
rect 0 667877 41657 668045
rect 0 667493 41713 667877
rect 0 667325 41657 667493
rect 41713 667381 42193 667437
rect 0 666849 41713 667325
rect 0 666681 41657 666849
rect 0 666205 41713 666681
rect 0 666037 41657 666205
rect 0 665653 41713 666037
rect 0 665485 41657 665653
rect 0 665009 41713 665485
rect 0 664841 41657 665009
rect 0 664365 41713 664841
rect 0 664197 41657 664365
rect 0 663813 41713 664197
rect 0 663645 41657 663813
rect 0 663169 41713 663645
rect 42260 663626 42288 670666
rect 41892 663598 42288 663626
rect 0 663001 41657 663169
rect 41892 663113 41920 663598
rect 41713 663057 42193 663113
rect 41722 663054 41920 663057
rect 0 662525 41713 663001
rect 0 662357 41657 662525
rect 0 661881 41713 662357
rect 0 661713 41657 661881
rect 41713 661769 42193 661825
rect 0 661329 41713 661713
rect 41800 661366 41828 661769
rect 0 661161 41657 661329
rect 41788 661302 41840 661366
rect 0 660685 41713 661161
rect 0 660517 41657 660685
rect 0 660041 41713 660517
rect 0 659873 41657 660041
rect 0 659489 41713 659873
rect 0 659321 41657 659489
rect 0 658845 41713 659321
rect 41788 659262 41840 659326
rect 0 658677 41657 658845
rect 41800 658789 41828 659262
rect 41713 658733 42193 658789
rect 0 658201 41713 658677
rect 0 658033 41657 658201
rect 42444 659326 42472 701626
rect 42536 661366 42564 704754
rect 42628 668778 42656 713050
rect 673564 683126 673592 728350
rect 673932 725286 673960 769626
rect 674012 761262 674064 761326
rect 673920 725222 673972 725286
rect 673644 717810 673696 717874
rect 673552 683062 673604 683126
rect 673552 680410 673604 680474
rect 42616 668714 42668 668778
rect 42524 661302 42576 661366
rect 42432 659262 42484 659326
rect 0 657649 41713 658033
rect 0 657481 41657 657649
rect 0 657005 41713 657481
rect 0 656837 41657 657005
rect 0 656361 41713 656837
rect 0 656193 41657 656361
rect 0 655809 41713 656193
rect 0 655641 41657 655809
rect 0 655442 41713 655641
rect 0 627973 41713 628183
rect 0 627805 41657 627973
rect 41713 627903 42193 627917
rect 41713 627875 42288 627903
rect 41713 627861 42193 627875
rect 0 627329 41713 627805
rect 0 627161 41657 627329
rect 0 626685 41713 627161
rect 0 626517 41657 626685
rect 41713 626573 42193 626629
rect 0 626133 41713 626517
rect 0 625965 41657 626133
rect 41722 626077 41828 626090
rect 41713 626021 42193 626077
rect 0 625489 41713 625965
rect 41800 625530 41828 626021
rect 0 625321 41657 625489
rect 41788 625466 41840 625530
rect 0 624845 41713 625321
rect 0 624677 41657 624845
rect 0 624293 41713 624677
rect 0 624125 41657 624293
rect 41713 624181 42193 624237
rect 0 623649 41713 624125
rect 0 623481 41657 623649
rect 0 623005 41713 623481
rect 0 622837 41657 623005
rect 0 622453 41713 622837
rect 0 622285 41657 622453
rect 0 621809 41713 622285
rect 0 621641 41657 621809
rect 0 621165 41713 621641
rect 0 620997 41657 621165
rect 0 620613 41713 620997
rect 0 620445 41657 620613
rect 0 619969 41713 620445
rect 42260 620378 42288 627875
rect 41892 620350 42288 620378
rect 0 619801 41657 619969
rect 41892 619913 41920 620350
rect 41713 619857 42193 619913
rect 0 619325 41713 619801
rect 0 619157 41657 619325
rect 0 618681 41713 619157
rect 0 618513 41657 618681
rect 41713 618569 42193 618625
rect 0 618129 41713 618513
rect 41800 618186 41828 618569
rect 0 617961 41657 618129
rect 41788 618122 41840 618186
rect 0 617485 41713 617961
rect 0 617317 41657 617485
rect 0 616841 41713 617317
rect 0 616673 41657 616841
rect 0 616289 41713 616673
rect 0 616121 41657 616289
rect 0 615645 41713 616121
rect 0 615477 41657 615645
rect 41713 615533 42193 615589
rect 0 615001 41713 615477
rect 41800 615058 41828 615533
rect 0 614833 41657 615001
rect 41788 614994 41840 615058
rect 0 614449 41713 614833
rect 42536 618186 42564 661302
rect 42628 625530 42656 668714
rect 42708 659262 42760 659326
rect 42616 625466 42668 625530
rect 42524 618122 42576 618186
rect 42248 614654 42300 614718
rect 0 614281 41657 614449
rect 0 613805 41713 614281
rect 0 613637 41657 613805
rect 0 613161 41713 613637
rect 0 612993 41657 613161
rect 0 612609 41713 612993
rect 0 612441 41657 612609
rect 0 612242 41713 612441
rect 0 584773 41713 584983
rect 42260 584882 42288 614654
rect 42260 584854 42380 584882
rect 0 584605 41657 584773
rect 41713 584703 42193 584717
rect 41713 584675 42288 584703
rect 41713 584661 42193 584675
rect 0 584129 41713 584605
rect 0 583961 41657 584129
rect 0 583485 41713 583961
rect 0 583317 41657 583485
rect 41713 583373 42193 583429
rect 0 582933 41713 583317
rect 41788 583238 41840 583302
rect 0 582765 41657 582933
rect 41800 582877 41828 583238
rect 41713 582821 42193 582877
rect 41722 582814 41828 582821
rect 0 582289 41713 582765
rect 0 582121 41657 582289
rect 0 581645 41713 582121
rect 0 581477 41657 581645
rect 0 581093 41713 581477
rect 0 580925 41657 581093
rect 41713 580981 42193 581037
rect 0 580449 41713 580925
rect 0 580281 41657 580449
rect 0 579805 41713 580281
rect 0 579637 41657 579805
rect 0 579253 41713 579637
rect 0 579085 41657 579253
rect 0 578609 41713 579085
rect 0 578441 41657 578609
rect 0 577965 41713 578441
rect 0 577797 41657 577965
rect 0 577413 41713 577797
rect 0 577245 41657 577413
rect 0 576769 41713 577245
rect 42260 576858 42288 584675
rect 41892 576830 42288 576858
rect 0 576601 41657 576769
rect 41892 576722 41920 576830
rect 41722 576713 41920 576722
rect 41713 576657 42193 576713
rect 0 576125 41713 576601
rect 0 575957 41657 576125
rect 0 575481 41713 575957
rect 41788 575894 41840 575958
rect 0 575313 41657 575481
rect 41800 575425 41828 575894
rect 41713 575369 42193 575425
rect 0 574929 41713 575313
rect 0 574761 41657 574929
rect 0 574285 41713 574761
rect 0 574117 41657 574285
rect 0 573641 41713 574117
rect 0 573473 41657 573641
rect 0 573089 41713 573473
rect 0 572921 41657 573089
rect 0 572445 41713 572921
rect 0 572277 41657 572445
rect 41713 572333 42193 572389
rect 0 571801 41713 572277
rect 41800 571878 41828 572333
rect 41788 571814 41840 571878
rect 0 571633 41657 571801
rect 42352 574094 42380 584854
rect 42536 575958 42564 618122
rect 42628 583302 42656 625466
rect 42720 615058 42748 659262
rect 673564 636342 673592 680410
rect 673656 673674 673684 717810
rect 673736 683062 673788 683126
rect 673644 673610 673696 673674
rect 673748 643094 673776 683062
rect 673932 680474 673960 725222
rect 674024 717874 674052 761262
rect 674012 717810 674064 717874
rect 673920 680410 673972 680474
rect 673656 643066 673776 643094
rect 673656 638926 673684 643066
rect 674012 673610 674064 673674
rect 673644 638862 673696 638926
rect 673552 636278 673604 636342
rect 673460 629410 673512 629474
rect 42708 614994 42760 615058
rect 673472 584186 673500 629410
rect 673564 591938 673592 636278
rect 673656 595202 673684 638862
rect 674024 629474 674052 673610
rect 674012 629410 674064 629474
rect 673644 595138 673696 595202
rect 673552 591874 673604 591938
rect 673460 584122 673512 584186
rect 42616 583238 42668 583302
rect 42524 575894 42576 575958
rect 42352 574066 42472 574094
rect 42444 571878 42472 574066
rect 42432 571814 42484 571878
rect 0 571249 41713 571633
rect 0 571081 41657 571249
rect 0 570605 41713 571081
rect 0 570437 41657 570605
rect 0 569961 41713 570437
rect 0 569793 41657 569961
rect 0 569409 41713 569793
rect 0 569241 41657 569409
rect 0 569042 41713 569241
rect 0 541573 41713 541783
rect 0 541405 41657 541573
rect 41713 541461 42193 541517
rect 0 540929 41713 541405
rect 41800 541362 41828 541461
rect 41800 541334 42288 541362
rect 0 540761 41657 540929
rect 0 540285 41713 540761
rect 0 540117 41657 540285
rect 41713 540173 42193 540229
rect 0 539733 41713 540117
rect 41788 540058 41840 540122
rect 0 539565 41657 539733
rect 41800 539677 41828 540058
rect 41713 539621 42193 539677
rect 0 539089 41713 539565
rect 0 538921 41657 539089
rect 0 538445 41713 538921
rect 0 538277 41657 538445
rect 0 537893 41713 538277
rect 0 537725 41657 537893
rect 41713 537781 42193 537837
rect 0 537249 41713 537725
rect 0 537081 41657 537249
rect 0 536605 41713 537081
rect 0 536437 41657 536605
rect 0 536053 41713 536437
rect 0 535885 41657 536053
rect 0 535409 41713 535885
rect 0 535241 41657 535409
rect 0 534765 41713 535241
rect 0 534597 41657 534765
rect 0 534213 41713 534597
rect 0 534045 41657 534213
rect 0 533569 41713 534045
rect 42260 533610 42288 541334
rect 41892 533582 42288 533610
rect 0 533401 41657 533569
rect 41892 533513 41920 533582
rect 41713 533457 42193 533513
rect 41722 533446 41920 533457
rect 0 532925 41713 533401
rect 0 532757 41657 532925
rect 0 532281 41713 532757
rect 0 532113 41657 532281
rect 41713 532169 42193 532225
rect 0 531729 41713 532113
rect 41800 531826 41828 532169
rect 41788 531762 41840 531826
rect 0 531561 41657 531729
rect 0 531085 41713 531561
rect 0 530917 41657 531085
rect 0 530441 41713 530917
rect 0 530273 41657 530441
rect 0 529889 41713 530273
rect 0 529721 41657 529889
rect 0 529245 41713 529721
rect 0 529077 41657 529245
rect 41713 529133 42193 529189
rect 0 528601 41713 529077
rect 41800 528698 41828 529133
rect 41788 528634 41840 528698
rect 0 528433 41657 528601
rect 42444 528698 42472 571814
rect 42536 531826 42564 575894
rect 42628 540122 42656 583238
rect 673564 548282 673592 591874
rect 673656 551410 673684 595138
rect 673920 584122 673972 584186
rect 673644 551346 673696 551410
rect 673552 548218 673604 548282
rect 42616 540058 42668 540122
rect 42524 531762 42576 531826
rect 42432 528634 42484 528698
rect 0 528049 41713 528433
rect 0 527881 41657 528049
rect 0 527405 41713 527881
rect 0 527237 41657 527405
rect 0 526761 41713 527237
rect 0 526593 41657 526761
rect 0 526209 41713 526593
rect 0 526041 41657 526209
rect 0 525842 41713 526041
rect 985 493478 40000 498258
rect 985 488279 39593 493478
rect 39616 488579 40000 488979
rect 985 483499 40000 488279
rect 985 483453 39593 483499
rect 7 456440 30281 458387
rect 30753 456200 31683 458428
rect 32033 456440 34915 458387
rect 7 456140 39593 456200
rect 7 452019 39600 456140
rect 7 451907 39593 452019
rect 7 445385 39600 451907
rect 7 445299 39593 445385
rect 7 441300 39600 445299
rect 7 441200 39593 441300
rect 30760 439005 31690 441200
rect 0 413773 41713 413983
rect 0 413605 41657 413773
rect 41713 413703 42193 413717
rect 41713 413675 42288 413703
rect 41713 413661 42193 413675
rect 0 413129 41713 413605
rect 0 412961 41657 413129
rect 0 412485 41713 412961
rect 0 412317 41657 412485
rect 41713 412373 42193 412429
rect 0 411933 41713 412317
rect 0 411765 41657 411933
rect 41722 411877 41828 411890
rect 41713 411821 42193 411877
rect 0 411289 41713 411765
rect 41800 411330 41828 411821
rect 0 411121 41657 411289
rect 41788 411266 41840 411330
rect 0 410645 41713 411121
rect 0 410477 41657 410645
rect 0 410093 41713 410477
rect 0 409925 41657 410093
rect 41713 409981 42193 410037
rect 0 409449 41713 409925
rect 0 409281 41657 409449
rect 0 408805 41713 409281
rect 0 408637 41657 408805
rect 0 408253 41713 408637
rect 0 408085 41657 408253
rect 0 407609 41713 408085
rect 0 407441 41657 407609
rect 0 406965 41713 407441
rect 0 406797 41657 406965
rect 0 406413 41713 406797
rect 0 406245 41657 406413
rect 0 405769 41713 406245
rect 42260 405770 42288 413675
rect 0 405601 41657 405769
rect 41892 405742 42288 405770
rect 41892 405713 41920 405742
rect 41713 405657 42193 405713
rect 0 405125 41713 405601
rect 0 404957 41657 405125
rect 0 404481 41713 404957
rect 41788 404874 41840 404938
rect 0 404313 41657 404481
rect 41800 404425 41828 404874
rect 41713 404369 42193 404425
rect 0 403929 41713 404313
rect 0 403761 41657 403929
rect 0 403285 41713 403761
rect 0 403117 41657 403285
rect 0 402641 41713 403117
rect 0 402473 41657 402641
rect 0 402089 41713 402473
rect 0 401921 41657 402089
rect 0 401445 41713 401921
rect 41788 401882 41840 401946
rect 0 401277 41657 401445
rect 41800 401389 41828 401882
rect 41713 401333 42193 401389
rect 0 400801 41713 401277
rect 0 400633 41657 400801
rect 42444 401946 42472 528634
rect 42628 419534 42656 540058
rect 42708 531762 42760 531826
rect 42536 419506 42656 419534
rect 42536 411330 42564 419506
rect 42524 411266 42576 411330
rect 42432 401882 42484 401946
rect 0 400249 41713 400633
rect 0 400081 41657 400249
rect 0 399605 41713 400081
rect 0 399437 41657 399605
rect 0 398961 41713 399437
rect 0 398793 41657 398961
rect 0 398409 41713 398793
rect 0 398241 41657 398409
rect 0 398042 41713 398241
rect 0 370573 41713 370783
rect 0 370405 41657 370573
rect 41713 370503 42193 370517
rect 41713 370475 42288 370503
rect 41713 370461 42193 370475
rect 0 369929 41713 370405
rect 0 369761 41657 369929
rect 0 369285 41713 369761
rect 0 369117 41657 369285
rect 41713 369173 42193 369229
rect 0 368733 41713 369117
rect 41788 369038 41840 369102
rect 0 368565 41657 368733
rect 41800 368677 41828 369038
rect 41713 368621 42193 368677
rect 41722 368614 41828 368621
rect 0 368089 41713 368565
rect 0 367921 41657 368089
rect 0 367445 41713 367921
rect 0 367277 41657 367445
rect 0 366893 41713 367277
rect 0 366725 41657 366893
rect 41713 366781 42193 366837
rect 0 366249 41713 366725
rect 0 366081 41657 366249
rect 0 365605 41713 366081
rect 0 365437 41657 365605
rect 0 365053 41713 365437
rect 0 364885 41657 365053
rect 0 364409 41713 364885
rect 0 364241 41657 364409
rect 0 363765 41713 364241
rect 0 363597 41657 363765
rect 0 363213 41713 363597
rect 0 363045 41657 363213
rect 0 362569 41713 363045
rect 42260 362658 42288 370475
rect 41800 362630 42288 362658
rect 0 362401 41657 362569
rect 41800 362522 41828 362630
rect 41722 362513 41828 362522
rect 41713 362457 42193 362513
rect 0 361925 41713 362401
rect 0 361757 41657 361925
rect 0 361281 41713 361757
rect 41788 361286 41840 361350
rect 0 361113 41657 361281
rect 41800 361225 41828 361286
rect 41713 361169 42193 361225
rect 0 360729 41713 361113
rect 0 360561 41657 360729
rect 0 360085 41713 360561
rect 0 359917 41657 360085
rect 0 359441 41713 359917
rect 0 359273 41657 359441
rect 0 358889 41713 359273
rect 0 358721 41657 358889
rect 0 358245 41713 358721
rect 0 358077 41657 358245
rect 41713 358133 42193 358189
rect 0 357601 41713 358077
rect 41800 357678 41828 358133
rect 41788 357614 41840 357678
rect 0 357433 41657 357601
rect 42444 357678 42472 401882
rect 42536 369102 42564 411266
rect 42720 404938 42748 531762
rect 42708 404874 42760 404938
rect 42720 400214 42748 404874
rect 42628 400186 42748 400214
rect 42524 369038 42576 369102
rect 42432 357614 42484 357678
rect 0 357049 41713 357433
rect 0 356881 41657 357049
rect 0 356405 41713 356881
rect 0 356237 41657 356405
rect 0 355761 41713 356237
rect 0 355593 41657 355761
rect 0 355209 41713 355593
rect 0 355041 41657 355209
rect 0 354842 41713 355041
rect 0 327173 41713 327383
rect 0 327005 41657 327173
rect 41713 327103 42193 327117
rect 41713 327075 42288 327103
rect 41713 327061 42193 327075
rect 0 326529 41713 327005
rect 0 326361 41657 326529
rect 0 325885 41713 326361
rect 0 325717 41657 325885
rect 41713 325773 42193 325829
rect 0 325333 41713 325717
rect 41788 325654 41840 325718
rect 0 325165 41657 325333
rect 41800 325277 41828 325654
rect 41713 325221 42193 325277
rect 0 324689 41713 325165
rect 0 324521 41657 324689
rect 0 324045 41713 324521
rect 0 323877 41657 324045
rect 0 323493 41713 323877
rect 0 323325 41657 323493
rect 41713 323381 42193 323437
rect 0 322849 41713 323325
rect 0 322681 41657 322849
rect 0 322205 41713 322681
rect 0 322037 41657 322205
rect 0 321653 41713 322037
rect 0 321485 41657 321653
rect 0 321009 41713 321485
rect 0 320841 41657 321009
rect 0 320365 41713 320841
rect 0 320197 41657 320365
rect 0 319813 41713 320197
rect 0 319645 41657 319813
rect 0 319169 41713 319645
rect 0 319001 41657 319169
rect 41713 319099 42193 319113
rect 42260 319099 42288 327075
rect 41713 319071 42288 319099
rect 41713 319057 42193 319071
rect 0 318525 41713 319001
rect 0 318357 41657 318525
rect 0 317881 41713 318357
rect 42536 325718 42564 369038
rect 42628 361350 42656 400186
rect 673932 540938 673960 584122
rect 673920 540874 673972 540938
rect 674760 422278 674788 996406
rect 678067 954065 716615 958947
rect 677600 953421 677984 953821
rect 678007 948978 716615 954065
rect 682788 944142 716615 948978
rect 685910 906400 686840 908595
rect 678007 906300 717593 906400
rect 678000 902301 717593 906300
rect 678007 902215 717593 902301
rect 678000 895693 717593 902215
rect 678007 895581 717593 895693
rect 678000 891460 717593 895581
rect 678007 891400 717593 891460
rect 682685 889213 685567 891160
rect 685917 889172 686847 891400
rect 687319 889213 717593 891160
rect 675887 862759 717600 862958
rect 675943 862591 717600 862759
rect 675887 862207 717600 862591
rect 675943 862039 717600 862207
rect 675887 861563 717600 862039
rect 675943 861395 717600 861563
rect 675887 860919 717600 861395
rect 675943 860751 717600 860919
rect 675887 860367 717600 860751
rect 675943 860199 717600 860367
rect 675887 859723 717600 860199
rect 675407 859639 675887 859667
rect 675404 859611 675887 859639
rect 675404 859178 675432 859611
rect 675943 859555 717600 859723
rect 675392 859114 675444 859178
rect 675887 859079 717600 859555
rect 675943 858911 717600 859079
rect 675887 858527 717600 858911
rect 675943 858359 717600 858527
rect 675887 857883 717600 858359
rect 675943 857715 717600 857883
rect 675887 857239 717600 857715
rect 675943 857071 717600 857239
rect 675887 856687 717600 857071
rect 675407 856596 675887 856631
rect 675404 856575 675887 856596
rect 675404 856118 675432 856575
rect 675943 856519 717600 856687
rect 675392 856054 675444 856118
rect 675887 856043 717600 856519
rect 675943 855875 717600 856043
rect 675887 855399 717600 855875
rect 675407 855329 675887 855343
rect 675312 855301 675887 855329
rect 675312 847325 675340 855301
rect 675407 855287 675887 855301
rect 675943 855231 717600 855399
rect 675887 854755 717600 855231
rect 675943 854587 717600 854755
rect 675887 854203 717600 854587
rect 675943 854035 717600 854203
rect 675887 853559 717600 854035
rect 675943 853391 717600 853559
rect 675887 852915 717600 853391
rect 675943 852747 717600 852915
rect 675887 852363 717600 852747
rect 675943 852195 717600 852363
rect 675887 851719 717600 852195
rect 675943 851551 717600 851719
rect 675887 851075 717600 851551
rect 675407 850963 675887 851019
rect 675943 850907 717600 851075
rect 675887 850523 717600 850907
rect 675943 850355 717600 850523
rect 675887 849879 717600 850355
rect 675392 849662 675444 849726
rect 675943 849711 717600 849879
rect 675404 849179 675432 849662
rect 675887 849235 717600 849711
rect 675404 849151 675887 849179
rect 675407 849123 675887 849151
rect 675943 849067 717600 849235
rect 675887 848683 717600 849067
rect 675407 848571 675887 848627
rect 675943 848515 717600 848683
rect 675887 848039 717600 848515
rect 675943 847871 717600 848039
rect 675887 847395 717600 847871
rect 675407 847325 675887 847339
rect 675312 847297 675887 847325
rect 675407 847283 675887 847297
rect 675943 847227 717600 847395
rect 675887 847017 717600 847227
rect 678007 818701 716615 818747
rect 677600 813921 716615 818701
rect 677600 813221 677984 813621
rect 678007 808722 716615 813921
rect 677600 803942 716615 808722
rect 675300 803762 675352 803826
rect 677598 803791 677654 803865
rect 677600 803762 677652 803791
rect 675208 767586 675260 767650
rect 675220 760238 675248 767586
rect 675208 760174 675260 760238
rect 675312 739694 675340 803762
rect 675887 775359 717600 775558
rect 675943 775191 717600 775359
rect 675887 774807 717600 775191
rect 675943 774639 717600 774807
rect 675887 774163 717600 774639
rect 675943 773995 717600 774163
rect 675887 773519 717600 773995
rect 675943 773351 717600 773519
rect 675887 772967 717600 773351
rect 675392 772754 675444 772818
rect 675943 772799 717600 772967
rect 675404 772267 675432 772754
rect 675887 772323 717600 772799
rect 675404 772239 675887 772267
rect 675407 772211 675887 772239
rect 675943 772155 717600 772323
rect 675887 771679 717600 772155
rect 675943 771511 717600 771679
rect 675887 771127 717600 771511
rect 675943 770959 717600 771127
rect 675887 770483 717600 770959
rect 675943 770315 717600 770483
rect 675887 769839 717600 770315
rect 675392 769626 675444 769690
rect 675943 769671 717600 769839
rect 675404 769231 675432 769626
rect 675887 769287 717600 769671
rect 675404 769203 675887 769231
rect 675407 769175 675887 769203
rect 675943 769119 717600 769287
rect 675887 768643 717600 769119
rect 675943 768475 717600 768643
rect 675887 767999 717600 768475
rect 675407 767924 675887 767943
rect 675404 767887 675887 767924
rect 675404 767650 675432 767887
rect 675943 767831 717600 767999
rect 675392 767586 675444 767650
rect 675887 767355 717600 767831
rect 675943 767187 717600 767355
rect 675887 766803 717600 767187
rect 675943 766635 717600 766803
rect 675887 766159 717600 766635
rect 675943 765991 717600 766159
rect 675887 765515 717600 765991
rect 675943 765347 717600 765515
rect 675887 764963 717600 765347
rect 675943 764795 717600 764963
rect 675887 764319 717600 764795
rect 675943 764151 717600 764319
rect 675887 763675 717600 764151
rect 675407 763563 675887 763619
rect 675943 763507 717600 763675
rect 675887 763123 717600 763507
rect 675943 762955 717600 763123
rect 675887 762479 717600 762955
rect 675943 762311 717600 762479
rect 675887 761835 717600 762311
rect 675407 761751 675887 761779
rect 675404 761723 675887 761751
rect 675404 761326 675432 761723
rect 675943 761667 717600 761835
rect 675392 761262 675444 761326
rect 675887 761283 717600 761667
rect 675407 761171 675887 761227
rect 675943 761115 717600 761283
rect 675887 760639 717600 761115
rect 675943 760471 717600 760639
rect 675392 760174 675444 760238
rect 675404 759939 675432 760174
rect 675887 759995 717600 760471
rect 675404 759900 675887 759939
rect 675407 759883 675887 759900
rect 675943 759827 717600 759995
rect 675887 759617 717600 759827
rect 675128 739666 675340 739694
rect 675128 709334 675156 739666
rect 675887 730959 717600 731158
rect 675943 730791 717600 730959
rect 675887 730407 717600 730791
rect 675943 730239 717600 730407
rect 675887 729763 717600 730239
rect 675943 729595 717600 729763
rect 675887 729119 717600 729595
rect 675943 728951 717600 729119
rect 675887 728567 717600 728951
rect 675392 728350 675444 728414
rect 675943 728399 717600 728567
rect 675404 727867 675432 728350
rect 675887 727923 717600 728399
rect 675404 727839 675887 727867
rect 675407 727811 675887 727839
rect 675943 727755 717600 727923
rect 675887 727279 717600 727755
rect 675943 727111 717600 727279
rect 675887 726727 717600 727111
rect 675943 726559 717600 726727
rect 675887 726083 717600 726559
rect 675943 725915 717600 726083
rect 675887 725439 717600 725915
rect 675392 725222 675444 725286
rect 675943 725271 717600 725439
rect 675404 724831 675432 725222
rect 675887 724887 717600 725271
rect 675404 724812 675887 724831
rect 675407 724775 675887 724812
rect 675943 724719 717600 724887
rect 675887 724243 717600 724719
rect 675943 724075 717600 724243
rect 675887 723599 717600 724075
rect 675407 723529 675887 723543
rect 675220 723501 675887 723529
rect 675220 715525 675248 723501
rect 675407 723487 675887 723501
rect 675943 723431 717600 723599
rect 675887 722955 717600 723431
rect 675943 722787 717600 722955
rect 675887 722403 717600 722787
rect 675943 722235 717600 722403
rect 675887 721759 717600 722235
rect 675943 721591 717600 721759
rect 675887 721115 717600 721591
rect 675943 720947 717600 721115
rect 675887 720563 717600 720947
rect 675943 720395 717600 720563
rect 675887 719919 717600 720395
rect 675943 719751 717600 719919
rect 675887 719275 717600 719751
rect 675407 719163 675887 719219
rect 675943 719107 717600 719275
rect 675887 718723 717600 719107
rect 675943 718555 717600 718723
rect 675887 718079 717600 718555
rect 675943 717911 717600 718079
rect 675392 717810 675444 717874
rect 675404 717379 675432 717810
rect 675887 717435 717600 717911
rect 675404 717332 675887 717379
rect 675407 717323 675887 717332
rect 675943 717267 717600 717435
rect 675887 716883 717600 717267
rect 675407 716771 675887 716827
rect 675943 716715 717600 716883
rect 675887 716239 717600 716715
rect 675943 716071 717600 716239
rect 675887 715595 717600 716071
rect 675407 715525 675887 715539
rect 675220 715497 675887 715525
rect 675407 715483 675887 715497
rect 675943 715427 717600 715595
rect 675887 715217 717600 715427
rect 675128 709306 675340 709334
rect 675312 690014 675340 709306
rect 675128 689986 675340 690014
rect 675128 670694 675156 689986
rect 675887 686759 717600 686958
rect 675943 686591 717600 686759
rect 675887 686207 717600 686591
rect 675943 686039 717600 686207
rect 675887 685563 717600 686039
rect 675943 685395 717600 685563
rect 675887 684919 717600 685395
rect 675943 684751 717600 684919
rect 675887 684367 717600 684751
rect 675943 684199 717600 684367
rect 675887 683723 717600 684199
rect 675407 683639 675887 683667
rect 675404 683611 675887 683639
rect 675404 683126 675432 683611
rect 675943 683555 717600 683723
rect 675392 683062 675444 683126
rect 675887 683079 717600 683555
rect 675943 682911 717600 683079
rect 675887 682527 717600 682911
rect 675943 682359 717600 682527
rect 675887 681883 717600 682359
rect 675943 681715 717600 681883
rect 675887 681239 717600 681715
rect 675943 681071 717600 681239
rect 675887 680687 717600 681071
rect 675407 680612 675887 680631
rect 675404 680575 675887 680612
rect 675404 680474 675432 680575
rect 675943 680519 717600 680687
rect 675392 680410 675444 680474
rect 675887 680043 717600 680519
rect 675943 679875 717600 680043
rect 675887 679399 717600 679875
rect 675407 679315 675887 679343
rect 675404 679287 675887 679315
rect 675404 678842 675432 679287
rect 675943 679231 717600 679399
rect 675208 678778 675260 678842
rect 675392 678778 675444 678842
rect 675220 671325 675248 678778
rect 675887 678755 717600 679231
rect 675943 678587 717600 678755
rect 675887 678203 717600 678587
rect 675943 678035 717600 678203
rect 675887 677559 717600 678035
rect 675943 677391 717600 677559
rect 675887 676915 717600 677391
rect 675943 676747 717600 676915
rect 675887 676363 717600 676747
rect 675943 676195 717600 676363
rect 675887 675719 717600 676195
rect 675943 675551 717600 675719
rect 675887 675075 717600 675551
rect 675407 674963 675887 675019
rect 675943 674907 717600 675075
rect 675887 674523 717600 674907
rect 675943 674355 717600 674523
rect 675887 673879 717600 674355
rect 675943 673711 717600 673879
rect 675392 673610 675444 673674
rect 675404 673179 675432 673610
rect 675887 673235 717600 673711
rect 675404 673132 675887 673179
rect 675407 673123 675887 673132
rect 675943 673067 717600 673235
rect 675887 672683 717600 673067
rect 675407 672571 675887 672627
rect 675943 672515 717600 672683
rect 675887 672039 717600 672515
rect 675943 671871 717600 672039
rect 675887 671395 717600 671871
rect 675407 671325 675887 671339
rect 675220 671297 675887 671325
rect 675407 671283 675887 671297
rect 675943 671227 717600 671395
rect 675887 671017 717600 671227
rect 675128 670666 675340 670694
rect 675312 651374 675340 670666
rect 675128 651346 675340 651374
rect 675128 623774 675156 651346
rect 675887 642559 717600 642758
rect 675943 642391 717600 642559
rect 675887 642007 717600 642391
rect 675943 641839 717600 642007
rect 675887 641363 717600 641839
rect 675943 641195 717600 641363
rect 675887 640719 717600 641195
rect 675943 640551 717600 640719
rect 675887 640167 717600 640551
rect 675943 639999 717600 640167
rect 675887 639523 717600 639999
rect 675407 639439 675887 639467
rect 675404 639411 675887 639439
rect 675404 638926 675432 639411
rect 675943 639355 717600 639523
rect 675392 638862 675444 638926
rect 675887 638879 717600 639355
rect 675943 638711 717600 638879
rect 675887 638327 717600 638711
rect 675943 638159 717600 638327
rect 675887 637683 717600 638159
rect 675943 637515 717600 637683
rect 675887 637039 717600 637515
rect 675943 636871 717600 637039
rect 675887 636487 717600 636871
rect 675407 636412 675887 636431
rect 675404 636375 675887 636412
rect 675404 636342 675432 636375
rect 675392 636278 675444 636342
rect 675943 636319 717600 636487
rect 675887 635843 717600 636319
rect 675943 635675 717600 635843
rect 675887 635199 717600 635675
rect 675407 635115 675887 635143
rect 675404 635087 675887 635115
rect 675404 634642 675432 635087
rect 675943 635031 717600 635199
rect 675208 634578 675260 634642
rect 675392 634578 675444 634642
rect 675220 627125 675248 634578
rect 675887 634555 717600 635031
rect 675943 634387 717600 634555
rect 675887 634003 717600 634387
rect 675943 633835 717600 634003
rect 675887 633359 717600 633835
rect 675943 633191 717600 633359
rect 675887 632715 717600 633191
rect 675943 632547 717600 632715
rect 675887 632163 717600 632547
rect 675943 631995 717600 632163
rect 675887 631519 717600 631995
rect 675943 631351 717600 631519
rect 675887 630875 717600 631351
rect 675407 630763 675887 630819
rect 675943 630707 717600 630875
rect 675887 630323 717600 630707
rect 675943 630155 717600 630323
rect 675887 629679 717600 630155
rect 675943 629511 717600 629679
rect 675392 629410 675444 629474
rect 675404 628979 675432 629410
rect 675887 629035 717600 629511
rect 675404 628932 675887 628979
rect 675407 628923 675887 628932
rect 675943 628867 717600 629035
rect 675887 628483 717600 628867
rect 675407 628371 675887 628427
rect 675943 628315 717600 628483
rect 675887 627839 717600 628315
rect 675943 627671 717600 627839
rect 675887 627195 717600 627671
rect 675407 627125 675887 627139
rect 675220 627097 675887 627125
rect 675407 627083 675887 627097
rect 675943 627027 717600 627195
rect 675887 626817 717600 627027
rect 675128 623746 675340 623774
rect 675312 590322 675340 623746
rect 675887 598159 717600 598358
rect 675943 597991 717600 598159
rect 675887 597607 717600 597991
rect 675943 597439 717600 597607
rect 675887 596963 717600 597439
rect 675943 596795 717600 596963
rect 675887 596319 717600 596795
rect 675943 596151 717600 596319
rect 675887 595767 717600 596151
rect 675943 595599 717600 595767
rect 675392 595138 675444 595202
rect 675404 595067 675432 595138
rect 675887 595123 717600 595599
rect 675404 595039 675887 595067
rect 675407 595011 675887 595039
rect 675943 594955 717600 595123
rect 675887 594479 717600 594955
rect 675943 594311 717600 594479
rect 675887 593927 717600 594311
rect 675943 593759 717600 593927
rect 675887 593283 717600 593759
rect 675943 593115 717600 593283
rect 675887 592639 717600 593115
rect 675943 592471 717600 592639
rect 675887 592087 717600 592471
rect 675407 592003 675887 592031
rect 675404 591975 675887 592003
rect 675404 591938 675432 591975
rect 675392 591874 675444 591938
rect 675943 591919 717600 592087
rect 675887 591443 717600 591919
rect 675943 591275 717600 591443
rect 675887 590799 717600 591275
rect 675407 590716 675887 590743
rect 675128 590294 675340 590322
rect 675404 590687 675887 590716
rect 675128 535454 675156 590294
rect 675404 590186 675432 590687
rect 675943 590631 717600 590799
rect 675312 590158 675432 590186
rect 675312 583250 675340 590158
rect 675887 590155 717600 590631
rect 675943 589987 717600 590155
rect 675887 589603 717600 589987
rect 675943 589435 717600 589603
rect 675887 588959 717600 589435
rect 675943 588791 717600 588959
rect 675887 588315 717600 588791
rect 675943 588147 717600 588315
rect 675887 587763 717600 588147
rect 675943 587595 717600 587763
rect 675887 587119 717600 587595
rect 675943 586951 717600 587119
rect 675887 586475 717600 586951
rect 675407 586363 675887 586419
rect 675943 586307 717600 586475
rect 675887 585923 717600 586307
rect 675943 585755 717600 585923
rect 675887 585279 717600 585755
rect 675943 585111 717600 585279
rect 675887 584635 717600 585111
rect 675407 584551 675887 584579
rect 675404 584523 675887 584551
rect 675404 584186 675432 584523
rect 675943 584467 717600 584635
rect 675392 584122 675444 584186
rect 675887 584083 717600 584467
rect 675407 583971 675887 584027
rect 675943 583915 717600 584083
rect 675887 583439 717600 583915
rect 675943 583271 717600 583439
rect 675312 583222 675432 583250
rect 675404 582739 675432 583222
rect 675887 582795 717600 583271
rect 675404 582692 675887 582739
rect 675407 582683 675887 582692
rect 675943 582627 717600 582795
rect 675887 582417 717600 582627
rect 675887 553959 717600 554158
rect 675943 553791 717600 553959
rect 675887 553407 717600 553791
rect 675943 553239 717600 553407
rect 675887 552763 717600 553239
rect 675943 552595 717600 552763
rect 675887 552119 717600 552595
rect 675943 551951 717600 552119
rect 675887 551567 717600 551951
rect 675392 551346 675444 551410
rect 675943 551399 717600 551567
rect 675404 550867 675432 551346
rect 675887 550923 717600 551399
rect 675404 550839 675887 550867
rect 675407 550811 675887 550839
rect 675943 550755 717600 550923
rect 675887 550279 717600 550755
rect 675943 550111 717600 550279
rect 675887 549727 717600 550111
rect 675943 549559 717600 549727
rect 675887 549083 717600 549559
rect 675943 548915 717600 549083
rect 675887 548439 717600 548915
rect 675392 548218 675444 548282
rect 675943 548271 717600 548439
rect 675404 547831 675432 548218
rect 675887 547887 717600 548271
rect 675404 547803 675887 547831
rect 675407 547775 675887 547803
rect 675943 547719 717600 547887
rect 675887 547243 717600 547719
rect 675943 547075 717600 547243
rect 675887 546599 717600 547075
rect 675407 546530 675887 546543
rect 675312 546502 675887 546530
rect 675312 539050 675340 546502
rect 675407 546487 675887 546502
rect 675943 546431 717600 546599
rect 675887 545955 717600 546431
rect 675943 545787 717600 545955
rect 675887 545403 717600 545787
rect 675943 545235 717600 545403
rect 675887 544759 717600 545235
rect 675943 544591 717600 544759
rect 675887 544115 717600 544591
rect 675943 543947 717600 544115
rect 675887 543563 717600 543947
rect 675943 543395 717600 543563
rect 675887 542919 717600 543395
rect 675943 542751 717600 542919
rect 675887 542275 717600 542751
rect 675407 542163 675887 542219
rect 675943 542107 717600 542275
rect 675887 541723 717600 542107
rect 675943 541555 717600 541723
rect 675887 541079 717600 541555
rect 675392 540874 675444 540938
rect 675943 540911 717600 541079
rect 675404 540379 675432 540874
rect 675887 540435 717600 540911
rect 675404 540351 675887 540379
rect 675407 540323 675887 540351
rect 675943 540267 717600 540435
rect 675887 539883 717600 540267
rect 675407 539771 675887 539827
rect 675943 539715 717600 539883
rect 675887 539239 717600 539715
rect 675943 539071 717600 539239
rect 675312 539022 675432 539050
rect 675404 538539 675432 539022
rect 675887 538595 717600 539071
rect 675404 538492 675887 538539
rect 675407 538483 675887 538492
rect 675943 538427 717600 538595
rect 675887 538217 717600 538427
rect 675128 535426 675340 535454
rect 675312 499526 675340 535426
rect 678007 509901 716615 509947
rect 677600 505121 716615 509901
rect 677600 504421 677984 504821
rect 678007 499922 716615 505121
rect 675300 499462 675352 499526
rect 676128 499462 676180 499526
rect 676140 494902 676168 499462
rect 677600 495142 716615 499922
rect 676128 494838 676180 494902
rect 677968 494873 678020 494902
rect 677966 494799 678022 494873
rect 685910 466600 686840 468795
rect 678007 466500 717593 466600
rect 678000 462501 717593 466500
rect 678007 462415 717593 462501
rect 678000 455893 717593 462415
rect 678007 455781 717593 455893
rect 678000 451660 717593 455781
rect 678007 451600 717593 451660
rect 682685 449413 685567 451360
rect 685917 449372 686847 451600
rect 687319 449413 717593 451360
rect 678007 423301 716615 423347
rect 674012 422214 674064 422278
rect 674748 422214 674800 422278
rect 674024 419937 674052 422214
rect 674010 419863 674066 419937
rect 674010 419183 674066 419257
rect 674012 419154 674064 419183
rect 677508 419154 677560 419218
rect 677520 418441 677548 419154
rect 677600 418521 716615 423301
rect 677506 418367 677562 418441
rect 677600 417821 677984 418221
rect 678007 413322 716615 418521
rect 677600 408542 716615 413322
rect 675887 379759 717600 379958
rect 675943 379591 717600 379759
rect 675887 379207 717600 379591
rect 675943 379039 717600 379207
rect 675887 378563 717600 379039
rect 675943 378395 717600 378563
rect 675887 377919 717600 378395
rect 675943 377751 717600 377919
rect 675887 377367 717600 377751
rect 673920 376110 673972 376174
rect 673736 373050 673788 373114
rect 42616 361286 42668 361350
rect 42524 325654 42576 325718
rect 42536 322934 42564 325654
rect 42444 322906 42564 322934
rect 0 317713 41657 317881
rect 41713 317769 42193 317825
rect 0 317329 41713 317713
rect 41800 317422 41828 317769
rect 41788 317358 41840 317422
rect 0 317161 41657 317329
rect 0 316685 41713 317161
rect 0 316517 41657 316685
rect 0 316041 41713 316517
rect 0 315873 41657 316041
rect 0 315489 41713 315873
rect 0 315321 41657 315489
rect 0 314845 41713 315321
rect 0 314677 41657 314845
rect 41713 314733 42193 314789
rect 0 314201 41713 314677
rect 41800 314294 41828 314733
rect 41788 314230 41840 314294
rect 0 314033 41657 314201
rect 0 313649 41713 314033
rect 0 313481 41657 313649
rect 0 313005 41713 313481
rect 42444 313018 42472 322906
rect 42628 317422 42656 361286
rect 42708 357614 42760 357678
rect 42616 317358 42668 317422
rect 42524 314230 42576 314294
rect 0 312837 41657 313005
rect 42260 312990 42472 313018
rect 0 312361 41713 312837
rect 0 312193 41657 312361
rect 0 311809 41713 312193
rect 0 311641 41657 311809
rect 0 311442 41713 311641
rect 0 283973 41713 284183
rect 42260 284050 42288 312990
rect 42260 284022 42472 284050
rect 0 283805 41657 283973
rect 41713 283914 42193 283917
rect 41713 283886 42288 283914
rect 41713 283861 42193 283886
rect 0 283329 41713 283805
rect 0 283161 41657 283329
rect 0 282685 41713 283161
rect 0 282517 41657 282685
rect 41713 282573 42193 282629
rect 0 282133 41713 282517
rect 0 281965 41657 282133
rect 41713 282021 42193 282077
rect 0 281489 41713 281965
rect 41800 281586 41828 282021
rect 41788 281522 41840 281586
rect 0 281321 41657 281489
rect 0 280845 41713 281321
rect 0 280677 41657 280845
rect 0 280293 41713 280677
rect 0 280125 41657 280293
rect 41713 280181 42193 280237
rect 0 279649 41713 280125
rect 0 279481 41657 279649
rect 0 279005 41713 279481
rect 0 278837 41657 279005
rect 0 278453 41713 278837
rect 0 278285 41657 278453
rect 0 277809 41713 278285
rect 0 277641 41657 277809
rect 0 277165 41713 277641
rect 0 276997 41657 277165
rect 0 276613 41713 276997
rect 0 276445 41657 276613
rect 0 275969 41713 276445
rect 42260 276026 42288 283886
rect 41800 275998 42288 276026
rect 0 275801 41657 275969
rect 41800 275913 41828 275998
rect 41713 275857 42193 275913
rect 0 275325 41713 275801
rect 42444 281586 42472 284022
rect 42432 281522 42484 281586
rect 0 275157 41657 275325
rect 0 274681 41713 275157
rect 0 274513 41657 274681
rect 41788 274654 41840 274718
rect 41800 274625 41828 274654
rect 41713 274569 42193 274625
rect 0 274129 41713 274513
rect 0 273961 41657 274129
rect 0 273485 41713 273961
rect 0 273317 41657 273485
rect 0 272841 41713 273317
rect 0 272673 41657 272841
rect 0 272289 41713 272673
rect 0 272121 41657 272289
rect 0 271645 41713 272121
rect 41788 272070 41840 272134
rect 0 271477 41657 271645
rect 41800 271589 41828 272070
rect 41713 271533 42193 271589
rect 0 271001 41713 271477
rect 0 270833 41657 271001
rect 42536 272134 42564 314230
rect 42628 274718 42656 317358
rect 42720 314294 42748 357614
rect 673748 334014 673776 373050
rect 673736 333950 673788 334014
rect 673932 331974 673960 376110
rect 675943 377199 717600 377367
rect 675887 376723 717600 377199
rect 675407 376652 675887 376667
rect 675404 376611 675887 376652
rect 675404 376174 675432 376611
rect 675943 376555 717600 376723
rect 675392 376110 675444 376174
rect 675887 376079 717600 376555
rect 675943 375911 717600 376079
rect 675887 375527 717600 375911
rect 675943 375359 717600 375527
rect 675887 374883 717600 375359
rect 675943 374715 717600 374883
rect 675887 374239 717600 374715
rect 675943 374071 717600 374239
rect 675887 373687 717600 374071
rect 675407 373603 675887 373631
rect 675404 373575 675887 373603
rect 675404 373114 675432 373575
rect 675943 373519 717600 373687
rect 675392 373050 675444 373114
rect 675887 373043 717600 373519
rect 675943 372875 717600 373043
rect 675887 372399 717600 372875
rect 675407 372314 675887 372343
rect 675312 372287 675887 372314
rect 675312 372286 675418 372287
rect 674012 365706 674064 365770
rect 673460 331910 673512 331974
rect 673920 331910 673972 331974
rect 42708 314230 42760 314294
rect 673472 288794 673500 331910
rect 673552 328850 673604 328914
rect 673460 288730 673512 288794
rect 42708 281522 42760 281586
rect 42616 274654 42668 274718
rect 42524 272070 42576 272134
rect 0 270449 41713 270833
rect 0 270281 41657 270449
rect 0 269805 41713 270281
rect 0 269637 41657 269805
rect 0 269161 41713 269637
rect 0 268993 41657 269161
rect 0 268609 41713 268993
rect 0 268441 41657 268609
rect 0 268242 41713 268441
rect 0 240773 41713 240983
rect 0 240605 41657 240773
rect 41713 240703 42193 240717
rect 41713 240675 42288 240703
rect 41713 240661 42193 240675
rect 0 240129 41713 240605
rect 0 239961 41657 240129
rect 0 239485 41713 239961
rect 0 239317 41657 239485
rect 41713 239373 42193 239429
rect 0 238933 41713 239317
rect 0 238765 41657 238933
rect 41713 238821 42193 238877
rect 0 238289 41713 238765
rect 41800 238338 41828 238821
rect 0 238121 41657 238289
rect 41788 238274 41840 238338
rect 0 237645 41713 238121
rect 0 237477 41657 237645
rect 41713 237533 42193 237589
rect 0 237093 41713 237477
rect 0 236925 41657 237093
rect 41713 236981 42193 237037
rect 0 236449 41713 236925
rect 0 236281 41657 236449
rect 0 235805 41713 236281
rect 0 235637 41657 235805
rect 41713 235693 42193 235749
rect 0 235253 41713 235637
rect 0 235085 41657 235253
rect 0 234609 41713 235085
rect 0 234441 41657 234609
rect 0 233965 41713 234441
rect 0 233797 41657 233965
rect 0 233413 41713 233797
rect 0 233245 41657 233413
rect 0 232769 41713 233245
rect 42260 232778 42288 240675
rect 0 232601 41657 232769
rect 41800 232750 42288 232778
rect 41800 232713 41828 232750
rect 41713 232657 42193 232713
rect 0 232125 41713 232601
rect 42432 238274 42484 238338
rect 0 231957 41657 232125
rect 0 231481 41713 231957
rect 41788 231882 41840 231946
rect 0 231313 41657 231481
rect 41800 231425 41828 231882
rect 41713 231369 42193 231425
rect 0 230929 41713 231313
rect 0 230761 41657 230929
rect 0 230285 41713 230761
rect 0 230117 41657 230285
rect 0 229641 41713 230117
rect 0 229473 41657 229641
rect 0 229089 41713 229473
rect 0 228921 41657 229089
rect 0 228445 41713 228921
rect 41788 228822 41840 228886
rect 0 228277 41657 228445
rect 41800 228389 41828 228822
rect 41713 228333 42193 228389
rect 0 227801 41713 228277
rect 0 227633 41657 227801
rect 0 227249 41713 227633
rect 0 227081 41657 227249
rect 0 226605 41713 227081
rect 0 226437 41657 226605
rect 0 225961 41713 226437
rect 0 225793 41657 225961
rect 0 225409 41713 225793
rect 0 225241 41657 225409
rect 0 225042 41713 225241
rect 0 197573 41713 197783
rect 0 197405 41657 197573
rect 41713 197503 42193 197517
rect 41713 197475 42288 197503
rect 41713 197461 42193 197475
rect 0 196929 41713 197405
rect 0 196761 41657 196929
rect 0 196285 41713 196761
rect 0 196117 41657 196285
rect 41713 196173 42193 196229
rect 0 195733 41713 196117
rect 0 195565 41657 195733
rect 41713 195621 42193 195677
rect 0 195089 41713 195565
rect 41800 195158 41828 195621
rect 41788 195094 41840 195158
rect 0 194921 41657 195089
rect 0 194445 41713 194921
rect 0 194277 41657 194445
rect 41713 194333 42193 194389
rect 0 193893 41713 194277
rect 0 193725 41657 193893
rect 41713 193781 42193 193837
rect 0 193249 41713 193725
rect 0 193081 41657 193249
rect 0 192605 41713 193081
rect 0 192437 41657 192605
rect 41713 192493 42193 192549
rect 0 192053 41713 192437
rect 0 191885 41657 192053
rect 0 191409 41713 191885
rect 0 191241 41657 191409
rect 0 190765 41713 191241
rect 0 190597 41657 190765
rect 0 190213 41713 190597
rect 0 190045 41657 190213
rect 0 189569 41713 190045
rect 0 189401 41657 189569
rect 42260 189530 42288 197475
rect 41708 189502 42288 189530
rect 41708 189485 42193 189502
rect 41713 189457 42193 189485
rect 0 188925 41713 189401
rect 42444 195158 42472 238274
rect 42536 228886 42564 272070
rect 42628 231946 42656 274654
rect 42720 238338 42748 281522
rect 673472 243778 673500 288730
rect 673564 285326 673592 328850
rect 673644 322458 673696 322522
rect 673552 285262 673604 285326
rect 673460 243714 673512 243778
rect 42708 238274 42760 238338
rect 42616 231882 42668 231946
rect 42628 231826 42656 231882
rect 42628 231798 42840 231826
rect 42524 228822 42576 228886
rect 42536 226334 42564 228822
rect 42536 226306 42748 226334
rect 42432 195094 42484 195158
rect 0 188757 41657 188925
rect 0 188281 41713 188757
rect 41788 188702 41840 188766
rect 0 188113 41657 188281
rect 41800 188225 41828 188702
rect 41713 188169 42193 188225
rect 0 187729 41713 188113
rect 0 187561 41657 187729
rect 0 187085 41713 187561
rect 0 186917 41657 187085
rect 0 186441 41713 186917
rect 0 186273 41657 186441
rect 0 185889 41713 186273
rect 0 185721 41657 185889
rect 0 185245 41713 185721
rect 41788 185642 41840 185706
rect 0 185077 41657 185245
rect 41800 185189 41828 185642
rect 41713 185133 42193 185189
rect 0 184601 41713 185077
rect 0 184433 41657 184601
rect 0 184049 41713 184433
rect 42248 184350 42300 184414
rect 0 183881 41657 184049
rect 0 183405 41713 183881
rect 0 183237 41657 183405
rect 0 182761 41713 183237
rect 0 182593 41657 182761
rect 0 182209 41713 182593
rect 0 182041 41657 182209
rect 0 181842 41713 182041
rect 985 120278 40000 125058
rect 985 115079 39593 120278
rect 39616 115379 40000 115779
rect 985 110299 40000 115079
rect 985 110253 39593 110299
rect 30753 83000 31683 85228
rect 31928 83049 32702 85239
rect 714 82940 39593 83000
rect 714 78819 39600 82940
rect 39670 80135 39726 80209
rect 714 78707 39593 78819
rect 714 72185 39600 78707
rect 39684 78305 39712 80135
rect 39670 78231 39726 78305
rect 714 72099 39593 72185
rect 714 68100 39600 72099
rect 714 68098 39593 68100
rect 42260 45694 42288 184350
rect 42248 45630 42300 45694
rect 42444 106078 42472 195094
rect 42524 188702 42576 188766
rect 42536 121514 42564 188702
rect 42720 185706 42748 226306
rect 42812 188766 42840 231798
rect 673472 199170 673500 243714
rect 673564 240310 673592 285262
rect 673656 277370 673684 322458
rect 674024 322522 674052 365706
rect 675312 364325 675340 372286
rect 675943 372231 717600 372399
rect 675887 371755 717600 372231
rect 675943 371587 717600 371755
rect 675887 371203 717600 371587
rect 675943 371035 717600 371203
rect 675887 370559 717600 371035
rect 675943 370391 717600 370559
rect 675887 369915 717600 370391
rect 675943 369747 717600 369915
rect 675887 369363 717600 369747
rect 675407 369251 675887 369307
rect 675943 369195 717600 369363
rect 675887 368719 717600 369195
rect 675943 368551 717600 368719
rect 675887 368075 717600 368551
rect 675407 367963 675887 368019
rect 675943 367907 717600 368075
rect 675887 367523 717600 367907
rect 675407 367411 675887 367467
rect 675943 367355 717600 367523
rect 675887 366879 717600 367355
rect 675943 366711 717600 366879
rect 675887 366235 717600 366711
rect 675407 366151 675887 366179
rect 675404 366123 675887 366151
rect 675404 365770 675432 366123
rect 675943 366067 717600 366235
rect 675392 365706 675444 365770
rect 675887 365683 717600 366067
rect 675407 365571 675887 365627
rect 675943 365515 717600 365683
rect 675887 365039 717600 365515
rect 675943 364871 717600 365039
rect 675887 364395 717600 364871
rect 675407 364325 675887 364339
rect 675312 364297 675887 364325
rect 675407 364283 675887 364297
rect 675943 364227 717600 364395
rect 675887 364017 717600 364227
rect 675887 335559 717600 335758
rect 675943 335391 717600 335559
rect 675887 335007 717600 335391
rect 675943 334839 717600 335007
rect 675887 334363 717600 334839
rect 675943 334195 717600 334363
rect 675208 333950 675260 334014
rect 675220 328914 675248 333950
rect 675887 333719 717600 334195
rect 675943 333551 717600 333719
rect 675887 333167 717600 333551
rect 675208 328850 675260 328914
rect 675943 332999 717600 333167
rect 675887 332523 717600 332999
rect 675407 332452 675887 332467
rect 675404 332411 675887 332452
rect 675404 331974 675432 332411
rect 675943 332355 717600 332523
rect 675392 331910 675444 331974
rect 675887 331879 717600 332355
rect 675943 331711 717600 331879
rect 675887 331327 717600 331711
rect 675943 331159 717600 331327
rect 675887 330683 717600 331159
rect 675943 330515 717600 330683
rect 675887 330039 717600 330515
rect 675943 329871 717600 330039
rect 675887 329487 717600 329871
rect 675407 329403 675887 329431
rect 675404 329375 675887 329403
rect 675404 328914 675432 329375
rect 675943 329319 717600 329487
rect 675392 328850 675444 328914
rect 675887 328843 717600 329319
rect 675943 328675 717600 328843
rect 675887 328199 717600 328675
rect 675407 328114 675887 328143
rect 675312 328087 675887 328114
rect 675312 328086 675418 328087
rect 674012 322458 674064 322522
rect 675312 320125 675340 328086
rect 675943 328031 717600 328199
rect 675887 327555 717600 328031
rect 675943 327387 717600 327555
rect 675887 327003 717600 327387
rect 675943 326835 717600 327003
rect 675887 326359 717600 326835
rect 675943 326191 717600 326359
rect 675887 325715 717600 326191
rect 675943 325547 717600 325715
rect 675887 325163 717600 325547
rect 675407 325051 675887 325107
rect 675943 324995 717600 325163
rect 675887 324519 717600 324995
rect 675943 324351 717600 324519
rect 675887 323875 717600 324351
rect 675407 323763 675887 323819
rect 675943 323707 717600 323875
rect 675887 323323 717600 323707
rect 675407 323211 675887 323267
rect 675943 323155 717600 323323
rect 675887 322679 717600 323155
rect 675392 322458 675444 322522
rect 675943 322511 717600 322679
rect 675404 321979 675432 322458
rect 675887 322035 717600 322511
rect 675404 321951 675887 321979
rect 675407 321923 675887 321951
rect 675943 321867 717600 322035
rect 675887 321483 717600 321867
rect 675407 321371 675887 321427
rect 675943 321315 717600 321483
rect 675887 320839 717600 321315
rect 675943 320671 717600 320839
rect 675887 320195 717600 320671
rect 675407 320125 675887 320139
rect 675312 320097 675887 320125
rect 675407 320083 675887 320097
rect 675943 320027 717600 320195
rect 675887 319817 717600 320027
rect 675887 291359 717600 291558
rect 675943 291191 717600 291359
rect 675887 290807 717600 291191
rect 675943 290639 717600 290807
rect 675887 290163 717600 290639
rect 675943 289995 717600 290163
rect 675887 289519 717600 289995
rect 675943 289351 717600 289519
rect 675887 288967 717600 289351
rect 675943 288799 717600 288967
rect 675392 288730 675444 288794
rect 675404 288267 675432 288730
rect 675887 288323 717600 288799
rect 675404 288252 675887 288267
rect 675407 288211 675887 288252
rect 675943 288155 717600 288323
rect 675887 287679 717600 288155
rect 675943 287511 717600 287679
rect 675887 287127 717600 287511
rect 675943 286959 717600 287127
rect 675887 286483 717600 286959
rect 675943 286315 717600 286483
rect 675887 285839 717600 286315
rect 675943 285671 717600 285839
rect 675392 285262 675444 285326
rect 675887 285287 717600 285671
rect 675404 285231 675432 285262
rect 675404 285203 675887 285231
rect 675407 285175 675887 285203
rect 675943 285119 717600 285287
rect 675887 284643 717600 285119
rect 675943 284475 717600 284643
rect 673644 277306 673696 277370
rect 673552 240246 673604 240310
rect 673460 199106 673512 199170
rect 42800 188702 42852 188766
rect 42708 185642 42760 185706
rect 42720 184414 42748 185642
rect 42708 184350 42760 184414
rect 673472 155990 673500 199106
rect 673564 197062 673592 240246
rect 673656 233918 673684 277306
rect 675887 283999 717600 284475
rect 675407 283914 675887 283943
rect 675312 283887 675887 283914
rect 675312 283886 675418 283887
rect 675312 275925 675340 283886
rect 675943 283831 717600 283999
rect 675887 283355 717600 283831
rect 675943 283187 717600 283355
rect 675887 282803 717600 283187
rect 675943 282635 717600 282803
rect 675887 282159 717600 282635
rect 675943 281991 717600 282159
rect 675887 281515 717600 281991
rect 675943 281347 717600 281515
rect 675887 280963 717600 281347
rect 675407 280851 675887 280907
rect 675943 280795 717600 280963
rect 675887 280319 717600 280795
rect 675943 280151 717600 280319
rect 675887 279675 717600 280151
rect 675407 279563 675887 279619
rect 675943 279507 717600 279675
rect 675887 279123 717600 279507
rect 675407 279011 675887 279067
rect 675943 278955 717600 279123
rect 675887 278479 717600 278955
rect 675943 278311 717600 278479
rect 675887 277835 717600 278311
rect 675407 277751 675887 277779
rect 675404 277723 675887 277751
rect 675404 277370 675432 277723
rect 675943 277667 717600 277835
rect 675392 277306 675444 277370
rect 675887 277283 717600 277667
rect 675407 277171 675887 277227
rect 675943 277115 717600 277283
rect 675887 276639 717600 277115
rect 675943 276471 717600 276639
rect 675887 275995 717600 276471
rect 675407 275925 675887 275939
rect 675312 275897 675887 275925
rect 675407 275883 675887 275897
rect 675943 275827 717600 275995
rect 675887 275617 717600 275827
rect 675887 246959 717600 247158
rect 675943 246791 717600 246959
rect 675887 246407 717600 246791
rect 675943 246239 717600 246407
rect 675887 245763 717600 246239
rect 675943 245595 717600 245763
rect 675887 245119 717600 245595
rect 675943 244951 717600 245119
rect 675887 244567 717600 244951
rect 675943 244399 717600 244567
rect 675887 243923 717600 244399
rect 675407 243839 675887 243867
rect 675404 243811 675887 243839
rect 675404 243778 675432 243811
rect 675392 243714 675444 243778
rect 675943 243755 717600 243923
rect 675887 243279 717600 243755
rect 675943 243111 717600 243279
rect 675887 242727 717600 243111
rect 675943 242559 717600 242727
rect 675887 242083 717600 242559
rect 675943 241915 717600 242083
rect 675887 241439 717600 241915
rect 675943 241271 717600 241439
rect 675887 240887 717600 241271
rect 675407 240788 675887 240831
rect 675404 240775 675887 240788
rect 675404 240310 675432 240775
rect 675943 240719 717600 240887
rect 675392 240246 675444 240310
rect 675887 240243 717600 240719
rect 675943 240075 717600 240243
rect 673644 233854 673696 233918
rect 673552 196998 673604 197062
rect 673460 155926 673512 155990
rect 673564 152862 673592 196998
rect 673656 189310 673684 233854
rect 675887 239599 717600 240075
rect 675407 239529 675887 239543
rect 675312 239501 675887 239529
rect 675312 231525 675340 239501
rect 675407 239487 675887 239501
rect 675943 239431 717600 239599
rect 675887 238955 717600 239431
rect 675943 238787 717600 238955
rect 675887 238403 717600 238787
rect 675943 238235 717600 238403
rect 675887 237759 717600 238235
rect 675943 237591 717600 237759
rect 675887 237115 717600 237591
rect 675943 236947 717600 237115
rect 675887 236563 717600 236947
rect 675407 236451 675887 236507
rect 675943 236395 717600 236563
rect 675887 235919 717600 236395
rect 675943 235751 717600 235919
rect 675887 235275 717600 235751
rect 675407 235163 675887 235219
rect 675943 235107 717600 235275
rect 675887 234723 717600 235107
rect 675407 234611 675887 234667
rect 675943 234555 717600 234723
rect 675887 234079 717600 234555
rect 675392 233854 675444 233918
rect 675943 233911 717600 234079
rect 675404 233379 675432 233854
rect 675887 233435 717600 233911
rect 675404 233351 675887 233379
rect 675407 233323 675887 233351
rect 675943 233267 717600 233435
rect 675887 232883 717600 233267
rect 675407 232771 675887 232827
rect 675943 232715 717600 232883
rect 675887 232239 717600 232715
rect 675943 232071 717600 232239
rect 675887 231595 717600 232071
rect 675407 231525 675887 231539
rect 675312 231497 675887 231525
rect 675407 231483 675887 231497
rect 675943 231427 717600 231595
rect 675887 231217 717600 231427
rect 675887 202759 717600 202958
rect 675943 202591 717600 202759
rect 675887 202207 717600 202591
rect 675943 202039 717600 202207
rect 675887 201563 717600 202039
rect 675943 201395 717600 201563
rect 675887 200919 717600 201395
rect 675943 200751 717600 200919
rect 675887 200367 717600 200751
rect 675943 200199 717600 200367
rect 675887 199723 717600 200199
rect 675407 199639 675887 199667
rect 675404 199611 675887 199639
rect 675404 199170 675432 199611
rect 675943 199555 717600 199723
rect 675392 199106 675444 199170
rect 675887 199079 717600 199555
rect 675943 198911 717600 199079
rect 675887 198527 717600 198911
rect 675943 198359 717600 198527
rect 675887 197883 717600 198359
rect 675943 197715 717600 197883
rect 675887 197239 717600 197715
rect 675943 197071 717600 197239
rect 675392 196998 675444 197062
rect 675404 196631 675432 196998
rect 675887 196687 717600 197071
rect 675404 196588 675887 196631
rect 675407 196575 675887 196588
rect 675943 196519 717600 196687
rect 675887 196043 717600 196519
rect 675943 195875 717600 196043
rect 673644 189246 673696 189310
rect 673552 152798 673604 152862
rect 42524 121450 42576 121514
rect 44180 121450 44232 121514
rect 44192 110537 44220 121450
rect 673460 111522 673512 111586
rect 44178 110463 44234 110537
rect 44822 110463 44878 110537
rect 44836 110414 44864 110463
rect 44836 110386 44956 110414
rect 42432 106014 42484 106078
rect 44180 106014 44232 106078
rect 44192 80209 44220 106014
rect 44178 80135 44234 80209
rect 44822 80135 44878 80209
rect 44836 46986 44864 80135
rect 44824 46922 44876 46986
rect 44928 45558 44956 110386
rect 143540 46854 143592 46918
rect 140964 45630 141016 45694
rect 44916 45494 44968 45558
rect 93768 41482 93820 41546
rect 93780 40225 93808 41482
rect 135168 40225 135220 40254
rect 93766 40151 93822 40225
rect 135166 40151 135222 40225
rect 140976 40202 141004 45630
rect 143552 40497 143580 46854
rect 151726 46815 151782 46889
rect 188526 46815 188582 46889
rect 200856 46854 200908 46918
rect 256240 46854 256292 46918
rect 297732 46854 297784 46918
rect 309416 46854 309468 46918
rect 352564 46854 352616 46918
rect 364248 46854 364300 46918
rect 407396 46854 407448 46918
rect 419080 46854 419132 46918
rect 462136 46854 462188 46918
rect 473820 46854 473872 46918
rect 516968 46854 517020 46918
rect 143538 40423 143594 40497
rect 143540 40225 143592 40254
rect 140976 40174 141036 40202
rect 141008 40118 141036 40174
rect 143078 40151 143134 40225
rect 143538 40151 143594 40225
rect 146300 41822 146352 41886
rect 143084 40118 143112 40151
rect 140996 40054 141048 40118
rect 143072 40054 143124 40118
rect 144552 40054 144604 40118
rect 141008 40000 141036 40054
rect 143084 40000 143112 40054
rect 144564 40000 144592 40054
rect 146312 40118 146340 41822
rect 151740 40497 151768 46815
rect 186688 45562 186740 45626
rect 186700 42193 186728 45562
rect 188540 44402 188568 46815
rect 194692 45562 194744 45626
rect 188528 44338 188580 44402
rect 192852 44338 192904 44402
rect 188540 42193 188568 44338
rect 192864 42193 192892 44338
rect 194704 42193 194732 45562
rect 195980 45494 196032 45558
rect 195992 44334 196020 45494
rect 195980 44270 196032 44334
rect 195992 42193 196020 44270
rect 200868 42193 200896 46854
rect 201500 44270 201552 44334
rect 201512 42193 201540 44270
rect 186683 41713 186739 42193
rect 187971 41713 188027 42193
rect 188523 41713 188579 42193
rect 189167 41834 189223 42193
rect 189264 41890 189316 41954
rect 189276 41834 189304 41890
rect 189167 41806 189304 41834
rect 189167 41713 189223 41806
rect 189811 41713 189867 42193
rect 190363 41713 190419 42193
rect 191007 41834 191063 42193
rect 191104 41890 191156 41954
rect 191116 41834 191144 41890
rect 191007 41806 191144 41834
rect 191007 41713 191063 41806
rect 191651 41713 191707 42193
rect 192203 41834 192259 42193
rect 192300 41890 192352 41954
rect 192312 41834 192340 41890
rect 192203 41806 192340 41834
rect 192203 41713 192259 41806
rect 192847 41713 192903 42193
rect 193491 41834 193547 42193
rect 193588 41890 193640 41954
rect 193600 41834 193628 41890
rect 193491 41806 193628 41834
rect 193491 41713 193547 41806
rect 194687 41713 194743 42193
rect 195975 41713 196031 42193
rect 196440 41890 196492 41954
rect 196452 41834 196480 41890
rect 196527 41834 196583 42193
rect 197171 41834 197227 42193
rect 197815 41834 197871 42193
rect 198367 41834 198423 42193
rect 198464 41890 198516 41954
rect 198476 41834 198504 41890
rect 199011 41834 199067 42193
rect 196452 41806 198504 41834
rect 198936 41818 199067 41834
rect 198924 41806 199067 41818
rect 196527 41713 196583 41806
rect 197171 41713 197227 41806
rect 197815 41713 197871 41806
rect 198367 41713 198423 41806
rect 198924 41754 198976 41806
rect 199011 41713 199067 41806
rect 200120 41890 200172 41954
rect 200132 41834 200160 41890
rect 200207 41834 200263 42193
rect 200851 41834 200907 42193
rect 200132 41806 200907 41834
rect 200207 41713 200263 41806
rect 200851 41713 200907 41806
rect 201495 41713 201551 42193
rect 202047 41713 202103 42193
rect 186417 41657 186627 41713
rect 186795 41657 187271 41713
rect 187439 41657 187915 41713
rect 188083 41657 188467 41713
rect 188635 41657 189111 41713
rect 189279 41657 189755 41713
rect 189923 41657 190307 41713
rect 190475 41657 190951 41713
rect 191119 41657 191595 41713
rect 191763 41657 192147 41713
rect 192315 41657 192791 41713
rect 192959 41657 193435 41713
rect 193603 41657 193987 41713
rect 194155 41657 194631 41713
rect 194799 41657 195275 41713
rect 195443 41657 195919 41713
rect 196087 41657 196471 41713
rect 196639 41657 197115 41713
rect 197283 41657 197759 41713
rect 197927 41657 198311 41713
rect 198479 41657 198955 41713
rect 199123 41657 199599 41713
rect 199767 41657 200151 41713
rect 200319 41657 200795 41713
rect 200963 41657 201439 41713
rect 201607 41657 201991 41713
rect 202159 41657 202358 41713
rect 151726 40423 151782 40497
rect 146300 40054 146352 40118
rect 78942 39593 83722 40000
rect 88221 39616 88621 40000
rect 88921 39593 93701 40000
rect 132617 39878 132897 40000
rect 132953 39934 133157 40000
rect 133213 39878 140940 40000
rect 132617 39816 140940 39878
rect 140996 39872 141048 40000
rect 141104 39878 141313 40000
rect 141369 39934 141499 40000
rect 141555 39878 141611 40000
rect 141667 39934 141813 40000
rect 141869 39878 141898 40000
rect 141954 39934 142084 40000
rect 142140 39878 143012 40000
rect 141104 39816 143012 39878
rect 78942 985 93747 39593
rect 132617 39204 143012 39816
rect 132617 39147 142955 39204
rect 143068 39151 143128 40000
rect 143184 39662 143299 40000
rect 143355 39718 143585 40000
rect 143641 39831 143762 40000
rect 143818 39887 144151 40000
rect 144207 39831 144517 40000
rect 144564 39916 144689 40000
rect 143641 39747 144517 39831
rect 144573 39803 144689 39916
rect 144745 39747 145035 40000
rect 143641 39662 145035 39747
rect 145199 39878 145765 40000
rect 145821 39934 145915 40000
rect 145971 39878 147532 40000
rect 143184 39650 145035 39662
rect 145199 39650 147532 39878
rect 143184 39369 147532 39650
rect 143184 39297 144495 39369
rect 145520 39341 147532 39369
rect 143184 39243 144441 39297
rect 144551 39285 145464 39313
rect 144551 39271 145530 39285
rect 145586 39275 147532 39341
rect 144551 39261 145436 39271
rect 143184 39207 144367 39243
rect 144551 39241 144623 39261
rect 144625 39241 144645 39261
rect 145414 39247 145461 39261
rect 145464 39247 145530 39271
rect 143244 39169 144367 39207
rect 144497 39233 144551 39241
rect 144571 39233 144625 39241
rect 144497 39205 144625 39233
rect 145414 39219 145530 39247
rect 145414 39214 145461 39219
rect 144497 39187 144551 39205
rect 144571 39187 144625 39205
rect 143068 39148 143188 39151
rect 132617 39076 141720 39147
rect 143011 39091 143188 39148
rect 143244 39147 144345 39169
rect 144423 39113 144571 39187
rect 144701 39185 145358 39205
rect 144681 39158 145358 39185
rect 145461 39191 145525 39214
rect 145530 39191 145599 39219
rect 145655 39206 147532 39275
rect 145461 39163 145599 39191
rect 144681 39131 145405 39158
rect 145461 39150 145525 39163
rect 145530 39150 145599 39163
rect 144401 39091 144497 39113
rect 132617 39010 141654 39076
rect 141776 39063 144497 39091
rect 141776 39049 141847 39063
rect 143068 39049 143128 39063
rect 144423 39049 144497 39063
rect 144627 39094 145405 39131
rect 145525 39135 145591 39150
rect 145599 39135 145653 39150
rect 144627 39057 145469 39094
rect 145525 39085 145653 39135
rect 145525 39084 145591 39085
rect 141776 39039 144497 39049
rect 141776 39020 141847 39039
rect 141850 39020 141869 39039
rect 144553 39028 145469 39057
rect 141710 39011 141776 39020
rect 141784 39011 141850 39020
rect 132617 37861 141628 39010
rect 141710 38969 141850 39011
rect 144553 38983 145545 39028
rect 141710 38954 141776 38969
rect 141784 38954 141850 38969
rect 141925 38964 145545 38983
rect 141684 38928 141710 38954
rect 141736 38928 141784 38954
rect 141684 38906 141784 38928
rect 132617 37823 141590 37861
rect 132617 36927 141538 37823
rect 141684 37805 141736 38906
rect 141906 38898 145545 38964
rect 141840 38850 145545 38898
rect 141646 37783 141736 37805
rect 141646 37767 141684 37783
rect 141720 37767 141736 37783
rect 141792 38284 145545 38850
rect 141792 38216 145477 38284
rect 145601 38228 145653 39085
rect 141792 38176 145437 38216
rect 145533 38178 145653 38228
rect 141792 38110 145371 38176
rect 145533 38160 145601 38178
rect 145607 38160 145653 38178
rect 145493 38150 145533 38160
rect 145567 38150 145607 38160
rect 145493 38136 145607 38150
rect 145493 38120 145533 38136
rect 145567 38120 145607 38136
rect 141594 37693 141720 37767
rect 141792 37711 145319 38110
rect 145427 38108 145493 38120
rect 145501 38108 145567 38120
rect 145427 38080 145567 38108
rect 145709 38104 147532 39206
rect 145427 38054 145493 38080
rect 145501 38054 145567 38080
rect 145663 38064 147532 38104
rect 132617 36860 141471 36927
rect 141594 36871 141646 37693
rect 141776 37637 145319 37711
rect 132617 35845 141419 36860
rect 141527 36821 141646 36871
rect 141527 36804 141594 36821
rect 141601 36804 141646 36821
rect 141475 36730 141601 36804
rect 141702 36748 145319 37637
rect 141475 35901 141527 36730
rect 141657 36674 145319 36748
rect 141583 35845 145319 36674
rect 132617 34484 145319 35845
rect 145375 37980 145501 38054
rect 145623 37998 147532 38064
rect 145375 34678 145427 37980
rect 145557 37924 147532 37998
rect 145483 34734 147532 37924
rect 145375 34540 145470 34678
rect 132617 34469 145362 34484
rect 132617 33839 145319 34469
rect 145418 34413 145470 34540
rect 145375 34371 145470 34413
rect 145375 34370 145418 34371
rect 145375 34275 145470 34370
rect 132617 33810 145290 33839
rect 132617 33765 145245 33810
rect 145375 33783 145427 34275
rect 145526 34219 147532 34734
rect 132617 32852 145240 33765
rect 145346 33754 145427 33783
rect 145301 33747 145346 33754
rect 145375 33747 145427 33754
rect 145301 33733 145427 33747
rect 145301 33709 145346 33733
rect 145375 33709 145427 33733
rect 145296 33704 145301 33709
rect 145348 33704 145375 33709
rect 145296 33682 145375 33704
rect 132617 32688 145114 32852
rect 145296 32796 145348 33682
rect 145483 33653 147532 34219
rect 145431 33626 147532 33653
rect 145170 32744 145348 32796
rect 145404 32688 147532 33626
rect 132617 158 147532 32688
rect 186417 0 202358 41657
rect 241260 39593 245381 39600
rect 245493 39593 252015 39600
rect 252101 39593 256100 39600
rect 238961 31928 241151 32702
rect 241200 31683 256100 39593
rect 256252 39545 256280 46854
rect 297088 44338 297140 44402
rect 295248 44270 295300 44334
rect 295260 42193 295288 44270
rect 297100 42193 297128 44338
rect 297744 42193 297772 46854
rect 299572 44338 299624 44402
rect 305736 44338 305788 44402
rect 299584 42193 299612 44338
rect 303252 44270 303304 44334
rect 303264 42193 303292 44270
rect 304540 44134 304592 44198
rect 304552 42193 304580 44134
rect 305748 42193 305776 44338
rect 309428 42193 309456 46854
rect 349988 44406 350040 44470
rect 350000 44198 350028 44406
rect 351920 44270 351972 44334
rect 349988 44134 350040 44198
rect 350080 44134 350132 44198
rect 350092 42193 350120 44134
rect 351932 42193 351960 44270
rect 352576 42193 352604 46854
rect 359372 44406 359424 44470
rect 354404 44270 354456 44334
rect 354416 42193 354444 44270
rect 358084 44134 358136 44198
rect 358096 42193 358124 44134
rect 359384 42193 359412 44406
rect 360568 44270 360620 44334
rect 360580 44198 360608 44270
rect 360568 44134 360620 44198
rect 360580 42193 360608 44134
rect 364260 42193 364288 46854
rect 404910 44231 404966 44305
rect 404924 42193 404952 44231
rect 406752 44202 406804 44266
rect 406764 42193 406792 44202
rect 407408 42193 407436 46854
rect 414204 44406 414256 44470
rect 412914 44231 412970 44305
rect 412928 42193 412956 44231
rect 414216 44198 414244 44406
rect 414204 44134 414256 44198
rect 414216 42193 414244 44134
rect 419092 42193 419120 46854
rect 459650 44231 459706 44305
rect 459664 42193 459692 44231
rect 461492 44202 461544 44266
rect 461504 42193 461532 44202
rect 462148 42193 462176 46854
rect 468944 44338 468996 44402
rect 467654 44231 467710 44305
rect 467668 42193 467696 44231
rect 468956 44198 468984 44338
rect 468944 44134 468996 44198
rect 468956 42193 468984 44134
rect 473832 42193 473860 46854
rect 514482 44231 514538 44305
rect 514496 42193 514524 44231
rect 516324 44202 516376 44266
rect 516336 42193 516364 44202
rect 516980 42193 517008 46854
rect 523776 45562 523828 45626
rect 518716 45494 518768 45558
rect 518728 44266 518756 45494
rect 522486 44367 522542 44441
rect 523788 44402 523816 45562
rect 518716 44202 518768 44266
rect 522500 42193 522528 44367
rect 523776 44338 523828 44402
rect 523788 42193 523816 44338
rect 673472 42770 673500 111522
rect 673564 108458 673592 152798
rect 673656 149054 673684 189246
rect 675887 195399 717600 195875
rect 675407 195329 675887 195343
rect 675312 195301 675887 195329
rect 675312 187325 675340 195301
rect 675407 195287 675887 195301
rect 675943 195231 717600 195399
rect 675887 194755 717600 195231
rect 675943 194587 717600 194755
rect 675887 194203 717600 194587
rect 675943 194035 717600 194203
rect 675887 193559 717600 194035
rect 675943 193391 717600 193559
rect 675887 192915 717600 193391
rect 675943 192747 717600 192915
rect 675887 192363 717600 192747
rect 675407 192251 675887 192307
rect 675943 192195 717600 192363
rect 675887 191719 717600 192195
rect 675943 191551 717600 191719
rect 675887 191075 717600 191551
rect 675407 190963 675887 191019
rect 675943 190907 717600 191075
rect 675887 190523 717600 190907
rect 675407 190411 675887 190467
rect 675943 190355 717600 190523
rect 675887 189879 717600 190355
rect 675943 189711 717600 189879
rect 675392 189246 675444 189310
rect 675404 189179 675432 189246
rect 675887 189235 717600 189711
rect 675404 189151 675887 189179
rect 675407 189123 675887 189151
rect 675943 189067 717600 189235
rect 675887 188683 717600 189067
rect 675407 188571 675887 188627
rect 675943 188515 717600 188683
rect 675887 188039 717600 188515
rect 675943 187871 717600 188039
rect 675887 187395 717600 187871
rect 675407 187325 675887 187339
rect 675312 187297 675887 187325
rect 675407 187283 675887 187297
rect 675943 187227 717600 187395
rect 675887 187017 717600 187227
rect 675887 158559 717600 158758
rect 675943 158391 717600 158559
rect 675887 158007 717600 158391
rect 675943 157839 717600 158007
rect 675887 157363 717600 157839
rect 675943 157195 717600 157363
rect 675887 156719 717600 157195
rect 675943 156551 717600 156719
rect 673920 155926 673972 155990
rect 673656 149026 673776 149054
rect 673748 144566 673776 149026
rect 673736 144502 673788 144566
rect 673552 108394 673604 108458
rect 673564 45626 673592 108394
rect 673748 100609 673776 144502
rect 673932 111586 673960 155926
rect 675887 156167 717600 156551
rect 675943 155999 717600 156167
rect 675392 155926 675444 155990
rect 675404 155467 675432 155926
rect 675887 155523 717600 155999
rect 675404 155439 675887 155467
rect 675407 155411 675887 155439
rect 675943 155355 717600 155523
rect 675887 154879 717600 155355
rect 675943 154711 717600 154879
rect 675887 154327 717600 154711
rect 675943 154159 717600 154327
rect 675887 153683 717600 154159
rect 675943 153515 717600 153683
rect 675887 153039 717600 153515
rect 675943 152871 717600 153039
rect 675392 152798 675444 152862
rect 675404 152431 675432 152798
rect 675887 152487 717600 152871
rect 675404 152388 675887 152431
rect 675407 152375 675887 152388
rect 675943 152319 717600 152487
rect 675887 151843 717600 152319
rect 675943 151675 717600 151843
rect 675887 151199 717600 151675
rect 675407 151129 675887 151143
rect 675312 151101 675887 151129
rect 675312 143125 675340 151101
rect 675407 151087 675887 151101
rect 675943 151031 717600 151199
rect 675887 150555 717600 151031
rect 675943 150387 717600 150555
rect 675887 150003 717600 150387
rect 675943 149835 717600 150003
rect 675887 149359 717600 149835
rect 675943 149191 717600 149359
rect 675887 148715 717600 149191
rect 675943 148547 717600 148715
rect 675887 148163 717600 148547
rect 675407 148051 675887 148107
rect 675943 147995 717600 148163
rect 675887 147519 717600 147995
rect 675943 147351 717600 147519
rect 675887 146875 717600 147351
rect 675407 146763 675887 146819
rect 675943 146707 717600 146875
rect 675887 146323 717600 146707
rect 675407 146211 675887 146267
rect 675943 146155 717600 146323
rect 675887 145679 717600 146155
rect 675943 145511 717600 145679
rect 675887 145035 717600 145511
rect 675407 144951 675887 144979
rect 675404 144923 675887 144951
rect 675404 144566 675432 144923
rect 675943 144867 717600 145035
rect 675392 144502 675444 144566
rect 675887 144483 717600 144867
rect 675407 144371 675887 144427
rect 675943 144315 717600 144483
rect 675887 143839 717600 144315
rect 675943 143671 717600 143839
rect 675887 143195 717600 143671
rect 675407 143125 675887 143139
rect 675312 143097 675887 143125
rect 675407 143083 675887 143097
rect 675943 143027 717600 143195
rect 675887 142817 717600 143027
rect 675887 114159 717600 114358
rect 675943 113991 717600 114159
rect 675887 113607 717600 113991
rect 675943 113439 717600 113607
rect 675887 112963 717600 113439
rect 675943 112795 717600 112963
rect 675887 112319 717600 112795
rect 675943 112151 717600 112319
rect 675887 111767 717600 112151
rect 673920 111522 673972 111586
rect 675943 111599 717600 111767
rect 675392 111522 675444 111586
rect 675404 111067 675432 111522
rect 675887 111123 717600 111599
rect 675404 111044 675887 111067
rect 675407 111011 675887 111044
rect 675943 110955 717600 111123
rect 675887 110479 717600 110955
rect 675943 110311 717600 110479
rect 675887 109927 717600 110311
rect 675943 109759 717600 109927
rect 675887 109283 717600 109759
rect 675943 109115 717600 109283
rect 675887 108639 717600 109115
rect 675943 108471 717600 108639
rect 675392 108394 675444 108458
rect 675404 108031 675432 108394
rect 675887 108087 717600 108471
rect 675404 108003 675887 108031
rect 675407 107975 675887 108003
rect 675943 107919 717600 108087
rect 675887 107443 717600 107919
rect 675943 107275 717600 107443
rect 675312 106814 675432 106842
rect 673734 100535 673790 100609
rect 673552 45562 673604 45626
rect 673748 45558 673776 100535
rect 675312 98725 675340 106814
rect 675404 106743 675432 106814
rect 675887 106799 717600 107275
rect 675404 106692 675887 106743
rect 675407 106687 675887 106692
rect 675943 106631 717600 106799
rect 675887 106155 717600 106631
rect 675943 105987 717600 106155
rect 675887 105603 717600 105987
rect 675943 105435 717600 105603
rect 675887 104959 717600 105435
rect 675943 104791 717600 104959
rect 675887 104315 717600 104791
rect 675943 104147 717600 104315
rect 675887 103763 717600 104147
rect 675407 103651 675887 103707
rect 675943 103595 717600 103763
rect 675887 103119 717600 103595
rect 675943 102951 717600 103119
rect 675887 102475 717600 102951
rect 675407 102363 675887 102419
rect 675943 102307 717600 102475
rect 675887 101923 717600 102307
rect 675407 101811 675887 101867
rect 675943 101755 717600 101923
rect 675887 101279 717600 101755
rect 675943 101111 717600 101279
rect 675887 100635 717600 101111
rect 675390 100579 675446 100609
rect 675390 100535 675887 100579
rect 675407 100523 675887 100535
rect 675943 100467 717600 100635
rect 675887 100083 717600 100467
rect 675407 99971 675887 100027
rect 675943 99915 717600 100083
rect 675887 99439 717600 99915
rect 675943 99271 717600 99439
rect 675887 98795 717600 99271
rect 675407 98725 675887 98739
rect 675312 98697 675887 98725
rect 675407 98683 675887 98697
rect 675943 98627 717600 98795
rect 675887 98417 717600 98627
rect 673736 45494 673788 45558
rect 579896 42706 579948 42770
rect 673460 42706 673512 42770
rect 295260 41806 295339 42193
rect 295283 41713 295339 41806
rect 295927 41713 295983 42193
rect 296571 41713 296627 42193
rect 297100 41806 297179 42193
rect 297744 41834 297823 42193
rect 297916 41890 297968 41954
rect 297928 41834 297956 41890
rect 297744 41806 297956 41834
rect 297123 41713 297179 41806
rect 297767 41713 297823 41806
rect 298411 41713 298467 42193
rect 298963 41713 299019 42193
rect 299584 41806 299663 42193
rect 299607 41713 299663 41806
rect 300251 41713 300307 42193
rect 300676 41890 300728 41954
rect 300688 41834 300716 41890
rect 300803 41834 300859 42193
rect 301447 41834 301503 42193
rect 302091 41834 302147 42193
rect 302240 41890 302292 41954
rect 302252 41834 302280 41890
rect 300688 41806 302280 41834
rect 300803 41713 300859 41806
rect 301447 41713 301503 41806
rect 302091 41713 302147 41806
rect 303264 41806 303343 42193
rect 304552 41806 304631 42193
rect 303287 41713 303343 41806
rect 304575 41713 304631 41806
rect 305127 41834 305183 42193
rect 305276 41890 305328 41954
rect 305288 41834 305316 41890
rect 305127 41806 305316 41834
rect 305748 41806 305827 42193
rect 305127 41713 305183 41806
rect 305771 41713 305827 41806
rect 306415 41834 306471 42193
rect 306564 41890 306616 41954
rect 306576 41834 306604 41890
rect 306415 41806 306604 41834
rect 306415 41713 306471 41806
rect 307611 41834 307667 42193
rect 307611 41818 307800 41834
rect 307611 41806 307812 41818
rect 308680 41890 308732 41954
rect 308692 41834 308720 41890
rect 308807 41834 308863 42193
rect 309428 41834 309507 42193
rect 308692 41806 309507 41834
rect 307611 41713 307667 41806
rect 307760 41754 307812 41806
rect 308807 41713 308863 41806
rect 309451 41713 309507 41806
rect 310647 41713 310703 42193
rect 350083 41713 350139 42193
rect 350727 41713 350783 42193
rect 351371 41713 351427 42193
rect 351923 41713 351979 42193
rect 352567 41970 352623 42193
rect 352567 41954 352696 41970
rect 352567 41942 352708 41954
rect 352567 41713 352623 41942
rect 352656 41890 352708 41942
rect 353211 41713 353267 42193
rect 353763 41713 353819 42193
rect 354407 41713 354463 42193
rect 355051 41713 355107 42193
rect 355508 41890 355560 41954
rect 355520 41834 355548 41890
rect 355603 41834 355659 42193
rect 356247 41834 356303 42193
rect 356891 41834 356947 42193
rect 356980 41890 357032 41954
rect 356992 41834 357020 41890
rect 355520 41806 357020 41834
rect 355603 41713 355659 41806
rect 356247 41713 356303 41806
rect 356891 41713 356947 41806
rect 358087 41713 358143 42193
rect 359375 41713 359431 42193
rect 359832 41890 359884 41954
rect 359844 41834 359872 41890
rect 359927 41834 359983 42193
rect 359844 41806 359983 41834
rect 359927 41713 359983 41806
rect 360571 41713 360627 42193
rect 361120 41890 361172 41954
rect 361132 41834 361160 41890
rect 361215 41834 361271 42193
rect 361132 41806 361271 41834
rect 361215 41713 361271 41806
rect 362411 41834 362467 42193
rect 362411 41818 362540 41834
rect 362411 41806 362552 41818
rect 362411 41713 362467 41806
rect 362500 41754 362552 41806
rect 363512 41890 363564 41954
rect 363524 41834 363552 41890
rect 363607 41834 363663 42193
rect 364251 41834 364307 42193
rect 363524 41806 364307 41834
rect 363607 41713 363663 41806
rect 364251 41713 364307 41806
rect 365447 41713 365503 42193
rect 404883 41820 404952 42193
rect 404883 41713 404939 41820
rect 406171 41713 406227 42193
rect 406723 41820 406792 42193
rect 407367 41970 407436 42193
rect 407367 41954 407528 41970
rect 407367 41942 407540 41954
rect 407367 41820 407436 41942
rect 407488 41890 407540 41942
rect 406723 41713 406779 41820
rect 407367 41713 407423 41820
rect 408011 41713 408067 42193
rect 408563 41713 408619 42193
rect 409851 41713 409907 42193
rect 410248 41890 410300 41954
rect 410260 41834 410288 41890
rect 410403 41834 410459 42193
rect 410260 41806 410459 41834
rect 410403 41713 410459 41806
rect 411536 41890 411588 41954
rect 411548 41834 411576 41890
rect 411691 41834 411747 42193
rect 411548 41806 411747 41834
rect 411691 41713 411747 41806
rect 412887 41820 412956 42193
rect 414175 41820 414244 42193
rect 414572 41890 414624 41954
rect 414584 41834 414612 41890
rect 414727 41834 414783 42193
rect 415860 41890 415912 41954
rect 412887 41713 412943 41820
rect 414175 41713 414231 41820
rect 414584 41806 414783 41834
rect 414727 41713 414783 41806
rect 415872 41834 415900 41890
rect 416015 41834 416071 42193
rect 415872 41806 416071 41834
rect 416015 41713 416071 41806
rect 417211 41834 417267 42193
rect 417211 41818 417372 41834
rect 418252 41890 418304 41954
rect 418264 41834 418292 41890
rect 418407 41834 418463 42193
rect 419051 41834 419120 42193
rect 418264 41820 419120 41834
rect 417211 41806 417384 41818
rect 417211 41713 417267 41806
rect 417332 41754 417384 41806
rect 418264 41806 419107 41820
rect 418407 41713 418463 41806
rect 419051 41713 419107 41806
rect 420247 41713 420303 42193
rect 459664 41806 459739 42193
rect 459683 41713 459739 41806
rect 460971 41713 461027 42193
rect 461504 41806 461579 42193
rect 462148 41834 462223 42193
rect 462320 41890 462372 41954
rect 462332 41834 462360 41890
rect 462148 41806 462360 41834
rect 461523 41713 461579 41806
rect 462167 41713 462223 41806
rect 462811 41713 462867 42193
rect 463363 41713 463419 42193
rect 464651 41713 464707 42193
rect 465080 41890 465132 41954
rect 465092 41834 465120 41890
rect 465203 41834 465259 42193
rect 465092 41806 465259 41834
rect 466368 41890 466420 41954
rect 466380 41834 466408 41890
rect 466491 41834 466547 42193
rect 466380 41806 466547 41834
rect 465203 41713 465259 41806
rect 466491 41713 466547 41806
rect 467668 41806 467743 42193
rect 468956 41806 469031 42193
rect 469404 41890 469456 41954
rect 469416 41834 469444 41890
rect 469527 41834 469583 42193
rect 470692 41890 470744 41954
rect 469416 41806 469583 41834
rect 467687 41713 467743 41806
rect 468975 41713 469031 41806
rect 469527 41713 469583 41806
rect 470704 41834 470732 41890
rect 470815 41834 470871 42193
rect 470704 41806 470871 41834
rect 470815 41713 470871 41806
rect 472011 41834 472067 42193
rect 472011 41818 472204 41834
rect 472011 41806 472216 41818
rect 473084 41890 473136 41954
rect 473096 41834 473124 41890
rect 473207 41834 473263 42193
rect 473832 41834 473907 42193
rect 473096 41806 473907 41834
rect 472011 41713 472067 41806
rect 472164 41754 472216 41806
rect 473207 41713 473263 41806
rect 473851 41713 473907 41806
rect 475047 41713 475103 42193
rect 514483 41713 514539 42193
rect 515771 41713 515827 42193
rect 516323 41713 516379 42193
rect 516967 41970 517023 42193
rect 516967 41954 517100 41970
rect 516967 41942 517112 41954
rect 516967 41713 517023 41942
rect 517060 41890 517112 41942
rect 517611 41713 517667 42193
rect 518163 41713 518219 42193
rect 519451 41713 519507 42193
rect 519912 41890 519964 41954
rect 519924 41834 519952 41890
rect 520003 41834 520059 42193
rect 519924 41806 520059 41834
rect 520003 41713 520059 41806
rect 521200 41890 521252 41954
rect 521212 41834 521240 41890
rect 521291 41834 521347 42193
rect 521212 41806 521347 41834
rect 521291 41713 521347 41806
rect 522487 41713 522543 42193
rect 523775 41713 523831 42193
rect 524236 41890 524288 41954
rect 524248 41834 524276 41890
rect 524327 41834 524383 42193
rect 524248 41806 524383 41834
rect 524327 41713 524383 41806
rect 525524 41890 525576 41954
rect 525536 41834 525564 41890
rect 525615 41834 525671 42193
rect 525536 41806 525671 41834
rect 525615 41713 525671 41806
rect 526811 41834 526867 42193
rect 526732 41818 526867 41834
rect 526720 41806 526867 41818
rect 526720 41754 526772 41806
rect 526811 41713 526867 41806
rect 527916 41890 527968 41954
rect 527928 41834 527956 41890
rect 528007 41834 528063 42193
rect 528651 41834 528707 42193
rect 527928 41806 528707 41834
rect 528007 41713 528063 41806
rect 528651 41713 528707 41806
rect 529847 41713 529903 42193
rect 579908 41886 579936 42706
rect 568856 41822 568908 41886
rect 579896 41822 579948 41886
rect 295017 41657 295227 41713
rect 295395 41657 295871 41713
rect 296039 41657 296515 41713
rect 296683 41657 297067 41713
rect 297235 41657 297711 41713
rect 297879 41657 298355 41713
rect 298523 41657 298907 41713
rect 299075 41657 299551 41713
rect 299719 41657 300195 41713
rect 300363 41657 300747 41713
rect 300915 41657 301391 41713
rect 301559 41657 302035 41713
rect 302203 41657 302587 41713
rect 302755 41657 303231 41713
rect 303399 41657 303875 41713
rect 304043 41657 304519 41713
rect 304687 41657 305071 41713
rect 305239 41657 305715 41713
rect 305883 41657 306359 41713
rect 306527 41657 306911 41713
rect 307079 41657 307555 41713
rect 307723 41657 308199 41713
rect 308367 41657 308751 41713
rect 308919 41657 309395 41713
rect 309563 41657 310039 41713
rect 310207 41657 310591 41713
rect 310759 41657 310958 41713
rect 256238 39471 256294 39545
rect 238972 30753 256100 31683
rect 241200 714 256100 30753
rect 295017 0 310958 41657
rect 349817 41657 350027 41713
rect 350195 41657 350671 41713
rect 350839 41657 351315 41713
rect 351483 41657 351867 41713
rect 352035 41657 352511 41713
rect 352679 41657 353155 41713
rect 353323 41657 353707 41713
rect 353875 41657 354351 41713
rect 354519 41657 354995 41713
rect 355163 41657 355547 41713
rect 355715 41657 356191 41713
rect 356359 41657 356835 41713
rect 357003 41657 357387 41713
rect 357555 41657 358031 41713
rect 358199 41657 358675 41713
rect 358843 41657 359319 41713
rect 359487 41657 359871 41713
rect 360039 41657 360515 41713
rect 360683 41657 361159 41713
rect 361327 41657 361711 41713
rect 361879 41657 362355 41713
rect 362523 41657 362999 41713
rect 363167 41657 363551 41713
rect 363719 41657 364195 41713
rect 364363 41657 364839 41713
rect 365007 41657 365391 41713
rect 365559 41657 365758 41713
rect 349817 0 365758 41657
rect 404617 41657 404827 41713
rect 404995 41657 405471 41713
rect 405639 41657 406115 41713
rect 406283 41657 406667 41713
rect 406835 41657 407311 41713
rect 407479 41657 407955 41713
rect 408123 41657 408507 41713
rect 408675 41657 409151 41713
rect 409319 41657 409795 41713
rect 409963 41657 410347 41713
rect 410515 41657 410991 41713
rect 411159 41657 411635 41713
rect 411803 41657 412187 41713
rect 412355 41657 412831 41713
rect 412999 41657 413475 41713
rect 413643 41657 414119 41713
rect 414287 41657 414671 41713
rect 414839 41657 415315 41713
rect 415483 41657 415959 41713
rect 416127 41657 416511 41713
rect 416679 41657 417155 41713
rect 417323 41657 417799 41713
rect 417967 41657 418351 41713
rect 418519 41657 418995 41713
rect 419163 41657 419639 41713
rect 419807 41657 420191 41713
rect 420359 41657 420558 41713
rect 404617 0 420558 41657
rect 459417 41657 459627 41713
rect 459795 41657 460271 41713
rect 460439 41657 460915 41713
rect 461083 41657 461467 41713
rect 461635 41657 462111 41713
rect 462279 41657 462755 41713
rect 462923 41657 463307 41713
rect 463475 41657 463951 41713
rect 464119 41657 464595 41713
rect 464763 41657 465147 41713
rect 465315 41657 465791 41713
rect 465959 41657 466435 41713
rect 466603 41657 466987 41713
rect 467155 41657 467631 41713
rect 467799 41657 468275 41713
rect 468443 41657 468919 41713
rect 469087 41657 469471 41713
rect 469639 41657 470115 41713
rect 470283 41657 470759 41713
rect 470927 41657 471311 41713
rect 471479 41657 471955 41713
rect 472123 41657 472599 41713
rect 472767 41657 473151 41713
rect 473319 41657 473795 41713
rect 473963 41657 474439 41713
rect 474607 41657 474991 41713
rect 475159 41657 475358 41713
rect 459417 0 475358 41657
rect 514217 41657 514427 41713
rect 514595 41657 515071 41713
rect 515239 41657 515715 41713
rect 515883 41657 516267 41713
rect 516435 41657 516911 41713
rect 517079 41657 517555 41713
rect 517723 41657 518107 41713
rect 518275 41657 518751 41713
rect 518919 41657 519395 41713
rect 519563 41657 519947 41713
rect 520115 41657 520591 41713
rect 520759 41657 521235 41713
rect 521403 41657 521787 41713
rect 521955 41657 522431 41713
rect 522599 41657 523075 41713
rect 523243 41657 523719 41713
rect 523887 41657 524271 41713
rect 524439 41657 524915 41713
rect 525083 41657 525559 41713
rect 525727 41657 526111 41713
rect 526279 41657 526755 41713
rect 526923 41657 527399 41713
rect 527567 41657 527951 41713
rect 528119 41657 528595 41713
rect 528763 41657 529239 41713
rect 529407 41657 529791 41713
rect 529959 41657 530158 41713
rect 514217 0 530158 41657
rect 568868 39681 568896 41822
rect 568854 39607 568910 39681
rect 569142 39593 573922 40000
rect 578421 39616 578821 40000
rect 579121 39593 583901 40000
rect 622942 39593 627722 40000
rect 632221 39616 632621 40000
rect 632921 39593 637701 40000
rect 569142 985 583947 39593
rect 622942 985 637747 39593
<< metal3 >>
rect 79944 997600 84944 1014070
rect 127944 997600 132944 1014070
rect 175944 997600 180944 1014070
rect 239478 997600 253800 1000737
rect 290878 997600 305200 1000737
rect 429744 997600 434744 1014070
rect 479144 997600 484144 1014070
rect 530744 997600 535744 1014070
rect 631944 997600 636944 1014070
rect 23530 960144 40000 965144
rect 677600 934600 680737 948922
rect 678000 461700 685920 466500
rect 31680 441300 39600 446100
rect 411069 44434 411135 44437
rect 465809 44434 465875 44437
rect 474457 44434 474523 44437
rect 411069 44432 419550 44434
rect 411069 44376 411074 44432
rect 411130 44376 419550 44432
rect 411069 44374 419550 44376
rect 411069 44371 411135 44374
rect 419490 44298 419550 44374
rect 465809 44432 474523 44434
rect 465809 44376 465814 44432
rect 465870 44376 474462 44432
rect 474518 44376 474523 44432
rect 465809 44374 474523 44376
rect 465809 44371 465875 44374
rect 474457 44371 474523 44374
rect 419717 44298 419783 44301
rect 419490 44296 419783 44298
rect 419490 44240 419722 44296
rect 419778 44240 419783 44296
rect 419490 44238 419783 44240
rect 419717 44235 419783 44238
rect 518801 44298 518867 44301
rect 524965 44298 525031 44301
rect 518801 44296 525031 44298
rect 518801 44240 518806 44296
rect 518862 44240 524970 44296
rect 525026 44240 525031 44296
rect 518801 44238 525031 44240
rect 518801 44235 518867 44238
rect 524965 44235 525031 44238
rect 141667 38031 141813 40000
rect 141667 37971 141873 38031
rect 141667 37911 141820 37971
rect 141873 37911 141966 37971
rect 141667 37818 141966 37911
rect 141820 37046 141966 37818
<< obsm3 >>
rect 75091 1014150 89850 1032263
rect 75091 1000581 79864 1014150
rect 85024 1000581 89850 1014150
rect 123091 1014150 137850 1032263
rect 123091 1000581 127864 1014150
rect 133024 1000581 137850 1014150
rect 171091 1014150 185850 1032263
rect 171091 1000581 175864 1014150
rect 181024 1000581 185850 1014150
rect 220000 1000817 253800 1037600
rect 271400 1000817 305200 1037600
rect 339448 1002850 354258 1037600
rect 424891 1014150 439650 1032263
rect 220000 997600 234279 1000737
rect 234359 999946 239398 1000817
rect 234359 998225 236898 999946
rect 234359 998145 234499 998225
rect 236859 998145 236898 998225
rect 234579 997600 236779 998145
rect 236978 997600 239178 999866
rect 239258 998145 239398 999946
rect 271400 997600 285679 1000737
rect 285759 999946 290798 1000817
rect 285759 998225 288298 999946
rect 285759 998145 285899 998225
rect 288259 998145 288298 998225
rect 285979 997600 288179 998145
rect 288378 997600 290578 999866
rect 290658 998145 290798 999946
rect 339499 997600 344279 1002770
rect 344359 998007 349398 1002850
rect 344579 997600 346779 998007
rect 346978 997600 349178 998007
rect 349478 997600 354258 1002770
rect 424891 1000581 429664 1014150
rect 434824 1000581 439650 1014150
rect 474291 1014150 489050 1032263
rect 474291 1000581 479064 1014150
rect 484224 1000581 489050 1014150
rect 525891 1014150 540650 1032263
rect 525891 1000581 530664 1014150
rect 535824 1000581 540650 1014150
rect 575648 1005032 590458 1036620
rect 627091 1014150 641850 1032263
rect 575648 1004183 585598 1005032
rect 575699 997600 580479 1004103
rect 580559 998007 585598 1004183
rect 580779 997600 582979 998007
rect 583178 997600 585378 998007
rect 585678 997600 590458 1004952
rect 627091 1000581 631864 1014150
rect 637024 1000581 641850 1014150
rect 339542 997117 339602 997600
rect 585734 997525 585794 997600
rect 585734 997462 585843 997525
rect 585777 997459 585843 997462
rect 339493 997054 339602 997117
rect 339493 997051 339559 997054
rect 5337 965224 37019 970050
rect 5337 960064 23450 965224
rect 5337 955291 37019 960064
rect 677600 954121 680737 968400
rect 680817 954041 717600 968400
rect 678145 953901 717600 954041
rect 677600 951621 678145 953821
rect 678225 951541 717600 953901
rect 678145 951502 717600 951541
rect 677600 949222 679866 951422
rect 679946 949142 717600 951502
rect 678145 949002 717600 949142
rect 680817 934600 717600 949002
rect 7 928240 4850 930187
rect 30753 928121 31683 930228
rect 33910 928240 34840 930187
rect 7 923071 38140 928000
rect 38220 923151 39600 927940
rect 7 922851 39593 923071
rect 7 920676 39600 922851
rect 7 920376 39593 920676
rect 7 918200 39600 920376
rect 7 917980 39593 918200
rect 7 913020 38140 917980
rect 38220 913100 39600 917900
rect 7 913000 39593 913020
rect 30760 910805 31690 912821
rect 685910 906579 686840 908595
rect 678007 906380 717593 906400
rect 678000 901500 679380 906300
rect 679460 901420 717593 906380
rect 678007 901200 717593 901420
rect 678000 899024 717593 901200
rect 678007 898724 717593 899024
rect 678000 896549 717593 898724
rect 678007 896329 717593 896549
rect 678000 891460 679380 896249
rect 679460 891400 717593 896329
rect 682760 889213 683690 891160
rect 685917 889172 686847 891279
rect 712750 889213 717593 891160
rect 44173 885866 44239 885869
rect 44817 885866 44883 885869
rect 44173 885806 44883 885866
rect 44173 885803 44239 885806
rect 44817 885803 44883 885806
rect 0 880798 35960 885658
rect 36040 880878 40000 885658
rect 0 880578 39593 880798
rect 0 878378 40000 880578
rect 0 878179 39593 878378
rect 0 875979 40000 878179
rect 0 875759 39593 875979
rect 0 870848 35960 875759
rect 36040 871042 40000 875679
rect 44173 871042 44239 871045
rect 36040 870982 44239 871042
rect 36040 870899 40000 870982
rect 44173 870979 44239 870982
rect 677338 847086 717600 862938
rect 980 838398 32568 843258
rect 32648 838478 40000 843258
rect 980 838178 39593 838398
rect 980 835978 40000 838178
rect 980 835779 39593 835978
rect 980 833579 40000 835779
rect 980 833359 39593 833579
rect 980 828448 33417 833359
rect 33497 828499 40000 833279
rect 677600 813921 680592 818701
rect 680672 813841 717600 818752
rect 678007 813621 717600 813841
rect 677600 811421 717600 813621
rect 678007 811222 717600 811421
rect 677600 809022 717600 811222
rect 678007 808802 717600 809022
rect 677600 803942 680592 808722
rect 680672 803942 717600 808802
rect 677593 803858 677659 803861
rect 677734 803858 677794 803942
rect 677593 803798 677794 803858
rect 677593 803795 677659 803798
rect 0 785262 40262 801114
rect 677338 759686 717600 775538
rect 0 742062 40262 757914
rect 677338 715286 717600 731138
rect 0 698862 40262 714714
rect 0 655462 40262 671314
rect 677338 671086 717600 686938
rect 0 612262 40262 628114
rect 677338 626886 717600 642738
rect 0 569062 40262 584914
rect 677338 582486 717600 598338
rect 0 525862 40262 541714
rect 677338 538286 717600 554138
rect 677600 505121 680592 509901
rect 680672 505041 717600 509952
rect 678007 504821 717600 505041
rect 677600 502621 717600 504821
rect 678007 502422 717600 502621
rect 677600 500222 717600 502422
rect 678007 500002 717600 500222
rect 0 493398 36928 498258
rect 37008 493478 40000 498258
rect 677600 495142 680592 499922
rect 680672 495142 717600 500002
rect 677918 494869 677978 495142
rect 677918 494806 678027 494869
rect 677961 494803 678027 494806
rect 0 493178 39593 493398
rect 0 490978 40000 493178
rect 0 490779 39593 490978
rect 0 488579 40000 490779
rect 0 488359 39593 488579
rect 0 483448 36928 488359
rect 37008 483499 40000 488279
rect 685910 466779 686840 468795
rect 678007 466580 717593 466600
rect 686000 461620 717593 466580
rect 678007 461400 717593 461620
rect 678000 459224 717593 461400
rect 678007 458924 717593 459224
rect 7 456440 4850 458387
rect 30753 456321 31683 458428
rect 33910 456440 34840 458387
rect 678000 456749 717593 458924
rect 678007 456529 717593 456749
rect 7 451271 31600 456200
rect 31680 451351 39600 456140
rect 678000 451660 685920 456449
rect 686000 451600 717593 456529
rect 7 451051 39593 451271
rect 7 448876 39600 451051
rect 682760 449413 683690 451360
rect 685917 449372 686847 451479
rect 712750 449413 717593 451360
rect 7 448576 39593 448876
rect 7 446400 39600 448576
rect 7 446180 39593 446400
rect 7 441220 31600 446180
rect 7 441200 39593 441220
rect 30760 439005 31690 441021
rect 673862 419930 673938 419932
rect 674005 419930 674071 419933
rect 673862 419870 674071 419930
rect 673862 419868 673938 419870
rect 674005 419867 674071 419870
rect 673862 419250 673938 419252
rect 674005 419250 674071 419253
rect 673862 419190 674071 419250
rect 673862 419188 673938 419190
rect 674005 419187 674071 419190
rect 677600 418521 684103 423301
rect 677501 418434 677567 418437
rect 677734 418434 677794 418521
rect 684183 418441 716620 423352
rect 677501 418374 677794 418434
rect 677501 418371 677567 418374
rect 678007 418221 716620 418441
rect 677600 416021 716620 418221
rect 678007 415822 716620 416021
rect 0 398062 40262 413914
rect 677600 413622 716620 415822
rect 678007 413402 716620 413622
rect 677600 408542 684952 413322
rect 685032 408542 716620 413402
rect 0 354862 40262 370714
rect 677338 364086 717600 379938
rect 0 311462 40262 327314
rect 677338 319886 717600 335738
rect 0 268262 40262 284114
rect 677338 275686 717600 291538
rect 0 225062 40262 240914
rect 677338 231286 717600 247138
rect 0 181862 40262 197714
rect 677338 187086 717600 202938
rect 677338 142886 717600 158738
rect 0 120198 35960 125058
rect 36040 120278 40000 125058
rect 0 119978 39593 120198
rect 0 117778 40000 119978
rect 0 117579 39593 117778
rect 0 115379 40000 117579
rect 0 115159 39593 115379
rect 0 110248 35960 115159
rect 36040 110530 40000 115079
rect 44173 110530 44239 110533
rect 44817 110530 44883 110533
rect 36040 110470 44883 110530
rect 36040 110299 40000 110470
rect 44173 110467 44239 110470
rect 44817 110467 44883 110470
rect 673729 100602 673795 100605
rect 675385 100602 675451 100605
rect 673729 100542 675451 100602
rect 673729 100539 673795 100542
rect 675385 100539 675451 100542
rect 677338 98486 717600 114338
rect 30753 83121 31683 85228
rect 31961 83088 32654 85228
rect 879 78071 38140 83000
rect 38220 78298 39600 82940
rect 39665 80202 39731 80205
rect 44173 80202 44239 80205
rect 44817 80202 44883 80205
rect 39665 80142 44883 80202
rect 39665 80139 39731 80142
rect 44173 80139 44239 80142
rect 44817 80139 44883 80142
rect 39665 78298 39731 78301
rect 38220 78238 39731 78298
rect 38220 78151 39600 78238
rect 39665 78235 39731 78238
rect 879 77851 39593 78071
rect 879 75676 39600 77851
rect 879 75376 39593 75676
rect 879 73200 39600 75376
rect 879 72980 39593 73200
rect 879 68098 38140 72980
rect 38220 68100 39600 72900
rect 151721 46882 151787 46885
rect 188521 46882 188587 46885
rect 151721 46822 188587 46882
rect 151721 46819 151787 46822
rect 188521 46819 188587 46822
rect 522481 44434 522547 44437
rect 404905 44298 404971 44301
rect 412909 44298 412975 44301
rect 404905 44238 412975 44298
rect 516090 44374 522547 44434
rect 404905 44235 404971 44238
rect 412909 44235 412975 44238
rect 459645 44298 459711 44301
rect 467649 44298 467715 44301
rect 459645 44238 467715 44298
rect 459645 44235 459711 44238
rect 467649 44235 467715 44238
rect 514477 44298 514543 44301
rect 516090 44298 516150 44374
rect 522481 44371 522547 44374
rect 514477 44238 516150 44298
rect 514477 44235 514543 44238
rect 143533 40490 143599 40493
rect 151721 40490 151787 40493
rect 143533 40430 151787 40490
rect 143533 40427 143599 40430
rect 145790 40354 145850 40430
rect 151721 40427 151787 40430
rect 145790 40294 145898 40354
rect 93761 40218 93827 40221
rect 135161 40218 135227 40221
rect 91142 40158 93827 40218
rect 91142 40000 91202 40158
rect 93761 40155 93827 40158
rect 133094 40158 135227 40218
rect 133094 40000 133154 40158
rect 135161 40155 135227 40158
rect 143073 40218 143139 40221
rect 143533 40218 143599 40221
rect 143073 40158 143458 40218
rect 143073 40155 143139 40158
rect 143398 40000 143458 40158
rect 143533 40158 144010 40218
rect 143533 40155 143599 40158
rect 143950 40000 144010 40158
rect 145838 40014 145898 40294
rect 145820 40000 145898 40014
rect 47600 32953 51202 36017
rect 51600 32953 55202 36017
rect 55600 32953 59202 36017
rect 59600 32953 63202 36017
rect 63600 32953 67202 36017
rect 67600 32953 71202 36017
rect 78942 32648 83722 40000
rect 84022 39593 86222 40000
rect 86421 39593 88621 40000
rect 83802 33417 88841 39593
rect 88921 33497 93701 40000
rect 83802 32568 93752 33417
rect 101400 32953 105002 36017
rect 105400 32953 109002 36017
rect 109400 32953 113002 36017
rect 113400 32953 117002 36017
rect 117400 32953 121002 36017
rect 121400 32953 125002 36017
rect 78942 980 93752 32568
rect 132660 30216 132868 39875
rect 132660 26680 132735 30216
rect 132948 30136 133162 40000
rect 132815 27080 133162 30136
rect 133242 37738 141587 39875
rect 141893 38746 143275 39875
rect 141893 38453 142982 38746
rect 143355 38666 143585 40000
rect 141893 38397 142926 38453
rect 141893 38111 142710 38397
rect 143062 38390 143585 38666
rect 143062 38373 143375 38390
rect 143388 38373 143585 38390
rect 143665 39293 143738 39875
rect 143818 39373 144151 40000
rect 144231 39293 145736 39875
rect 143006 38360 143062 38373
rect 143079 38360 143388 38373
rect 143006 38330 143388 38360
rect 143006 38317 143315 38330
rect 143332 38317 143388 38330
rect 141953 38051 142710 38111
rect 133242 36966 141740 37738
rect 142046 37467 142710 38051
rect 142790 38300 143006 38317
rect 143019 38300 143332 38317
rect 142790 38004 143332 38300
rect 143665 38293 145736 39293
rect 143468 38237 145736 38293
rect 142790 37547 143019 38004
rect 143412 37924 145736 38237
rect 143099 37467 145736 37924
rect 142046 36966 145736 37467
rect 133242 36603 145736 36966
rect 145816 36843 145920 40000
rect 146000 36923 147407 39875
rect 146042 36881 147407 36923
rect 145816 36801 145962 36843
rect 145816 36711 146052 36801
rect 146132 36791 147407 36881
rect 145816 36683 145934 36711
rect 145936 36683 146142 36711
rect 146222 36701 147407 36791
rect 145934 36621 146142 36683
rect 133242 36511 145854 36603
rect 145934 36591 146245 36621
rect 133242 36396 145946 36511
rect 146026 36476 146245 36591
rect 133242 33821 146061 36396
rect 133242 33704 145944 33821
rect 146141 33741 146245 36476
rect 133242 33561 145801 33704
rect 146024 33639 146245 33741
rect 146024 33624 146155 33639
rect 146170 33624 146245 33639
rect 145881 33609 146024 33624
rect 146027 33609 146170 33624
rect 133242 33444 145684 33561
rect 145881 33489 146170 33609
rect 146325 33544 147407 36701
rect 145881 33481 146024 33489
rect 146027 33481 146170 33489
rect 145764 33459 145881 33481
rect 145889 33459 146027 33481
rect 133242 33401 145641 33444
rect 133242 33095 143065 33401
rect 145764 33369 146027 33459
rect 146250 33401 147407 33544
rect 145764 33364 145885 33369
rect 145910 33364 146027 33369
rect 145721 33339 145764 33364
rect 145769 33339 145910 33364
rect 145721 33321 145910 33339
rect 143145 33261 145910 33321
rect 146107 33284 147407 33401
rect 143145 33260 145777 33261
rect 145806 33260 145910 33261
rect 143145 33175 145806 33260
rect 145990 33180 147407 33284
rect 145886 33095 147407 33180
rect 133242 27160 147407 33095
rect 155200 32953 158802 36017
rect 159200 32953 162802 36017
rect 163200 32953 166802 36017
rect 167200 32953 170802 36017
rect 171200 32953 174802 36017
rect 175200 32953 178802 36017
rect 132815 26760 133482 27080
rect 133562 26840 147407 27160
rect 132660 26360 133082 26680
rect 133162 26480 133762 26760
rect 133842 26560 147407 26840
rect 133162 26450 133949 26480
rect 133162 26440 133482 26450
rect 133502 26440 133949 26450
rect 132660 26103 133402 26360
rect 133482 26293 133949 26440
rect 134029 26373 147407 26560
rect 133482 26270 133942 26293
rect 133949 26270 134122 26293
rect 133482 26210 134122 26270
rect 133482 26183 133739 26210
rect 133742 26183 134122 26210
rect 134202 26200 147407 26373
rect 133739 26120 134122 26183
rect 132660 25913 133659 26103
rect 133739 26000 134392 26120
rect 133739 25993 133929 26000
rect 133952 25993 134392 26000
rect 132660 25720 133849 25913
rect 133929 25850 134392 25993
rect 134472 25930 147407 26200
rect 133929 25820 134628 25850
rect 133929 25800 134122 25820
rect 134132 25800 134628 25820
rect 132660 25478 134042 25720
rect 134122 25584 134628 25800
rect 134122 25558 134364 25584
rect 134368 25558 134628 25584
rect 134364 25520 134628 25558
rect 132660 25440 134284 25478
rect 132660 20991 134322 25440
rect 134402 21071 134628 25520
rect 134708 20991 147407 25930
rect 132660 0 147407 20991
rect 186486 0 202338 40262
rect 210000 32953 213602 36017
rect 214000 32953 217602 36017
rect 218000 32953 221602 36017
rect 222000 32953 225602 36017
rect 226000 32953 229602 36017
rect 230000 32953 233602 36017
rect 238972 31961 241112 32654
rect 238972 30753 241079 31683
rect 241260 31680 246049 39600
rect 246349 39593 248524 39600
rect 248824 39593 251000 39600
rect 246129 31600 251220 39593
rect 251300 39538 256100 39600
rect 256233 39538 256299 39541
rect 251300 39478 256299 39538
rect 251300 31680 256100 39478
rect 256233 39475 256299 39478
rect 263800 32953 267402 36017
rect 267800 32953 271402 36017
rect 271800 32953 275402 36017
rect 275800 32953 279402 36017
rect 279800 32953 283402 36017
rect 283800 32953 287402 36017
rect 241200 879 256100 31600
rect 295086 0 310938 40262
rect 318600 32953 322202 36017
rect 322600 32953 326202 36017
rect 326600 32953 330202 36017
rect 330600 32953 334202 36017
rect 334600 32953 338202 36017
rect 338600 32953 342202 36017
rect 349886 0 365738 40262
rect 373400 32953 377002 36017
rect 377400 32953 381002 36017
rect 381400 32953 385002 36017
rect 385400 32953 389002 36017
rect 389400 32953 393002 36017
rect 393400 32953 397002 36017
rect 404686 0 420538 40262
rect 428200 32953 431802 36017
rect 432200 32953 435802 36017
rect 436200 32953 439802 36017
rect 440200 32953 443802 36017
rect 444200 32953 447802 36017
rect 448200 32953 451802 36017
rect 459486 0 475338 40262
rect 483000 32953 486602 36017
rect 487000 32953 490602 36017
rect 491000 32953 494602 36017
rect 495000 32953 498602 36017
rect 499000 32953 502602 36017
rect 503000 32953 506602 36017
rect 514286 0 530138 40262
rect 568849 39674 568915 39677
rect 569142 39674 573922 40000
rect 568849 39614 573922 39674
rect 568849 39611 568915 39614
rect 537800 32953 541402 36017
rect 541800 32953 545402 36017
rect 545800 32953 549402 36017
rect 549800 32953 553402 36017
rect 553800 32953 557402 36017
rect 557800 32953 561402 36017
rect 569142 34830 573922 39614
rect 574222 39593 576422 40000
rect 576621 39593 578821 40000
rect 574002 34750 579041 39593
rect 579121 34830 583901 40000
rect 622942 37008 627722 40000
rect 628022 39593 630222 40000
rect 630421 39593 632621 40000
rect 627802 36928 632841 39593
rect 632921 37008 637701 40000
rect 569142 0 583952 34750
rect 591600 32953 595202 36017
rect 595600 32953 599202 36017
rect 599600 32953 603202 36017
rect 603600 32953 607202 36017
rect 607600 32953 611202 36017
rect 611600 32953 615202 36017
rect 622942 0 637752 36928
rect 645400 32953 649002 36017
rect 649400 32953 653002 36017
rect 653400 32953 657002 36017
rect 657400 32953 661002 36017
rect 661400 32953 665002 36017
rect 665400 32953 669002 36017
<< metal4 >>
rect 7 456200 4843 456493
rect 0 455946 4843 456200
rect 28653 407418 28719 526322
rect 32933 455946 33623 483654
rect 36323 456007 37013 483593
rect 37293 455946 38223 483654
rect 38503 455946 39593 483654
rect 679377 423146 680307 451854
rect 680587 423207 681277 451793
rect 688881 423146 688947 544782
rect 93607 36323 132793 37013
rect 93546 31674 132854 31683
rect 93546 30762 132869 31674
rect 93546 30753 132854 30762
rect 93546 28653 192982 28719
<< obsm4 >>
rect 0 1032677 40466 1037600
rect 40546 1032757 75254 1037600
rect 0 1016680 40549 1032677
rect 40800 1016680 75000 1032757
rect 75334 1032677 89666 1037600
rect 89746 1032757 123254 1037600
rect 75193 1016680 89807 1032677
rect 90000 1016680 123000 1032757
rect 123334 1032677 137666 1037600
rect 137746 1032757 171254 1037600
rect 123193 1016680 137807 1032677
rect 138000 1016680 171000 1032757
rect 171334 1032677 185666 1037600
rect 185746 1032757 229641 1037600
rect 171193 1016680 185807 1032677
rect 186000 1016680 220000 1032757
rect 229721 1032677 245097 1037600
rect 245177 1032757 281041 1037600
rect 229448 1016680 245177 1032677
rect 253800 1016680 271400 1032757
rect 281121 1032677 296497 1037600
rect 296577 1032757 339654 1037600
rect 280848 1016680 296577 1032677
rect 305200 1016680 339400 1032757
rect 339734 1032677 354066 1037600
rect 354146 1032757 425054 1037600
rect 339593 1016680 354207 1032677
rect 354400 1016680 388600 1032757
rect 389600 1016680 424800 1032757
rect 425134 1032677 439466 1037600
rect 439546 1032757 474454 1037600
rect 424993 1016680 439607 1032677
rect 439800 1016680 474200 1032757
rect 474534 1032677 488866 1037600
rect 488946 1032757 526054 1037600
rect 474393 1016680 489007 1032677
rect 489200 1016680 525800 1032757
rect 526134 1032677 540466 1037600
rect 540546 1032757 575854 1037600
rect 525993 1016680 540607 1032677
rect 540800 1016680 575600 1032757
rect 575934 1032677 590266 1037600
rect 590346 1032757 627254 1037600
rect 575793 1016680 590407 1032677
rect 590600 1016680 627000 1032757
rect 627334 1032677 641666 1037600
rect 641746 1032757 677887 1037600
rect 642000 1032677 677600 1032757
rect 677967 1032677 717600 1037600
rect 627193 1016680 641807 1032677
rect 642000 1016680 717600 1032677
rect 0 1011527 40349 1016680
rect 40429 1011607 75254 1016600
rect 75334 1011527 89666 1016680
rect 89746 1011607 123254 1016600
rect 123334 1011527 137666 1016680
rect 137746 1011607 171254 1016600
rect 171334 1011527 185666 1016680
rect 185746 1011607 229543 1016600
rect 229623 1011527 245097 1016680
rect 245177 1011607 280943 1016600
rect 281023 1011527 296497 1016680
rect 296577 1011607 339654 1016600
rect 339734 1011527 354066 1016680
rect 354146 1011607 425054 1016600
rect 425134 1011527 439466 1016680
rect 439546 1011607 474454 1016600
rect 474534 1011527 488866 1016680
rect 488946 1011607 526054 1016600
rect 526134 1011527 540466 1016680
rect 540546 1011607 575854 1016600
rect 575934 1011527 590266 1016680
rect 590346 1011607 627254 1016600
rect 627334 1011527 641666 1016680
rect 641746 1011607 678129 1016600
rect 678209 1011527 717600 1016680
rect 0 1011387 40549 1011527
rect 40800 1011387 75000 1011527
rect 75193 1011387 89807 1011527
rect 90000 1011387 123000 1011527
rect 123193 1011387 137807 1011527
rect 138000 1011387 171000 1011527
rect 171193 1011387 185807 1011527
rect 186000 1011387 220000 1011527
rect 229448 1011387 245177 1011527
rect 253800 1011387 271400 1011527
rect 280848 1011387 296577 1011527
rect 305200 1011387 339400 1011527
rect 339593 1011387 354207 1011527
rect 354400 1011387 388600 1011527
rect 389600 1011387 424800 1011527
rect 424993 1011387 439607 1011527
rect 439800 1011387 474200 1011527
rect 474393 1011387 489007 1011527
rect 489200 1011387 525800 1011527
rect 525993 1011387 540607 1011527
rect 540800 1011387 575600 1011527
rect 575793 1011387 590407 1011527
rect 590600 1011387 627000 1011527
rect 627193 1011387 641807 1011527
rect 642000 1011387 717600 1011527
rect 0 1010337 40466 1011387
rect 40546 1010417 75254 1011307
rect 75334 1010337 89666 1011387
rect 89746 1010417 123254 1011307
rect 123334 1010337 137666 1011387
rect 137746 1010417 171254 1011307
rect 171334 1010337 185666 1011387
rect 185746 1010417 229543 1011307
rect 229623 1010337 245097 1011387
rect 245177 1010417 280943 1011307
rect 281023 1010337 296497 1011387
rect 296577 1010417 339654 1011307
rect 339734 1010337 354066 1011387
rect 354146 1010417 425054 1011307
rect 425134 1010337 439466 1011387
rect 439546 1010417 474454 1011307
rect 474534 1010337 488866 1011387
rect 488946 1010417 526054 1011307
rect 526134 1010337 540466 1011387
rect 540546 1010417 575854 1011307
rect 575934 1010337 590266 1011387
rect 590346 1010417 627254 1011307
rect 627334 1010337 641666 1011387
rect 641746 1010417 677896 1011307
rect 677976 1010337 717600 1011387
rect 0 1010217 40549 1010337
rect 40800 1010217 75000 1010337
rect 75193 1010217 89807 1010337
rect 90000 1010217 123000 1010337
rect 123193 1010217 137807 1010337
rect 138000 1010217 171000 1010337
rect 171193 1010217 185807 1010337
rect 186000 1010217 220000 1010337
rect 229448 1010217 245177 1010337
rect 253800 1010217 271400 1010337
rect 280848 1010217 296577 1010337
rect 305200 1010217 339400 1010337
rect 339593 1010217 354207 1010337
rect 354400 1010217 388600 1010337
rect 389600 1010217 424800 1010337
rect 424993 1010217 439607 1010337
rect 439800 1010217 474200 1010337
rect 474393 1010217 489007 1010337
rect 489200 1010217 525800 1010337
rect 525993 1010217 540607 1010337
rect 540800 1010217 575600 1010337
rect 575793 1010217 590407 1010337
rect 590600 1010217 627000 1010337
rect 627193 1010217 641807 1010337
rect 642000 1010217 717600 1010337
rect 0 1009167 40466 1010217
rect 40546 1009247 75254 1010137
rect 75334 1009167 89666 1010217
rect 89746 1009247 123254 1010137
rect 123334 1009167 137666 1010217
rect 137746 1009247 171254 1010137
rect 171334 1009167 185666 1010217
rect 185746 1009247 229543 1010137
rect 229623 1009167 245097 1010217
rect 245177 1009247 280943 1010137
rect 281023 1009167 296497 1010217
rect 296577 1009247 339654 1010137
rect 339734 1009167 354066 1010217
rect 354146 1009247 425054 1010137
rect 425134 1009167 439466 1010217
rect 439546 1009247 474454 1010137
rect 474534 1009167 488866 1010217
rect 488946 1009247 526054 1010137
rect 526134 1009167 540466 1010217
rect 540546 1009247 575854 1010137
rect 575934 1009167 590266 1010217
rect 590346 1009247 627254 1010137
rect 627334 1009167 641666 1010217
rect 641746 1009247 677925 1010137
rect 678005 1009167 717600 1010217
rect 0 1009027 40549 1009167
rect 40800 1009027 75000 1009167
rect 75193 1009027 89807 1009167
rect 90000 1009027 123000 1009167
rect 123193 1009027 137807 1009167
rect 138000 1009027 171000 1009167
rect 171193 1009027 185807 1009167
rect 186000 1009027 220000 1009167
rect 229448 1009027 245177 1009167
rect 253800 1009027 271400 1009167
rect 280848 1009027 296577 1009167
rect 305200 1009027 339400 1009167
rect 339593 1009027 354207 1009167
rect 354400 1009027 388600 1009167
rect 389600 1009027 424800 1009167
rect 424993 1009027 439607 1009167
rect 439800 1009027 474200 1009167
rect 474393 1009027 489007 1009167
rect 489200 1009027 525800 1009167
rect 525993 1009027 540607 1009167
rect 540800 1009027 575600 1009167
rect 575793 1009027 590407 1009167
rect 590600 1009027 627000 1009167
rect 627193 1009027 641807 1009167
rect 642000 1009027 717600 1009167
rect 0 1008801 35285 1009027
rect 35365 1008881 388600 1008947
rect 389600 1008881 575854 1008947
rect 575934 1008901 590266 1009027
rect 590346 1008881 682235 1008947
rect 0 1008145 35338 1008801
rect 35418 1008225 682182 1008821
rect 682315 1008801 717600 1009027
rect 0 1007849 36409 1008145
rect 36489 1007929 75254 1008165
rect 75334 1007949 89666 1008145
rect 89746 1007929 123254 1008165
rect 123334 1007949 137666 1008145
rect 137746 1007929 171254 1008165
rect 171334 1007949 185666 1008145
rect 185746 1007929 229448 1008165
rect 229528 1007949 245097 1008145
rect 245177 1007929 280848 1008165
rect 280928 1007949 296497 1008145
rect 296577 1007929 339654 1008165
rect 339734 1007949 354066 1008145
rect 354146 1007929 388600 1008165
rect 389600 1007929 425054 1008165
rect 425134 1007949 439466 1008145
rect 439546 1007929 474454 1008165
rect 474534 1007949 488866 1008145
rect 488946 1007929 526054 1008165
rect 526134 1007949 540466 1008145
rect 540546 1007929 575854 1008165
rect 575934 1007949 590266 1008145
rect 590346 1007929 627254 1008165
rect 627334 1007949 641666 1008145
rect 641746 1007929 681910 1008165
rect 682262 1008145 717600 1008801
rect 0 1007293 36545 1007849
rect 0 1007067 36005 1007293
rect 36625 1007273 681787 1007869
rect 681990 1007849 717600 1008145
rect 36085 1007147 388600 1007213
rect 389600 1007147 575854 1007213
rect 575934 1007067 590266 1007193
rect 590346 1007147 681515 1007213
rect 681867 1007193 717600 1007849
rect 681595 1007067 717600 1007193
rect 0 1006927 40549 1007067
rect 75193 1006927 89807 1007067
rect 123193 1006927 137807 1007067
rect 171193 1006927 185807 1007067
rect 229448 1006927 245177 1007067
rect 280848 1006927 296577 1007067
rect 339593 1006927 354207 1007067
rect 424993 1006927 439607 1007067
rect 474393 1006927 489007 1007067
rect 525993 1006927 540607 1007067
rect 575793 1006927 590407 1007067
rect 627193 1006927 641807 1007067
rect 677600 1006927 717600 1007067
rect 0 1005837 40466 1006927
rect 40546 1005917 75254 1006847
rect 75334 1005837 89666 1006927
rect 89746 1005917 123254 1006847
rect 123334 1005837 137666 1006927
rect 137746 1005917 171254 1006847
rect 171334 1005837 185666 1006927
rect 185746 1005917 229450 1006847
rect 229530 1005837 245097 1006927
rect 245177 1005917 280850 1006847
rect 280930 1005837 296497 1006927
rect 296577 1005917 339654 1006847
rect 339734 1005837 354066 1006927
rect 354146 1005917 389600 1006847
rect 390600 1005917 425054 1006847
rect 425134 1005837 439466 1006927
rect 439546 1005917 474454 1006847
rect 474534 1005837 488866 1006927
rect 488946 1005917 526054 1006847
rect 526134 1005837 540466 1006927
rect 540546 1005917 575854 1006847
rect 575934 1005837 590266 1006927
rect 590346 1005917 627254 1006847
rect 627334 1005837 641666 1006927
rect 641746 1005917 677895 1006847
rect 677975 1005837 717600 1006927
rect 0 1005717 40549 1005837
rect 75193 1005717 89807 1005837
rect 123193 1005717 137807 1005837
rect 171193 1005717 185807 1005837
rect 229448 1005717 245177 1005837
rect 280848 1005717 296577 1005837
rect 339593 1005717 354207 1005837
rect 424993 1005717 439607 1005837
rect 474393 1005717 489007 1005837
rect 525993 1005717 540607 1005837
rect 575793 1005717 590407 1005837
rect 627193 1005717 641807 1005837
rect 677600 1005717 717600 1005837
rect 0 1004867 40466 1005717
rect 40546 1004947 75254 1005637
rect 75334 1004867 89666 1005717
rect 89746 1004947 123254 1005637
rect 123334 1004867 137666 1005717
rect 137746 1004947 171254 1005637
rect 171334 1004867 185666 1005717
rect 185746 1004947 229543 1005637
rect 229623 1004867 245097 1005717
rect 245177 1004947 280943 1005637
rect 281023 1004867 296497 1005717
rect 296577 1004947 339654 1005637
rect 339734 1004867 354066 1005717
rect 354146 1004947 388600 1005637
rect 389600 1004947 425054 1005637
rect 425134 1004867 439466 1005717
rect 439546 1004947 474454 1005637
rect 474534 1004867 488866 1005717
rect 488946 1004947 526054 1005637
rect 526134 1004867 540466 1005717
rect 540546 1004947 575854 1005637
rect 575934 1004867 590266 1005717
rect 590346 1004947 627254 1005637
rect 627334 1004867 641666 1005717
rect 641746 1004947 677867 1005637
rect 677947 1004867 717600 1005717
rect 0 1004747 40549 1004867
rect 75193 1004747 89807 1004867
rect 123193 1004747 137807 1004867
rect 171193 1004747 185807 1004867
rect 229448 1004747 245177 1004867
rect 280848 1004747 296577 1004867
rect 339593 1004747 354207 1004867
rect 424993 1004747 439607 1004867
rect 474393 1004747 489007 1004867
rect 525993 1004747 540607 1004867
rect 575793 1004747 590407 1004867
rect 627193 1004747 641807 1004867
rect 677600 1004747 717600 1004867
rect 0 1003897 40466 1004747
rect 40546 1003977 75254 1004667
rect 75334 1003897 89666 1004747
rect 89746 1003977 123254 1004667
rect 123334 1003897 137666 1004747
rect 137746 1003977 171254 1004667
rect 171334 1003897 185666 1004747
rect 185746 1003977 229543 1004667
rect 229623 1003897 245097 1004747
rect 245177 1003977 280943 1004667
rect 281023 1003897 296497 1004747
rect 296577 1003977 339654 1004667
rect 339734 1003897 354066 1004747
rect 354146 1003977 425054 1004667
rect 425134 1003897 439466 1004747
rect 439546 1003977 474454 1004667
rect 474534 1003897 488866 1004747
rect 488946 1003977 526054 1004667
rect 526134 1003897 540466 1004747
rect 540546 1003977 575854 1004667
rect 575934 1003897 590266 1004747
rect 590346 1003977 627254 1004667
rect 627334 1003897 641666 1004747
rect 641746 1003977 677877 1004667
rect 677957 1003897 717600 1004747
rect 0 1003777 40549 1003897
rect 75193 1003777 89807 1003897
rect 123193 1003777 137807 1003897
rect 171193 1003777 185807 1003897
rect 229448 1003777 245177 1003897
rect 280848 1003777 296577 1003897
rect 339593 1003777 354207 1003897
rect 424993 1003777 439607 1003897
rect 474393 1003777 489007 1003897
rect 525993 1003777 540607 1003897
rect 575793 1003777 590407 1003897
rect 627193 1003777 641807 1003897
rect 677600 1003777 717600 1003897
rect 0 1002687 40466 1003777
rect 40546 1002767 75254 1003697
rect 75334 1002687 89666 1003777
rect 89746 1002767 123254 1003697
rect 123334 1002687 137666 1003777
rect 137746 1002767 171254 1003697
rect 171334 1002687 185666 1003777
rect 185746 1002767 229543 1003697
rect 229623 1002687 245097 1003777
rect 245177 1002767 280943 1003697
rect 281023 1002687 296497 1003777
rect 296577 1002767 339654 1003697
rect 339734 1002687 354066 1003777
rect 354146 1002767 425054 1003697
rect 425134 1002687 439466 1003777
rect 439546 1002767 474454 1003697
rect 474534 1002687 488866 1003777
rect 488946 1002767 526054 1003697
rect 526134 1002687 540466 1003777
rect 540546 1002767 575854 1003697
rect 575934 1002687 590266 1003777
rect 590346 1002767 627254 1003697
rect 627334 1002687 641666 1003777
rect 641746 1002767 677920 1003697
rect 678000 1002687 717600 1003777
rect 0 1002567 40549 1002687
rect 75193 1002567 89807 1002687
rect 123193 1002567 137807 1002687
rect 171193 1002567 185807 1002687
rect 229448 1002567 245177 1002687
rect 280848 1002567 296577 1002687
rect 339593 1002567 354207 1002687
rect 424993 1002567 439607 1002687
rect 474393 1002567 489007 1002687
rect 525993 1002567 540607 1002687
rect 575793 1002567 590407 1002687
rect 627193 1002567 641807 1002687
rect 677600 1002567 717600 1002687
rect 0 1002315 40466 1002567
rect 0 998209 28573 1002315
rect 28799 1002262 40466 1002315
rect 0 997967 20920 998209
rect 0 997600 4843 997887
rect 4923 997600 20920 997967
rect 0 970200 20920 997600
rect 0 969946 4843 970200
rect 4923 969866 20920 970007
rect 21000 969946 25993 998129
rect 26073 998005 28573 998209
rect 26073 997976 27383 998005
rect 26073 970200 26213 997976
rect 26073 969866 26213 970007
rect 26293 969946 27183 997896
rect 27263 970200 27383 997976
rect 27263 969866 27383 970007
rect 27463 969946 28353 997925
rect 28433 970200 28573 998005
rect 28433 969866 28573 970007
rect 0 955534 28573 969866
rect 0 955200 4843 955454
rect 4923 955393 20920 955534
rect 0 928000 20920 955200
rect 0 927957 4850 928000
rect 0 927746 4843 927957
rect 4923 927666 20920 928000
rect 21000 927746 25993 955454
rect 26073 955393 26213 955534
rect 26073 927666 26213 955200
rect 26293 927746 27183 955454
rect 27263 955393 27383 955534
rect 27263 927666 27383 955200
rect 27463 927746 28353 955454
rect 28433 955393 28573 955534
rect 28433 927666 28573 955200
rect 0 913334 28573 927666
rect 0 913000 4843 913254
rect 4923 913000 20920 913334
rect 0 885800 20920 913000
rect 0 885546 4843 885800
rect 4923 885466 20920 885607
rect 21000 885546 25993 913254
rect 26073 885800 26213 913334
rect 26073 885466 26213 885607
rect 26293 885546 27183 913254
rect 27263 885800 27383 913334
rect 27263 885466 27383 885607
rect 27463 885546 28353 913254
rect 28433 885800 28573 913334
rect 28433 885466 28573 885607
rect 0 871134 28573 885466
rect 0 870800 4843 871054
rect 4923 870993 20920 871134
rect 0 843400 20920 870800
rect 0 843146 4843 843400
rect 4923 843066 20920 843207
rect 21000 843146 25993 871054
rect 26073 870993 26213 871134
rect 26073 843400 26213 870800
rect 26073 843066 26213 843207
rect 26293 843146 27183 871054
rect 27263 870993 27383 871134
rect 27263 843400 27383 870800
rect 27263 843066 27383 843207
rect 27463 843146 28353 871054
rect 28433 870993 28573 871134
rect 28433 843400 28573 870800
rect 28433 843066 28573 843207
rect 28653 843146 28719 1002235
rect 0 828734 28699 843066
rect 0 828400 4843 828654
rect 4923 828593 20920 828734
rect 0 801200 20920 828400
rect 0 800946 4843 801200
rect 4923 800866 20920 800994
rect 21000 800946 25993 828654
rect 26073 828593 26213 828734
rect 26073 801200 26213 828400
rect 26073 800866 26213 800994
rect 26293 800946 27183 828654
rect 27263 828593 27383 828734
rect 27263 801200 27383 828400
rect 27263 800866 27383 800994
rect 27463 800946 28353 828654
rect 28433 828593 28573 828734
rect 28433 801200 28573 828400
rect 28433 800866 28573 800994
rect 0 794538 28573 800866
rect 28653 794618 28719 828654
rect 0 792872 28699 794538
rect 28779 792952 29375 1002182
rect 29455 1001990 40466 1002262
rect 29435 969946 29671 1001910
rect 29751 1001867 40466 1001990
rect 29455 955534 29651 969866
rect 29435 927746 29671 955454
rect 29455 913334 29651 927666
rect 29435 885546 29671 913254
rect 29455 871134 29651 885466
rect 29435 843146 29671 871054
rect 29455 828734 29651 843066
rect 29435 800946 29671 828654
rect 29455 796013 29651 800866
rect 29731 796093 30327 1001787
rect 30407 1001595 40466 1001867
rect 30387 843146 30453 1001515
rect 30533 1001477 40466 1001595
rect 40546 1001557 75254 1002487
rect 75334 1001477 89666 1002567
rect 89746 1001557 123254 1002487
rect 123334 1001477 137666 1002567
rect 137746 1001557 171254 1002487
rect 171334 1001477 185666 1002567
rect 185746 1001557 229543 1002487
rect 229623 1001477 244161 1002567
rect 244241 1001557 280943 1002487
rect 281023 1001477 295561 1002567
rect 295641 1001557 339654 1002487
rect 339734 1001477 354066 1002567
rect 354146 1001557 425054 1002487
rect 425134 1001477 439466 1002567
rect 439546 1001557 474454 1002487
rect 474534 1001477 488866 1002567
rect 488946 1001557 526054 1002487
rect 526134 1001477 540466 1002567
rect 540546 1001557 575854 1002487
rect 575934 1001477 590266 1002567
rect 590346 1001557 627254 1002487
rect 627334 1001477 641666 1002567
rect 641746 1001557 677905 1002487
rect 677985 1002315 717600 1002567
rect 677985 1002262 688801 1002315
rect 677985 1001595 688145 1002262
rect 677985 1001477 687067 1001595
rect 30533 1001357 40549 1001477
rect 75193 1001357 89807 1001477
rect 123193 1001357 137807 1001477
rect 171193 1001357 185807 1001477
rect 229448 1001357 245177 1001477
rect 280848 1001357 296577 1001477
rect 339593 1001357 354207 1001477
rect 424993 1001357 439607 1001477
rect 474393 1001357 489007 1001477
rect 525993 1001357 540607 1001477
rect 575793 1001357 590407 1001477
rect 627193 1001357 641807 1001477
rect 677600 1001357 687067 1001477
rect 30533 1000507 40469 1001357
rect 40549 1000587 75193 1001277
rect 75273 1000507 89727 1001357
rect 89807 1000587 123193 1001277
rect 123273 1000507 137727 1001357
rect 137807 1000587 171193 1001277
rect 171273 1000507 185727 1001357
rect 185807 1000587 229543 1001277
rect 229623 1000507 244161 1001357
rect 244241 1000587 280943 1001277
rect 281023 1000507 295561 1001357
rect 295641 1000587 339593 1001277
rect 339673 1000507 354127 1001357
rect 354207 1000587 388600 1001277
rect 389600 1000587 424993 1001277
rect 425073 1000507 439527 1001357
rect 439607 1000587 474393 1001277
rect 474473 1000507 488927 1001357
rect 489007 1000587 525993 1001277
rect 526073 1000507 540527 1001357
rect 540607 1000587 575793 1001277
rect 575873 1000507 590327 1001357
rect 590407 1000587 627193 1001277
rect 627273 1000507 641727 1001357
rect 641807 1000587 677894 1001277
rect 677974 1000507 687067 1001357
rect 30533 1000387 40549 1000507
rect 75193 1000387 89807 1000507
rect 123193 1000387 137807 1000507
rect 171193 1000387 185807 1000507
rect 229448 1000387 245177 1000507
rect 280848 1000387 296577 1000507
rect 339593 1000387 354207 1000507
rect 424993 1000387 439607 1000507
rect 474393 1000387 489007 1000507
rect 525993 1000387 540607 1000507
rect 575793 1000387 590407 1000507
rect 627193 1000387 641807 1000507
rect 677600 1000387 687067 1000507
rect 30533 999297 40466 1000387
rect 40546 999377 75254 1000307
rect 75334 999297 89666 1000387
rect 89746 999377 123254 1000307
rect 123334 999297 137666 1000387
rect 137746 999377 171254 1000307
rect 171334 999297 185666 1000387
rect 185746 999377 229543 1000307
rect 229623 999297 245097 1000387
rect 245177 999377 280943 1000307
rect 281023 999297 296497 1000387
rect 296577 999377 339654 1000307
rect 339734 999297 354066 1000387
rect 354146 999377 389600 1000307
rect 390600 999377 425054 1000307
rect 425134 999297 439466 1000387
rect 439546 999377 474454 1000307
rect 474534 999297 488866 1000387
rect 488946 999377 526054 1000307
rect 526134 999297 540466 1000387
rect 540546 999377 575854 1000307
rect 575934 999297 590266 1000387
rect 590346 999377 627254 1000307
rect 627334 999297 641666 1000387
rect 641746 999377 678357 1000307
rect 678437 999297 687067 1000387
rect 30533 999177 40549 999297
rect 75193 999177 89807 999297
rect 123193 999177 137807 999297
rect 171193 999177 185807 999297
rect 229448 999177 245177 999297
rect 280848 999177 296577 999297
rect 339593 999177 354207 999297
rect 424993 999177 439607 999297
rect 474393 999177 489007 999297
rect 525993 999177 540607 999297
rect 575793 999177 590407 999297
rect 627193 999177 641807 999297
rect 677600 999177 687067 999297
rect 30533 998437 40466 999177
rect 30533 998000 37213 998437
rect 30533 997975 33823 998000
rect 30533 997600 30673 997975
rect 31763 997957 33823 997975
rect 31763 997947 32853 997957
rect 30533 969866 30673 970007
rect 30753 969946 31683 997895
rect 31763 997600 31883 997947
rect 31763 969866 31883 970007
rect 31963 969946 32653 997867
rect 32733 997600 32853 997947
rect 32733 969866 32853 970007
rect 32933 969946 33623 997877
rect 33703 997600 33823 997957
rect 34913 997985 37213 998000
rect 33703 969866 33823 970007
rect 33903 969946 34833 997920
rect 34913 997600 35033 997985
rect 36123 997974 37213 997985
rect 34913 969866 35033 970007
rect 35113 969946 36043 997905
rect 36123 997600 36243 997974
rect 36323 970007 37013 997894
rect 37093 997600 37213 997974
rect 36123 969927 36243 970007
rect 37093 969927 37213 970007
rect 37293 969946 38223 998357
rect 38303 998150 40466 998437
rect 38303 997600 38423 998150
rect 36123 969866 37213 969927
rect 38303 969866 38423 970007
rect 38503 969946 39593 998070
rect 39673 997927 40466 998150
rect 40546 998007 75254 999097
rect 75334 998007 89666 999177
rect 89746 998007 123254 999097
rect 123334 998007 137666 999177
rect 137746 998007 171254 999097
rect 171334 998007 185666 999177
rect 185746 998007 229543 999097
rect 229623 998007 245097 999177
rect 245177 998007 280943 999097
rect 281023 998007 296497 999177
rect 296577 998007 339654 999097
rect 339734 998007 354066 999177
rect 354146 998007 425054 999097
rect 425134 998007 439466 999177
rect 439546 998007 474454 999097
rect 474534 998007 488866 999177
rect 488946 998007 526054 999097
rect 526134 998007 540466 999177
rect 540546 998007 575854 999097
rect 575934 998007 590266 999177
rect 590346 998007 627254 999097
rect 627334 998007 641666 999177
rect 641746 998007 678070 999097
rect 678150 997927 687067 999177
rect 39673 997600 40549 997927
rect 677600 997134 687067 997927
rect 677600 997051 677927 997134
rect 30533 955534 39593 969866
rect 678007 958857 679097 997054
rect 679177 997051 679297 997134
rect 680387 997131 681477 997134
rect 679177 958777 679297 958952
rect 679377 958857 680307 997054
rect 680387 997051 680507 997131
rect 681357 997051 681477 997131
rect 680387 958777 680507 958952
rect 680587 958857 681277 997051
rect 681357 958777 681477 958952
rect 681557 958857 682487 997054
rect 682567 997051 682687 997134
rect 682567 958777 682687 958952
rect 682767 958857 683697 997054
rect 683777 997051 683897 997134
rect 683777 958777 683897 958952
rect 683977 958857 684667 997054
rect 684747 997051 684867 997134
rect 684747 958777 684867 958952
rect 684947 958857 685637 997054
rect 685717 997051 685837 997134
rect 685717 958870 685837 958952
rect 685917 958950 686847 997054
rect 686927 997051 687067 997134
rect 686927 958870 687067 958952
rect 685717 958777 687067 958870
rect 30533 955393 30673 955534
rect 30533 927666 30673 928000
rect 30753 927746 31683 955454
rect 31763 955393 31883 955534
rect 31763 927666 31883 928000
rect 31963 927746 32653 955454
rect 32733 955393 32853 955534
rect 32733 927666 32853 928000
rect 32933 927746 33623 955454
rect 33703 955393 33823 955534
rect 33903 930187 34833 955454
rect 34913 955393 35033 955534
rect 36123 955473 37213 955534
rect 33703 927666 33823 928000
rect 33903 927987 34840 930187
rect 33903 927746 34833 927987
rect 34913 927666 35033 928000
rect 35113 927746 36043 955454
rect 36123 955393 36243 955473
rect 37093 955393 37213 955473
rect 36123 927727 36243 928000
rect 36323 927807 37013 955393
rect 37093 927727 37213 928000
rect 37293 927746 38223 955454
rect 38303 955393 38423 955534
rect 36123 927666 37213 927727
rect 38303 927666 38423 928000
rect 38503 927746 39593 955454
rect 678007 944239 687067 958777
rect 678007 943303 680507 944239
rect 679177 943223 679297 943303
rect 680387 943223 680507 943303
rect 30533 913334 39593 927666
rect 30533 913000 30673 913334
rect 30753 913014 31683 913254
rect 30753 910805 31690 913014
rect 31763 913000 31883 913334
rect 30533 885466 30673 885607
rect 30753 885546 31683 910805
rect 31763 885466 31883 885607
rect 31963 885546 32653 913254
rect 32733 913000 32853 913334
rect 32733 885466 32853 885607
rect 32933 885546 33623 913254
rect 33703 913000 33823 913334
rect 33703 885466 33823 885607
rect 33903 885546 34833 913254
rect 34913 913000 35033 913334
rect 36123 913273 37213 913334
rect 34913 885466 35033 885607
rect 35113 885546 36043 913254
rect 36123 913000 36243 913273
rect 36323 885607 37013 913193
rect 37093 913000 37213 913273
rect 36123 885527 36243 885607
rect 37093 885527 37213 885607
rect 37293 885546 38223 913254
rect 38303 913000 38423 913334
rect 36123 885466 37213 885527
rect 38303 885466 38423 885607
rect 38503 885546 39593 913254
rect 678007 906146 679097 943223
rect 679177 906066 679297 906400
rect 679377 906146 680307 943223
rect 680387 906127 680507 906400
rect 680587 906207 681277 944159
rect 681357 943223 681477 944239
rect 681357 906127 681477 906400
rect 681557 906146 682487 944159
rect 682567 943303 687067 944239
rect 682567 943223 682687 943303
rect 683777 943223 683897 943303
rect 684747 943223 684867 943303
rect 685717 943223 685837 943303
rect 686927 943223 687067 943303
rect 680387 906066 681477 906127
rect 682567 906066 682687 906400
rect 682767 906146 683697 943223
rect 683777 906066 683897 906400
rect 683977 906146 684667 943223
rect 684747 906066 684867 906400
rect 684947 906146 685637 943223
rect 685917 908595 686847 943223
rect 685717 906066 685837 906400
rect 685910 906386 686847 908595
rect 685917 906146 686847 906386
rect 686927 906066 687067 906400
rect 678007 891734 687067 906066
rect 30533 871134 39593 885466
rect 30533 870993 30673 871134
rect 30533 843066 30673 843207
rect 30753 843146 31683 871054
rect 31763 870993 31883 871134
rect 31763 843066 31883 843207
rect 31963 843146 32653 871054
rect 32733 870993 32853 871134
rect 32733 843066 32853 843207
rect 32933 843146 33623 871054
rect 33703 870993 33823 871134
rect 33703 843066 33823 843207
rect 33903 843146 34833 871054
rect 34913 870993 35033 871134
rect 36123 871073 37213 871134
rect 34913 843066 35033 843207
rect 35113 843146 36043 871054
rect 36123 870993 36243 871073
rect 37093 870993 37213 871073
rect 36323 843207 37013 870993
rect 36123 843127 36243 843207
rect 37093 843127 37213 843207
rect 37293 843146 38223 871054
rect 38303 870993 38423 871134
rect 36123 843066 37213 843127
rect 38303 843066 38423 843207
rect 38503 843146 39593 871054
rect 677707 862666 677927 862807
rect 678007 862746 679097 891654
rect 679177 891400 679297 891734
rect 680387 891673 681477 891734
rect 679177 862666 679297 862807
rect 679377 862746 680307 891654
rect 680387 891400 680507 891673
rect 680587 862807 681277 891593
rect 681357 891400 681477 891673
rect 680387 862727 680507 862807
rect 681357 862727 681477 862807
rect 681557 862746 682487 891654
rect 682567 891400 682687 891734
rect 682767 891413 683697 891654
rect 682760 889213 683697 891413
rect 683777 891400 683897 891734
rect 680387 862666 681477 862727
rect 682567 862666 682687 862807
rect 682767 862746 683697 889213
rect 683777 862666 683897 862807
rect 683977 862746 684667 891654
rect 684747 891400 684867 891734
rect 684747 862666 684867 862807
rect 684947 862746 685637 891654
rect 685717 891400 685837 891734
rect 685717 862666 685837 862807
rect 685917 862746 686847 891654
rect 686927 891400 687067 891734
rect 686927 862666 687067 862807
rect 677707 862398 687067 862666
rect 687147 862478 687213 1001515
rect 687293 1001191 688145 1001595
rect 687293 1001055 687849 1001191
rect 677707 853662 687193 862398
rect 677707 847334 687067 853662
rect 677707 847206 677927 847334
rect 30407 828734 39593 843066
rect 29455 795709 30307 796013
rect 29455 792872 29651 795709
rect 0 792568 29651 792872
rect 0 785802 28699 792568
rect 0 785534 28573 785802
rect 0 785200 4843 785454
rect 4923 785393 20920 785534
rect 0 758000 20920 785200
rect 0 757746 4843 758000
rect 4923 757666 20920 757794
rect 21000 757746 25993 785454
rect 26073 785393 26213 785534
rect 26073 758000 26213 785200
rect 26073 757666 26213 757794
rect 26293 757746 27183 785454
rect 27263 785393 27383 785534
rect 27263 758000 27383 785200
rect 27263 757666 27383 757794
rect 27463 757746 28353 785454
rect 28433 785393 28573 785534
rect 28433 758000 28573 785200
rect 28433 757666 28573 757794
rect 0 751338 28573 757666
rect 28653 751418 28719 785722
rect 0 749672 28699 751338
rect 28779 749752 29375 792488
rect 29455 785534 29651 792568
rect 29435 757746 29671 785454
rect 29455 752813 29651 757666
rect 29731 752893 30327 795629
rect 30387 794618 30453 828654
rect 30533 828593 30673 828734
rect 30533 800866 30673 800994
rect 30753 800946 31683 828654
rect 31763 828593 31883 828734
rect 31763 800866 31883 800994
rect 31963 800946 32653 828654
rect 32733 828593 32853 828734
rect 32733 800866 32853 800994
rect 32933 800946 33623 828654
rect 33703 828593 33823 828734
rect 33703 800866 33823 800994
rect 33903 800946 34833 828654
rect 34913 828593 35033 828734
rect 36123 828673 37213 828734
rect 34913 800866 35033 800994
rect 35113 800946 36043 828654
rect 36123 828593 36243 828673
rect 37093 828593 37213 828673
rect 36323 800994 37013 828593
rect 36123 800914 36243 800994
rect 37093 800914 37213 800994
rect 37293 800946 38223 828654
rect 38303 828593 38423 828734
rect 36123 800866 37213 800914
rect 38303 800866 38423 800994
rect 38503 800946 39593 828654
rect 678007 818546 679097 847254
rect 679177 847206 679297 847334
rect 680387 847286 681477 847334
rect 679177 818466 679297 818607
rect 679377 818546 680307 847254
rect 680387 847206 680507 847286
rect 681357 847206 681477 847286
rect 680587 818607 681277 847206
rect 680387 818527 680507 818607
rect 681357 818527 681477 818607
rect 681557 818546 682487 847254
rect 682567 847206 682687 847334
rect 680387 818466 681477 818527
rect 682567 818466 682687 818607
rect 682767 818546 683697 847254
rect 683777 847206 683897 847334
rect 683777 818466 683897 818607
rect 683977 818546 684667 847254
rect 684747 847206 684867 847334
rect 684747 818466 684867 818607
rect 684947 818546 685637 847254
rect 685717 847206 685837 847334
rect 685717 818466 685837 818607
rect 685917 818546 686847 847254
rect 686927 847206 687067 847334
rect 686927 818466 687067 818607
rect 678007 804134 687067 818466
rect 39673 800866 39893 800994
rect 30533 794538 39893 800866
rect 30407 785802 39893 794538
rect 29455 752509 30307 752813
rect 29455 749672 29651 752509
rect 0 749368 29651 749672
rect 0 742602 28699 749368
rect 0 742334 28573 742602
rect 0 742000 4843 742254
rect 4923 742193 20920 742334
rect 0 714800 20920 742000
rect 0 714546 4843 714800
rect 4923 714466 20920 714594
rect 21000 714546 25993 742254
rect 26073 742193 26213 742334
rect 26073 714800 26213 742000
rect 26073 714466 26213 714594
rect 26293 714546 27183 742254
rect 27263 742193 27383 742334
rect 27263 714800 27383 742000
rect 27263 714466 27383 714594
rect 27463 714546 28353 742254
rect 28433 742193 28573 742334
rect 28433 714800 28573 742000
rect 28433 714466 28573 714594
rect 0 708138 28573 714466
rect 28653 708218 28719 742522
rect 0 706472 28699 708138
rect 28779 706552 29375 749288
rect 29455 742334 29651 749368
rect 29435 714546 29671 742254
rect 29455 709613 29651 714466
rect 29731 709693 30327 752429
rect 30387 751418 30453 785722
rect 30533 785534 39893 785802
rect 30533 785393 30673 785534
rect 30533 757666 30673 757794
rect 30753 757746 31683 785454
rect 31763 785393 31883 785534
rect 31763 757666 31883 757794
rect 31963 757746 32653 785454
rect 32733 785393 32853 785534
rect 32733 757666 32853 757794
rect 32933 757746 33623 785454
rect 33703 785393 33823 785534
rect 33703 757666 33823 757794
rect 33903 757746 34833 785454
rect 34913 785393 35033 785534
rect 36123 785473 37213 785534
rect 34913 757666 35033 757794
rect 35113 757746 36043 785454
rect 36123 785393 36243 785473
rect 37093 785393 37213 785473
rect 36323 757794 37013 785393
rect 36123 757714 36243 757794
rect 37093 757714 37213 757794
rect 37293 757746 38223 785454
rect 38303 785393 38423 785534
rect 36123 757666 37213 757714
rect 38303 757666 38423 757794
rect 38503 757746 39593 785454
rect 39673 785393 39893 785534
rect 677707 775266 677927 775407
rect 678007 775346 679097 804054
rect 679177 803993 679297 804134
rect 680387 804073 681477 804134
rect 679177 775266 679297 775407
rect 679377 775346 680307 804054
rect 680387 803993 680507 804073
rect 681357 803993 681477 804073
rect 680587 775407 681277 803993
rect 680387 775327 680507 775407
rect 681357 775327 681477 775407
rect 681557 775346 682487 804054
rect 682567 803993 682687 804134
rect 680387 775266 681477 775327
rect 682567 775266 682687 775407
rect 682767 775346 683697 804054
rect 683777 803993 683897 804134
rect 683777 775266 683897 775407
rect 683977 775346 684667 804054
rect 684747 803993 684867 804134
rect 684747 775266 684867 775407
rect 684947 775346 685637 804054
rect 685717 803993 685837 804134
rect 685717 775266 685837 775407
rect 685917 775346 686847 804054
rect 686927 803993 687067 804134
rect 686927 775266 687067 775407
rect 677707 774998 687067 775266
rect 687147 775078 687213 853582
rect 687273 852571 687869 1000975
rect 687929 958952 688165 1001111
rect 687949 943303 688145 958872
rect 687929 906146 688165 943223
rect 687949 891734 688145 906066
rect 687929 862746 688165 891654
rect 687949 855632 688145 862666
rect 688225 855712 688821 1002182
rect 688881 862478 688947 1002235
rect 689027 997251 717600 1002315
rect 689027 997134 691527 997251
rect 689027 997051 689167 997134
rect 689027 968400 689167 996800
rect 689027 958777 689167 958952
rect 689247 958857 690137 997054
rect 690217 997051 690337 997134
rect 690217 968400 690337 996800
rect 690217 958777 690337 958952
rect 690417 958857 691307 997054
rect 691387 997051 691527 997134
rect 691387 968400 691527 996800
rect 691387 958777 691527 958952
rect 691607 958857 696600 997171
rect 696680 997134 717600 997251
rect 696680 997051 712677 997134
rect 712757 996800 717600 997054
rect 696680 968400 717600 996800
rect 696680 958777 712677 958952
rect 689027 958679 712677 958777
rect 712757 958759 717600 968400
rect 689027 943303 717600 958679
rect 689027 943223 689167 943303
rect 690217 943223 690337 943303
rect 691387 943223 691527 943303
rect 696680 943223 712677 943303
rect 689027 906066 689167 934600
rect 689247 906146 690137 943223
rect 690217 906066 690337 934600
rect 690417 906146 691307 943223
rect 691387 906066 691527 934600
rect 691607 906146 696600 943223
rect 712757 934600 717600 943223
rect 696680 906400 717600 934600
rect 696680 906066 712677 906400
rect 712757 906146 717600 906400
rect 689027 891734 717600 906066
rect 689027 863000 689167 891734
rect 689027 862666 689167 862807
rect 689247 862746 690137 891654
rect 690217 863000 690337 891734
rect 690217 862666 690337 862807
rect 690417 862746 691307 891654
rect 691387 863000 691527 891734
rect 691387 862666 691527 862807
rect 691607 862746 696600 891654
rect 696680 891400 712677 891734
rect 712757 891443 717600 891654
rect 712750 891400 717600 891443
rect 696680 863000 717600 891400
rect 696680 862666 712677 862807
rect 712757 862746 717600 863000
rect 689027 862398 717600 862666
rect 688901 855632 717600 862398
rect 687949 855328 717600 855632
rect 687949 852491 688145 855328
rect 687293 852187 688145 852491
rect 677707 766262 687193 774998
rect 677707 759934 687067 766262
rect 677707 759806 677927 759934
rect 39673 757666 39893 757794
rect 30533 751338 39893 757666
rect 30407 742602 39893 751338
rect 29455 709309 30307 709613
rect 29455 706472 29651 709309
rect 0 706168 29651 706472
rect 0 699402 28699 706168
rect 0 699134 28573 699402
rect 0 698800 4843 699054
rect 4923 698993 20920 699134
rect 0 671400 20920 698800
rect 0 671146 4843 671400
rect 4923 671066 20920 671194
rect 21000 671146 25993 699054
rect 26073 698993 26213 699134
rect 26073 671400 26213 698800
rect 26073 671066 26213 671194
rect 26293 671146 27183 699054
rect 27263 698993 27383 699134
rect 27263 671400 27383 698800
rect 27263 671066 27383 671194
rect 27463 671146 28353 699054
rect 28433 698993 28573 699134
rect 28433 671400 28573 698800
rect 28433 671066 28573 671194
rect 0 664738 28573 671066
rect 28653 664818 28719 699322
rect 0 663072 28699 664738
rect 28779 663152 29375 706088
rect 29455 699134 29651 706168
rect 29435 671146 29671 699054
rect 29455 666213 29651 671066
rect 29731 666293 30327 709229
rect 30387 708218 30453 742522
rect 30533 742334 39893 742602
rect 30533 742193 30673 742334
rect 30533 714466 30673 714594
rect 30753 714546 31683 742254
rect 31763 742193 31883 742334
rect 31763 714466 31883 714594
rect 31963 714546 32653 742254
rect 32733 742193 32853 742334
rect 32733 714466 32853 714594
rect 32933 714546 33623 742254
rect 33703 742193 33823 742334
rect 33703 714466 33823 714594
rect 33903 714546 34833 742254
rect 34913 742193 35033 742334
rect 36123 742273 37213 742334
rect 34913 714466 35033 714594
rect 35113 714546 36043 742254
rect 36123 742193 36243 742273
rect 37093 742193 37213 742273
rect 36323 714594 37013 742193
rect 36123 714514 36243 714594
rect 37093 714514 37213 714594
rect 37293 714546 38223 742254
rect 38303 742193 38423 742334
rect 36123 714466 37213 714514
rect 38303 714466 38423 714594
rect 38503 714546 39593 742254
rect 39673 742193 39893 742334
rect 677707 730866 677927 731007
rect 678007 730946 679097 759854
rect 679177 759806 679297 759934
rect 680387 759886 681477 759934
rect 679177 730866 679297 731007
rect 679377 730946 680307 759854
rect 680387 759806 680507 759886
rect 681357 759806 681477 759886
rect 680587 731007 681277 759806
rect 680387 730927 680507 731007
rect 681357 730927 681477 731007
rect 681557 730946 682487 759854
rect 682567 759806 682687 759934
rect 680387 730866 681477 730927
rect 682567 730866 682687 731007
rect 682767 730946 683697 759854
rect 683777 759806 683897 759934
rect 683777 730866 683897 731007
rect 683977 730946 684667 759854
rect 684747 759806 684867 759934
rect 684747 730866 684867 731007
rect 684947 730946 685637 759854
rect 685717 759806 685837 759934
rect 685717 730866 685837 731007
rect 685917 730946 686847 759854
rect 686927 759806 687067 759934
rect 686927 730866 687067 731007
rect 677707 730598 687067 730866
rect 687147 730678 687213 766182
rect 687273 765171 687869 852107
rect 687949 847334 688145 852187
rect 687929 818546 688165 847254
rect 687949 804134 688145 818466
rect 687929 775346 688165 804054
rect 687949 768232 688145 775266
rect 688225 768312 688821 855248
rect 688901 853662 717600 855328
rect 688881 775078 688947 853582
rect 689027 847334 717600 853662
rect 689027 847206 689167 847334
rect 689027 818800 689167 847000
rect 689027 818466 689167 818607
rect 689247 818546 690137 847254
rect 690217 847206 690337 847334
rect 690217 818800 690337 847000
rect 690217 818466 690337 818607
rect 690417 818546 691307 847254
rect 691387 847206 691527 847334
rect 691387 818800 691527 847000
rect 691387 818466 691527 818607
rect 691607 818546 696600 847254
rect 696680 847206 712677 847334
rect 712757 847000 717600 847254
rect 696680 818800 717600 847000
rect 696680 818466 712677 818607
rect 712757 818546 717600 818800
rect 689027 804134 717600 818466
rect 689027 803993 689167 804134
rect 689027 775600 689167 803800
rect 689027 775266 689167 775407
rect 689247 775346 690137 804054
rect 690217 803993 690337 804134
rect 690217 775600 690337 803800
rect 690217 775266 690337 775407
rect 690417 775346 691307 804054
rect 691387 803993 691527 804134
rect 691387 775600 691527 803800
rect 691387 775266 691527 775407
rect 691607 775346 696600 804054
rect 696680 803993 712677 804134
rect 712757 803800 717600 804054
rect 696680 775600 717600 803800
rect 696680 775266 712677 775407
rect 712757 775346 717600 775600
rect 689027 774998 717600 775266
rect 688901 768232 717600 774998
rect 687949 767928 717600 768232
rect 687949 765091 688145 767928
rect 687293 764787 688145 765091
rect 677707 721862 687193 730598
rect 677707 715534 687067 721862
rect 677707 715406 677927 715534
rect 39673 714466 39893 714594
rect 30533 708138 39893 714466
rect 30407 699402 39893 708138
rect 29455 665909 30307 666213
rect 29455 663072 29651 665909
rect 0 662768 29651 663072
rect 0 656002 28699 662768
rect 0 655734 28573 656002
rect 0 655400 4843 655654
rect 4923 655593 20920 655734
rect 0 628200 20920 655400
rect 0 627946 4843 628200
rect 4923 627866 20920 627994
rect 21000 627946 25993 655654
rect 26073 655593 26213 655734
rect 26073 628200 26213 655400
rect 26073 627866 26213 627994
rect 26293 627946 27183 655654
rect 27263 655593 27383 655734
rect 27263 628200 27383 655400
rect 27263 627866 27383 627994
rect 27463 627946 28353 655654
rect 28433 655593 28573 655734
rect 28433 628200 28573 655400
rect 28433 627866 28573 627994
rect 0 621538 28573 627866
rect 28653 621618 28719 655922
rect 0 619872 28699 621538
rect 28779 619952 29375 662688
rect 29455 655734 29651 662768
rect 29435 627946 29671 655654
rect 29455 623013 29651 627866
rect 29731 623093 30327 665829
rect 30387 664818 30453 699322
rect 30533 699134 39893 699402
rect 30533 698993 30673 699134
rect 30533 671066 30673 671194
rect 30753 671146 31683 699054
rect 31763 698993 31883 699134
rect 31763 671066 31883 671194
rect 31963 671146 32653 699054
rect 32733 698993 32853 699134
rect 32733 671066 32853 671194
rect 32933 671146 33623 699054
rect 33703 698993 33823 699134
rect 33703 671066 33823 671194
rect 33903 671146 34833 699054
rect 34913 698993 35033 699134
rect 36123 699073 37213 699134
rect 34913 671066 35033 671194
rect 35113 671146 36043 699054
rect 36123 698993 36243 699073
rect 37093 698993 37213 699073
rect 36323 671194 37013 698993
rect 36123 671114 36243 671194
rect 37093 671114 37213 671194
rect 37293 671146 38223 699054
rect 38303 698993 38423 699134
rect 36123 671066 37213 671114
rect 38303 671066 38423 671194
rect 38503 671146 39593 699054
rect 39673 698993 39893 699134
rect 677707 686666 677927 686807
rect 678007 686746 679097 715454
rect 679177 715406 679297 715534
rect 680387 715486 681477 715534
rect 679177 686666 679297 686807
rect 679377 686746 680307 715454
rect 680387 715406 680507 715486
rect 681357 715406 681477 715486
rect 680587 686807 681277 715406
rect 680387 686727 680507 686807
rect 681357 686727 681477 686807
rect 681557 686746 682487 715454
rect 682567 715406 682687 715534
rect 680387 686666 681477 686727
rect 682567 686666 682687 686807
rect 682767 686746 683697 715454
rect 683777 715406 683897 715534
rect 683777 686666 683897 686807
rect 683977 686746 684667 715454
rect 684747 715406 684867 715534
rect 684747 686666 684867 686807
rect 684947 686746 685637 715454
rect 685717 715406 685837 715534
rect 685717 686666 685837 686807
rect 685917 686746 686847 715454
rect 686927 715406 687067 715534
rect 686927 686666 687067 686807
rect 677707 686398 687067 686666
rect 687147 686478 687213 721782
rect 687273 720771 687869 764707
rect 687949 759934 688145 764787
rect 687929 730946 688165 759854
rect 687949 723832 688145 730866
rect 688225 723912 688821 767848
rect 688901 766262 717600 767928
rect 688881 730678 688947 766182
rect 689027 759934 717600 766262
rect 689027 759806 689167 759934
rect 689027 731200 689167 759600
rect 689027 730866 689167 731007
rect 689247 730946 690137 759854
rect 690217 759806 690337 759934
rect 690217 731200 690337 759600
rect 690217 730866 690337 731007
rect 690417 730946 691307 759854
rect 691387 759806 691527 759934
rect 691387 731200 691527 759600
rect 691387 730866 691527 731007
rect 691607 730946 696600 759854
rect 696680 759806 712677 759934
rect 712757 759600 717600 759854
rect 696680 731200 717600 759600
rect 696680 730866 712677 731007
rect 712757 730946 717600 731200
rect 689027 730598 717600 730866
rect 688901 723832 717600 730598
rect 687949 723528 717600 723832
rect 687949 720691 688145 723528
rect 687293 720387 688145 720691
rect 677707 677662 687193 686398
rect 677707 671334 687067 677662
rect 677707 671206 677927 671334
rect 39673 671066 39893 671194
rect 30533 664738 39893 671066
rect 30407 656002 39893 664738
rect 29455 622709 30307 623013
rect 29455 619872 29651 622709
rect 0 619568 29651 619872
rect 0 612802 28699 619568
rect 0 612534 28573 612802
rect 0 612200 4843 612454
rect 4923 612393 20920 612534
rect 0 585000 20920 612200
rect 0 584746 4843 585000
rect 4923 584666 20920 584794
rect 21000 584746 25993 612454
rect 26073 612393 26213 612534
rect 26073 585000 26213 612200
rect 26073 584666 26213 584794
rect 26293 584746 27183 612454
rect 27263 612393 27383 612534
rect 27263 585000 27383 612200
rect 27263 584666 27383 584794
rect 27463 584746 28353 612454
rect 28433 612393 28573 612534
rect 28433 585000 28573 612200
rect 28433 584666 28573 584794
rect 0 578338 28573 584666
rect 28653 578418 28719 612722
rect 0 576672 28699 578338
rect 28779 576752 29375 619488
rect 29455 612534 29651 619568
rect 29435 584746 29671 612454
rect 29455 579813 29651 584666
rect 29731 579893 30327 622629
rect 30387 621618 30453 655922
rect 30533 655734 39893 656002
rect 30533 655593 30673 655734
rect 30533 627866 30673 627994
rect 30753 627946 31683 655654
rect 31763 655593 31883 655734
rect 31763 627866 31883 627994
rect 31963 627946 32653 655654
rect 32733 655593 32853 655734
rect 32733 627866 32853 627994
rect 32933 627946 33623 655654
rect 33703 655593 33823 655734
rect 33703 627866 33823 627994
rect 33903 627946 34833 655654
rect 34913 655593 35033 655734
rect 36123 655673 37213 655734
rect 34913 627866 35033 627994
rect 35113 627946 36043 655654
rect 36123 655593 36243 655673
rect 37093 655593 37213 655673
rect 36323 627994 37013 655593
rect 36123 627914 36243 627994
rect 37093 627914 37213 627994
rect 37293 627946 38223 655654
rect 38303 655593 38423 655734
rect 36123 627866 37213 627914
rect 38303 627866 38423 627994
rect 38503 627946 39593 655654
rect 39673 655593 39893 655734
rect 677707 642466 677927 642607
rect 678007 642546 679097 671254
rect 679177 671206 679297 671334
rect 680387 671286 681477 671334
rect 679177 642466 679297 642607
rect 679377 642546 680307 671254
rect 680387 671206 680507 671286
rect 681357 671206 681477 671286
rect 680587 642607 681277 671206
rect 680387 642527 680507 642607
rect 681357 642527 681477 642607
rect 681557 642546 682487 671254
rect 682567 671206 682687 671334
rect 680387 642466 681477 642527
rect 682567 642466 682687 642607
rect 682767 642546 683697 671254
rect 683777 671206 683897 671334
rect 683777 642466 683897 642607
rect 683977 642546 684667 671254
rect 684747 671206 684867 671334
rect 684747 642466 684867 642607
rect 684947 642546 685637 671254
rect 685717 671206 685837 671334
rect 685717 642466 685837 642607
rect 685917 642546 686847 671254
rect 686927 671206 687067 671334
rect 686927 642466 687067 642607
rect 677707 642198 687067 642466
rect 687147 642278 687213 677582
rect 687273 676571 687869 720307
rect 687949 715534 688145 720387
rect 687929 686746 688165 715454
rect 687949 679632 688145 686666
rect 688225 679712 688821 723448
rect 688901 721862 717600 723528
rect 688881 686478 688947 721782
rect 689027 715534 717600 721862
rect 689027 715406 689167 715534
rect 689027 687000 689167 715200
rect 689027 686666 689167 686807
rect 689247 686746 690137 715454
rect 690217 715406 690337 715534
rect 690217 687000 690337 715200
rect 690217 686666 690337 686807
rect 690417 686746 691307 715454
rect 691387 715406 691527 715534
rect 691387 687000 691527 715200
rect 691387 686666 691527 686807
rect 691607 686746 696600 715454
rect 696680 715406 712677 715534
rect 712757 715200 717600 715454
rect 696680 687000 717600 715200
rect 696680 686666 712677 686807
rect 712757 686746 717600 687000
rect 689027 686398 717600 686666
rect 688901 679632 717600 686398
rect 687949 679328 717600 679632
rect 687949 676491 688145 679328
rect 687293 676187 688145 676491
rect 677707 633462 687193 642198
rect 39673 627866 39893 627994
rect 30533 621538 39893 627866
rect 677707 627134 687067 633462
rect 677707 627006 677927 627134
rect 30407 612802 39893 621538
rect 29455 579509 30307 579813
rect 29455 576672 29651 579509
rect 0 576368 29651 576672
rect 0 569602 28699 576368
rect 0 569334 28573 569602
rect 0 569000 4843 569254
rect 4923 569193 20920 569334
rect 0 541800 20920 569000
rect 0 541546 4843 541800
rect 4923 541466 20920 541594
rect 21000 541546 25993 569254
rect 26073 569193 26213 569334
rect 26073 541800 26213 569000
rect 26073 541466 26213 541594
rect 26293 541546 27183 569254
rect 27263 569193 27383 569334
rect 27263 541800 27383 569000
rect 27263 541466 27383 541594
rect 27463 541546 28353 569254
rect 28433 569193 28573 569334
rect 28433 541800 28573 569000
rect 28433 541466 28573 541594
rect 0 535138 28573 541466
rect 28653 535218 28719 569522
rect 0 533472 28699 535138
rect 28779 533552 29375 576288
rect 29455 569334 29651 576368
rect 29435 541546 29671 569254
rect 29455 536613 29651 541466
rect 29731 536693 30327 579429
rect 30387 578418 30453 612722
rect 30533 612534 39893 612802
rect 30533 612393 30673 612534
rect 30533 584666 30673 584794
rect 30753 584746 31683 612454
rect 31763 612393 31883 612534
rect 31763 584666 31883 584794
rect 31963 584746 32653 612454
rect 32733 612393 32853 612534
rect 32733 584666 32853 584794
rect 32933 584746 33623 612454
rect 33703 612393 33823 612534
rect 33703 584666 33823 584794
rect 33903 584746 34833 612454
rect 34913 612393 35033 612534
rect 36123 612473 37213 612534
rect 34913 584666 35033 584794
rect 35113 584746 36043 612454
rect 36123 612393 36243 612473
rect 37093 612393 37213 612473
rect 36323 584794 37013 612393
rect 36123 584714 36243 584794
rect 37093 584714 37213 584794
rect 37293 584746 38223 612454
rect 38303 612393 38423 612534
rect 36123 584666 37213 584714
rect 38303 584666 38423 584794
rect 38503 584746 39593 612454
rect 39673 612393 39893 612534
rect 677707 598066 677927 598207
rect 678007 598146 679097 627054
rect 679177 627006 679297 627134
rect 680387 627086 681477 627134
rect 679177 598066 679297 598207
rect 679377 598146 680307 627054
rect 680387 627006 680507 627086
rect 681357 627006 681477 627086
rect 680587 598207 681277 627006
rect 680387 598127 680507 598207
rect 681357 598127 681477 598207
rect 681557 598146 682487 627054
rect 682567 627006 682687 627134
rect 680387 598066 681477 598127
rect 682567 598066 682687 598207
rect 682767 598146 683697 627054
rect 683777 627006 683897 627134
rect 683777 598066 683897 598207
rect 683977 598146 684667 627054
rect 684747 627006 684867 627134
rect 684747 598066 684867 598207
rect 684947 598146 685637 627054
rect 685717 627006 685837 627134
rect 685717 598066 685837 598207
rect 685917 598146 686847 627054
rect 686927 627006 687067 627134
rect 686927 598066 687067 598207
rect 677707 597798 687067 598066
rect 687147 597878 687213 633382
rect 687273 632371 687869 676107
rect 687949 671334 688145 676187
rect 687929 642546 688165 671254
rect 687949 635432 688145 642466
rect 688225 635512 688821 679248
rect 688901 677662 717600 679328
rect 688881 642278 688947 677582
rect 689027 671334 717600 677662
rect 689027 671206 689167 671334
rect 689027 642800 689167 671000
rect 689027 642466 689167 642607
rect 689247 642546 690137 671254
rect 690217 671206 690337 671334
rect 690217 642800 690337 671000
rect 690217 642466 690337 642607
rect 690417 642546 691307 671254
rect 691387 671206 691527 671334
rect 691387 642800 691527 671000
rect 691387 642466 691527 642607
rect 691607 642546 696600 671254
rect 696680 671206 712677 671334
rect 712757 671000 717600 671254
rect 696680 642800 717600 671000
rect 696680 642466 712677 642607
rect 712757 642546 717600 642800
rect 689027 642198 717600 642466
rect 688901 635432 717600 642198
rect 687949 635128 717600 635432
rect 687949 632291 688145 635128
rect 687293 631987 688145 632291
rect 677707 589062 687193 597798
rect 39673 584666 39893 584794
rect 30533 578338 39893 584666
rect 677707 582734 687067 589062
rect 677707 582606 677927 582734
rect 30407 569602 39893 578338
rect 29455 536309 30307 536613
rect 29455 533472 29651 536309
rect 0 533168 29651 533472
rect 0 526402 28699 533168
rect 0 526134 28573 526402
rect 0 525800 4843 526054
rect 4923 525993 20920 526134
rect 0 498400 20920 525800
rect 0 498146 4843 498400
rect 4923 498066 20920 498207
rect 21000 498146 25993 526054
rect 26073 525993 26213 526134
rect 26073 498400 26213 525800
rect 26073 498066 26213 498207
rect 26293 498146 27183 526054
rect 27263 525993 27383 526134
rect 27263 498400 27383 525800
rect 27263 498066 27383 498207
rect 27463 498146 28353 526054
rect 28433 525993 28573 526134
rect 28433 498400 28573 525800
rect 28433 498066 28573 498207
rect 0 483734 28573 498066
rect 0 483400 4843 483654
rect 4923 483593 20920 483734
rect 0 456493 20920 483400
rect 0 456200 7 456493
rect 4843 456200 20920 456493
rect 4843 456157 4850 456200
rect 4923 455866 20920 456200
rect 21000 455946 25993 483654
rect 26073 483593 26213 483734
rect 26073 455866 26213 483400
rect 26293 455946 27183 483654
rect 27263 483593 27383 483734
rect 27263 455866 27383 483400
rect 27463 455946 28353 483654
rect 28433 483593 28573 483734
rect 28433 455866 28573 483400
rect 0 441534 28573 455866
rect 0 441200 4843 441454
rect 4923 441200 20920 441534
rect 0 414000 20920 441200
rect 0 413746 4843 414000
rect 4923 413666 20920 413794
rect 21000 413746 25993 441454
rect 26073 414000 26213 441534
rect 26073 413666 26213 413794
rect 26293 413746 27183 441454
rect 27263 414000 27383 441534
rect 27263 413666 27383 413794
rect 27463 413746 28353 441454
rect 28433 414000 28573 441534
rect 28433 413666 28573 413794
rect 0 407338 28573 413666
rect 0 405672 28699 407338
rect 28779 405752 29375 533088
rect 29455 526134 29651 533168
rect 29435 498146 29671 526054
rect 29455 483734 29651 498066
rect 29435 455946 29671 483654
rect 29455 441534 29651 455866
rect 29435 413746 29671 441454
rect 29455 408813 29651 413666
rect 29731 408893 30327 536229
rect 30387 535218 30453 569522
rect 30533 569334 39893 569602
rect 30533 569193 30673 569334
rect 30533 541466 30673 541594
rect 30753 541546 31683 569254
rect 31763 569193 31883 569334
rect 31763 541466 31883 541594
rect 31963 541546 32653 569254
rect 32733 569193 32853 569334
rect 32733 541466 32853 541594
rect 32933 541546 33623 569254
rect 33703 569193 33823 569334
rect 33703 541466 33823 541594
rect 33903 541546 34833 569254
rect 34913 569193 35033 569334
rect 36123 569273 37213 569334
rect 34913 541466 35033 541594
rect 35113 541546 36043 569254
rect 36123 569193 36243 569273
rect 37093 569193 37213 569273
rect 36323 541594 37013 569193
rect 36123 541514 36243 541594
rect 37093 541514 37213 541594
rect 37293 541546 38223 569254
rect 38303 569193 38423 569334
rect 36123 541466 37213 541514
rect 38303 541466 38423 541594
rect 38503 541546 39593 569254
rect 39673 569193 39893 569334
rect 677707 553866 677927 554007
rect 678007 553946 679097 582654
rect 679177 582606 679297 582734
rect 680387 582686 681477 582734
rect 679177 553866 679297 554007
rect 679377 553946 680307 582654
rect 680387 582606 680507 582686
rect 681357 582606 681477 582686
rect 680587 554007 681277 582606
rect 680387 553927 680507 554007
rect 681357 553927 681477 554007
rect 681557 553946 682487 582654
rect 682567 582606 682687 582734
rect 680387 553866 681477 553927
rect 682567 553866 682687 554007
rect 682767 553946 683697 582654
rect 683777 582606 683897 582734
rect 683777 553866 683897 554007
rect 683977 553946 684667 582654
rect 684747 582606 684867 582734
rect 684747 553866 684867 554007
rect 684947 553946 685637 582654
rect 685717 582606 685837 582734
rect 685717 553866 685837 554007
rect 685917 553946 686847 582654
rect 686927 582606 687067 582734
rect 686927 553866 687067 554007
rect 677707 553598 687067 553866
rect 687147 553678 687213 588982
rect 687273 587971 687869 631907
rect 687949 627134 688145 631987
rect 687929 598146 688165 627054
rect 687949 591032 688145 598066
rect 688225 591112 688821 635048
rect 688901 633462 717600 635128
rect 688881 597878 688947 633382
rect 689027 627134 717600 633462
rect 689027 627006 689167 627134
rect 689027 598400 689167 626800
rect 689027 598066 689167 598207
rect 689247 598146 690137 627054
rect 690217 627006 690337 627134
rect 690217 598400 690337 626800
rect 690217 598066 690337 598207
rect 690417 598146 691307 627054
rect 691387 627006 691527 627134
rect 691387 598400 691527 626800
rect 691387 598066 691527 598207
rect 691607 598146 696600 627054
rect 696680 627006 712677 627134
rect 712757 626800 717600 627054
rect 696680 598400 717600 626800
rect 696680 598066 712677 598207
rect 712757 598146 717600 598400
rect 689027 597798 717600 598066
rect 688901 591032 717600 597798
rect 687949 590728 717600 591032
rect 687949 587891 688145 590728
rect 687293 587587 688145 587891
rect 677707 544862 687193 553598
rect 39673 541466 39893 541594
rect 30533 535138 39893 541466
rect 677707 538534 687067 544862
rect 677707 538406 677927 538534
rect 30407 526402 39893 535138
rect 29455 408509 30307 408813
rect 29455 405672 29651 408509
rect 0 405368 29651 405672
rect 0 398602 28699 405368
rect 0 398334 28573 398602
rect 0 398000 4843 398254
rect 4923 398193 20920 398334
rect 0 370800 20920 398000
rect 0 370546 4843 370800
rect 4923 370466 20920 370594
rect 21000 370546 25993 398254
rect 26073 398193 26213 398334
rect 26073 370800 26213 398000
rect 26073 370466 26213 370594
rect 26293 370546 27183 398254
rect 27263 398193 27383 398334
rect 27263 370800 27383 398000
rect 27263 370466 27383 370594
rect 27463 370546 28353 398254
rect 28433 398193 28573 398334
rect 28433 370800 28573 398000
rect 28433 370466 28573 370594
rect 0 364138 28573 370466
rect 28653 364218 28719 398522
rect 0 362472 28699 364138
rect 28779 362552 29375 405288
rect 29455 398334 29651 405368
rect 29435 370546 29671 398254
rect 29455 365613 29651 370466
rect 29731 365693 30327 408429
rect 30387 407418 30453 526322
rect 30533 526134 39893 526402
rect 30533 525993 30673 526134
rect 30533 498066 30673 498207
rect 30753 498146 31683 526054
rect 31763 525993 31883 526134
rect 31763 498066 31883 498207
rect 31963 498146 32653 526054
rect 32733 525993 32853 526134
rect 32733 498066 32853 498207
rect 32933 498146 33623 526054
rect 33703 525993 33823 526134
rect 33703 498066 33823 498207
rect 33903 498146 34833 526054
rect 34913 525993 35033 526134
rect 36123 526073 37213 526134
rect 34913 498066 35033 498207
rect 35113 498146 36043 526054
rect 36123 525993 36243 526073
rect 37093 525993 37213 526073
rect 36323 498207 37013 525993
rect 36123 498127 36243 498207
rect 37093 498127 37213 498207
rect 37293 498146 38223 526054
rect 38303 525993 38423 526134
rect 36123 498066 37213 498127
rect 38303 498066 38423 498207
rect 38503 498146 39593 526054
rect 39673 525993 39893 526134
rect 678007 509746 679097 538454
rect 679177 538406 679297 538534
rect 680387 538486 681477 538534
rect 679177 509666 679297 509807
rect 679377 509746 680307 538454
rect 680387 538406 680507 538486
rect 681357 538406 681477 538486
rect 680587 509807 681277 538406
rect 680387 509727 680507 509807
rect 681357 509727 681477 509807
rect 681557 509746 682487 538454
rect 682567 538406 682687 538534
rect 680387 509666 681477 509727
rect 682567 509666 682687 509807
rect 682767 509746 683697 538454
rect 683777 538406 683897 538534
rect 683777 509666 683897 509807
rect 683977 509746 684667 538454
rect 684747 538406 684867 538534
rect 684747 509666 684867 509807
rect 684947 509746 685637 538454
rect 685717 538406 685837 538534
rect 685717 509666 685837 509807
rect 685917 509746 686847 538454
rect 686927 538406 687067 538534
rect 686927 509666 687067 509807
rect 30533 483734 39593 498066
rect 678007 495334 687067 509666
rect 30533 483593 30673 483734
rect 30533 455866 30673 456200
rect 30753 455946 31683 483654
rect 31763 483593 31883 483734
rect 31763 455866 31883 456200
rect 31963 455946 32653 483654
rect 32733 483593 32853 483734
rect 32733 455866 32853 456200
rect 33703 483593 33823 483734
rect 33903 458387 34833 483654
rect 34913 483593 35033 483734
rect 36123 483673 37213 483734
rect 33703 455866 33823 456200
rect 33903 456187 34840 458387
rect 33903 455946 34833 456187
rect 34913 455866 35033 456200
rect 35113 455946 36043 483654
rect 36123 483593 36243 483673
rect 37093 483593 37213 483673
rect 36123 455927 36243 456200
rect 37093 455927 37213 456200
rect 38303 483593 38423 483734
rect 36123 455866 37213 455927
rect 38303 455866 38423 456200
rect 678007 466346 679097 495254
rect 679177 495193 679297 495334
rect 680387 495273 681477 495334
rect 679177 466266 679297 466600
rect 679377 466346 680307 495254
rect 680387 495193 680507 495273
rect 681357 495193 681477 495273
rect 680387 466327 680507 466600
rect 680587 466407 681277 495193
rect 681357 466327 681477 466600
rect 681557 466346 682487 495254
rect 682567 495193 682687 495334
rect 680387 466266 681477 466327
rect 682567 466266 682687 466600
rect 682767 466346 683697 495254
rect 683777 495193 683897 495334
rect 683777 466266 683897 466600
rect 683977 466346 684667 495254
rect 684747 495193 684867 495334
rect 684747 466266 684867 466600
rect 684947 466346 685637 495254
rect 685717 495193 685837 495334
rect 685917 468795 686847 495254
rect 686927 495193 687067 495334
rect 685717 466266 685837 466600
rect 685910 466586 686847 468795
rect 685917 466346 686847 466586
rect 686927 466266 687067 466600
rect 30533 441534 39593 455866
rect 678007 451934 687067 466266
rect 30533 441200 30673 441534
rect 30753 441214 31683 441454
rect 30753 439005 31690 441214
rect 31763 441200 31883 441534
rect 30533 413666 30673 413794
rect 30753 413746 31683 439005
rect 31763 413666 31883 413794
rect 31963 413746 32653 441454
rect 32733 441200 32853 441534
rect 32733 413666 32853 413794
rect 32933 413746 33623 441454
rect 33703 441200 33823 441534
rect 33703 413666 33823 413794
rect 33903 413746 34833 441454
rect 34913 441200 35033 441534
rect 36123 441473 37213 441534
rect 34913 413666 35033 413794
rect 35113 413746 36043 441454
rect 36123 441200 36243 441473
rect 36323 413794 37013 441393
rect 37093 441200 37213 441473
rect 36123 413714 36243 413794
rect 37093 413714 37213 413794
rect 37293 413746 38223 441454
rect 38303 441200 38423 441534
rect 36123 413666 37213 413714
rect 38303 413666 38423 413794
rect 38503 413746 39593 441454
rect 678007 423146 679097 451854
rect 679177 451600 679297 451934
rect 680387 451873 681477 451934
rect 679177 423066 679297 423207
rect 680387 451600 680507 451873
rect 681357 451600 681477 451873
rect 680387 423127 680507 423207
rect 681357 423127 681477 423207
rect 681557 423146 682487 451854
rect 682567 451600 682687 451934
rect 682767 451613 683697 451854
rect 682760 449413 683697 451613
rect 683777 451600 683897 451934
rect 680387 423066 681477 423127
rect 682567 423066 682687 423207
rect 682767 423146 683697 449413
rect 683777 423066 683897 423207
rect 683977 423146 684667 451854
rect 684747 451600 684867 451934
rect 684747 423066 684867 423207
rect 684947 423146 685637 451854
rect 685717 451600 685837 451934
rect 685717 423066 685837 423207
rect 685917 423146 686847 451854
rect 686927 451600 687067 451934
rect 686927 423066 687067 423207
rect 687147 423146 687213 544782
rect 687273 543771 687869 587507
rect 687949 582734 688145 587587
rect 687929 553946 688165 582654
rect 687949 546832 688145 553866
rect 688225 546912 688821 590648
rect 688901 589062 717600 590728
rect 688881 553678 688947 588982
rect 689027 582734 717600 589062
rect 689027 582606 689167 582734
rect 689027 554200 689167 582400
rect 689027 553866 689167 554007
rect 689247 553946 690137 582654
rect 690217 582606 690337 582734
rect 690217 554200 690337 582400
rect 690217 553866 690337 554007
rect 690417 553946 691307 582654
rect 691387 582606 691527 582734
rect 691387 554200 691527 582400
rect 691387 553866 691527 554007
rect 691607 553946 696600 582654
rect 696680 582606 712677 582734
rect 712757 582400 717600 582654
rect 696680 554200 717600 582400
rect 696680 553866 712677 554007
rect 712757 553946 717600 554200
rect 689027 553598 717600 553866
rect 688901 546832 717600 553598
rect 687949 546528 717600 546832
rect 687949 543691 688145 546528
rect 687293 543387 688145 543691
rect 673867 419930 673933 419933
rect 673867 419870 674114 419930
rect 673867 419867 673933 419870
rect 673867 419250 673933 419253
rect 674054 419250 674114 419870
rect 673867 419190 674114 419250
rect 673867 419187 673933 419190
rect 39673 413666 39893 413794
rect 30533 407338 39893 413666
rect 678007 408734 687193 423066
rect 30407 398602 39893 407338
rect 29455 365309 30307 365613
rect 29455 362472 29651 365309
rect 0 362168 29651 362472
rect 0 355402 28699 362168
rect 0 355134 28573 355402
rect 0 354800 4843 355054
rect 4923 354993 20920 355134
rect 0 327400 20920 354800
rect 0 327146 4843 327400
rect 4923 327066 20920 327194
rect 21000 327146 25993 355054
rect 26073 354993 26213 355134
rect 26073 327400 26213 354800
rect 26073 327066 26213 327194
rect 26293 327146 27183 355054
rect 27263 354993 27383 355134
rect 27263 327400 27383 354800
rect 27263 327066 27383 327194
rect 27463 327146 28353 355054
rect 28433 354993 28573 355134
rect 28433 327400 28573 354800
rect 28433 327066 28573 327194
rect 0 320738 28573 327066
rect 28653 320818 28719 355322
rect 0 319072 28699 320738
rect 28779 319152 29375 362088
rect 29455 355134 29651 362168
rect 29435 327146 29671 355054
rect 29455 322213 29651 327066
rect 29731 322293 30327 365229
rect 30387 364218 30453 398522
rect 30533 398334 39893 398602
rect 30533 398193 30673 398334
rect 30533 370466 30673 370594
rect 30753 370546 31683 398254
rect 31763 398193 31883 398334
rect 31763 370466 31883 370594
rect 31963 370546 32653 398254
rect 32733 398193 32853 398334
rect 32733 370466 32853 370594
rect 32933 370546 33623 398254
rect 33703 398193 33823 398334
rect 33703 370466 33823 370594
rect 33903 370546 34833 398254
rect 34913 398193 35033 398334
rect 36123 398273 37213 398334
rect 34913 370466 35033 370594
rect 35113 370546 36043 398254
rect 36123 398193 36243 398273
rect 37093 398193 37213 398273
rect 36323 370594 37013 398193
rect 36123 370514 36243 370594
rect 37093 370514 37213 370594
rect 37293 370546 38223 398254
rect 38303 398193 38423 398334
rect 36123 370466 37213 370514
rect 38303 370466 38423 370594
rect 38503 370546 39593 398254
rect 39673 398193 39893 398334
rect 677707 379666 677927 379807
rect 678007 379746 679097 408654
rect 679177 408593 679297 408734
rect 680387 408673 681477 408734
rect 679177 379666 679297 379807
rect 679377 379746 680307 408654
rect 680387 408593 680507 408673
rect 681357 408593 681477 408673
rect 680587 379807 681277 408593
rect 680387 379727 680507 379807
rect 681357 379727 681477 379807
rect 681557 379746 682487 408654
rect 682567 408593 682687 408734
rect 680387 379666 681477 379727
rect 682567 379666 682687 379807
rect 682767 379746 683697 408654
rect 683777 408593 683897 408734
rect 683777 379666 683897 379807
rect 683977 379746 684667 408654
rect 684747 408593 684867 408734
rect 684747 379666 684867 379807
rect 684947 379746 685637 408654
rect 685717 408593 685837 408734
rect 685717 379666 685837 379807
rect 685917 379746 686847 408654
rect 686927 408593 687067 408734
rect 686927 379666 687067 379807
rect 677707 379398 687067 379666
rect 687147 379478 687213 408654
rect 677707 370662 687193 379398
rect 39673 370466 39893 370594
rect 30533 364138 39893 370466
rect 677707 364334 687067 370662
rect 677707 364206 677927 364334
rect 30407 355402 39893 364138
rect 29455 321909 30307 322213
rect 29455 319072 29651 321909
rect 0 318768 29651 319072
rect 0 312002 28699 318768
rect 0 311734 28573 312002
rect 0 311400 4843 311654
rect 4923 311593 20920 311734
rect 0 284200 20920 311400
rect 0 283946 4843 284200
rect 4923 283866 20920 283994
rect 21000 283946 25993 311654
rect 26073 311593 26213 311734
rect 26073 284200 26213 311400
rect 26073 283866 26213 283994
rect 26293 283946 27183 311654
rect 27263 311593 27383 311734
rect 27263 284200 27383 311400
rect 27263 283866 27383 283994
rect 27463 283946 28353 311654
rect 28433 311593 28573 311734
rect 28433 284200 28573 311400
rect 28433 283866 28573 283994
rect 0 277538 28573 283866
rect 28653 277618 28719 311922
rect 0 275872 28699 277538
rect 28779 275952 29375 318688
rect 29455 311734 29651 318768
rect 29435 283946 29671 311654
rect 29455 279013 29651 283866
rect 29731 279093 30327 321829
rect 30387 320818 30453 355322
rect 30533 355134 39893 355402
rect 30533 354993 30673 355134
rect 30533 327066 30673 327194
rect 30753 327146 31683 355054
rect 31763 354993 31883 355134
rect 31763 327066 31883 327194
rect 31963 327146 32653 355054
rect 32733 354993 32853 355134
rect 32733 327066 32853 327194
rect 32933 327146 33623 355054
rect 33703 354993 33823 355134
rect 33703 327066 33823 327194
rect 33903 327146 34833 355054
rect 34913 354993 35033 355134
rect 36123 355073 37213 355134
rect 34913 327066 35033 327194
rect 35113 327146 36043 355054
rect 36123 354993 36243 355073
rect 37093 354993 37213 355073
rect 36323 327194 37013 354993
rect 36123 327114 36243 327194
rect 37093 327114 37213 327194
rect 37293 327146 38223 355054
rect 38303 354993 38423 355134
rect 36123 327066 37213 327114
rect 38303 327066 38423 327194
rect 38503 327146 39593 355054
rect 39673 354993 39893 355134
rect 677707 335466 677927 335607
rect 678007 335546 679097 364254
rect 679177 364206 679297 364334
rect 680387 364286 681477 364334
rect 679177 335466 679297 335607
rect 679377 335546 680307 364254
rect 680387 364206 680507 364286
rect 681357 364206 681477 364286
rect 680587 335607 681277 364206
rect 680387 335527 680507 335607
rect 681357 335527 681477 335607
rect 681557 335546 682487 364254
rect 682567 364206 682687 364334
rect 680387 335466 681477 335527
rect 682567 335466 682687 335607
rect 682767 335546 683697 364254
rect 683777 364206 683897 364334
rect 683777 335466 683897 335607
rect 683977 335546 684667 364254
rect 684747 364206 684867 364334
rect 684747 335466 684867 335607
rect 684947 335546 685637 364254
rect 685717 364206 685837 364334
rect 685717 335466 685837 335607
rect 685917 335546 686847 364254
rect 686927 364206 687067 364334
rect 686927 335466 687067 335607
rect 677707 335198 687067 335466
rect 687147 335278 687213 370582
rect 687273 369571 687869 543307
rect 687949 538534 688145 543387
rect 687929 509746 688165 538454
rect 687949 495334 688145 509666
rect 687929 466346 688165 495254
rect 687949 451934 688145 466266
rect 687929 423146 688165 451854
rect 687949 408734 688145 423066
rect 687929 379746 688165 408654
rect 687949 372632 688145 379666
rect 688225 372712 688821 546448
rect 688901 544862 717600 546528
rect 689027 538534 717600 544862
rect 689027 538406 689167 538534
rect 689027 510000 689167 538200
rect 689027 509666 689167 509807
rect 689247 509746 690137 538454
rect 690217 538406 690337 538534
rect 690217 510000 690337 538200
rect 690217 509666 690337 509807
rect 690417 509746 691307 538454
rect 691387 538406 691527 538534
rect 691387 510000 691527 538200
rect 691387 509666 691527 509807
rect 691607 509746 696600 538454
rect 696680 538406 712677 538534
rect 712757 538200 717600 538454
rect 696680 510000 717600 538200
rect 696680 509666 712677 509807
rect 712757 509746 717600 510000
rect 689027 495334 717600 509666
rect 689027 495193 689167 495334
rect 689027 466266 689167 495000
rect 689247 466346 690137 495254
rect 690217 495193 690337 495334
rect 690217 466266 690337 495000
rect 690417 466346 691307 495254
rect 691387 495193 691527 495334
rect 691387 466266 691527 495000
rect 691607 466346 696600 495254
rect 696680 495193 712677 495334
rect 712757 495000 717600 495254
rect 696680 466600 717600 495000
rect 696680 466266 712677 466600
rect 712757 466346 717600 466600
rect 689027 451934 717600 466266
rect 689027 423400 689167 451934
rect 689027 423066 689167 423207
rect 689247 423146 690137 451854
rect 690217 423400 690337 451934
rect 690217 423066 690337 423207
rect 690417 423146 691307 451854
rect 691387 423400 691527 451934
rect 691387 423066 691527 423207
rect 691607 423146 696600 451854
rect 696680 451600 712677 451934
rect 712757 451643 717600 451854
rect 712750 451600 717600 451643
rect 696680 423400 717600 451600
rect 696680 423066 712677 423207
rect 712757 423146 717600 423400
rect 688901 408734 717600 423066
rect 688881 379478 688947 408654
rect 689027 408593 689167 408734
rect 689027 380000 689167 408400
rect 689027 379666 689167 379807
rect 689247 379746 690137 408654
rect 690217 408593 690337 408734
rect 690217 380000 690337 408400
rect 690217 379666 690337 379807
rect 690417 379746 691307 408654
rect 691387 408593 691527 408734
rect 691387 380000 691527 408400
rect 691387 379666 691527 379807
rect 691607 379746 696600 408654
rect 696680 408593 712677 408734
rect 712757 408400 717600 408654
rect 696680 380000 717600 408400
rect 696680 379666 712677 379807
rect 712757 379746 717600 380000
rect 689027 379398 717600 379666
rect 688901 372632 717600 379398
rect 687949 372328 717600 372632
rect 687949 369491 688145 372328
rect 687293 369187 688145 369491
rect 39673 327066 39893 327194
rect 30533 320738 39893 327066
rect 30407 312002 39893 320738
rect 677707 326462 687193 335198
rect 677707 320134 687067 326462
rect 677707 320006 677927 320134
rect 29455 278709 30307 279013
rect 29455 275872 29651 278709
rect 0 275568 29651 275872
rect 0 268802 28699 275568
rect 0 268534 28573 268802
rect 0 268200 4843 268454
rect 4923 268393 20920 268534
rect 0 241000 20920 268200
rect 0 240746 4843 241000
rect 4923 240666 20920 240794
rect 21000 240746 25993 268454
rect 26073 268393 26213 268534
rect 26073 241000 26213 268200
rect 26073 240666 26213 240794
rect 26293 240746 27183 268454
rect 27263 268393 27383 268534
rect 27263 241000 27383 268200
rect 27263 240666 27383 240794
rect 27463 240746 28353 268454
rect 28433 268393 28573 268534
rect 28433 241000 28573 268200
rect 28433 240666 28573 240794
rect 0 234338 28573 240666
rect 28653 234418 28719 268722
rect 0 232672 28699 234338
rect 28779 232752 29375 275488
rect 29455 268534 29651 275568
rect 29435 240746 29671 268454
rect 29455 235813 29651 240666
rect 29731 235893 30327 278629
rect 30387 277618 30453 311922
rect 30533 311734 39893 312002
rect 30533 311593 30673 311734
rect 30533 283866 30673 283994
rect 30753 283946 31683 311654
rect 31763 311593 31883 311734
rect 31763 283866 31883 283994
rect 31963 283946 32653 311654
rect 32733 311593 32853 311734
rect 32733 283866 32853 283994
rect 32933 283946 33623 311654
rect 33703 311593 33823 311734
rect 33703 283866 33823 283994
rect 33903 283946 34833 311654
rect 34913 311593 35033 311734
rect 36123 311673 37213 311734
rect 34913 283866 35033 283994
rect 35113 283946 36043 311654
rect 36123 311593 36243 311673
rect 37093 311593 37213 311673
rect 36323 283994 37013 311593
rect 36123 283914 36243 283994
rect 37093 283914 37213 283994
rect 37293 283946 38223 311654
rect 38303 311593 38423 311734
rect 36123 283866 37213 283914
rect 38303 283866 38423 283994
rect 38503 283946 39593 311654
rect 39673 311593 39893 311734
rect 677707 291266 677927 291407
rect 678007 291346 679097 320054
rect 679177 320006 679297 320134
rect 680387 320086 681477 320134
rect 679177 291266 679297 291407
rect 679377 291346 680307 320054
rect 680387 320006 680507 320086
rect 681357 320006 681477 320086
rect 680587 291407 681277 320006
rect 680387 291327 680507 291407
rect 681357 291327 681477 291407
rect 681557 291346 682487 320054
rect 682567 320006 682687 320134
rect 680387 291266 681477 291327
rect 682567 291266 682687 291407
rect 682767 291346 683697 320054
rect 683777 320006 683897 320134
rect 683777 291266 683897 291407
rect 683977 291346 684667 320054
rect 684747 320006 684867 320134
rect 684747 291266 684867 291407
rect 684947 291346 685637 320054
rect 685717 320006 685837 320134
rect 685717 291266 685837 291407
rect 685917 291346 686847 320054
rect 686927 320006 687067 320134
rect 686927 291266 687067 291407
rect 677707 290998 687067 291266
rect 687147 291078 687213 326382
rect 687273 325371 687869 369107
rect 687949 364334 688145 369187
rect 687929 335546 688165 364254
rect 687949 328432 688145 335466
rect 688225 328512 688821 372248
rect 688901 370662 717600 372328
rect 688881 335278 688947 370582
rect 689027 364334 717600 370662
rect 689027 364206 689167 364334
rect 689027 335800 689167 364000
rect 689027 335466 689167 335607
rect 689247 335546 690137 364254
rect 690217 364206 690337 364334
rect 690217 335800 690337 364000
rect 690217 335466 690337 335607
rect 690417 335546 691307 364254
rect 691387 364206 691527 364334
rect 691387 335800 691527 364000
rect 691387 335466 691527 335607
rect 691607 335546 696600 364254
rect 696680 364206 712677 364334
rect 712757 364000 717600 364254
rect 696680 335800 717600 364000
rect 696680 335466 712677 335607
rect 712757 335546 717600 335800
rect 689027 335198 717600 335466
rect 688901 328432 717600 335198
rect 687949 328128 717600 328432
rect 687949 325291 688145 328128
rect 687293 324987 688145 325291
rect 39673 283866 39893 283994
rect 30533 277538 39893 283866
rect 30407 268802 39893 277538
rect 677707 282262 687193 290998
rect 677707 275934 687067 282262
rect 677707 275806 677927 275934
rect 29455 235509 30307 235813
rect 29455 232672 29651 235509
rect 0 232368 29651 232672
rect 0 225602 28699 232368
rect 0 225334 28573 225602
rect 0 225000 4843 225254
rect 4923 225193 20920 225334
rect 0 197800 20920 225000
rect 0 197546 4843 197800
rect 4923 197466 20920 197594
rect 21000 197546 25993 225254
rect 26073 225193 26213 225334
rect 26073 197800 26213 225000
rect 26073 197466 26213 197594
rect 26293 197546 27183 225254
rect 27263 225193 27383 225334
rect 27263 197800 27383 225000
rect 27263 197466 27383 197594
rect 27463 197546 28353 225254
rect 28433 225193 28573 225334
rect 28433 197800 28573 225000
rect 28433 197466 28573 197594
rect 0 191138 28573 197466
rect 28653 191218 28719 225522
rect 0 189472 28699 191138
rect 28779 189552 29375 232288
rect 29455 225334 29651 232368
rect 29435 197546 29671 225254
rect 29455 192613 29651 197466
rect 29731 192693 30327 235429
rect 30387 234418 30453 268722
rect 30533 268534 39893 268802
rect 30533 268393 30673 268534
rect 30533 240666 30673 240794
rect 30753 240746 31683 268454
rect 31763 268393 31883 268534
rect 31763 240666 31883 240794
rect 31963 240746 32653 268454
rect 32733 268393 32853 268534
rect 32733 240666 32853 240794
rect 32933 240746 33623 268454
rect 33703 268393 33823 268534
rect 33703 240666 33823 240794
rect 33903 240746 34833 268454
rect 34913 268393 35033 268534
rect 36123 268473 37213 268534
rect 34913 240666 35033 240794
rect 35113 240746 36043 268454
rect 36123 268393 36243 268473
rect 37093 268393 37213 268473
rect 36323 240794 37013 268393
rect 36123 240714 36243 240794
rect 37093 240714 37213 240794
rect 37293 240746 38223 268454
rect 38303 268393 38423 268534
rect 36123 240666 37213 240714
rect 38303 240666 38423 240794
rect 38503 240746 39593 268454
rect 39673 268393 39893 268534
rect 677707 246866 677927 247007
rect 678007 246946 679097 275854
rect 679177 275806 679297 275934
rect 680387 275886 681477 275934
rect 679177 246866 679297 247007
rect 679377 246946 680307 275854
rect 680387 275806 680507 275886
rect 681357 275806 681477 275886
rect 680587 247007 681277 275806
rect 680387 246927 680507 247007
rect 681357 246927 681477 247007
rect 681557 246946 682487 275854
rect 682567 275806 682687 275934
rect 680387 246866 681477 246927
rect 682567 246866 682687 247007
rect 682767 246946 683697 275854
rect 683777 275806 683897 275934
rect 683777 246866 683897 247007
rect 683977 246946 684667 275854
rect 684747 275806 684867 275934
rect 684747 246866 684867 247007
rect 684947 246946 685637 275854
rect 685717 275806 685837 275934
rect 685717 246866 685837 247007
rect 685917 246946 686847 275854
rect 686927 275806 687067 275934
rect 686927 246866 687067 247007
rect 677707 246598 687067 246866
rect 687147 246678 687213 282182
rect 687273 281171 687869 324907
rect 687949 320134 688145 324987
rect 687929 291346 688165 320054
rect 687949 284232 688145 291266
rect 688225 284312 688821 328048
rect 688901 326462 717600 328128
rect 688881 291078 688947 326382
rect 689027 320134 717600 326462
rect 689027 320006 689167 320134
rect 689027 291600 689167 319800
rect 689027 291266 689167 291407
rect 689247 291346 690137 320054
rect 690217 320006 690337 320134
rect 690217 291600 690337 319800
rect 690217 291266 690337 291407
rect 690417 291346 691307 320054
rect 691387 320006 691527 320134
rect 691387 291600 691527 319800
rect 691387 291266 691527 291407
rect 691607 291346 696600 320054
rect 696680 320006 712677 320134
rect 712757 319800 717600 320054
rect 696680 291600 717600 319800
rect 696680 291266 712677 291407
rect 712757 291346 717600 291600
rect 689027 290998 717600 291266
rect 688901 284232 717600 290998
rect 687949 283928 717600 284232
rect 687949 281091 688145 283928
rect 687293 280787 688145 281091
rect 39673 240666 39893 240794
rect 30533 234338 39893 240666
rect 30407 225602 39893 234338
rect 677707 237862 687193 246598
rect 677707 231534 687067 237862
rect 677707 231406 677927 231534
rect 29455 192309 30307 192613
rect 29455 189472 29651 192309
rect 0 189168 29651 189472
rect 0 182402 28699 189168
rect 0 182134 28573 182402
rect 0 181800 4843 182054
rect 4923 181993 20920 182134
rect 0 153400 20920 181800
rect 0 152400 4843 153400
rect 0 125200 20920 152400
rect 0 124946 4843 125200
rect 4923 124866 20920 125007
rect 21000 124946 25993 182054
rect 26073 181993 26213 182134
rect 26073 153400 26213 181800
rect 26073 125200 26213 152400
rect 26073 124866 26213 125007
rect 26293 124946 27183 182054
rect 27263 181993 27383 182134
rect 27263 153400 27383 181800
rect 27263 125200 27383 152400
rect 27263 124866 27383 125007
rect 27463 124946 28353 182054
rect 28433 181993 28573 182134
rect 28433 153400 28573 181800
rect 28653 153400 28719 182322
rect 28433 125200 28573 152400
rect 28433 124866 28573 125007
rect 0 110534 28573 124866
rect 0 110200 4843 110454
rect 4923 110393 20920 110534
rect 0 83000 20920 110200
rect 0 82746 4843 83000
rect 4923 82666 20920 83000
rect 21000 82746 25993 110454
rect 26073 110393 26213 110534
rect 26073 82666 26213 110200
rect 26293 82746 27183 110454
rect 27263 110393 27383 110534
rect 27263 82666 27383 110200
rect 27463 82746 28353 110454
rect 28433 110393 28573 110534
rect 28433 82666 28573 110200
rect 0 68334 28573 82666
rect 0 68000 4843 68254
rect 4923 68193 20920 68334
rect 0 40800 20920 68000
rect 0 40546 4843 40800
rect 4923 40466 20920 40549
rect 0 40349 20920 40466
rect 21000 40429 25993 68254
rect 26073 68193 26213 68334
rect 26073 40800 26213 68000
rect 26073 40466 26213 40549
rect 26293 40546 27183 68254
rect 27263 68193 27383 68334
rect 27263 40800 27383 68000
rect 27263 40466 27383 40549
rect 27463 40546 28353 68254
rect 28433 68193 28573 68334
rect 28433 40800 28573 68000
rect 28433 40466 28573 40549
rect 26073 40349 28573 40466
rect 0 35285 28573 40349
rect 28653 35365 28719 152400
rect 28779 35418 29375 189088
rect 29455 182134 29651 189168
rect 29435 153400 29671 182054
rect 29435 124946 29671 152400
rect 29455 110534 29651 124866
rect 29435 82746 29671 110454
rect 29455 68334 29651 82666
rect 29435 36489 29671 68254
rect 29731 36625 30327 192229
rect 30387 191218 30453 225522
rect 30533 225334 39893 225602
rect 30533 225193 30673 225334
rect 30533 197466 30673 197594
rect 30753 197546 31683 225254
rect 31763 225193 31883 225334
rect 31763 197466 31883 197594
rect 31963 197546 32653 225254
rect 32733 225193 32853 225334
rect 32733 197466 32853 197594
rect 32933 197546 33623 225254
rect 33703 225193 33823 225334
rect 33703 197466 33823 197594
rect 33903 197546 34833 225254
rect 34913 225193 35033 225334
rect 36123 225273 37213 225334
rect 34913 197466 35033 197594
rect 35113 197546 36043 225254
rect 36123 225193 36243 225273
rect 37093 225193 37213 225273
rect 36323 197594 37013 225193
rect 36123 197514 36243 197594
rect 37093 197514 37213 197594
rect 37293 197546 38223 225254
rect 38303 225193 38423 225334
rect 36123 197466 37213 197514
rect 38303 197466 38423 197594
rect 38503 197546 39593 225254
rect 39673 225193 39893 225334
rect 677707 202666 677927 202807
rect 678007 202746 679097 231454
rect 679177 231406 679297 231534
rect 680387 231486 681477 231534
rect 679177 202666 679297 202807
rect 679377 202746 680307 231454
rect 680387 231406 680507 231486
rect 681357 231406 681477 231486
rect 680587 202807 681277 231406
rect 680387 202727 680507 202807
rect 681357 202727 681477 202807
rect 681557 202746 682487 231454
rect 682567 231406 682687 231534
rect 680387 202666 681477 202727
rect 682567 202666 682687 202807
rect 682767 202746 683697 231454
rect 683777 231406 683897 231534
rect 683777 202666 683897 202807
rect 683977 202746 684667 231454
rect 684747 231406 684867 231534
rect 684747 202666 684867 202807
rect 684947 202746 685637 231454
rect 685717 231406 685837 231534
rect 685717 202666 685837 202807
rect 685917 202746 686847 231454
rect 686927 231406 687067 231534
rect 686927 202666 687067 202807
rect 677707 202398 687067 202666
rect 687147 202478 687213 237782
rect 687273 236771 687869 280707
rect 687949 275934 688145 280787
rect 687929 246946 688165 275854
rect 687949 239832 688145 246866
rect 688225 239912 688821 283848
rect 688901 282262 717600 283928
rect 688881 246678 688947 282182
rect 689027 275934 717600 282262
rect 689027 275806 689167 275934
rect 689027 247200 689167 275600
rect 689027 246866 689167 247007
rect 689247 246946 690137 275854
rect 690217 275806 690337 275934
rect 690217 247200 690337 275600
rect 690217 246866 690337 247007
rect 690417 246946 691307 275854
rect 691387 275806 691527 275934
rect 691387 247200 691527 275600
rect 691387 246866 691527 247007
rect 691607 246946 696600 275854
rect 696680 275806 712677 275934
rect 712757 275600 717600 275854
rect 696680 247200 717600 275600
rect 696680 246866 712677 247007
rect 712757 246946 717600 247200
rect 689027 246598 717600 246866
rect 688901 239832 717600 246598
rect 687949 239528 717600 239832
rect 687949 236691 688145 239528
rect 687293 236387 688145 236691
rect 39673 197466 39893 197594
rect 30533 191138 39893 197466
rect 30407 182402 39893 191138
rect 677707 193662 687193 202398
rect 677707 187334 687067 193662
rect 677707 187206 677927 187334
rect 30387 153400 30453 182322
rect 30533 182134 39893 182402
rect 30533 181993 30673 182134
rect 30753 154400 31683 182054
rect 31763 181993 31883 182134
rect 31963 153400 32653 182054
rect 32733 181993 32853 182134
rect 29751 36409 30307 36545
rect 29455 36005 30307 36409
rect 30387 36085 30453 152400
rect 30533 124866 30673 125007
rect 30753 124946 31683 153400
rect 31763 124866 31883 125007
rect 31963 124946 32653 152400
rect 32733 124866 32853 125007
rect 32933 124946 33623 182054
rect 33703 181993 33823 182134
rect 33703 124866 33823 125007
rect 33903 124946 34833 182054
rect 34913 181993 35033 182134
rect 36123 182073 37213 182134
rect 34913 124866 35033 125007
rect 35113 124946 36043 182054
rect 36123 181993 36243 182073
rect 37093 181993 37213 182073
rect 36323 153400 37013 181993
rect 37293 154400 38223 182054
rect 38303 181993 38423 182134
rect 36323 125007 37013 152400
rect 36123 124927 36243 125007
rect 37093 124927 37213 125007
rect 37293 124946 38223 153400
rect 36123 124866 37213 124927
rect 38303 124866 38423 125007
rect 38503 124946 39593 182054
rect 39673 181993 39893 182134
rect 677707 158466 677927 158607
rect 678007 158546 679097 187254
rect 679177 187206 679297 187334
rect 680387 187286 681477 187334
rect 679177 158466 679297 158607
rect 679377 158546 680307 187254
rect 680387 187206 680507 187286
rect 681357 187206 681477 187286
rect 680587 158607 681277 187206
rect 680387 158527 680507 158607
rect 681357 158527 681477 158607
rect 681557 158546 682487 187254
rect 682567 187206 682687 187334
rect 680387 158466 681477 158527
rect 682567 158466 682687 158607
rect 682767 158546 683697 187254
rect 683777 187206 683897 187334
rect 683777 158466 683897 158607
rect 683977 158546 684667 187254
rect 684747 187206 684867 187334
rect 684747 158466 684867 158607
rect 684947 158546 685637 187254
rect 685717 187206 685837 187334
rect 685717 158466 685837 158607
rect 685917 158546 686847 187254
rect 686927 187206 687067 187334
rect 686927 158466 687067 158607
rect 677707 158198 687067 158466
rect 687147 158278 687213 193582
rect 687273 192571 687869 236307
rect 687949 231534 688145 236387
rect 687929 202746 688165 231454
rect 687949 195632 688145 202666
rect 688225 195712 688821 239448
rect 688901 237862 717600 239528
rect 688881 202478 688947 237782
rect 689027 231534 717600 237862
rect 689027 231406 689167 231534
rect 689027 203000 689167 231200
rect 689027 202666 689167 202807
rect 689247 202746 690137 231454
rect 690217 231406 690337 231534
rect 690217 203000 690337 231200
rect 690217 202666 690337 202807
rect 690417 202746 691307 231454
rect 691387 231406 691527 231534
rect 691387 203000 691527 231200
rect 691387 202666 691527 202807
rect 691607 202746 696600 231454
rect 696680 231406 712677 231534
rect 712757 231200 717600 231454
rect 696680 203000 717600 231200
rect 696680 202666 712677 202807
rect 712757 202746 717600 203000
rect 689027 202398 717600 202666
rect 688901 195632 717600 202398
rect 687949 195328 717600 195632
rect 687949 192491 688145 195328
rect 687293 192187 688145 192491
rect 677707 149462 687193 158198
rect 677707 143134 687067 149462
rect 677707 143006 677927 143134
rect 30533 110534 39593 124866
rect 677707 114066 677927 114207
rect 678007 114146 679097 143054
rect 679177 143006 679297 143134
rect 680387 143086 681477 143134
rect 679177 114066 679297 114207
rect 679377 114146 680307 143054
rect 680387 143006 680507 143086
rect 681357 143006 681477 143086
rect 680587 114207 681277 143006
rect 680387 114127 680507 114207
rect 681357 114127 681477 114207
rect 681557 114146 682487 143054
rect 682567 143006 682687 143134
rect 680387 114066 681477 114127
rect 682567 114066 682687 114207
rect 682767 114146 683697 143054
rect 683777 143006 683897 143134
rect 683777 114066 683897 114207
rect 683977 114146 684667 143054
rect 684747 143006 684867 143134
rect 684747 114066 684867 114207
rect 684947 114146 685637 143054
rect 685717 143006 685837 143134
rect 685717 114066 685837 114207
rect 685917 114146 686847 143054
rect 686927 143006 687067 143134
rect 686927 114066 687067 114207
rect 677707 113798 687067 114066
rect 687147 113878 687213 149382
rect 687273 148371 687869 192107
rect 687949 187334 688145 192187
rect 687929 158546 688165 187254
rect 687949 151432 688145 158466
rect 688225 151512 688821 195248
rect 688901 193662 717600 195328
rect 688881 158278 688947 193582
rect 689027 187334 717600 193662
rect 689027 187206 689167 187334
rect 689027 158800 689167 187000
rect 689027 158466 689167 158607
rect 689247 158546 690137 187254
rect 690217 187206 690337 187334
rect 690217 158800 690337 187000
rect 690217 158466 690337 158607
rect 690417 158546 691307 187254
rect 691387 187206 691527 187334
rect 691387 158800 691527 187000
rect 691387 158466 691527 158607
rect 691607 158546 696600 187254
rect 696680 187206 712677 187334
rect 712757 187000 717600 187254
rect 696680 158800 717600 187000
rect 696680 158466 712677 158607
rect 712757 158546 717600 158800
rect 689027 158198 717600 158466
rect 688901 151432 717600 158198
rect 687949 151128 717600 151432
rect 687949 148291 688145 151128
rect 687293 147987 688145 148291
rect 30533 110393 30673 110534
rect 30533 82666 30673 83000
rect 30753 82746 31683 110454
rect 31763 110393 31883 110534
rect 31763 82666 31883 83000
rect 31963 82746 32653 110454
rect 32733 110393 32853 110534
rect 32733 82666 32853 83000
rect 32933 82746 33623 110454
rect 33703 110393 33823 110534
rect 33703 82666 33823 83000
rect 33903 82746 34833 110454
rect 34913 110393 35033 110534
rect 36123 110473 37213 110534
rect 34913 82666 35033 83000
rect 35113 82746 36043 110454
rect 36123 110393 36243 110473
rect 37093 110393 37213 110473
rect 36123 82727 36243 83000
rect 36323 82807 37013 110393
rect 37093 82727 37213 83000
rect 37293 82746 38223 110454
rect 38303 110393 38423 110534
rect 36123 82666 37213 82727
rect 38303 82666 38423 83000
rect 38503 82746 39593 110454
rect 677707 105062 687193 113798
rect 677707 98734 687067 105062
rect 677707 98606 677927 98734
rect 30533 68334 39593 82666
rect 30533 68193 30673 68334
rect 30533 40466 30673 40549
rect 30753 40546 31683 68254
rect 31763 68193 31883 68334
rect 31763 40466 31883 40549
rect 31963 40546 32653 68254
rect 32733 68193 32853 68334
rect 32733 40466 32853 40549
rect 32933 40546 33623 68254
rect 33703 68193 33823 68334
rect 33703 40466 33823 40549
rect 33903 40546 34833 68254
rect 34913 68193 35033 68334
rect 36123 68273 37213 68334
rect 34913 40466 35033 40549
rect 35113 40546 36043 68254
rect 36123 68193 36243 68273
rect 37093 68193 37213 68273
rect 36323 40549 37013 68193
rect 36123 40469 36243 40549
rect 37093 40469 37213 40549
rect 37293 40546 38223 68254
rect 38303 68193 38423 68334
rect 36123 40466 37213 40469
rect 38303 40466 38423 40549
rect 38503 40546 39593 68254
rect 39673 40466 40000 40549
rect 30533 39673 40000 40466
rect 186606 39673 202207 39893
rect 295206 39673 310807 39893
rect 350006 39673 365607 39893
rect 404806 39673 420407 39893
rect 459606 39673 475207 39893
rect 514406 39673 530007 39893
rect 677051 39673 677927 40000
rect 30533 38423 39450 39673
rect 39530 38503 79054 39593
rect 79134 38423 93466 39593
rect 93546 38503 132854 39593
rect 132934 38423 147266 39593
rect 147346 38503 186654 39593
rect 186734 38423 202066 39673
rect 202146 38503 241454 39593
rect 241534 38423 255866 39593
rect 255946 38503 295254 39593
rect 295334 38423 310666 39673
rect 310746 38503 350054 39593
rect 350134 38423 365466 39673
rect 365546 38503 404854 39593
rect 404934 38423 420266 39673
rect 420346 38503 459654 39593
rect 459734 38423 475066 39673
rect 475146 38503 514454 39593
rect 514534 38423 529866 39673
rect 529946 38503 569254 39593
rect 569334 38423 583666 39593
rect 583746 38503 623054 39593
rect 623134 38423 637466 39593
rect 637546 38503 677054 39593
rect 677134 39450 677927 39673
rect 678007 39530 679097 98654
rect 679177 98606 679297 98734
rect 680387 98686 681477 98734
rect 679377 70200 680307 98654
rect 680387 98606 680507 98686
rect 681357 98606 681477 98686
rect 680587 69200 681277 98606
rect 679177 39450 679297 40000
rect 677134 39163 679297 39450
rect 679377 39243 680307 69200
rect 680387 39626 680507 40000
rect 680587 39706 681277 68200
rect 681357 39626 681477 40000
rect 681557 39695 682487 98654
rect 682567 98606 682687 98734
rect 680387 39615 681477 39626
rect 682567 39615 682687 40000
rect 682767 39680 683697 98654
rect 683777 98606 683897 98734
rect 680387 39600 682687 39615
rect 683777 39643 683897 40000
rect 683977 39723 684667 98654
rect 684747 98606 684867 98734
rect 684947 69200 685637 98654
rect 685717 98606 685837 98734
rect 685917 70200 686847 98654
rect 686927 98606 687067 98734
rect 687147 69200 687213 104982
rect 687273 103971 687869 147907
rect 687949 143134 688145 147987
rect 687929 114146 688165 143054
rect 687949 107032 688145 114066
rect 688225 107112 688821 151048
rect 688901 149462 717600 151128
rect 688881 113878 688947 149382
rect 689027 143134 717600 149462
rect 689027 143006 689167 143134
rect 689027 114400 689167 142800
rect 689027 114066 689167 114207
rect 689247 114146 690137 143054
rect 690217 143006 690337 143134
rect 690217 114400 690337 142800
rect 690217 114066 690337 114207
rect 690417 114146 691307 143054
rect 691387 143006 691527 143134
rect 691387 114400 691527 142800
rect 691387 114066 691527 114207
rect 691607 114146 696600 143054
rect 696680 143006 712677 143134
rect 712757 142800 717600 143054
rect 696680 114400 717600 142800
rect 696680 114066 712677 114207
rect 712757 114146 717600 114400
rect 689027 113798 717600 114066
rect 688901 107032 717600 113798
rect 687949 106728 717600 107032
rect 687949 103891 688145 106728
rect 687293 103587 688145 103891
rect 684747 39653 684867 40000
rect 684947 39733 685637 68200
rect 685717 39653 685837 40000
rect 685917 39705 686847 69200
rect 684747 39643 685837 39653
rect 683777 39625 685837 39643
rect 686927 39625 687067 40000
rect 683777 39600 687067 39625
rect 680387 39163 687067 39600
rect 677134 38423 687067 39163
rect 30533 38303 40000 38423
rect 78993 38303 93607 38423
rect 132793 38303 147407 38423
rect 186606 38303 202207 38423
rect 241200 38303 256007 38423
rect 295206 38303 310807 38423
rect 350006 38303 365607 38423
rect 404806 38303 420407 38423
rect 459606 38303 475207 38423
rect 514406 38303 530007 38423
rect 569193 38303 583807 38423
rect 622993 38303 637607 38423
rect 677051 38303 687067 38423
rect 30533 37213 39163 38303
rect 39243 37293 79054 38223
rect 79134 37213 93466 38303
rect 93546 37293 132854 38223
rect 132934 37213 147266 38303
rect 147346 37293 186654 38223
rect 186734 37213 202066 38303
rect 202146 37293 241454 38223
rect 241534 37213 255866 38303
rect 255946 37293 295254 38223
rect 295334 37213 310666 38303
rect 310746 37293 350054 38223
rect 350134 37213 365466 38303
rect 365546 37293 404854 38223
rect 404934 37213 420266 38303
rect 420346 37293 459654 38223
rect 459734 37213 475066 38303
rect 475146 37293 514454 38223
rect 514534 37213 529866 38303
rect 529946 37293 569254 38223
rect 569334 37213 583666 38303
rect 583746 37293 623054 38223
rect 623134 37213 637466 38303
rect 637546 37293 677054 38223
rect 677134 37213 687067 38303
rect 30533 37093 40000 37213
rect 78993 37093 93607 37213
rect 132793 37093 147407 37213
rect 186606 37093 202207 37213
rect 241200 37093 256007 37213
rect 295206 37093 310807 37213
rect 350006 37093 365607 37213
rect 404806 37093 420407 37213
rect 459606 37093 475207 37213
rect 514406 37093 530007 37213
rect 569193 37093 583807 37213
rect 622993 37093 637607 37213
rect 677051 37093 687067 37213
rect 30533 36243 39626 37093
rect 39706 36323 78993 37013
rect 79073 36243 93527 37093
rect 132873 36243 147327 37093
rect 147407 36323 186606 37013
rect 186686 36243 202127 37093
rect 202207 36323 241393 37013
rect 241473 36243 255927 37093
rect 256007 36323 295206 37013
rect 295286 36243 310727 37093
rect 310807 36323 350006 37013
rect 350086 36243 365527 37093
rect 365607 36323 404806 37013
rect 404886 36243 420327 37093
rect 420407 36323 459606 37013
rect 459686 36243 475127 37093
rect 475207 36323 514406 37013
rect 514486 36243 529927 37093
rect 530007 36323 569193 37013
rect 569273 36243 583727 37093
rect 583807 36323 622993 37013
rect 623073 36243 637527 37093
rect 637607 36323 677051 37013
rect 677131 36243 687067 37093
rect 30533 36123 40000 36243
rect 78993 36123 93607 36243
rect 132793 36123 147407 36243
rect 186606 36123 202207 36243
rect 241200 36123 256007 36243
rect 295206 36123 310807 36243
rect 350006 36123 365607 36243
rect 404806 36123 420407 36243
rect 459606 36123 475207 36243
rect 514406 36123 530007 36243
rect 569193 36123 583807 36243
rect 622993 36123 637607 36243
rect 677051 36123 687067 36243
rect 30533 36005 39615 36123
rect 29455 35338 39615 36005
rect 28799 35285 39615 35338
rect 0 35033 39615 35285
rect 39695 35113 79054 36043
rect 79134 35033 93466 36123
rect 93546 35113 132854 36043
rect 132934 35033 147266 36123
rect 147346 35113 186654 36043
rect 186734 35033 202066 36123
rect 202146 35113 241454 36043
rect 241534 35033 255866 36123
rect 255946 35113 295254 36043
rect 295334 35033 310666 36123
rect 310746 35113 350054 36043
rect 350134 35033 365466 36123
rect 365546 35113 404854 36043
rect 404934 35033 420266 36123
rect 420346 35113 459654 36043
rect 459734 35033 475066 36123
rect 475146 35113 514454 36043
rect 514534 35033 529866 36123
rect 529946 35113 569254 36043
rect 569334 35033 583666 36123
rect 583746 35113 623054 36043
rect 623134 35033 637466 36123
rect 637546 35113 677054 36043
rect 677134 36005 687067 36123
rect 687147 36085 687213 68200
rect 677134 35733 687193 36005
rect 687273 35813 687869 103507
rect 687949 98734 688145 103587
rect 687929 69200 688165 98654
rect 677134 35610 687849 35733
rect 687929 35690 688165 68200
rect 677134 35338 688145 35610
rect 688225 35418 688821 106648
rect 688901 105062 717600 106728
rect 688881 69200 688947 104982
rect 689027 98734 717600 105062
rect 689027 98606 689167 98734
rect 689027 69200 689167 98400
rect 688881 35365 688947 68200
rect 689027 39595 689167 68200
rect 689247 39675 690137 98654
rect 690217 98606 690337 98734
rect 690217 69200 690337 98400
rect 690217 39624 690337 68200
rect 690417 39704 691307 98654
rect 691387 98606 691527 98734
rect 691387 69200 691527 98400
rect 691387 39624 691527 68200
rect 690217 39595 691527 39624
rect 689027 39391 691527 39595
rect 691607 39471 696600 98654
rect 696680 98606 712677 98734
rect 712757 98400 717600 98654
rect 696680 69200 717600 98400
rect 712757 68200 717600 69200
rect 696680 40000 717600 68200
rect 696680 39633 712677 40000
rect 712757 39713 717600 40000
rect 696680 39391 717600 39633
rect 677134 35285 688801 35338
rect 689027 35285 717600 39391
rect 677134 35033 717600 35285
rect 0 34913 40000 35033
rect 78993 34913 93607 35033
rect 132793 34913 147407 35033
rect 186606 34913 202207 35033
rect 241200 34913 256007 35033
rect 295206 34913 310807 35033
rect 350006 34913 365607 35033
rect 404806 34913 420407 35033
rect 459606 34913 475207 35033
rect 514406 34913 530007 35033
rect 569193 34913 583807 35033
rect 622993 34913 637607 35033
rect 677051 34913 717600 35033
rect 0 33823 39600 34913
rect 39680 33903 79054 34833
rect 79134 33823 93466 34913
rect 93546 33903 132854 34833
rect 132934 33823 147266 34913
rect 147346 33903 186654 34833
rect 186734 33823 202066 34913
rect 202146 33903 241454 34833
rect 241534 33823 255866 34913
rect 255946 33903 295254 34833
rect 295334 33823 310666 34913
rect 310746 33903 350054 34833
rect 350134 33823 365466 34913
rect 365546 33903 404854 34833
rect 404934 33823 420266 34913
rect 420346 33903 459654 34833
rect 459734 33823 475066 34913
rect 475146 33903 514454 34833
rect 514534 33823 529866 34913
rect 529946 33903 569254 34833
rect 569334 33823 583666 34913
rect 583746 33903 623054 34833
rect 623134 33823 637466 34913
rect 637546 33903 677054 34833
rect 677134 33823 717600 34913
rect 0 33703 40000 33823
rect 78993 33703 93607 33823
rect 132793 33703 147407 33823
rect 186606 33703 202207 33823
rect 241200 33703 256007 33823
rect 295206 33703 310807 33823
rect 350006 33703 365607 33823
rect 404806 33703 420407 33823
rect 459606 33703 475207 33823
rect 514406 33703 530007 33823
rect 569193 33703 583807 33823
rect 622993 33703 637607 33823
rect 677051 33703 717600 33823
rect 0 32853 39643 33703
rect 39723 32933 79054 33623
rect 79134 32853 93466 33703
rect 93546 32933 132854 33623
rect 132934 32853 147266 33703
rect 147346 32933 186654 33623
rect 186734 32853 202066 33703
rect 202146 32933 241454 33623
rect 241534 32853 255866 33703
rect 255946 32933 295254 33623
rect 295334 32853 310666 33703
rect 310746 32933 350054 33623
rect 350134 32853 365466 33703
rect 365546 32933 404854 33623
rect 404934 32853 420266 33703
rect 420346 32933 459654 33623
rect 459734 32853 475066 33703
rect 475146 32933 514454 33623
rect 514534 32853 529866 33703
rect 529946 32933 569254 33623
rect 569334 32853 583666 33703
rect 583746 32933 623054 33623
rect 623134 32853 637466 33703
rect 637546 32933 677054 33623
rect 677134 32853 717600 33703
rect 0 32733 40000 32853
rect 78993 32733 93607 32853
rect 132793 32733 147407 32853
rect 186606 32733 202207 32853
rect 241200 32733 256007 32853
rect 295206 32733 310807 32853
rect 350006 32733 365607 32853
rect 404806 32733 420407 32853
rect 459606 32733 475207 32853
rect 514406 32733 530007 32853
rect 569193 32733 583807 32853
rect 622993 32733 637607 32853
rect 677051 32733 717600 32853
rect 0 31883 39653 32733
rect 39733 31963 79054 32653
rect 79134 31883 93466 32733
rect 93546 31963 132854 32653
rect 132934 31883 147266 32733
rect 147346 31963 186654 32653
rect 186734 31883 202066 32733
rect 202146 31963 241454 32653
rect 241534 31883 255866 32733
rect 255946 31963 295254 32653
rect 295334 31883 310666 32733
rect 310746 31963 350054 32653
rect 350134 31883 365466 32733
rect 365546 31963 404854 32653
rect 404934 31883 420266 32733
rect 420346 31963 459654 32653
rect 459734 31883 475066 32733
rect 475146 31963 514454 32653
rect 514534 31883 529866 32733
rect 529946 31963 569254 32653
rect 569334 31883 583666 32733
rect 583746 31963 623054 32653
rect 623134 31883 637466 32733
rect 637546 31963 677054 32653
rect 677134 31883 717600 32733
rect 0 31763 40000 31883
rect 78993 31763 93607 31883
rect 132793 31763 147407 31883
rect 186606 31763 202207 31883
rect 241200 31763 256007 31883
rect 295206 31763 310807 31883
rect 350006 31763 365607 31883
rect 404806 31763 420407 31883
rect 459606 31763 475207 31883
rect 514406 31763 530007 31883
rect 569193 31763 583807 31883
rect 622993 31763 637607 31883
rect 677051 31763 717600 31883
rect 0 30673 39625 31763
rect 39705 30753 79054 31683
rect 79134 30673 93466 31763
rect 132934 31754 147266 31763
rect 132949 30682 147266 31754
rect 147346 30753 186654 31683
rect 132934 30673 147266 30682
rect 186734 30673 202066 31763
rect 202146 30753 241454 31683
rect 241534 30673 255866 31763
rect 255946 30753 295254 31683
rect 295334 30673 310666 31763
rect 310746 30753 350054 31683
rect 350134 30673 365466 31763
rect 365546 30753 404854 31683
rect 404934 30673 420266 31763
rect 420346 30753 459654 31683
rect 459734 30673 475066 31763
rect 475146 30753 514454 31683
rect 514534 30673 529866 31763
rect 529946 30753 569254 31683
rect 569334 30673 583666 31763
rect 583746 30753 623054 31683
rect 623134 30673 637466 31763
rect 637546 30753 677054 31683
rect 677134 30673 717600 31763
rect 0 30533 40000 30673
rect 78993 30533 93607 30673
rect 132793 30533 147407 30673
rect 186606 30533 202207 30673
rect 241200 30533 256007 30673
rect 295206 30533 310807 30673
rect 350006 30533 365607 30673
rect 404806 30533 420407 30673
rect 459606 30533 475207 30673
rect 514406 30533 530007 30673
rect 569193 30533 583807 30673
rect 622993 30533 637607 30673
rect 677051 30533 717600 30673
rect 0 30407 36005 30533
rect 0 29751 35733 30407
rect 36085 30387 79054 30453
rect 79134 30407 93466 30533
rect 93546 30387 192982 30453
rect 193062 30407 201798 30533
rect 201878 30387 301582 30453
rect 301662 30407 310398 30533
rect 310478 30387 356382 30453
rect 356462 30407 365198 30533
rect 365278 30387 411182 30453
rect 411262 30407 419998 30533
rect 420078 30387 465982 30453
rect 466062 30407 474798 30533
rect 474878 30387 520782 30453
rect 520862 30407 529598 30533
rect 529678 30387 681515 30453
rect 0 29455 35610 29751
rect 35813 29731 191507 30327
rect 0 28799 35338 29455
rect 35690 29435 79054 29671
rect 79134 29455 93466 29651
rect 93546 29435 132854 29671
rect 132934 29455 147266 29651
rect 147346 29435 186654 29671
rect 191587 29651 191891 30307
rect 191971 29731 300107 30327
rect 186734 29455 202066 29651
rect 0 28573 35285 28799
rect 35418 28779 194648 29375
rect 35365 28653 79054 28719
rect 79134 28573 93466 28699
rect 194728 28699 195032 29455
rect 202146 29435 241454 29671
rect 241534 29455 255866 29651
rect 255946 29435 295254 29671
rect 300187 29651 300491 30307
rect 300571 29731 354907 30327
rect 295334 29455 310666 29651
rect 195112 28779 303248 29375
rect 193062 28573 201798 28699
rect 201878 28653 301582 28719
rect 303328 28699 303632 29455
rect 310746 29435 350054 29671
rect 354987 29651 355291 30307
rect 355371 29731 409707 30327
rect 350134 29455 365466 29651
rect 303712 28779 358048 29375
rect 301662 28573 310398 28699
rect 310478 28653 356382 28719
rect 358128 28699 358432 29455
rect 365546 29435 404854 29671
rect 409787 29651 410091 30307
rect 410171 29731 464507 30327
rect 404934 29455 420266 29651
rect 358512 28779 412848 29375
rect 356462 28573 365198 28699
rect 365278 28653 411182 28719
rect 412928 28699 413232 29455
rect 420346 29435 459654 29671
rect 464587 29651 464891 30307
rect 464971 29731 519307 30327
rect 459734 29455 475066 29651
rect 413312 28779 467648 29375
rect 411262 28573 419998 28699
rect 420078 28653 465982 28719
rect 467728 28699 468032 29455
rect 475146 29435 514454 29671
rect 519387 29651 519691 30307
rect 519771 29731 680975 30327
rect 681595 30307 717600 30533
rect 681055 29751 717600 30307
rect 514534 29455 529866 29651
rect 468112 28779 522448 29375
rect 466062 28573 474798 28699
rect 474878 28653 520782 28719
rect 522528 28699 522832 29455
rect 529946 29435 569254 29671
rect 569334 29455 583666 29651
rect 583746 29435 623054 29671
rect 623134 29455 637466 29651
rect 637546 29435 681111 29671
rect 681191 29455 717600 29751
rect 522912 28779 682182 29375
rect 682262 28799 717600 29455
rect 520862 28573 529598 28699
rect 529678 28653 682235 28719
rect 682315 28573 717600 28799
rect 0 28433 78800 28573
rect 78993 28433 93607 28573
rect 93800 28433 132600 28573
rect 132793 28433 147407 28573
rect 147600 28433 186400 28573
rect 186606 28433 202207 28573
rect 202400 28433 256007 28573
rect 256200 28433 295000 28573
rect 295206 28433 310807 28573
rect 311000 28433 349800 28573
rect 350006 28433 365607 28573
rect 365800 28433 404600 28573
rect 404806 28433 420407 28573
rect 420600 28433 459400 28573
rect 459606 28433 475207 28573
rect 475400 28433 514200 28573
rect 514406 28433 530007 28573
rect 530200 28433 569000 28573
rect 569193 28433 583807 28573
rect 584000 28433 622800 28573
rect 622993 28433 637607 28573
rect 637800 28433 676800 28573
rect 677051 28433 717600 28573
rect 0 27383 39595 28433
rect 39675 27463 79054 28353
rect 79134 27383 93466 28433
rect 93546 27463 132854 28353
rect 132934 27383 147266 28433
rect 147346 27463 186654 28353
rect 186734 27383 202066 28433
rect 202146 27463 241454 28353
rect 241534 27383 255866 28433
rect 255946 27463 295254 28353
rect 295334 27383 310666 28433
rect 310746 27463 350054 28353
rect 350134 27383 365466 28433
rect 365546 27463 404854 28353
rect 404934 27383 420266 28433
rect 420346 27463 459654 28353
rect 459734 27383 475066 28433
rect 475146 27463 514454 28353
rect 514534 27383 529866 28433
rect 529946 27463 569254 28353
rect 569334 27383 583666 28433
rect 583746 27463 623054 28353
rect 623134 27383 637466 28433
rect 637546 27463 677054 28353
rect 677134 27383 717600 28433
rect 0 27263 78800 27383
rect 78993 27263 93607 27383
rect 93800 27263 132600 27383
rect 132793 27263 147407 27383
rect 147600 27263 186400 27383
rect 186606 27263 202207 27383
rect 202400 27263 256007 27383
rect 256200 27263 295000 27383
rect 295206 27263 310807 27383
rect 311000 27263 349800 27383
rect 350006 27263 365607 27383
rect 365800 27263 404600 27383
rect 404806 27263 420407 27383
rect 420600 27263 459400 27383
rect 459606 27263 475207 27383
rect 475400 27263 514200 27383
rect 514406 27263 530007 27383
rect 530200 27263 569000 27383
rect 569193 27263 583807 27383
rect 584000 27263 622800 27383
rect 622993 27263 637607 27383
rect 637800 27263 676800 27383
rect 677051 27263 717600 27383
rect 0 26213 39624 27263
rect 39704 26293 79054 27183
rect 79134 26213 93466 27263
rect 93546 26293 132854 27183
rect 132934 26213 147266 27263
rect 147346 26293 186654 27183
rect 186734 26213 202066 27263
rect 202146 26293 241454 27183
rect 241534 26213 255866 27263
rect 255946 26293 295254 27183
rect 295334 26213 310666 27263
rect 310746 26293 350054 27183
rect 350134 26213 365466 27263
rect 365546 26293 404854 27183
rect 404934 26213 420266 27263
rect 420346 26293 459654 27183
rect 459734 26213 475066 27263
rect 475146 26293 514454 27183
rect 514534 26213 529866 27263
rect 529946 26293 569254 27183
rect 569334 26213 583666 27263
rect 583746 26293 623054 27183
rect 623134 26213 637466 27263
rect 637546 26293 677054 27183
rect 677134 26213 717600 27263
rect 0 26073 78800 26213
rect 78993 26073 93607 26213
rect 93800 26073 132600 26213
rect 132793 26073 147407 26213
rect 147600 26073 186400 26213
rect 186606 26073 202207 26213
rect 202400 26073 256007 26213
rect 256200 26073 295000 26213
rect 295206 26073 310807 26213
rect 311000 26073 349800 26213
rect 350006 26073 365607 26213
rect 365800 26073 404600 26213
rect 404806 26073 420407 26213
rect 420600 26073 459400 26213
rect 459606 26073 475207 26213
rect 475400 26073 514200 26213
rect 514406 26073 530007 26213
rect 530200 26073 569000 26213
rect 569193 26073 583807 26213
rect 584000 26073 622800 26213
rect 622993 26073 637607 26213
rect 637800 26073 676800 26213
rect 677051 26073 717600 26213
rect 0 20920 39391 26073
rect 39471 21000 79054 25993
rect 79134 20920 93466 26073
rect 93546 21000 132854 25993
rect 132934 20920 147266 26073
rect 147346 21000 186654 25993
rect 186734 20920 202066 26073
rect 202146 21000 241454 25993
rect 241534 20920 255866 26073
rect 255946 21000 295254 25993
rect 295334 20920 310666 26073
rect 310746 21000 350054 25993
rect 350134 20920 365466 26073
rect 365546 21000 404854 25993
rect 404934 20920 420266 26073
rect 420346 21000 459654 25993
rect 459734 20920 475066 26073
rect 475146 21000 514454 25993
rect 514534 20920 529866 26073
rect 529946 21000 569254 25993
rect 569334 20920 583666 26073
rect 583746 21000 623054 25993
rect 623134 20920 637466 26073
rect 637546 21000 677171 25993
rect 677251 20920 717600 26073
rect 0 4923 78800 20920
rect 78993 4923 93607 20920
rect 0 0 39633 4923
rect 40000 4843 78800 4923
rect 39713 0 79054 4843
rect 79134 0 93466 4923
rect 93800 4843 132600 20920
rect 132793 4923 147407 20920
rect 93546 0 132854 4843
rect 132934 0 147266 4923
rect 147600 4843 186400 20920
rect 186606 4923 202207 20920
rect 202400 4923 256007 20920
rect 147346 0 186654 4843
rect 186734 0 202066 4923
rect 202400 4843 241200 4923
rect 202146 0 241454 4843
rect 241534 0 255866 4923
rect 256200 4843 295000 20920
rect 295206 4923 310807 20920
rect 255946 0 295254 4843
rect 295334 0 310666 4923
rect 311000 4843 349800 20920
rect 350006 4923 365607 20920
rect 310746 0 350054 4843
rect 350134 0 365466 4923
rect 365800 4843 404600 20920
rect 404806 4923 420407 20920
rect 365546 0 404854 4843
rect 404934 0 420266 4923
rect 420600 4843 459400 20920
rect 459606 4923 475207 20920
rect 420346 0 459654 4843
rect 459734 0 475066 4923
rect 475400 4843 514200 20920
rect 514406 4923 530007 20920
rect 475146 0 514454 4843
rect 514534 0 529866 4923
rect 530200 4843 569000 20920
rect 569193 4923 583807 20920
rect 529946 0 569254 4843
rect 569334 0 583666 4923
rect 584000 4843 622800 20920
rect 622993 4923 637607 20920
rect 583746 0 623054 4843
rect 623134 0 637466 4923
rect 637800 4843 676800 20920
rect 677051 4923 717600 20920
rect 637546 0 677054 4843
rect 677134 0 717600 4923
<< metal5 >>
rect 76410 1018624 88578 1030789
rect 124410 1018624 136578 1030789
rect 172410 1018624 184578 1030789
rect 230810 1018624 242978 1030789
rect 282210 1018624 294378 1030789
rect 340810 1018624 352978 1030789
rect 426210 1018624 438378 1030789
rect 475610 1018624 487778 1030789
rect 527210 1018624 539378 1030789
rect 577010 1018624 589178 1030789
rect 628410 1018624 640578 1030789
rect 6811 956610 18976 968778
rect 698624 945422 710789 957590
rect 6167 915054 19620 925934
rect 697980 893466 711433 904346
rect 6811 872210 18976 884378
rect 698512 848240 711002 860780
rect 6811 829810 18976 841978
rect 698624 805222 710789 817390
rect 6598 787420 19088 799960
rect 698512 760840 711002 773380
rect 6598 744220 19088 756760
rect 698512 716440 711002 728980
rect 6598 701020 19088 713560
rect 698512 672240 711002 684780
rect 6598 657620 19088 670160
rect 698512 628040 711002 640580
rect 6598 614420 19088 626960
rect 6598 571220 19088 583760
rect 698512 583640 711002 596180
rect 6598 528020 19088 540560
rect 698512 539440 711002 551980
rect 6811 484810 18976 496978
rect 698624 496422 710789 508590
rect 6167 443254 19620 454134
rect 697980 453666 711433 464546
rect 6598 400220 19088 412760
rect 698624 409822 710789 421990
rect 6598 357020 19088 369560
rect 698512 365240 711002 377780
rect 6598 313620 19088 326160
rect 698512 321040 711002 333580
rect 6598 270420 19088 282960
rect 698512 276840 711002 289380
rect 6598 227220 19088 239760
rect 698512 232440 711002 244980
rect 6598 184020 19088 196560
rect 698512 188240 711002 200780
rect 698512 144040 711002 156580
rect 6811 111610 18976 123778
rect 698512 99640 711002 112180
rect 6167 70054 19620 80934
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19620
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
<< obsm5 >>
rect 0 1032757 75254 1037600
rect 0 1016917 40800 1032757
rect 75574 1032437 89426 1037600
rect 89746 1032757 123254 1037600
rect 123574 1032437 137426 1037600
rect 137746 1032757 171254 1037600
rect 171574 1032437 185426 1037600
rect 185746 1032757 425054 1037600
rect 75000 1031109 90000 1032437
rect 75000 1018304 76090 1031109
rect 88898 1018304 90000 1031109
rect 75000 1016917 90000 1018304
rect 123000 1031109 138000 1032437
rect 123000 1018304 124090 1031109
rect 136898 1018304 138000 1031109
rect 123000 1016917 138000 1018304
rect 171000 1031109 186000 1032437
rect 171000 1018304 172090 1031109
rect 184898 1018304 186000 1031109
rect 171000 1016917 186000 1018304
rect 220000 1031109 253800 1032757
rect 220000 1018304 230490 1031109
rect 243298 1018304 253800 1031109
rect 220000 1016917 253800 1018304
rect 271400 1031109 305200 1032757
rect 271400 1018304 281890 1031109
rect 294698 1018304 305200 1031109
rect 271400 1016917 305200 1018304
rect 339400 1031109 354400 1032757
rect 425374 1032437 439226 1037600
rect 439546 1032757 474454 1037600
rect 474774 1032437 488626 1037600
rect 488946 1032757 526054 1037600
rect 526374 1032437 540226 1037600
rect 540546 1032757 627254 1037600
rect 339400 1018304 340490 1031109
rect 353298 1018304 354400 1031109
rect 339400 1016917 354400 1018304
rect 424800 1031109 439800 1032437
rect 424800 1018304 425890 1031109
rect 438698 1018304 439800 1031109
rect 424800 1016917 439800 1018304
rect 474200 1031109 489200 1032437
rect 474200 1018304 475290 1031109
rect 488098 1018304 489200 1031109
rect 474200 1016917 489200 1018304
rect 525800 1031109 540800 1032437
rect 525800 1018304 526890 1031109
rect 539698 1018304 540800 1031109
rect 525800 1016917 540800 1018304
rect 575600 1031109 590600 1032757
rect 627574 1032437 641426 1037600
rect 641746 1032757 717600 1037600
rect 575600 1018304 576690 1031109
rect 589498 1018304 590600 1031109
rect 575600 1016917 590600 1018304
rect 627000 1031109 642000 1032437
rect 627000 1018304 628090 1031109
rect 640898 1018304 642000 1031109
rect 627000 1016917 642000 1018304
rect 677600 1016917 717600 1032757
rect 0 1011287 40109 1016917
rect 40429 1011607 75254 1016597
rect 0 1009267 40226 1011287
rect 40546 1010437 75254 1011287
rect 40546 1009267 75254 1010117
rect 0 1006827 35049 1009267
rect 35369 1007147 75254 1008947
rect 0 1002551 40226 1006827
rect 40546 1005937 75254 1006827
rect 40546 1004968 75254 1005617
rect 75574 1004968 89426 1016917
rect 89746 1011607 123254 1016597
rect 89746 1010437 123254 1011287
rect 89746 1009267 123254 1010117
rect 89746 1007147 123254 1008947
rect 89746 1005937 123254 1006827
rect 89746 1004968 123254 1005617
rect 123574 1004968 137426 1016917
rect 137746 1011607 171254 1016597
rect 137746 1010437 171254 1011287
rect 137746 1009267 171254 1010117
rect 137746 1007147 171254 1008947
rect 137746 1005937 171254 1006827
rect 137746 1004968 171254 1005617
rect 171574 1004968 185426 1016917
rect 185746 1011607 229543 1016597
rect 185746 1010437 229543 1011287
rect 185746 1009267 229543 1010117
rect 229863 1008947 244857 1016917
rect 245177 1011607 280943 1016597
rect 245177 1010437 280943 1011287
rect 245177 1009267 280943 1010117
rect 281263 1008947 296257 1016917
rect 296577 1011607 339654 1016597
rect 296577 1010437 339654 1011287
rect 296577 1009267 339654 1010117
rect 185746 1007147 229448 1008947
rect 229768 1007147 244857 1008947
rect 245177 1007147 280848 1008947
rect 281168 1007147 296257 1008947
rect 296577 1007147 339654 1008947
rect 185746 1005937 229543 1006827
rect 185746 1004968 229543 1005617
rect 40800 1004967 229543 1004968
rect 40546 1003997 75254 1004647
rect 40546 1002787 75254 1003677
rect 0 998449 28333 1002551
rect 0 997600 20683 998449
rect 26313 998245 28333 998449
rect 26313 998216 27163 998245
rect 0 969946 4843 997600
rect 5163 969626 20683 970200
rect 21003 969946 25993 998129
rect 26313 969946 27163 997896
rect 27483 969946 28333 997925
rect 28653 969946 30453 1002231
rect 30773 1001257 40226 1002551
rect 40546 1001577 75254 1002467
rect 75574 1001257 89426 1004967
rect 89746 1003997 123254 1004647
rect 89746 1002787 123254 1003677
rect 89746 1001577 123254 1002467
rect 123574 1001257 137426 1004967
rect 137746 1003997 171254 1004647
rect 137746 1002787 171254 1003677
rect 137746 1001577 171254 1002467
rect 171574 1001257 185426 1004967
rect 185746 1003997 229543 1004647
rect 185746 1002787 229543 1003677
rect 185746 1001577 229543 1002467
rect 229863 1001577 244857 1007147
rect 245177 1005937 280943 1006827
rect 245177 1004967 280943 1005617
rect 245177 1003997 280943 1004647
rect 245177 1002787 280943 1003677
rect 245177 1001577 280943 1002467
rect 281263 1001577 296257 1007147
rect 296577 1005937 339654 1006827
rect 296577 1004968 339654 1005617
rect 339974 1004968 353826 1016917
rect 354146 1011607 425054 1016597
rect 354146 1010437 425054 1011287
rect 354146 1009267 425054 1010117
rect 354146 1007147 388600 1008947
rect 389600 1007147 425054 1008947
rect 354146 1005937 389600 1006827
rect 390600 1005937 425054 1006827
rect 354146 1004968 388600 1005617
rect 296577 1004967 388600 1004968
rect 389600 1004968 425054 1005617
rect 425374 1004968 439226 1016917
rect 439546 1011607 474454 1016597
rect 439546 1010437 474454 1011287
rect 439546 1009267 474454 1010117
rect 439546 1007147 474454 1008947
rect 439546 1005937 474454 1006827
rect 439546 1004968 474454 1005617
rect 474774 1004968 488626 1016917
rect 488946 1011607 526054 1016597
rect 488946 1010437 526054 1011287
rect 488946 1009267 526054 1010117
rect 488946 1007147 526054 1008947
rect 488946 1005937 526054 1006827
rect 488946 1004968 526054 1005617
rect 526374 1004968 540226 1016917
rect 540546 1011607 575854 1016597
rect 540546 1010437 575854 1011287
rect 540546 1009267 575854 1010117
rect 540546 1007147 575854 1008947
rect 540546 1005937 575854 1006827
rect 540546 1004968 575854 1005617
rect 576174 1004968 590026 1016917
rect 590346 1011607 627254 1016597
rect 590346 1010437 627254 1011287
rect 590346 1009267 627254 1010117
rect 590346 1007147 627254 1008947
rect 590346 1005937 627254 1006827
rect 590346 1004968 627254 1005617
rect 627574 1004968 641426 1016917
rect 641746 1011607 678129 1016597
rect 678449 1011287 717600 1016917
rect 641746 1010437 677896 1011287
rect 678216 1010437 717600 1011287
rect 641746 1009267 677925 1010117
rect 678245 1009267 717600 1010437
rect 641746 1007147 682231 1008947
rect 682551 1006827 717600 1009267
rect 641746 1005937 677895 1006827
rect 678215 1005617 717600 1006827
rect 641746 1004968 677867 1005617
rect 389600 1004967 677867 1004968
rect 678187 1004967 717600 1005617
rect 296577 1003997 339654 1004647
rect 296577 1002787 339654 1003677
rect 296577 1001577 339654 1002467
rect 30773 1000607 40229 1001257
rect 40549 1000607 75193 1001257
rect 75513 1000607 89487 1001257
rect 89807 1000607 123193 1001257
rect 123513 1000607 137487 1001257
rect 137807 1000607 171193 1001257
rect 171513 1000607 185487 1001257
rect 185807 1000607 229543 1001257
rect 30773 998677 40226 1000607
rect 40546 999397 75254 1000287
rect 30773 998240 36993 998677
rect 38523 998390 40226 998677
rect 30773 998215 33603 998240
rect 35133 998225 36993 998240
rect 31983 998197 33603 998215
rect 36343 998214 36993 998225
rect 31983 998187 32633 998197
rect 30773 969946 31663 997895
rect 31983 969946 32633 997867
rect 32953 969946 33603 997877
rect 33923 969946 34813 997920
rect 35133 969946 36023 997905
rect 36343 970007 36993 997894
rect 37313 969946 38203 998357
rect 38523 969946 39573 998070
rect 39893 997707 40226 998390
rect 40546 998027 75254 999077
rect 75574 998027 89426 1000607
rect 89746 999397 123254 1000287
rect 89746 998027 123254 999077
rect 123574 998027 137426 1000607
rect 137746 999397 171254 1000287
rect 137746 998027 171254 999077
rect 171574 998027 185426 1000607
rect 229863 1000287 243921 1001577
rect 244241 1000607 280943 1001257
rect 281263 1000287 295321 1001577
rect 339974 1001257 353826 1004967
rect 354146 1003997 425054 1004647
rect 354146 1002787 425054 1003677
rect 354146 1001577 425054 1002467
rect 425374 1001257 439226 1004967
rect 439546 1003997 474454 1004647
rect 439546 1002787 474454 1003677
rect 439546 1001577 474454 1002467
rect 474774 1001257 488626 1004967
rect 488946 1003997 526054 1004647
rect 488946 1002787 526054 1003677
rect 488946 1001577 526054 1002467
rect 526374 1001257 540226 1004967
rect 540546 1003997 575854 1004647
rect 540546 1002787 575854 1003677
rect 540546 1001577 575854 1002467
rect 576174 1001257 590026 1004967
rect 590346 1003997 627254 1004647
rect 590346 1002787 627254 1003677
rect 590346 1001577 627254 1002467
rect 627574 1001257 641426 1004967
rect 641746 1003997 677877 1004647
rect 678197 1003997 717600 1004967
rect 641746 1002787 677920 1003677
rect 678240 1002551 717600 1003997
rect 678240 1002467 686827 1002551
rect 641746 1001577 677905 1002467
rect 678225 1001257 686827 1002467
rect 295641 1000607 339593 1001257
rect 339913 1000607 353887 1001257
rect 354207 1000607 388600 1001257
rect 389600 1000607 424993 1001257
rect 425313 1000607 439287 1001257
rect 439607 1000607 474393 1001257
rect 474713 1000607 488687 1001257
rect 489007 1000607 525993 1001257
rect 526313 1000607 540287 1001257
rect 540607 1000607 575793 1001257
rect 576113 1000607 590087 1001257
rect 590407 1000607 627193 1001257
rect 627513 1000607 641487 1001257
rect 641807 1000607 677894 1001257
rect 678214 1000607 686827 1001257
rect 185746 999397 229543 1000287
rect 185746 998027 229543 999077
rect 229863 998027 244857 1000287
rect 245177 999397 280943 1000287
rect 245177 998027 280943 999077
rect 281263 998027 296257 1000287
rect 296577 999397 339654 1000287
rect 296577 998027 339654 999077
rect 339974 998027 353826 1000607
rect 354146 999397 389600 1000287
rect 390600 999397 425054 1000287
rect 354146 998027 425054 999077
rect 425374 998027 439226 1000607
rect 439546 999397 474454 1000287
rect 439546 998027 474454 999077
rect 474774 998027 488626 1000607
rect 488946 999397 526054 1000287
rect 488946 998027 526054 999077
rect 526374 998027 540226 1000607
rect 540546 999397 575854 1000287
rect 540546 998027 575854 999077
rect 576174 998027 590026 1000607
rect 590346 999397 627254 1000287
rect 590346 998027 627254 999077
rect 627574 998027 641426 1000607
rect 641746 999397 678357 1000287
rect 678677 999077 686827 1000607
rect 641746 998027 678070 999077
rect 678390 997707 686827 999077
rect 39893 997600 40800 997707
rect 677600 997374 686827 997707
rect 677600 996800 677707 997374
rect 680607 997371 681257 997374
rect 32632 969626 32633 969946
rect 36343 969626 36993 969687
rect 0 969098 39573 969626
rect 0 956290 6491 969098
rect 19296 956290 39573 969098
rect 678027 958857 679077 997054
rect 679397 958857 680287 997054
rect 680607 958857 681257 997051
rect 681577 958857 682467 997054
rect 682787 958857 683677 997054
rect 683997 958857 684647 997054
rect 684968 996800 685617 997054
rect 684967 958857 685617 996800
rect 685937 958857 686827 997054
rect 687147 958952 688947 1002231
rect 689267 997491 717600 1002551
rect 689267 997374 691287 997491
rect 689267 958857 690117 997054
rect 690437 958857 691287 997054
rect 691607 958857 696597 997171
rect 696917 996800 717600 997491
rect 712757 968400 717600 996800
rect 687147 958537 688947 958632
rect 696917 958537 717600 968400
rect 0 955774 39573 956290
rect 678027 957910 717600 958537
rect 0 928000 4843 955454
rect 5163 955200 20683 955774
rect 32632 955454 32633 955774
rect 36343 955713 36993 955774
rect 0 927426 20683 928000
rect 21003 927746 25993 955454
rect 26313 927746 27163 955454
rect 27483 927746 28333 955454
rect 28653 927746 30453 955454
rect 30773 927746 31663 955454
rect 31983 928000 32633 955454
rect 31983 927746 32632 928000
rect 32953 927746 33603 955454
rect 33923 927746 34813 955454
rect 35133 927746 36023 955454
rect 36343 927807 36993 955393
rect 37313 927746 38203 955454
rect 38523 927746 39573 955454
rect 678027 945102 698304 957910
rect 711109 945102 717600 957910
rect 678027 944479 717600 945102
rect 678027 943543 680287 944479
rect 36343 927426 36993 927487
rect 0 926254 39573 927426
rect 0 914734 5847 926254
rect 19940 914734 39573 926254
rect 0 913574 39573 914734
rect 0 913000 20683 913574
rect 36343 913513 36993 913574
rect 0 885800 4843 913000
rect 0 885226 20683 885800
rect 21003 885546 25993 913254
rect 26313 885546 27163 913254
rect 27483 885546 28333 913254
rect 28653 885546 30453 913254
rect 30773 885546 31663 913254
rect 31983 913000 32632 913254
rect 31983 885546 32633 913000
rect 32953 885546 33603 913254
rect 33923 885546 34813 913254
rect 35133 885546 36023 913254
rect 36343 885607 36993 913193
rect 37313 885546 38203 913254
rect 38523 885546 39573 913254
rect 678027 906146 679077 943223
rect 679397 906146 680287 943223
rect 680607 906207 681257 944159
rect 681577 943543 717600 944479
rect 681577 906146 682467 943223
rect 682787 906146 683677 943223
rect 683997 906146 684647 943223
rect 684967 906400 685617 943223
rect 684968 906146 685617 906400
rect 685937 906146 686827 943223
rect 687147 906146 688947 943223
rect 689267 906146 690117 943223
rect 690437 906146 691287 943223
rect 691607 906146 696597 943223
rect 696917 934600 717600 943543
rect 712757 906400 717600 934600
rect 680607 905826 681257 905887
rect 696917 905826 717600 906400
rect 678027 904666 717600 905826
rect 678027 893146 697660 904666
rect 711753 893146 717600 904666
rect 678027 891974 717600 893146
rect 680607 891913 681257 891974
rect 32632 885226 32633 885546
rect 36343 885226 36993 885287
rect 0 884698 39573 885226
rect 0 871890 6491 884698
rect 19296 871890 39573 884698
rect 0 871374 39573 871890
rect 0 870800 20683 871374
rect 32632 871054 32633 871374
rect 36343 871313 36993 871374
rect 0 843400 4843 870800
rect 0 842826 20683 843400
rect 21003 843146 25993 871054
rect 26313 843146 27163 871054
rect 27483 843146 28333 871054
rect 28653 843146 30453 871054
rect 30773 843146 31663 871054
rect 31983 843146 32633 871054
rect 32953 843146 33603 871054
rect 33923 843146 34813 871054
rect 35133 843146 36023 871054
rect 36343 843207 36993 870993
rect 37313 843146 38203 871054
rect 38523 843146 39573 871054
rect 678027 862746 679077 891654
rect 679397 862746 680287 891654
rect 680607 862807 681257 891593
rect 681577 862746 682467 891654
rect 682787 862746 683677 891654
rect 683997 862746 684647 891654
rect 684968 891400 685617 891654
rect 684967 863000 685617 891400
rect 684968 862746 685617 863000
rect 685937 862746 686827 891654
rect 687147 862746 688947 891654
rect 689267 862746 690117 891654
rect 690437 862746 691287 891654
rect 691607 862746 696597 891654
rect 696917 891400 717600 891974
rect 712757 863000 717600 891400
rect 680607 862426 681257 862487
rect 696917 862426 717600 863000
rect 678027 861100 717600 862426
rect 678027 847920 698192 861100
rect 711322 847920 717600 861100
rect 678027 847574 717600 847920
rect 680607 847526 681257 847574
rect 32632 842826 32633 843146
rect 36343 842826 36993 842887
rect 0 842298 39573 842826
rect 0 829490 6491 842298
rect 19296 829490 39573 842298
rect 0 828974 39573 829490
rect 0 828400 20683 828974
rect 32632 828654 32633 828974
rect 36343 828913 36993 828974
rect 0 801200 4843 828400
rect 0 800626 20683 801200
rect 21003 800946 25993 828654
rect 26313 800946 27163 828654
rect 27483 800946 28333 828654
rect 28653 800946 30453 828654
rect 30773 800946 31663 828654
rect 31983 801200 32633 828654
rect 31983 800946 32632 801200
rect 32953 800946 33603 828654
rect 33923 800946 34813 828654
rect 35133 800946 36023 828654
rect 36343 800994 36993 828593
rect 37313 800946 38203 828654
rect 38523 800946 39573 828654
rect 678027 818546 679077 847254
rect 679397 818546 680287 847254
rect 680607 818607 681257 847206
rect 681577 818546 682467 847254
rect 682787 818546 683677 847254
rect 683997 818546 684647 847254
rect 684968 847000 685617 847254
rect 684967 818546 685617 847000
rect 685937 818546 686827 847254
rect 687147 818546 688947 847254
rect 689267 818546 690117 847254
rect 690437 818546 691287 847254
rect 691607 818546 696597 847254
rect 696917 847000 717600 847574
rect 712757 818800 717600 847000
rect 680607 818226 681257 818287
rect 684967 818226 684968 818546
rect 696917 818226 717600 818800
rect 678027 817710 717600 818226
rect 678027 804902 698304 817710
rect 711109 804902 717600 817710
rect 678027 804374 717600 804902
rect 680607 804313 681257 804374
rect 684967 804054 684968 804374
rect 36343 800626 36993 800674
rect 0 800280 39573 800626
rect 0 787100 6278 800280
rect 19408 787100 39573 800280
rect 0 785774 39573 787100
rect 0 785200 20683 785774
rect 36343 785713 36993 785774
rect 0 758000 4843 785200
rect 0 757426 20683 758000
rect 21003 757746 25993 785454
rect 26313 757746 27163 785454
rect 27483 757746 28333 785454
rect 28653 757746 30453 785454
rect 30773 757746 31663 785454
rect 31983 785200 32632 785454
rect 31983 758000 32633 785200
rect 31983 757746 32632 758000
rect 32953 757746 33603 785454
rect 33923 757746 34813 785454
rect 35133 757746 36023 785454
rect 36343 757794 36993 785393
rect 37313 757746 38203 785454
rect 38523 757746 39573 785454
rect 678027 775346 679077 804054
rect 679397 775346 680287 804054
rect 680607 775407 681257 803993
rect 681577 775346 682467 804054
rect 682787 775346 683677 804054
rect 683997 775346 684647 804054
rect 684967 775600 685617 804054
rect 684968 775346 685617 775600
rect 685937 775346 686827 804054
rect 687147 775346 688947 804054
rect 689267 775346 690117 804054
rect 690437 775346 691287 804054
rect 691607 775346 696597 804054
rect 696917 803800 717600 804374
rect 712757 775600 717600 803800
rect 680607 775026 681257 775087
rect 696917 775026 717600 775600
rect 678027 773700 717600 775026
rect 678027 760520 698192 773700
rect 711322 760520 717600 773700
rect 678027 760174 717600 760520
rect 680607 760126 681257 760174
rect 36343 757426 36993 757474
rect 0 757080 39573 757426
rect 0 743900 6278 757080
rect 19408 743900 39573 757080
rect 0 742574 39573 743900
rect 0 742000 20683 742574
rect 36343 742513 36993 742574
rect 0 714800 4843 742000
rect 0 714226 20683 714800
rect 21003 714546 25993 742254
rect 26313 714546 27163 742254
rect 27483 714546 28333 742254
rect 28653 714546 30453 742254
rect 30773 714546 31663 742254
rect 31983 742000 32632 742254
rect 31983 714800 32633 742000
rect 31983 714546 32632 714800
rect 32953 714546 33603 742254
rect 33923 714546 34813 742254
rect 35133 714546 36023 742254
rect 36343 714594 36993 742193
rect 37313 714546 38203 742254
rect 38523 714546 39573 742254
rect 678027 730946 679077 759854
rect 679397 730946 680287 759854
rect 680607 731007 681257 759806
rect 681577 730946 682467 759854
rect 682787 730946 683677 759854
rect 683997 730946 684647 759854
rect 684968 759600 685617 759854
rect 684967 731200 685617 759600
rect 684968 730946 685617 731200
rect 685937 730946 686827 759854
rect 687147 730946 688947 759854
rect 689267 730946 690117 759854
rect 690437 730946 691287 759854
rect 691607 730946 696597 759854
rect 696917 759600 717600 760174
rect 712757 731200 717600 759600
rect 680607 730626 681257 730687
rect 696917 730626 717600 731200
rect 678027 729300 717600 730626
rect 678027 716120 698192 729300
rect 711322 716120 717600 729300
rect 678027 715774 717600 716120
rect 680607 715726 681257 715774
rect 36343 714226 36993 714274
rect 0 713880 39573 714226
rect 0 700700 6278 713880
rect 19408 700700 39573 713880
rect 0 699374 39573 700700
rect 0 698800 20683 699374
rect 36343 699313 36993 699374
rect 0 671400 4843 698800
rect 0 670826 20683 671400
rect 21003 671146 25993 699054
rect 26313 671146 27163 699054
rect 27483 671146 28333 699054
rect 28653 671146 30453 699054
rect 30773 671146 31663 699054
rect 31983 698800 32632 699054
rect 31983 671400 32633 698800
rect 31983 671146 32632 671400
rect 32953 671146 33603 699054
rect 33923 671146 34813 699054
rect 35133 671146 36023 699054
rect 36343 671194 36993 698993
rect 37313 671146 38203 699054
rect 38523 671146 39573 699054
rect 678027 686746 679077 715454
rect 679397 686746 680287 715454
rect 680607 686807 681257 715406
rect 681577 686746 682467 715454
rect 682787 686746 683677 715454
rect 683997 686746 684647 715454
rect 684968 715200 685617 715454
rect 684967 687000 685617 715200
rect 684968 686746 685617 687000
rect 685937 686746 686827 715454
rect 687147 686746 688947 715454
rect 689267 686746 690117 715454
rect 690437 686746 691287 715454
rect 691607 686746 696597 715454
rect 696917 715200 717600 715774
rect 712757 687000 717600 715200
rect 680607 686426 681257 686487
rect 696917 686426 717600 687000
rect 678027 685100 717600 686426
rect 678027 671920 698192 685100
rect 711322 671920 717600 685100
rect 678027 671574 717600 671920
rect 680607 671526 681257 671574
rect 36343 670826 36993 670874
rect 0 670480 39573 670826
rect 0 657300 6278 670480
rect 19408 657300 39573 670480
rect 0 655974 39573 657300
rect 0 655400 20683 655974
rect 36343 655913 36993 655974
rect 0 628200 4843 655400
rect 0 627626 20683 628200
rect 21003 627946 25993 655654
rect 26313 627946 27163 655654
rect 27483 627946 28333 655654
rect 28653 627946 30453 655654
rect 30773 627946 31663 655654
rect 31983 655400 32632 655654
rect 31983 628200 32633 655400
rect 31983 627946 32632 628200
rect 32953 627946 33603 655654
rect 33923 627946 34813 655654
rect 35133 627946 36023 655654
rect 36343 627994 36993 655593
rect 37313 627946 38203 655654
rect 38523 627946 39573 655654
rect 678027 642546 679077 671254
rect 679397 642546 680287 671254
rect 680607 642607 681257 671206
rect 681577 642546 682467 671254
rect 682787 642546 683677 671254
rect 683997 642546 684647 671254
rect 684968 671000 685617 671254
rect 684967 642800 685617 671000
rect 684968 642546 685617 642800
rect 685937 642546 686827 671254
rect 687147 642546 688947 671254
rect 689267 642546 690117 671254
rect 690437 642546 691287 671254
rect 691607 642546 696597 671254
rect 696917 671000 717600 671574
rect 712757 642800 717600 671000
rect 680607 642226 681257 642287
rect 696917 642226 717600 642800
rect 678027 640900 717600 642226
rect 678027 627720 698192 640900
rect 711322 627720 717600 640900
rect 36343 627626 36993 627674
rect 0 627280 39573 627626
rect 678027 627374 717600 627720
rect 680607 627326 681257 627374
rect 0 614100 6278 627280
rect 19408 614100 39573 627280
rect 0 612774 39573 614100
rect 0 612200 20683 612774
rect 36343 612713 36993 612774
rect 0 585000 4843 612200
rect 0 584426 20683 585000
rect 21003 584746 25993 612454
rect 26313 584746 27163 612454
rect 27483 584746 28333 612454
rect 28653 584746 30453 612454
rect 30773 584746 31663 612454
rect 31983 612200 32632 612454
rect 31983 585000 32633 612200
rect 31983 584746 32632 585000
rect 32953 584746 33603 612454
rect 33923 584746 34813 612454
rect 35133 584746 36023 612454
rect 36343 584794 36993 612393
rect 37313 584746 38203 612454
rect 38523 584746 39573 612454
rect 678027 598146 679077 627054
rect 679397 598146 680287 627054
rect 680607 598207 681257 627006
rect 681577 598146 682467 627054
rect 682787 598146 683677 627054
rect 683997 598146 684647 627054
rect 684968 626800 685617 627054
rect 684967 598400 685617 626800
rect 684968 598146 685617 598400
rect 685937 598146 686827 627054
rect 687147 598146 688947 627054
rect 689267 598146 690117 627054
rect 690437 598146 691287 627054
rect 691607 598146 696597 627054
rect 696917 626800 717600 627374
rect 712757 598400 717600 626800
rect 680607 597826 681257 597887
rect 696917 597826 717600 598400
rect 678027 596500 717600 597826
rect 36343 584426 36993 584474
rect 0 584080 39573 584426
rect 0 570900 6278 584080
rect 19408 570900 39573 584080
rect 678027 583320 698192 596500
rect 711322 583320 717600 596500
rect 678027 582974 717600 583320
rect 680607 582926 681257 582974
rect 0 569574 39573 570900
rect 0 569000 20683 569574
rect 36343 569513 36993 569574
rect 0 541800 4843 569000
rect 0 541226 20683 541800
rect 21003 541546 25993 569254
rect 26313 541546 27163 569254
rect 27483 541546 28333 569254
rect 28653 541546 30453 569254
rect 30773 541546 31663 569254
rect 31983 569000 32632 569254
rect 31983 541800 32633 569000
rect 31983 541546 32632 541800
rect 32953 541546 33603 569254
rect 33923 541546 34813 569254
rect 35133 541546 36023 569254
rect 36343 541594 36993 569193
rect 37313 541546 38203 569254
rect 38523 541546 39573 569254
rect 678027 553946 679077 582654
rect 679397 553946 680287 582654
rect 680607 554007 681257 582606
rect 681577 553946 682467 582654
rect 682787 553946 683677 582654
rect 683997 553946 684647 582654
rect 684968 582400 685617 582654
rect 684967 554200 685617 582400
rect 684968 553946 685617 554200
rect 685937 553946 686827 582654
rect 687147 553946 688947 582654
rect 689267 553946 690117 582654
rect 690437 553946 691287 582654
rect 691607 553946 696597 582654
rect 696917 582400 717600 582974
rect 712757 554200 717600 582400
rect 680607 553626 681257 553687
rect 696917 553626 717600 554200
rect 678027 552300 717600 553626
rect 36343 541226 36993 541274
rect 0 540880 39573 541226
rect 0 527700 6278 540880
rect 19408 527700 39573 540880
rect 678027 539120 698192 552300
rect 711322 539120 717600 552300
rect 678027 538774 717600 539120
rect 680607 538726 681257 538774
rect 0 526374 39573 527700
rect 0 525800 20683 526374
rect 36343 526313 36993 526374
rect 0 498400 4843 525800
rect 0 497826 20683 498400
rect 21003 498146 25993 526054
rect 26313 498146 27163 526054
rect 27483 498146 28333 526054
rect 28653 498146 30453 526054
rect 30773 498146 31663 526054
rect 31983 525800 32632 526054
rect 31983 498146 32633 525800
rect 32953 498146 33603 526054
rect 33923 498146 34813 526054
rect 35133 498146 36023 526054
rect 36343 498207 36993 525993
rect 37313 498146 38203 526054
rect 38523 498146 39573 526054
rect 678027 509746 679077 538454
rect 679397 509746 680287 538454
rect 680607 509807 681257 538406
rect 681577 509746 682467 538454
rect 682787 509746 683677 538454
rect 683997 509746 684647 538454
rect 684968 538200 685617 538454
rect 684967 509746 685617 538200
rect 685937 509746 686827 538454
rect 687147 509746 688947 538454
rect 689267 509746 690117 538454
rect 690437 509746 691287 538454
rect 691607 509746 696597 538454
rect 696917 538200 717600 538774
rect 712757 510000 717600 538200
rect 680607 509426 681257 509487
rect 684967 509426 684968 509746
rect 696917 509426 717600 510000
rect 678027 508910 717600 509426
rect 32632 497826 32633 498146
rect 36343 497826 36993 497887
rect 0 497298 39573 497826
rect 0 484490 6491 497298
rect 19296 484490 39573 497298
rect 678027 496102 698304 508910
rect 711109 496102 717600 508910
rect 678027 495574 717600 496102
rect 680607 495513 681257 495574
rect 684967 495254 684968 495574
rect 0 483974 39573 484490
rect 0 483400 20683 483974
rect 32632 483654 32633 483974
rect 36343 483913 36993 483974
rect 0 456200 4843 483400
rect 0 455626 20683 456200
rect 21003 455946 25993 483654
rect 26313 455946 27163 483654
rect 27483 455946 28333 483654
rect 28653 455946 30453 483654
rect 30773 455946 31663 483654
rect 31983 456200 32633 483654
rect 31983 455946 32632 456200
rect 32953 455946 33603 483654
rect 33923 455946 34813 483654
rect 35133 455946 36023 483654
rect 36343 456007 36993 483593
rect 37313 455946 38203 483654
rect 38523 455946 39573 483654
rect 678027 466346 679077 495254
rect 679397 466346 680287 495254
rect 680607 466407 681257 495193
rect 681577 466346 682467 495254
rect 682787 466346 683677 495254
rect 683997 466346 684647 495254
rect 684967 466600 685617 495254
rect 684968 466346 685617 466600
rect 685937 466346 686827 495254
rect 687147 466346 688947 495254
rect 689267 466346 690117 495254
rect 690437 466346 691287 495254
rect 691607 466346 696597 495254
rect 696917 495000 717600 495574
rect 712757 466600 717600 495000
rect 680607 466026 681257 466087
rect 696917 466026 717600 466600
rect 678027 464866 717600 466026
rect 36343 455626 36993 455687
rect 0 454454 39573 455626
rect 0 442934 5847 454454
rect 19940 442934 39573 454454
rect 678027 453346 697660 464866
rect 711753 453346 717600 464866
rect 678027 452174 717600 453346
rect 680607 452113 681257 452174
rect 0 441774 39573 442934
rect 0 441200 20683 441774
rect 36343 441713 36993 441774
rect 0 414000 4843 441200
rect 0 413426 20683 414000
rect 21003 413746 25993 441454
rect 26313 413746 27163 441454
rect 27483 413746 28333 441454
rect 28653 413746 30453 441454
rect 30773 413746 31663 441454
rect 31983 441200 32632 441454
rect 31983 414000 32633 441200
rect 31983 413746 32632 414000
rect 32953 413746 33603 441454
rect 33923 413746 34813 441454
rect 35133 413746 36023 441454
rect 36343 413794 36993 441393
rect 37313 413746 38203 441454
rect 38523 413746 39573 441454
rect 678027 423146 679077 451854
rect 679397 423146 680287 451854
rect 680607 423207 681257 451793
rect 681577 423146 682467 451854
rect 682787 423146 683677 451854
rect 683997 423146 684647 451854
rect 684968 451600 685617 451854
rect 684967 423146 685617 451600
rect 685937 423146 686827 451854
rect 687147 423146 688947 451854
rect 689267 423146 690117 451854
rect 690437 423146 691287 451854
rect 691607 423146 696597 451854
rect 696917 451600 717600 452174
rect 712757 423400 717600 451600
rect 680607 422826 681257 422887
rect 684967 422826 684968 423146
rect 696917 422826 717600 423400
rect 678027 422310 717600 422826
rect 36343 413426 36993 413474
rect 0 413080 39573 413426
rect 0 399900 6278 413080
rect 19408 399900 39573 413080
rect 678027 409502 698304 422310
rect 711109 409502 717600 422310
rect 678027 408974 717600 409502
rect 680607 408913 681257 408974
rect 684967 408654 684968 408974
rect 0 398574 39573 399900
rect 0 398000 20683 398574
rect 36343 398513 36993 398574
rect 0 370800 4843 398000
rect 0 370226 20683 370800
rect 21003 370546 25993 398254
rect 26313 370546 27163 398254
rect 27483 370546 28333 398254
rect 28653 370546 30453 398254
rect 30773 370546 31663 398254
rect 31983 398000 32632 398254
rect 31983 370800 32633 398000
rect 31983 370546 32632 370800
rect 32953 370546 33603 398254
rect 33923 370546 34813 398254
rect 35133 370546 36023 398254
rect 36343 370594 36993 398193
rect 37313 370546 38203 398254
rect 38523 370546 39573 398254
rect 678027 379746 679077 408654
rect 679397 379746 680287 408654
rect 680607 379807 681257 408593
rect 681577 379746 682467 408654
rect 682787 379746 683677 408654
rect 683997 379746 684647 408654
rect 684967 380000 685617 408654
rect 684968 379746 685617 380000
rect 685937 379746 686827 408654
rect 687147 379746 688947 408654
rect 689267 379746 690117 408654
rect 690437 379746 691287 408654
rect 691607 379746 696597 408654
rect 696917 408400 717600 408974
rect 712757 380000 717600 408400
rect 680607 379426 681257 379487
rect 696917 379426 717600 380000
rect 678027 378100 717600 379426
rect 36343 370226 36993 370274
rect 0 369880 39573 370226
rect 0 356700 6278 369880
rect 19408 356700 39573 369880
rect 678027 364920 698192 378100
rect 711322 364920 717600 378100
rect 678027 364574 717600 364920
rect 680607 364526 681257 364574
rect 0 355374 39573 356700
rect 0 354800 20683 355374
rect 36343 355313 36993 355374
rect 0 327400 4843 354800
rect 0 326826 20683 327400
rect 21003 327146 25993 355054
rect 26313 327146 27163 355054
rect 27483 327146 28333 355054
rect 28653 327146 30453 355054
rect 30773 327146 31663 355054
rect 31983 354800 32632 355054
rect 31983 327400 32633 354800
rect 31983 327146 32632 327400
rect 32953 327146 33603 355054
rect 33923 327146 34813 355054
rect 35133 327146 36023 355054
rect 36343 327194 36993 354993
rect 37313 327146 38203 355054
rect 38523 327146 39573 355054
rect 678027 335546 679077 364254
rect 679397 335546 680287 364254
rect 680607 335607 681257 364206
rect 681577 335546 682467 364254
rect 682787 335546 683677 364254
rect 683997 335546 684647 364254
rect 684968 364000 685617 364254
rect 684967 335800 685617 364000
rect 684968 335546 685617 335800
rect 685937 335546 686827 364254
rect 687147 335546 688947 364254
rect 689267 335546 690117 364254
rect 690437 335546 691287 364254
rect 691607 335546 696597 364254
rect 696917 364000 717600 364574
rect 712757 335800 717600 364000
rect 680607 335226 681257 335287
rect 696917 335226 717600 335800
rect 678027 333900 717600 335226
rect 36343 326826 36993 326874
rect 0 326480 39573 326826
rect 0 313300 6278 326480
rect 19408 313300 39573 326480
rect 678027 320720 698192 333900
rect 711322 320720 717600 333900
rect 678027 320374 717600 320720
rect 680607 320326 681257 320374
rect 0 311974 39573 313300
rect 0 311400 20683 311974
rect 36343 311913 36993 311974
rect 0 284200 4843 311400
rect 0 283626 20683 284200
rect 21003 283946 25993 311654
rect 26313 283946 27163 311654
rect 27483 283946 28333 311654
rect 28653 283946 30453 311654
rect 30773 283946 31663 311654
rect 31983 311400 32632 311654
rect 31983 284200 32633 311400
rect 31983 283946 32632 284200
rect 32953 283946 33603 311654
rect 33923 283946 34813 311654
rect 35133 283946 36023 311654
rect 36343 283994 36993 311593
rect 37313 283946 38203 311654
rect 38523 283946 39573 311654
rect 678027 291346 679077 320054
rect 679397 291346 680287 320054
rect 680607 291407 681257 320006
rect 681577 291346 682467 320054
rect 682787 291346 683677 320054
rect 683997 291346 684647 320054
rect 684968 319800 685617 320054
rect 684967 291600 685617 319800
rect 684968 291346 685617 291600
rect 685937 291346 686827 320054
rect 687147 291346 688947 320054
rect 689267 291346 690117 320054
rect 690437 291346 691287 320054
rect 691607 291346 696597 320054
rect 696917 319800 717600 320374
rect 712757 291600 717600 319800
rect 680607 291026 681257 291087
rect 696917 291026 717600 291600
rect 678027 289700 717600 291026
rect 36343 283626 36993 283674
rect 0 283280 39573 283626
rect 0 270100 6278 283280
rect 19408 270100 39573 283280
rect 678027 276520 698192 289700
rect 711322 276520 717600 289700
rect 678027 276174 717600 276520
rect 680607 276126 681257 276174
rect 0 268774 39573 270100
rect 0 268200 20683 268774
rect 36343 268713 36993 268774
rect 0 241000 4843 268200
rect 0 240426 20683 241000
rect 21003 240746 25993 268454
rect 26313 240746 27163 268454
rect 27483 240746 28333 268454
rect 28653 240746 30453 268454
rect 30773 240746 31663 268454
rect 31983 268200 32632 268454
rect 31983 241000 32633 268200
rect 31983 240746 32632 241000
rect 32953 240746 33603 268454
rect 33923 240746 34813 268454
rect 35133 240746 36023 268454
rect 36343 240794 36993 268393
rect 37313 240746 38203 268454
rect 38523 240746 39573 268454
rect 678027 246946 679077 275854
rect 679397 246946 680287 275854
rect 680607 247007 681257 275806
rect 681577 246946 682467 275854
rect 682787 246946 683677 275854
rect 683997 246946 684647 275854
rect 684968 275600 685617 275854
rect 684967 247200 685617 275600
rect 684968 246946 685617 247200
rect 685937 246946 686827 275854
rect 687147 246946 688947 275854
rect 689267 246946 690117 275854
rect 690437 246946 691287 275854
rect 691607 246946 696597 275854
rect 696917 275600 717600 276174
rect 712757 247200 717600 275600
rect 680607 246626 681257 246687
rect 696917 246626 717600 247200
rect 678027 245300 717600 246626
rect 36343 240426 36993 240474
rect 0 240080 39573 240426
rect 0 226900 6278 240080
rect 19408 226900 39573 240080
rect 678027 232120 698192 245300
rect 711322 232120 717600 245300
rect 678027 231774 717600 232120
rect 680607 231726 681257 231774
rect 0 225574 39573 226900
rect 0 225000 20683 225574
rect 36343 225513 36993 225574
rect 0 197800 4843 225000
rect 0 197226 20683 197800
rect 21003 197546 25993 225254
rect 26313 197546 27163 225254
rect 27483 197546 28333 225254
rect 28653 197546 30453 225254
rect 30773 197546 31663 225254
rect 31983 225000 32632 225254
rect 31983 197800 32633 225000
rect 31983 197546 32632 197800
rect 32953 197546 33603 225254
rect 33923 197546 34813 225254
rect 35133 197546 36023 225254
rect 36343 197594 36993 225193
rect 37313 197546 38203 225254
rect 38523 197546 39573 225254
rect 678027 202746 679077 231454
rect 679397 202746 680287 231454
rect 680607 202807 681257 231406
rect 681577 202746 682467 231454
rect 682787 202746 683677 231454
rect 683997 202746 684647 231454
rect 684968 231200 685617 231454
rect 684967 203000 685617 231200
rect 684968 202746 685617 203000
rect 685937 202746 686827 231454
rect 687147 202746 688947 231454
rect 689267 202746 690117 231454
rect 690437 202746 691287 231454
rect 691607 202746 696597 231454
rect 696917 231200 717600 231774
rect 712757 203000 717600 231200
rect 680607 202426 681257 202487
rect 696917 202426 717600 203000
rect 678027 201100 717600 202426
rect 36343 197226 36993 197274
rect 0 196880 39573 197226
rect 0 183700 6278 196880
rect 19408 183700 39573 196880
rect 678027 187920 698192 201100
rect 711322 187920 717600 201100
rect 678027 187574 717600 187920
rect 680607 187526 681257 187574
rect 0 182374 39573 183700
rect 0 181800 20683 182374
rect 36343 182313 36993 182374
rect 0 125200 4843 181800
rect 0 124626 20683 125200
rect 21003 124946 25993 182054
rect 26313 124946 27163 182054
rect 27483 124946 28333 182054
rect 28653 153400 30453 182054
rect 30773 154400 31663 182054
rect 31983 181800 32632 182054
rect 31983 153400 32633 181800
rect 28653 124946 30453 152400
rect 30773 124946 31663 153400
rect 31983 124946 32633 152400
rect 32953 124946 33603 182054
rect 33923 124946 34813 182054
rect 35133 124946 36023 182054
rect 36343 153400 36993 181993
rect 37313 154400 38203 182054
rect 36343 125007 36993 152400
rect 37313 124946 38203 153400
rect 38523 124946 39573 182054
rect 678027 158546 679077 187254
rect 679397 158546 680287 187254
rect 680607 158607 681257 187206
rect 681577 158546 682467 187254
rect 682787 158546 683677 187254
rect 683997 158546 684647 187254
rect 684968 187000 685617 187254
rect 684967 158800 685617 187000
rect 684968 158546 685617 158800
rect 685937 158546 686827 187254
rect 687147 158546 688947 187254
rect 689267 158546 690117 187254
rect 690437 158546 691287 187254
rect 691607 158546 696597 187254
rect 696917 187000 717600 187574
rect 712757 158800 717600 187000
rect 680607 158226 681257 158287
rect 696917 158226 717600 158800
rect 678027 156900 717600 158226
rect 678027 143720 698192 156900
rect 711322 143720 717600 156900
rect 678027 143374 717600 143720
rect 680607 143326 681257 143374
rect 32632 124626 32633 124946
rect 36343 124626 36993 124687
rect 0 124098 39573 124626
rect 0 111290 6491 124098
rect 19296 111290 39573 124098
rect 678027 114146 679077 143054
rect 679397 114146 680287 143054
rect 680607 114207 681257 143006
rect 681577 114146 682467 143054
rect 682787 114146 683677 143054
rect 683997 114146 684647 143054
rect 684968 142800 685617 143054
rect 684967 114400 685617 142800
rect 684968 114146 685617 114400
rect 685937 114146 686827 143054
rect 687147 114146 688947 143054
rect 689267 114146 690117 143054
rect 690437 114146 691287 143054
rect 691607 114146 696597 143054
rect 696917 142800 717600 143374
rect 712757 114400 717600 142800
rect 680607 113826 681257 113887
rect 696917 113826 717600 114400
rect 0 110774 39573 111290
rect 678027 112500 717600 113826
rect 0 110200 20683 110774
rect 32632 110454 32633 110774
rect 36343 110713 36993 110774
rect 0 83000 4843 110200
rect 0 82426 20683 83000
rect 21003 82746 25993 110454
rect 26313 82746 27163 110454
rect 27483 82746 28333 110454
rect 28653 82746 30453 110454
rect 30773 82746 31663 110454
rect 31983 82746 32633 110454
rect 32953 82746 33603 110454
rect 33923 82746 34813 110454
rect 35133 82746 36023 110454
rect 36343 82807 36993 110393
rect 37313 82746 38203 110454
rect 38523 82746 39573 110454
rect 678027 99320 698192 112500
rect 711322 99320 717600 112500
rect 678027 98974 717600 99320
rect 680607 98926 681257 98974
rect 32632 82426 32633 82746
rect 36343 82426 36993 82487
rect 0 81254 39573 82426
rect 0 69734 5847 81254
rect 19940 69734 39573 81254
rect 0 68574 39573 69734
rect 0 68000 20683 68574
rect 32632 68254 32633 68574
rect 36343 68513 36993 68574
rect 0 40800 4843 68000
rect 0 40109 20683 40800
rect 21003 40429 25993 68254
rect 26313 40546 27163 68254
rect 27483 40546 28333 68254
rect 26313 40109 28333 40226
rect 0 35049 28333 40109
rect 28653 35369 30453 68254
rect 30773 40546 31663 68254
rect 31983 40800 32633 68254
rect 31983 40546 32632 40800
rect 32953 40546 33603 68254
rect 33923 40546 34813 68254
rect 35133 40546 36023 68254
rect 36343 40549 36993 68193
rect 37313 40546 38203 68254
rect 38523 40546 39573 68254
rect 36343 40226 36993 40229
rect 39893 40226 40000 40800
rect 30773 39893 40000 40226
rect 676800 39893 677707 40000
rect 30773 38523 39210 39893
rect 39530 38523 79054 39573
rect 30773 36993 38923 38523
rect 47400 38203 71400 38523
rect 39243 37313 79054 38203
rect 79374 36993 93226 39573
rect 93546 38523 132854 39573
rect 101200 38203 125200 38523
rect 93546 37313 132854 38203
rect 133174 36993 147026 39573
rect 147346 38523 186654 39573
rect 155000 38203 179000 38523
rect 147346 37313 186654 38203
rect 186974 36993 201826 39573
rect 202146 38523 241454 39573
rect 209800 38203 233800 38523
rect 202146 37313 241454 38203
rect 241774 36993 255626 39573
rect 255946 38523 295254 39573
rect 263600 38203 287600 38523
rect 255946 37313 295254 38203
rect 295574 36993 310426 39573
rect 310746 38523 350054 39573
rect 318400 38203 342400 38523
rect 310746 37313 350054 38203
rect 350374 36993 365226 39573
rect 365546 38523 404854 39573
rect 373200 38203 397200 38523
rect 365546 37313 404854 38203
rect 405174 36993 420026 39573
rect 420346 38523 459654 39573
rect 428000 38203 452000 38523
rect 420346 37313 459654 38203
rect 459974 36993 474826 39573
rect 475146 38523 514454 39573
rect 482800 38203 506800 38523
rect 475146 37313 514454 38203
rect 514774 36993 529626 39573
rect 529946 38523 569254 39573
rect 537600 38203 561600 38523
rect 529946 37313 569254 38203
rect 569574 36993 583426 39573
rect 583746 38523 623054 39573
rect 591400 38203 615400 38523
rect 583746 37313 623054 38203
rect 623374 36993 637226 39573
rect 637546 38523 677054 39573
rect 677374 39210 677707 39893
rect 678027 39530 679077 98654
rect 679397 70200 680287 98654
rect 680607 69200 681257 98606
rect 679397 39243 680287 69200
rect 680607 39706 681257 68200
rect 681577 39695 682467 98654
rect 682787 39680 683677 98654
rect 683997 39723 684647 98654
rect 684968 98400 685617 98654
rect 684967 69200 685617 98400
rect 685937 70200 686827 98654
rect 687147 69200 688947 98654
rect 684967 39733 685617 68200
rect 685937 39705 686827 69200
rect 684967 39403 685617 39413
rect 680607 39375 681257 39386
rect 683997 39385 685617 39403
rect 680607 39360 682467 39375
rect 683997 39360 686827 39385
rect 677374 38923 679077 39210
rect 680607 38923 686827 39360
rect 645200 38203 669200 38523
rect 637546 37313 677054 38203
rect 677374 36993 686827 38923
rect 30773 36343 39386 36993
rect 39706 36343 78993 36993
rect 79313 36343 93287 36993
rect 93607 36343 132793 36993
rect 133113 36343 147087 36993
rect 147407 36343 186606 36993
rect 186926 36343 201887 36993
rect 202207 36343 241393 36993
rect 241713 36343 255687 36993
rect 256007 36343 295206 36993
rect 295526 36343 310487 36993
rect 310807 36343 350006 36993
rect 350326 36343 365287 36993
rect 365607 36343 404806 36993
rect 405126 36343 420087 36993
rect 420407 36343 459606 36993
rect 459926 36343 474887 36993
rect 475207 36343 514406 36993
rect 514726 36343 529687 36993
rect 530007 36343 569193 36993
rect 569513 36343 583487 36993
rect 583807 36343 622993 36993
rect 623313 36343 637287 36993
rect 637607 36343 677051 36993
rect 677371 36343 686827 36993
rect 30773 35133 39375 36343
rect 39695 35133 79054 36023
rect 30773 35049 39360 35133
rect 0 33603 39360 35049
rect 39680 33923 79054 34813
rect 0 32633 39403 33603
rect 39723 32953 79054 33603
rect 79374 32633 93226 36343
rect 93546 35133 132854 36023
rect 93546 33923 132854 34813
rect 93546 32953 132854 33603
rect 0 31983 39413 32633
rect 39733 32632 132600 32633
rect 39733 31983 79054 32632
rect 0 30773 39385 31983
rect 39705 30773 79054 31663
rect 0 28333 35049 30773
rect 35369 28653 79054 30453
rect 0 27163 39355 28333
rect 39675 27483 79054 28333
rect 0 26313 39384 27163
rect 39704 26313 79054 27163
rect 0 20683 39151 26313
rect 39471 21003 79054 25993
rect 79374 20683 93226 32632
rect 93546 31983 132854 32632
rect 93546 30773 132854 31663
rect 93546 28653 132854 30453
rect 93546 27483 132854 28333
rect 93546 26313 132854 27163
rect 93546 21003 132854 25993
rect 133174 20683 147026 36343
rect 147346 35133 186654 36023
rect 147346 33923 186654 34813
rect 147346 32953 186654 33603
rect 147600 32632 186400 32633
rect 147346 31983 186654 32632
rect 147346 30773 186654 31663
rect 147346 28653 186654 30453
rect 147346 27483 186654 28333
rect 147346 26313 186654 27163
rect 147346 21003 186654 25993
rect 186974 20683 201826 36343
rect 202146 35133 241454 36023
rect 202146 33923 241454 34813
rect 202146 32953 241454 33603
rect 241774 32633 255626 36343
rect 255946 35133 295254 36023
rect 255946 33923 295254 34813
rect 255946 32953 295254 33603
rect 202400 32632 295000 32633
rect 202146 31983 241454 32632
rect 202146 30773 241454 31663
rect 202146 28653 241454 30453
rect 202146 27483 241454 28333
rect 202146 26313 241454 27163
rect 202146 21003 241454 25993
rect 241774 20683 255626 32632
rect 255946 31983 295254 32632
rect 255946 30773 295254 31663
rect 255946 28653 295254 30453
rect 255946 27483 295254 28333
rect 255946 26313 295254 27163
rect 255946 21003 295254 25993
rect 295574 20683 310426 36343
rect 310746 35133 350054 36023
rect 310746 33923 350054 34813
rect 310746 32953 350054 33603
rect 311000 32632 349800 32633
rect 310746 31983 350054 32632
rect 310746 30773 350054 31663
rect 310746 28653 350054 30453
rect 310746 27483 350054 28333
rect 310746 26313 350054 27163
rect 310746 21003 350054 25993
rect 350374 20683 365226 36343
rect 365546 35133 404854 36023
rect 365546 33923 404854 34813
rect 365546 32953 404854 33603
rect 365800 32632 404600 32633
rect 365546 31983 404854 32632
rect 365546 30773 404854 31663
rect 365546 28653 404854 30453
rect 365546 27483 404854 28333
rect 365546 26313 404854 27163
rect 365546 21003 404854 25993
rect 405174 20683 420026 36343
rect 420346 35133 459654 36023
rect 420346 33923 459654 34813
rect 420346 32953 459654 33603
rect 420600 32632 459400 32633
rect 420346 31983 459654 32632
rect 420346 30773 459654 31663
rect 420346 28653 459654 30453
rect 420346 27483 459654 28333
rect 420346 26313 459654 27163
rect 420346 21003 459654 25993
rect 459974 20683 474826 36343
rect 475146 35133 514454 36023
rect 475146 33923 514454 34813
rect 475146 32953 514454 33603
rect 475400 32632 514200 32633
rect 475146 31983 514454 32632
rect 475146 30773 514454 31663
rect 475146 28653 514454 30453
rect 475146 27483 514454 28333
rect 475146 26313 514454 27163
rect 475146 21003 514454 25993
rect 514774 20683 529626 36343
rect 529946 35133 569254 36023
rect 529946 33923 569254 34813
rect 529946 32953 569254 33603
rect 569574 32633 583426 36343
rect 583746 35133 623054 36023
rect 583746 33923 623054 34813
rect 583746 32953 623054 33603
rect 623374 32633 637226 36343
rect 637546 35133 677054 36023
rect 677374 35049 686827 36343
rect 687147 35369 688947 68200
rect 689267 39675 690117 98654
rect 690437 39704 691287 98654
rect 691607 39471 696597 98654
rect 696917 98400 717600 98974
rect 712757 40000 717600 98400
rect 690437 39355 691287 39384
rect 689267 39151 691287 39355
rect 696917 39151 717600 40000
rect 689267 35049 717600 39151
rect 637546 33923 677054 34813
rect 637546 32953 677054 33603
rect 530200 32632 676800 32633
rect 529946 31983 569254 32632
rect 529946 30773 569254 31663
rect 529946 28653 569254 30453
rect 529946 27483 569254 28333
rect 529946 26313 569254 27163
rect 529946 21003 569254 25993
rect 569574 20683 583426 32632
rect 583746 31983 623054 32632
rect 583746 30773 623054 31663
rect 583746 28653 623054 30453
rect 583746 27483 623054 28333
rect 583746 26313 623054 27163
rect 583746 21003 623054 25993
rect 623374 20683 637226 32632
rect 637546 31983 677054 32632
rect 637546 30773 677054 31663
rect 677374 30773 717600 35049
rect 637546 28653 682231 30453
rect 682551 28333 717600 30773
rect 637546 27483 677054 28333
rect 637546 26313 677054 27163
rect 677374 26313 717600 28333
rect 637546 21003 677171 25993
rect 677491 20683 717600 26313
rect 0 4843 40000 20683
rect 78800 19296 93800 20683
rect 78800 6491 79902 19296
rect 92710 6491 93800 19296
rect 78800 4843 93800 6491
rect 132600 18629 147600 20683
rect 132600 6823 136393 18629
rect 144470 6823 147600 18629
rect 132600 5163 147600 6823
rect 186400 19408 202400 20683
rect 186400 6278 187320 19408
rect 200500 6278 202400 19408
rect 0 0 132854 4843
rect 133174 0 147026 5163
rect 186400 4843 202400 6278
rect 241200 19940 256200 20683
rect 241200 5847 242946 19940
rect 254466 5847 256200 19940
rect 241200 4843 256200 5847
rect 295000 19408 311000 20683
rect 295000 6278 295920 19408
rect 309100 6278 311000 19408
rect 295000 4843 311000 6278
rect 349800 19408 365800 20683
rect 349800 6278 350720 19408
rect 363900 6278 365800 19408
rect 349800 4843 365800 6278
rect 404600 19408 420600 20683
rect 404600 6278 405520 19408
rect 418700 6278 420600 19408
rect 404600 4843 420600 6278
rect 459400 19408 475400 20683
rect 459400 6278 460320 19408
rect 473500 6278 475400 19408
rect 459400 4843 475400 6278
rect 514200 19408 530200 20683
rect 514200 6278 515120 19408
rect 528300 6278 530200 19408
rect 514200 4843 530200 6278
rect 569000 19296 584000 20683
rect 569000 6491 570102 19296
rect 582910 6491 584000 19296
rect 569000 4843 584000 6491
rect 622800 19296 637800 20683
rect 622800 6491 623902 19296
rect 636710 6491 637800 19296
rect 622800 4843 637800 6491
rect 676800 4843 717600 20683
rect 147346 0 717600 4843
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 1 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 2 nsew signal output
rlabel metal2 s 194043 41713 194099 42193 6 por
port 3 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 4 nsew signal output
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 5 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 6 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 7 nsew signal input
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 8 nsew signal output
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 9 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 10 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 11 nsew signal input
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 12 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 13 nsew signal output
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 14 nsew signal input
rlabel metal2 s 415371 41713 415427 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41754 415268 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41806 415427 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412364 41754 412416 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41713 412299 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41806 412416 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409328 41754 409380 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41713 409263 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41806 409380 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415228 41818 415427 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41818 412404 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41818 409368 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415371 41834 415427 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41834 412299 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41834 409263 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 415216 41760 415268 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 412364 41760 412416 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 409328 41760 409380 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41760 415274 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41760 412422 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41760 409386 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41772 415274 41800 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41800 415274 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41800 412422 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41800 409386 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal3 s 419717 44235 419783 44238 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 419490 44238 419783 44298 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 419717 44298 419783 44301 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 419490 44298 419550 44374 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44371 411135 44374 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44374 419550 44434 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal3 s 411069 44434 411135 44437 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via2 s 419722 44240 419778 44296 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via2 s 411074 44376 411130 44432 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419695 41713 419751 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41713 411103 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419695 41820 419764 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41820 411116 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419736 42193 419764 44231 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419722 44231 419778 44305 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411088 42193 411116 44367 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411074 44367 411130 44441 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 17 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 18 nsew signal output
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 19 nsew signal input
rlabel metal2 s 470171 41713 470227 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41754 470100 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41806 470227 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467196 41754 467248 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41713 467099 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41806 467248 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464160 41754 464212 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41713 464063 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41806 464212 41818 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470060 41818 470227 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41818 467236 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41818 464200 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470171 41834 470227 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41834 467099 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41834 464063 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 470048 41760 470100 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 467196 41760 467248 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 464160 41760 464212 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41760 470106 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41760 467254 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41760 464218 41772 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41772 470106 41800 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41800 470106 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41800 467254 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41800 464218 41812 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal3 s 474457 44371 474523 44374 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44371 465875 44374 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44374 474523 44434 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 474457 44434 474523 44437 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44434 465875 44437 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 474462 44376 474518 44432 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 465814 44376 465870 44432 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474495 41713 474551 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465847 41713 465903 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 41806 474551 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 41806 465903 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 42193 474504 44367 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 42193 465856 44367 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474462 44367 474518 44441 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465814 44367 465870 44441 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 22 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 23 nsew signal output
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 24 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 25 nsew signal input
rlabel metal3 s 524965 44235 525031 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44235 518867 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44238 525031 44298 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 524965 44298 525031 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44298 518867 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 524970 44240 525026 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 518806 44240 518862 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518807 41713 518863 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524984 42193 525012 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518820 42193 518848 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524970 44231 525026 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518806 44231 518862 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 27 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 28 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd_pad
port 29 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda_pad
port 30 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio_pad
port 31 nsew signal bidirectional
rlabel metal5 s 6811 872210 18976 884378 6 vddio_pad2
port 32 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa_pad
port 33 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd_pad
port 34 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio_pad
port 35 nsew signal bidirectional
rlabel metal5 s 340810 1018624 352978 1030789 6 vssio_pad2
port 36 nsew signal bidirectional
rlabel metal5 s 698512 99640 711002 112180 6 mprj_io[0]
port 37 nsew signal bidirectional
rlabel metal2 s 675407 104203 675887 104259 6 mprj_io_analog_en[0]
port 38 nsew signal input
rlabel metal2 s 675407 105491 675887 105547 6 mprj_io_analog_pol[0]
port 39 nsew signal input
rlabel metal2 s 675407 108527 675887 108583 6 mprj_io_analog_sel[0]
port 40 nsew signal input
rlabel metal2 s 675407 104847 675887 104903 6 mprj_io_dm[0]
port 41 nsew signal input
rlabel metal2 s 675407 103007 675887 103063 6 mprj_io_dm[1]
port 42 nsew signal input
rlabel metal2 s 675407 109171 675887 109227 6 mprj_io_dm[2]
port 43 nsew signal input
rlabel metal2 s 675407 109815 675887 109871 6 mprj_io_holdover[0]
port 44 nsew signal input
rlabel metal2 s 675407 112851 675887 112907 6 mprj_io_ib_mode_sel[0]
port 45 nsew signal input
rlabel metal2 s 675407 106043 675887 106099 6 mprj_io_inp_dis[0]
port 46 nsew signal input
rlabel metal2 s 675407 113495 675887 113551 6 mprj_io_oeb[0]
port 47 nsew signal input
rlabel metal2 s 675407 110367 675887 110423 6 mprj_io_out[0]
port 48 nsew signal input
rlabel metal2 s 675407 101167 675887 101223 6 mprj_io_slow_sel[0]
port 49 nsew signal input
rlabel metal2 s 675407 112207 675887 112263 6 mprj_io_vtrip_sel[0]
port 50 nsew signal input
rlabel metal2 s 675407 99327 675887 99383 6 mprj_io_in[0]
port 51 nsew signal output
rlabel metal2 s 675407 114047 675887 114103 6 mprj_io_in_3v3[0]
port 52 nsew signal output
rlabel metal2 s 675407 674411 675887 674467 6 mprj_gpio_analog[3]
port 53 nsew signal bidirectional
rlabel metal2 s 675407 676251 675887 676307 6 mprj_gpio_noesd[3]
port 54 nsew signal bidirectional
rlabel metal5 s 698512 672240 711002 684780 6 mprj_io[10]
port 55 nsew signal bidirectional
rlabel metal2 s 675407 676803 675887 676859 6 mprj_io_analog_en[10]
port 56 nsew signal input
rlabel metal2 s 675407 678091 675887 678147 6 mprj_io_analog_pol[10]
port 57 nsew signal input
rlabel metal2 s 675407 681127 675887 681183 6 mprj_io_analog_sel[10]
port 58 nsew signal input
rlabel metal2 s 675407 677447 675887 677503 6 mprj_io_dm[30]
port 59 nsew signal input
rlabel metal2 s 675407 675607 675887 675663 6 mprj_io_dm[31]
port 60 nsew signal input
rlabel metal2 s 675407 681771 675887 681827 6 mprj_io_dm[32]
port 61 nsew signal input
rlabel metal2 s 675407 682415 675887 682471 6 mprj_io_holdover[10]
port 62 nsew signal input
rlabel metal2 s 675407 685451 675887 685507 6 mprj_io_ib_mode_sel[10]
port 63 nsew signal input
rlabel metal2 s 675407 678643 675887 678699 6 mprj_io_inp_dis[10]
port 64 nsew signal input
rlabel metal2 s 675407 686095 675887 686151 6 mprj_io_oeb[10]
port 65 nsew signal input
rlabel metal2 s 675407 682967 675887 683023 6 mprj_io_out[10]
port 66 nsew signal input
rlabel metal2 s 675407 673767 675887 673823 6 mprj_io_slow_sel[10]
port 67 nsew signal input
rlabel metal2 s 675407 684807 675887 684863 6 mprj_io_vtrip_sel[10]
port 68 nsew signal input
rlabel metal2 s 675407 671927 675887 671983 6 mprj_io_in[10]
port 69 nsew signal output
rlabel metal2 s 675407 686647 675887 686703 6 mprj_io_in_3v3[10]
port 70 nsew signal output
rlabel metal2 s 675407 718611 675887 718667 6 mprj_gpio_analog[4]
port 71 nsew signal bidirectional
rlabel metal2 s 675407 720451 675887 720507 6 mprj_gpio_noesd[4]
port 72 nsew signal bidirectional
rlabel metal5 s 698512 716440 711002 728980 6 mprj_io[11]
port 73 nsew signal bidirectional
rlabel metal2 s 675407 721003 675887 721059 6 mprj_io_analog_en[11]
port 74 nsew signal input
rlabel metal2 s 675407 722291 675887 722347 6 mprj_io_analog_pol[11]
port 75 nsew signal input
rlabel metal2 s 675407 725327 675887 725383 6 mprj_io_analog_sel[11]
port 76 nsew signal input
rlabel metal2 s 675407 721647 675887 721703 6 mprj_io_dm[33]
port 77 nsew signal input
rlabel metal2 s 675407 719807 675887 719863 6 mprj_io_dm[34]
port 78 nsew signal input
rlabel metal2 s 675407 725971 675887 726027 6 mprj_io_dm[35]
port 79 nsew signal input
rlabel metal2 s 675407 726615 675887 726671 6 mprj_io_holdover[11]
port 80 nsew signal input
rlabel metal2 s 675407 729651 675887 729707 6 mprj_io_ib_mode_sel[11]
port 81 nsew signal input
rlabel metal2 s 675407 722843 675887 722899 6 mprj_io_inp_dis[11]
port 82 nsew signal input
rlabel metal2 s 675407 730295 675887 730351 6 mprj_io_oeb[11]
port 83 nsew signal input
rlabel metal2 s 675407 727167 675887 727223 6 mprj_io_out[11]
port 84 nsew signal input
rlabel metal2 s 675407 717967 675887 718023 6 mprj_io_slow_sel[11]
port 85 nsew signal input
rlabel metal2 s 675407 729007 675887 729063 6 mprj_io_vtrip_sel[11]
port 86 nsew signal input
rlabel metal2 s 675407 716127 675887 716183 6 mprj_io_in[11]
port 87 nsew signal output
rlabel metal2 s 675407 730847 675887 730903 6 mprj_io_in_3v3[11]
port 88 nsew signal output
rlabel metal2 s 675407 763011 675887 763067 6 mprj_gpio_analog[5]
port 89 nsew signal bidirectional
rlabel metal2 s 675407 764851 675887 764907 6 mprj_gpio_noesd[5]
port 90 nsew signal bidirectional
rlabel metal5 s 698512 760840 711002 773380 6 mprj_io[12]
port 91 nsew signal bidirectional
rlabel metal2 s 675407 765403 675887 765459 6 mprj_io_analog_en[12]
port 92 nsew signal input
rlabel metal2 s 675407 766691 675887 766747 6 mprj_io_analog_pol[12]
port 93 nsew signal input
rlabel metal2 s 675407 769727 675887 769783 6 mprj_io_analog_sel[12]
port 94 nsew signal input
rlabel metal2 s 675407 766047 675887 766103 6 mprj_io_dm[36]
port 95 nsew signal input
rlabel metal2 s 675407 764207 675887 764263 6 mprj_io_dm[37]
port 96 nsew signal input
rlabel metal2 s 675407 770371 675887 770427 6 mprj_io_dm[38]
port 97 nsew signal input
rlabel metal2 s 675407 771015 675887 771071 6 mprj_io_holdover[12]
port 98 nsew signal input
rlabel metal2 s 675407 774051 675887 774107 6 mprj_io_ib_mode_sel[12]
port 99 nsew signal input
rlabel metal2 s 675407 767243 675887 767299 6 mprj_io_inp_dis[12]
port 100 nsew signal input
rlabel metal2 s 675407 774695 675887 774751 6 mprj_io_oeb[12]
port 101 nsew signal input
rlabel metal2 s 675407 771567 675887 771623 6 mprj_io_out[12]
port 102 nsew signal input
rlabel metal2 s 675407 762367 675887 762423 6 mprj_io_slow_sel[12]
port 103 nsew signal input
rlabel metal2 s 675407 773407 675887 773463 6 mprj_io_vtrip_sel[12]
port 104 nsew signal input
rlabel metal2 s 675407 760527 675887 760583 6 mprj_io_in[12]
port 105 nsew signal output
rlabel metal2 s 675407 775247 675887 775303 6 mprj_io_in_3v3[12]
port 106 nsew signal output
rlabel metal2 s 675407 850411 675887 850467 6 mprj_gpio_analog[6]
port 107 nsew signal bidirectional
rlabel metal2 s 675407 852251 675887 852307 6 mprj_gpio_noesd[6]
port 108 nsew signal bidirectional
rlabel metal5 s 698512 848240 711002 860780 6 mprj_io[13]
port 109 nsew signal bidirectional
rlabel metal2 s 675407 852803 675887 852859 6 mprj_io_analog_en[13]
port 110 nsew signal input
rlabel metal2 s 675407 854091 675887 854147 6 mprj_io_analog_pol[13]
port 111 nsew signal input
rlabel metal2 s 675407 857127 675887 857183 6 mprj_io_analog_sel[13]
port 112 nsew signal input
rlabel metal2 s 675407 853447 675887 853503 6 mprj_io_dm[39]
port 113 nsew signal input
rlabel metal2 s 675407 851607 675887 851663 6 mprj_io_dm[40]
port 114 nsew signal input
rlabel metal2 s 675407 857771 675887 857827 6 mprj_io_dm[41]
port 115 nsew signal input
rlabel metal2 s 675407 858415 675887 858471 6 mprj_io_holdover[13]
port 116 nsew signal input
rlabel metal2 s 675407 861451 675887 861507 6 mprj_io_ib_mode_sel[13]
port 117 nsew signal input
rlabel metal2 s 675407 854643 675887 854699 6 mprj_io_inp_dis[13]
port 118 nsew signal input
rlabel metal2 s 675407 862095 675887 862151 6 mprj_io_oeb[13]
port 119 nsew signal input
rlabel metal2 s 675407 858967 675887 859023 6 mprj_io_out[13]
port 120 nsew signal input
rlabel metal2 s 675407 849767 675887 849823 6 mprj_io_slow_sel[13]
port 121 nsew signal input
rlabel metal2 s 675407 860807 675887 860863 6 mprj_io_vtrip_sel[13]
port 122 nsew signal input
rlabel metal2 s 675407 847927 675887 847983 6 mprj_io_in[13]
port 123 nsew signal output
rlabel metal2 s 675407 862647 675887 862703 6 mprj_io_in_3v3[13]
port 124 nsew signal output
rlabel metal5 s 698512 144040 711002 156580 6 mprj_io[1]
port 125 nsew signal bidirectional
rlabel metal2 s 675407 148603 675887 148659 6 mprj_io_analog_en[1]
port 126 nsew signal input
rlabel metal2 s 675407 149891 675887 149947 6 mprj_io_analog_pol[1]
port 127 nsew signal input
rlabel metal2 s 675407 152927 675887 152983 6 mprj_io_analog_sel[1]
port 128 nsew signal input
rlabel metal2 s 675407 149247 675887 149303 6 mprj_io_dm[3]
port 129 nsew signal input
rlabel metal2 s 675407 147407 675887 147463 6 mprj_io_dm[4]
port 130 nsew signal input
rlabel metal2 s 675407 153571 675887 153627 6 mprj_io_dm[5]
port 131 nsew signal input
rlabel metal2 s 675407 154215 675887 154271 6 mprj_io_holdover[1]
port 132 nsew signal input
rlabel metal2 s 675407 157251 675887 157307 6 mprj_io_ib_mode_sel[1]
port 133 nsew signal input
rlabel metal2 s 675407 150443 675887 150499 6 mprj_io_inp_dis[1]
port 134 nsew signal input
rlabel metal2 s 675407 157895 675887 157951 6 mprj_io_oeb[1]
port 135 nsew signal input
rlabel metal2 s 675407 154767 675887 154823 6 mprj_io_out[1]
port 136 nsew signal input
rlabel metal2 s 675407 145567 675887 145623 6 mprj_io_slow_sel[1]
port 137 nsew signal input
rlabel metal2 s 675407 156607 675887 156663 6 mprj_io_vtrip_sel[1]
port 138 nsew signal input
rlabel metal2 s 675407 143727 675887 143783 6 mprj_io_in[1]
port 139 nsew signal output
rlabel metal2 s 675407 158447 675887 158503 6 mprj_io_in_3v3[1]
port 140 nsew signal output
rlabel metal5 s 698512 188240 711002 200780 6 mprj_io[2]
port 141 nsew signal bidirectional
rlabel metal2 s 675407 192803 675887 192859 6 mprj_io_analog_en[2]
port 142 nsew signal input
rlabel metal2 s 675407 194091 675887 194147 6 mprj_io_analog_pol[2]
port 143 nsew signal input
rlabel metal2 s 675407 197127 675887 197183 6 mprj_io_analog_sel[2]
port 144 nsew signal input
rlabel metal2 s 675407 193447 675887 193503 6 mprj_io_dm[6]
port 145 nsew signal input
rlabel metal2 s 675407 191607 675887 191663 6 mprj_io_dm[7]
port 146 nsew signal input
rlabel metal2 s 675407 197771 675887 197827 6 mprj_io_dm[8]
port 147 nsew signal input
rlabel metal2 s 675407 198415 675887 198471 6 mprj_io_holdover[2]
port 148 nsew signal input
rlabel metal2 s 675407 201451 675887 201507 6 mprj_io_ib_mode_sel[2]
port 149 nsew signal input
rlabel metal2 s 675407 194643 675887 194699 6 mprj_io_inp_dis[2]
port 150 nsew signal input
rlabel metal2 s 675407 202095 675887 202151 6 mprj_io_oeb[2]
port 151 nsew signal input
rlabel metal2 s 675407 198967 675887 199023 6 mprj_io_out[2]
port 152 nsew signal input
rlabel metal2 s 675407 189767 675887 189823 6 mprj_io_slow_sel[2]
port 153 nsew signal input
rlabel metal2 s 675407 200807 675887 200863 6 mprj_io_vtrip_sel[2]
port 154 nsew signal input
rlabel metal2 s 675407 187927 675887 187983 6 mprj_io_in[2]
port 155 nsew signal output
rlabel metal2 s 675407 202647 675887 202703 6 mprj_io_in_3v3[2]
port 156 nsew signal output
rlabel metal5 s 698512 232440 711002 244980 6 mprj_io[3]
port 157 nsew signal bidirectional
rlabel metal2 s 675407 237003 675887 237059 6 mprj_io_analog_en[3]
port 158 nsew signal input
rlabel metal2 s 675407 238291 675887 238347 6 mprj_io_analog_pol[3]
port 159 nsew signal input
rlabel metal2 s 675407 241327 675887 241383 6 mprj_io_analog_sel[3]
port 160 nsew signal input
rlabel metal2 s 675407 235807 675887 235863 6 mprj_io_dm[10]
port 161 nsew signal input
rlabel metal2 s 675407 241971 675887 242027 6 mprj_io_dm[11]
port 162 nsew signal input
rlabel metal2 s 675407 237647 675887 237703 6 mprj_io_dm[9]
port 163 nsew signal input
rlabel metal2 s 675407 242615 675887 242671 6 mprj_io_holdover[3]
port 164 nsew signal input
rlabel metal2 s 675407 245651 675887 245707 6 mprj_io_ib_mode_sel[3]
port 165 nsew signal input
rlabel metal2 s 675407 238843 675887 238899 6 mprj_io_inp_dis[3]
port 166 nsew signal input
rlabel metal2 s 675407 246295 675887 246351 6 mprj_io_oeb[3]
port 167 nsew signal input
rlabel metal2 s 675407 243167 675887 243223 6 mprj_io_out[3]
port 168 nsew signal input
rlabel metal2 s 675407 233967 675887 234023 6 mprj_io_slow_sel[3]
port 169 nsew signal input
rlabel metal2 s 675407 245007 675887 245063 6 mprj_io_vtrip_sel[3]
port 170 nsew signal input
rlabel metal2 s 675407 232127 675887 232183 6 mprj_io_in[3]
port 171 nsew signal output
rlabel metal2 s 675407 246847 675887 246903 6 mprj_io_in_3v3[3]
port 172 nsew signal output
rlabel metal5 s 698512 276840 711002 289380 6 mprj_io[4]
port 173 nsew signal bidirectional
rlabel metal2 s 675407 281403 675887 281459 6 mprj_io_analog_en[4]
port 174 nsew signal input
rlabel metal2 s 675407 282691 675887 282747 6 mprj_io_analog_pol[4]
port 175 nsew signal input
rlabel metal2 s 675407 285727 675887 285783 6 mprj_io_analog_sel[4]
port 176 nsew signal input
rlabel metal2 s 675407 282047 675887 282103 6 mprj_io_dm[12]
port 177 nsew signal input
rlabel metal2 s 675407 280207 675887 280263 6 mprj_io_dm[13]
port 178 nsew signal input
rlabel metal2 s 675407 286371 675887 286427 6 mprj_io_dm[14]
port 179 nsew signal input
rlabel metal2 s 675407 287015 675887 287071 6 mprj_io_holdover[4]
port 180 nsew signal input
rlabel metal2 s 675407 290051 675887 290107 6 mprj_io_ib_mode_sel[4]
port 181 nsew signal input
rlabel metal2 s 675407 283243 675887 283299 6 mprj_io_inp_dis[4]
port 182 nsew signal input
rlabel metal2 s 675407 290695 675887 290751 6 mprj_io_oeb[4]
port 183 nsew signal input
rlabel metal2 s 675407 287567 675887 287623 6 mprj_io_out[4]
port 184 nsew signal input
rlabel metal2 s 675407 278367 675887 278423 6 mprj_io_slow_sel[4]
port 185 nsew signal input
rlabel metal2 s 675407 289407 675887 289463 6 mprj_io_vtrip_sel[4]
port 186 nsew signal input
rlabel metal2 s 675407 276527 675887 276583 6 mprj_io_in[4]
port 187 nsew signal output
rlabel metal2 s 675407 291247 675887 291303 6 mprj_io_in_3v3[4]
port 188 nsew signal output
rlabel metal5 s 698512 321040 711002 333580 6 mprj_io[5]
port 189 nsew signal bidirectional
rlabel metal2 s 675407 325603 675887 325659 6 mprj_io_analog_en[5]
port 190 nsew signal input
rlabel metal2 s 675407 326891 675887 326947 6 mprj_io_analog_pol[5]
port 191 nsew signal input
rlabel metal2 s 675407 329927 675887 329983 6 mprj_io_analog_sel[5]
port 192 nsew signal input
rlabel metal2 s 675407 326247 675887 326303 6 mprj_io_dm[15]
port 193 nsew signal input
rlabel metal2 s 675407 324407 675887 324463 6 mprj_io_dm[16]
port 194 nsew signal input
rlabel metal2 s 675407 330571 675887 330627 6 mprj_io_dm[17]
port 195 nsew signal input
rlabel metal2 s 675407 331215 675887 331271 6 mprj_io_holdover[5]
port 196 nsew signal input
rlabel metal2 s 675407 334251 675887 334307 6 mprj_io_ib_mode_sel[5]
port 197 nsew signal input
rlabel metal2 s 675407 327443 675887 327499 6 mprj_io_inp_dis[5]
port 198 nsew signal input
rlabel metal2 s 675407 334895 675887 334951 6 mprj_io_oeb[5]
port 199 nsew signal input
rlabel metal2 s 675407 331767 675887 331823 6 mprj_io_out[5]
port 200 nsew signal input
rlabel metal2 s 675407 322567 675887 322623 6 mprj_io_slow_sel[5]
port 201 nsew signal input
rlabel metal2 s 675407 333607 675887 333663 6 mprj_io_vtrip_sel[5]
port 202 nsew signal input
rlabel metal2 s 675407 320727 675887 320783 6 mprj_io_in[5]
port 203 nsew signal output
rlabel metal2 s 675407 335447 675887 335503 6 mprj_io_in_3v3[5]
port 204 nsew signal output
rlabel metal5 s 698512 365240 711002 377780 6 mprj_io[6]
port 205 nsew signal bidirectional
rlabel metal2 s 675407 369803 675887 369859 6 mprj_io_analog_en[6]
port 206 nsew signal input
rlabel metal2 s 675407 371091 675887 371147 6 mprj_io_analog_pol[6]
port 207 nsew signal input
rlabel metal2 s 675407 374127 675887 374183 6 mprj_io_analog_sel[6]
port 208 nsew signal input
rlabel metal2 s 675407 370447 675887 370503 6 mprj_io_dm[18]
port 209 nsew signal input
rlabel metal2 s 675407 368607 675887 368663 6 mprj_io_dm[19]
port 210 nsew signal input
rlabel metal2 s 675407 374771 675887 374827 6 mprj_io_dm[20]
port 211 nsew signal input
rlabel metal2 s 675407 375415 675887 375471 6 mprj_io_holdover[6]
port 212 nsew signal input
rlabel metal2 s 675407 378451 675887 378507 6 mprj_io_ib_mode_sel[6]
port 213 nsew signal input
rlabel metal2 s 675407 371643 675887 371699 6 mprj_io_inp_dis[6]
port 214 nsew signal input
rlabel metal2 s 675407 379095 675887 379151 6 mprj_io_oeb[6]
port 215 nsew signal input
rlabel metal2 s 675407 375967 675887 376023 6 mprj_io_out[6]
port 216 nsew signal input
rlabel metal2 s 675407 366767 675887 366823 6 mprj_io_slow_sel[6]
port 217 nsew signal input
rlabel metal2 s 675407 377807 675887 377863 6 mprj_io_vtrip_sel[6]
port 218 nsew signal input
rlabel metal2 s 675407 364927 675887 364983 6 mprj_io_in[6]
port 219 nsew signal output
rlabel metal2 s 675407 379647 675887 379703 6 mprj_io_in_3v3[6]
port 220 nsew signal output
rlabel metal2 s 675407 541611 675887 541667 6 mprj_gpio_analog[0]
port 221 nsew signal bidirectional
rlabel metal2 s 675407 543451 675887 543507 6 mprj_gpio_noesd[0]
port 222 nsew signal bidirectional
rlabel metal5 s 698512 539440 711002 551980 6 mprj_io[7]
port 223 nsew signal bidirectional
rlabel metal2 s 675407 544003 675887 544059 6 mprj_io_analog_en[7]
port 224 nsew signal input
rlabel metal2 s 675407 545291 675887 545347 6 mprj_io_analog_pol[7]
port 225 nsew signal input
rlabel metal2 s 675407 548327 675887 548383 6 mprj_io_analog_sel[7]
port 226 nsew signal input
rlabel metal2 s 675407 544647 675887 544703 6 mprj_io_dm[21]
port 227 nsew signal input
rlabel metal2 s 675407 542807 675887 542863 6 mprj_io_dm[22]
port 228 nsew signal input
rlabel metal2 s 675407 548971 675887 549027 6 mprj_io_dm[23]
port 229 nsew signal input
rlabel metal2 s 675407 549615 675887 549671 6 mprj_io_holdover[7]
port 230 nsew signal input
rlabel metal2 s 675407 552651 675887 552707 6 mprj_io_ib_mode_sel[7]
port 231 nsew signal input
rlabel metal2 s 675407 545843 675887 545899 6 mprj_io_inp_dis[7]
port 232 nsew signal input
rlabel metal2 s 675407 553295 675887 553351 6 mprj_io_oeb[7]
port 233 nsew signal input
rlabel metal2 s 675407 550167 675887 550223 6 mprj_io_out[7]
port 234 nsew signal input
rlabel metal2 s 675407 540967 675887 541023 6 mprj_io_slow_sel[7]
port 235 nsew signal input
rlabel metal2 s 675407 552007 675887 552063 6 mprj_io_vtrip_sel[7]
port 236 nsew signal input
rlabel metal2 s 675407 539127 675887 539183 6 mprj_io_in[7]
port 237 nsew signal output
rlabel metal2 s 675407 553847 675887 553903 6 mprj_io_in_3v3[7]
port 238 nsew signal output
rlabel metal2 s 675407 585811 675887 585867 6 mprj_gpio_analog[1]
port 239 nsew signal bidirectional
rlabel metal2 s 675407 587651 675887 587707 6 mprj_gpio_noesd[1]
port 240 nsew signal bidirectional
rlabel metal5 s 698512 583640 711002 596180 6 mprj_io[8]
port 241 nsew signal bidirectional
rlabel metal2 s 675407 588203 675887 588259 6 mprj_io_analog_en[8]
port 242 nsew signal input
rlabel metal2 s 675407 589491 675887 589547 6 mprj_io_analog_pol[8]
port 243 nsew signal input
rlabel metal2 s 675407 592527 675887 592583 6 mprj_io_analog_sel[8]
port 244 nsew signal input
rlabel metal2 s 675407 588847 675887 588903 6 mprj_io_dm[24]
port 245 nsew signal input
rlabel metal2 s 675407 587007 675887 587063 6 mprj_io_dm[25]
port 246 nsew signal input
rlabel metal2 s 675407 593171 675887 593227 6 mprj_io_dm[26]
port 247 nsew signal input
rlabel metal2 s 675407 593815 675887 593871 6 mprj_io_holdover[8]
port 248 nsew signal input
rlabel metal2 s 675407 596851 675887 596907 6 mprj_io_ib_mode_sel[8]
port 249 nsew signal input
rlabel metal2 s 675407 590043 675887 590099 6 mprj_io_inp_dis[8]
port 250 nsew signal input
rlabel metal2 s 675407 597495 675887 597551 6 mprj_io_oeb[8]
port 251 nsew signal input
rlabel metal2 s 675407 594367 675887 594423 6 mprj_io_out[8]
port 252 nsew signal input
rlabel metal2 s 675407 585167 675887 585223 6 mprj_io_slow_sel[8]
port 253 nsew signal input
rlabel metal2 s 675407 596207 675887 596263 6 mprj_io_vtrip_sel[8]
port 254 nsew signal input
rlabel metal2 s 675407 583327 675887 583383 6 mprj_io_in[8]
port 255 nsew signal output
rlabel metal2 s 675407 598047 675887 598103 6 mprj_io_in_3v3[8]
port 256 nsew signal output
rlabel metal2 s 675407 630211 675887 630267 6 mprj_gpio_analog[2]
port 257 nsew signal bidirectional
rlabel metal2 s 675407 632051 675887 632107 6 mprj_gpio_noesd[2]
port 258 nsew signal bidirectional
rlabel metal5 s 698512 628040 711002 640580 6 mprj_io[9]
port 259 nsew signal bidirectional
rlabel metal2 s 675407 632603 675887 632659 6 mprj_io_analog_en[9]
port 260 nsew signal input
rlabel metal2 s 675407 633891 675887 633947 6 mprj_io_analog_pol[9]
port 261 nsew signal input
rlabel metal2 s 675407 636927 675887 636983 6 mprj_io_analog_sel[9]
port 262 nsew signal input
rlabel metal2 s 675407 633247 675887 633303 6 mprj_io_dm[27]
port 263 nsew signal input
rlabel metal2 s 675407 631407 675887 631463 6 mprj_io_dm[28]
port 264 nsew signal input
rlabel metal2 s 675407 637571 675887 637627 6 mprj_io_dm[29]
port 265 nsew signal input
rlabel metal2 s 675407 638215 675887 638271 6 mprj_io_holdover[9]
port 266 nsew signal input
rlabel metal2 s 675407 641251 675887 641307 6 mprj_io_ib_mode_sel[9]
port 267 nsew signal input
rlabel metal2 s 675407 634443 675887 634499 6 mprj_io_inp_dis[9]
port 268 nsew signal input
rlabel metal2 s 675407 641895 675887 641951 6 mprj_io_oeb[9]
port 269 nsew signal input
rlabel metal2 s 675407 638767 675887 638823 6 mprj_io_out[9]
port 270 nsew signal input
rlabel metal2 s 675407 629567 675887 629623 6 mprj_io_slow_sel[9]
port 271 nsew signal input
rlabel metal2 s 675407 640607 675887 640663 6 mprj_io_vtrip_sel[9]
port 272 nsew signal input
rlabel metal2 s 675407 627727 675887 627783 6 mprj_io_in[9]
port 273 nsew signal output
rlabel metal2 s 675407 642447 675887 642503 6 mprj_io_in_3v3[9]
port 274 nsew signal output
rlabel metal2 s 41713 797733 42193 797789 6 mprj_gpio_analog[7]
port 275 nsew signal bidirectional
rlabel metal2 s 41713 795893 42193 795949 6 mprj_gpio_noesd[7]
port 276 nsew signal bidirectional
rlabel metal5 s 6598 787420 19088 799960 6 mprj_io[25]
port 277 nsew signal bidirectional
rlabel metal2 s 41713 795341 42193 795397 6 mprj_io_analog_en[14]
port 278 nsew signal input
rlabel metal2 s 41713 794053 42193 794109 6 mprj_io_analog_pol[14]
port 279 nsew signal input
rlabel metal2 s 41713 791017 42193 791073 6 mprj_io_analog_sel[14]
port 280 nsew signal input
rlabel metal2 s 41713 794697 42193 794753 6 mprj_io_dm[42]
port 281 nsew signal input
rlabel metal2 s 41713 796537 42193 796593 6 mprj_io_dm[43]
port 282 nsew signal input
rlabel metal2 s 41713 790373 42193 790429 6 mprj_io_dm[44]
port 283 nsew signal input
rlabel metal2 s 41713 789729 42193 789785 6 mprj_io_holdover[14]
port 284 nsew signal input
rlabel metal2 s 41713 786693 42193 786749 6 mprj_io_ib_mode_sel[14]
port 285 nsew signal input
rlabel metal2 s 41713 793501 42193 793557 6 mprj_io_inp_dis[14]
port 286 nsew signal input
rlabel metal2 s 41713 786049 42193 786105 6 mprj_io_oeb[14]
port 287 nsew signal input
rlabel metal2 s 41713 789177 42193 789233 6 mprj_io_out[14]
port 288 nsew signal input
rlabel metal2 s 41713 798377 42193 798433 6 mprj_io_slow_sel[14]
port 289 nsew signal input
rlabel metal2 s 41713 787337 42193 787393 6 mprj_io_vtrip_sel[14]
port 290 nsew signal input
rlabel metal2 s 41713 800217 42193 800273 6 mprj_io_in[14]
port 291 nsew signal output
rlabel metal2 s 41713 785497 42193 785553 6 mprj_io_in_3v3[14]
port 292 nsew signal output
rlabel metal2 s 41713 280733 42193 280789 6 mprj_gpio_analog[17]
port 293 nsew signal bidirectional
rlabel metal2 s 41713 278893 42193 278949 6 mprj_gpio_noesd[17]
port 294 nsew signal bidirectional
rlabel metal5 s 6598 270420 19088 282960 6 mprj_io[35]
port 295 nsew signal bidirectional
rlabel metal2 s 41713 278341 42193 278397 6 mprj_io_analog_en[24]
port 296 nsew signal input
rlabel metal2 s 41713 277053 42193 277109 6 mprj_io_analog_pol[24]
port 297 nsew signal input
rlabel metal2 s 41713 274017 42193 274073 6 mprj_io_analog_sel[24]
port 298 nsew signal input
rlabel metal2 s 41713 277697 42193 277753 6 mprj_io_dm[72]
port 299 nsew signal input
rlabel metal2 s 41713 279537 42193 279593 6 mprj_io_dm[73]
port 300 nsew signal input
rlabel metal2 s 41713 273373 42193 273429 6 mprj_io_dm[74]
port 301 nsew signal input
rlabel metal2 s 41713 272729 42193 272785 6 mprj_io_holdover[24]
port 302 nsew signal input
rlabel metal2 s 41713 269693 42193 269749 6 mprj_io_ib_mode_sel[24]
port 303 nsew signal input
rlabel metal2 s 41713 276501 42193 276557 6 mprj_io_inp_dis[24]
port 304 nsew signal input
rlabel metal2 s 41713 269049 42193 269105 6 mprj_io_oeb[24]
port 305 nsew signal input
rlabel metal2 s 41713 272177 42193 272233 6 mprj_io_out[24]
port 306 nsew signal input
rlabel metal2 s 41713 281377 42193 281433 6 mprj_io_slow_sel[24]
port 307 nsew signal input
rlabel metal2 s 41713 270337 42193 270393 6 mprj_io_vtrip_sel[24]
port 308 nsew signal input
rlabel metal2 s 41713 283217 42193 283273 6 mprj_io_in[24]
port 309 nsew signal output
rlabel metal2 s 41713 268497 42193 268553 6 mprj_io_in_3v3[24]
port 310 nsew signal output
rlabel metal5 s 6598 227220 19088 239760 6 mprj_io[36]
port 311 nsew signal bidirectional
rlabel metal2 s 41713 235141 42193 235197 6 mprj_io_analog_en[25]
port 312 nsew signal input
rlabel metal2 s 41713 233853 42193 233909 6 mprj_io_analog_pol[25]
port 313 nsew signal input
rlabel metal2 s 41713 230817 42193 230873 6 mprj_io_analog_sel[25]
port 314 nsew signal input
rlabel metal2 s 41713 234497 42193 234553 6 mprj_io_dm[75]
port 315 nsew signal input
rlabel metal2 s 41713 236337 42193 236393 6 mprj_io_dm[76]
port 316 nsew signal input
rlabel metal2 s 41713 230173 42193 230229 6 mprj_io_dm[77]
port 317 nsew signal input
rlabel metal2 s 41713 229529 42193 229585 6 mprj_io_holdover[25]
port 318 nsew signal input
rlabel metal2 s 41713 226493 42193 226549 6 mprj_io_ib_mode_sel[25]
port 319 nsew signal input
rlabel metal2 s 41713 233301 42193 233357 6 mprj_io_inp_dis[25]
port 320 nsew signal input
rlabel metal2 s 41713 225849 42193 225905 6 mprj_io_oeb[25]
port 321 nsew signal input
rlabel metal2 s 41713 228977 42193 229033 6 mprj_io_out[25]
port 322 nsew signal input
rlabel metal2 s 41713 238177 42193 238233 6 mprj_io_slow_sel[25]
port 323 nsew signal input
rlabel metal2 s 41713 227137 42193 227193 6 mprj_io_vtrip_sel[25]
port 324 nsew signal input
rlabel metal2 s 41713 240017 42193 240073 6 mprj_io_in[25]
port 325 nsew signal output
rlabel metal2 s 41713 225297 42193 225353 6 mprj_io_in_3v3[25]
port 326 nsew signal output
rlabel metal5 s 6598 184020 19088 196560 6 mprj_io[37]
port 327 nsew signal bidirectional
rlabel metal2 s 41713 191941 42193 191997 6 mprj_io_analog_en[26]
port 328 nsew signal input
rlabel metal2 s 41713 190653 42193 190709 6 mprj_io_analog_pol[26]
port 329 nsew signal input
rlabel metal2 s 41713 187617 42193 187673 6 mprj_io_analog_sel[26]
port 330 nsew signal input
rlabel metal2 s 41713 191297 42193 191353 6 mprj_io_dm[78]
port 331 nsew signal input
rlabel metal2 s 41713 193137 42193 193193 6 mprj_io_dm[79]
port 332 nsew signal input
rlabel metal2 s 41713 186973 42193 187029 6 mprj_io_dm[80]
port 333 nsew signal input
rlabel metal2 s 41713 186329 42193 186385 6 mprj_io_holdover[26]
port 334 nsew signal input
rlabel metal2 s 41713 183293 42193 183349 6 mprj_io_ib_mode_sel[26]
port 335 nsew signal input
rlabel metal2 s 41713 190101 42193 190157 6 mprj_io_inp_dis[26]
port 336 nsew signal input
rlabel metal2 s 41713 182649 42193 182705 6 mprj_io_oeb[26]
port 337 nsew signal input
rlabel metal2 s 41713 185777 42193 185833 6 mprj_io_out[26]
port 338 nsew signal input
rlabel metal2 s 41713 194977 42193 195033 6 mprj_io_slow_sel[26]
port 339 nsew signal input
rlabel metal2 s 41713 183937 42193 183993 6 mprj_io_vtrip_sel[26]
port 340 nsew signal input
rlabel metal2 s 41713 196817 42193 196873 6 mprj_io_in[26]
port 341 nsew signal output
rlabel metal2 s 41713 182097 42193 182153 6 mprj_io_in_3v3[26]
port 342 nsew signal output
rlabel metal2 s 41713 754533 42193 754589 6 mprj_gpio_analog[8]
port 343 nsew signal bidirectional
rlabel metal2 s 41713 752693 42193 752749 6 mprj_gpio_noesd[8]
port 344 nsew signal bidirectional
rlabel metal5 s 6598 744220 19088 756760 6 mprj_io[26]
port 345 nsew signal bidirectional
rlabel metal2 s 41713 752141 42193 752197 6 mprj_io_analog_en[15]
port 346 nsew signal input
rlabel metal2 s 41713 750853 42193 750909 6 mprj_io_analog_pol[15]
port 347 nsew signal input
rlabel metal2 s 41713 747817 42193 747873 6 mprj_io_analog_sel[15]
port 348 nsew signal input
rlabel metal2 s 41713 751497 42193 751553 6 mprj_io_dm[45]
port 349 nsew signal input
rlabel metal2 s 41713 753337 42193 753393 6 mprj_io_dm[46]
port 350 nsew signal input
rlabel metal2 s 41713 747173 42193 747229 6 mprj_io_dm[47]
port 351 nsew signal input
rlabel metal2 s 41713 746529 42193 746585 6 mprj_io_holdover[15]
port 352 nsew signal input
rlabel metal2 s 41713 743493 42193 743549 6 mprj_io_ib_mode_sel[15]
port 353 nsew signal input
rlabel metal2 s 41713 750301 42193 750357 6 mprj_io_inp_dis[15]
port 354 nsew signal input
rlabel metal2 s 41713 742849 42193 742905 6 mprj_io_oeb[15]
port 355 nsew signal input
rlabel metal2 s 41713 745977 42193 746033 6 mprj_io_out[15]
port 356 nsew signal input
rlabel metal2 s 41713 755177 42193 755233 6 mprj_io_slow_sel[15]
port 357 nsew signal input
rlabel metal2 s 41713 744137 42193 744193 6 mprj_io_vtrip_sel[15]
port 358 nsew signal input
rlabel metal2 s 41713 757017 42193 757073 6 mprj_io_in[15]
port 359 nsew signal output
rlabel metal2 s 41713 742297 42193 742353 6 mprj_io_in_3v3[15]
port 360 nsew signal output
rlabel metal2 s 41713 711333 42193 711389 6 mprj_gpio_analog[9]
port 361 nsew signal bidirectional
rlabel metal2 s 41713 709493 42193 709549 6 mprj_gpio_noesd[9]
port 362 nsew signal bidirectional
rlabel metal5 s 6598 701020 19088 713560 6 mprj_io[27]
port 363 nsew signal bidirectional
rlabel metal2 s 41713 708941 42193 708997 6 mprj_io_analog_en[16]
port 364 nsew signal input
rlabel metal2 s 41713 707653 42193 707709 6 mprj_io_analog_pol[16]
port 365 nsew signal input
rlabel metal2 s 41713 704617 42193 704673 6 mprj_io_analog_sel[16]
port 366 nsew signal input
rlabel metal2 s 41713 708297 42193 708353 6 mprj_io_dm[48]
port 367 nsew signal input
rlabel metal2 s 41713 710137 42193 710193 6 mprj_io_dm[49]
port 368 nsew signal input
rlabel metal2 s 41713 703973 42193 704029 6 mprj_io_dm[50]
port 369 nsew signal input
rlabel metal2 s 41713 703329 42193 703385 6 mprj_io_holdover[16]
port 370 nsew signal input
rlabel metal2 s 41713 700293 42193 700349 6 mprj_io_ib_mode_sel[16]
port 371 nsew signal input
rlabel metal2 s 41713 707101 42193 707157 6 mprj_io_inp_dis[16]
port 372 nsew signal input
rlabel metal2 s 41713 699649 42193 699705 6 mprj_io_oeb[16]
port 373 nsew signal input
rlabel metal2 s 41713 702777 42193 702833 6 mprj_io_out[16]
port 374 nsew signal input
rlabel metal2 s 41713 711977 42193 712033 6 mprj_io_slow_sel[16]
port 375 nsew signal input
rlabel metal2 s 41713 700937 42193 700993 6 mprj_io_vtrip_sel[16]
port 376 nsew signal input
rlabel metal2 s 41713 713817 42193 713873 6 mprj_io_in[16]
port 377 nsew signal output
rlabel metal2 s 41713 699097 42193 699153 6 mprj_io_in_3v3[16]
port 378 nsew signal output
rlabel metal2 s 41713 667933 42193 667989 6 mprj_gpio_analog[10]
port 379 nsew signal bidirectional
rlabel metal2 s 41713 666093 42193 666149 6 mprj_gpio_noesd[10]
port 380 nsew signal bidirectional
rlabel metal5 s 6598 657620 19088 670160 6 mprj_io[28]
port 381 nsew signal bidirectional
rlabel metal2 s 41713 665541 42193 665597 6 mprj_io_analog_en[17]
port 382 nsew signal input
rlabel metal2 s 41713 664253 42193 664309 6 mprj_io_analog_pol[17]
port 383 nsew signal input
rlabel metal2 s 41713 661217 42193 661273 6 mprj_io_analog_sel[17]
port 384 nsew signal input
rlabel metal2 s 41713 664897 42193 664953 6 mprj_io_dm[51]
port 385 nsew signal input
rlabel metal2 s 41713 666737 42193 666793 6 mprj_io_dm[52]
port 386 nsew signal input
rlabel metal2 s 41713 660573 42193 660629 6 mprj_io_dm[53]
port 387 nsew signal input
rlabel metal2 s 41713 659929 42193 659985 6 mprj_io_holdover[17]
port 388 nsew signal input
rlabel metal2 s 41713 656893 42193 656949 6 mprj_io_ib_mode_sel[17]
port 389 nsew signal input
rlabel metal2 s 41713 663701 42193 663757 6 mprj_io_inp_dis[17]
port 390 nsew signal input
rlabel metal2 s 41713 656249 42193 656305 6 mprj_io_oeb[17]
port 391 nsew signal input
rlabel metal2 s 41713 659377 42193 659433 6 mprj_io_out[17]
port 392 nsew signal input
rlabel metal2 s 41713 668577 42193 668633 6 mprj_io_slow_sel[17]
port 393 nsew signal input
rlabel metal2 s 41713 657537 42193 657593 6 mprj_io_vtrip_sel[17]
port 394 nsew signal input
rlabel metal2 s 41713 670417 42193 670473 6 mprj_io_in[17]
port 395 nsew signal output
rlabel metal2 s 41713 655697 42193 655753 6 mprj_io_in_3v3[17]
port 396 nsew signal output
rlabel metal2 s 41713 624733 42193 624789 6 mprj_gpio_analog[11]
port 397 nsew signal bidirectional
rlabel metal2 s 41713 622893 42193 622949 6 mprj_gpio_noesd[11]
port 398 nsew signal bidirectional
rlabel metal5 s 6598 614420 19088 626960 6 mprj_io[29]
port 399 nsew signal bidirectional
rlabel metal2 s 41713 622341 42193 622397 6 mprj_io_analog_en[18]
port 400 nsew signal input
rlabel metal2 s 41713 621053 42193 621109 6 mprj_io_analog_pol[18]
port 401 nsew signal input
rlabel metal2 s 41713 618017 42193 618073 6 mprj_io_analog_sel[18]
port 402 nsew signal input
rlabel metal2 s 41713 621697 42193 621753 6 mprj_io_dm[54]
port 403 nsew signal input
rlabel metal2 s 41713 623537 42193 623593 6 mprj_io_dm[55]
port 404 nsew signal input
rlabel metal2 s 41713 617373 42193 617429 6 mprj_io_dm[56]
port 405 nsew signal input
rlabel metal2 s 41713 616729 42193 616785 6 mprj_io_holdover[18]
port 406 nsew signal input
rlabel metal2 s 41713 613693 42193 613749 6 mprj_io_ib_mode_sel[18]
port 407 nsew signal input
rlabel metal2 s 41713 620501 42193 620557 6 mprj_io_inp_dis[18]
port 408 nsew signal input
rlabel metal2 s 41713 613049 42193 613105 6 mprj_io_oeb[18]
port 409 nsew signal input
rlabel metal2 s 41713 616177 42193 616233 6 mprj_io_out[18]
port 410 nsew signal input
rlabel metal2 s 41713 625377 42193 625433 6 mprj_io_slow_sel[18]
port 411 nsew signal input
rlabel metal2 s 41713 614337 42193 614393 6 mprj_io_vtrip_sel[18]
port 412 nsew signal input
rlabel metal2 s 41713 627217 42193 627273 6 mprj_io_in[18]
port 413 nsew signal output
rlabel metal2 s 41713 612497 42193 612553 6 mprj_io_in_3v3[18]
port 414 nsew signal output
rlabel metal2 s 41713 581533 42193 581589 6 mprj_gpio_analog[12]
port 415 nsew signal bidirectional
rlabel metal2 s 41713 579693 42193 579749 6 mprj_gpio_noesd[12]
port 416 nsew signal bidirectional
rlabel metal5 s 6598 571220 19088 583760 6 mprj_io[30]
port 417 nsew signal bidirectional
rlabel metal2 s 41713 579141 42193 579197 6 mprj_io_analog_en[19]
port 418 nsew signal input
rlabel metal2 s 41713 577853 42193 577909 6 mprj_io_analog_pol[19]
port 419 nsew signal input
rlabel metal2 s 41713 574817 42193 574873 6 mprj_io_analog_sel[19]
port 420 nsew signal input
rlabel metal2 s 41713 578497 42193 578553 6 mprj_io_dm[57]
port 421 nsew signal input
rlabel metal2 s 41713 580337 42193 580393 6 mprj_io_dm[58]
port 422 nsew signal input
rlabel metal2 s 41713 574173 42193 574229 6 mprj_io_dm[59]
port 423 nsew signal input
rlabel metal2 s 41713 573529 42193 573585 6 mprj_io_holdover[19]
port 424 nsew signal input
rlabel metal2 s 41713 570493 42193 570549 6 mprj_io_ib_mode_sel[19]
port 425 nsew signal input
rlabel metal2 s 41713 577301 42193 577357 6 mprj_io_inp_dis[19]
port 426 nsew signal input
rlabel metal2 s 41713 569849 42193 569905 6 mprj_io_oeb[19]
port 427 nsew signal input
rlabel metal2 s 41713 572977 42193 573033 6 mprj_io_out[19]
port 428 nsew signal input
rlabel metal2 s 41713 582177 42193 582233 6 mprj_io_slow_sel[19]
port 429 nsew signal input
rlabel metal2 s 41713 571137 42193 571193 6 mprj_io_vtrip_sel[19]
port 430 nsew signal input
rlabel metal2 s 41713 584017 42193 584073 6 mprj_io_in[19]
port 431 nsew signal output
rlabel metal2 s 41713 569297 42193 569353 6 mprj_io_in_3v3[19]
port 432 nsew signal output
rlabel metal2 s 41713 538333 42193 538389 6 mprj_gpio_analog[13]
port 433 nsew signal bidirectional
rlabel metal2 s 41713 536493 42193 536549 6 mprj_gpio_noesd[13]
port 434 nsew signal bidirectional
rlabel metal5 s 6598 528020 19088 540560 6 mprj_io[31]
port 435 nsew signal bidirectional
rlabel metal2 s 41713 535941 42193 535997 6 mprj_io_analog_en[20]
port 436 nsew signal input
rlabel metal2 s 41713 534653 42193 534709 6 mprj_io_analog_pol[20]
port 437 nsew signal input
rlabel metal2 s 41713 531617 42193 531673 6 mprj_io_analog_sel[20]
port 438 nsew signal input
rlabel metal2 s 41713 535297 42193 535353 6 mprj_io_dm[60]
port 439 nsew signal input
rlabel metal2 s 41713 537137 42193 537193 6 mprj_io_dm[61]
port 440 nsew signal input
rlabel metal2 s 41713 530973 42193 531029 6 mprj_io_dm[62]
port 441 nsew signal input
rlabel metal2 s 41713 530329 42193 530385 6 mprj_io_holdover[20]
port 442 nsew signal input
rlabel metal2 s 41713 527293 42193 527349 6 mprj_io_ib_mode_sel[20]
port 443 nsew signal input
rlabel metal2 s 41713 534101 42193 534157 6 mprj_io_inp_dis[20]
port 444 nsew signal input
rlabel metal2 s 41713 526649 42193 526705 6 mprj_io_oeb[20]
port 445 nsew signal input
rlabel metal2 s 41713 529777 42193 529833 6 mprj_io_out[20]
port 446 nsew signal input
rlabel metal2 s 41713 538977 42193 539033 6 mprj_io_slow_sel[20]
port 447 nsew signal input
rlabel metal2 s 41713 527937 42193 527993 6 mprj_io_vtrip_sel[20]
port 448 nsew signal input
rlabel metal2 s 41713 540817 42193 540873 6 mprj_io_in[20]
port 449 nsew signal output
rlabel metal2 s 41713 526097 42193 526153 6 mprj_io_in_3v3[20]
port 450 nsew signal output
rlabel metal2 s 41713 410533 42193 410589 6 mprj_gpio_analog[14]
port 451 nsew signal bidirectional
rlabel metal2 s 41713 408693 42193 408749 6 mprj_gpio_noesd[14]
port 452 nsew signal bidirectional
rlabel metal5 s 6598 400220 19088 412760 6 mprj_io[32]
port 453 nsew signal bidirectional
rlabel metal2 s 41713 408141 42193 408197 6 mprj_io_analog_en[21]
port 454 nsew signal input
rlabel metal2 s 41713 406853 42193 406909 6 mprj_io_analog_pol[21]
port 455 nsew signal input
rlabel metal2 s 41713 403817 42193 403873 6 mprj_io_analog_sel[21]
port 456 nsew signal input
rlabel metal2 s 41713 407497 42193 407553 6 mprj_io_dm[63]
port 457 nsew signal input
rlabel metal2 s 41713 409337 42193 409393 6 mprj_io_dm[64]
port 458 nsew signal input
rlabel metal2 s 41713 403173 42193 403229 6 mprj_io_dm[65]
port 459 nsew signal input
rlabel metal2 s 41713 402529 42193 402585 6 mprj_io_holdover[21]
port 460 nsew signal input
rlabel metal2 s 41713 399493 42193 399549 6 mprj_io_ib_mode_sel[21]
port 461 nsew signal input
rlabel metal2 s 41713 406301 42193 406357 6 mprj_io_inp_dis[21]
port 462 nsew signal input
rlabel metal2 s 41713 398849 42193 398905 6 mprj_io_oeb[21]
port 463 nsew signal input
rlabel metal2 s 41713 401977 42193 402033 6 mprj_io_out[21]
port 464 nsew signal input
rlabel metal2 s 41713 411177 42193 411233 6 mprj_io_slow_sel[21]
port 465 nsew signal input
rlabel metal2 s 41713 400137 42193 400193 6 mprj_io_vtrip_sel[21]
port 466 nsew signal input
rlabel metal2 s 41713 413017 42193 413073 6 mprj_io_in[21]
port 467 nsew signal output
rlabel metal2 s 41713 398297 42193 398353 6 mprj_io_in_3v3[21]
port 468 nsew signal output
rlabel metal2 s 41713 367333 42193 367389 6 mprj_gpio_analog[15]
port 469 nsew signal bidirectional
rlabel metal2 s 41713 365493 42193 365549 6 mprj_gpio_noesd[15]
port 470 nsew signal bidirectional
rlabel metal5 s 6598 357020 19088 369560 6 mprj_io[33]
port 471 nsew signal bidirectional
rlabel metal2 s 41713 364941 42193 364997 6 mprj_io_analog_en[22]
port 472 nsew signal input
rlabel metal2 s 41713 363653 42193 363709 6 mprj_io_analog_pol[22]
port 473 nsew signal input
rlabel metal2 s 41713 360617 42193 360673 6 mprj_io_analog_sel[22]
port 474 nsew signal input
rlabel metal2 s 41713 364297 42193 364353 6 mprj_io_dm[66]
port 475 nsew signal input
rlabel metal2 s 41713 366137 42193 366193 6 mprj_io_dm[67]
port 476 nsew signal input
rlabel metal2 s 41713 359973 42193 360029 6 mprj_io_dm[68]
port 477 nsew signal input
rlabel metal2 s 41713 359329 42193 359385 6 mprj_io_holdover[22]
port 478 nsew signal input
rlabel metal2 s 41713 356293 42193 356349 6 mprj_io_ib_mode_sel[22]
port 479 nsew signal input
rlabel metal2 s 41713 363101 42193 363157 6 mprj_io_inp_dis[22]
port 480 nsew signal input
rlabel metal2 s 41713 355649 42193 355705 6 mprj_io_oeb[22]
port 481 nsew signal input
rlabel metal2 s 41713 358777 42193 358833 6 mprj_io_out[22]
port 482 nsew signal input
rlabel metal2 s 41713 367977 42193 368033 6 mprj_io_slow_sel[22]
port 483 nsew signal input
rlabel metal2 s 41713 356937 42193 356993 6 mprj_io_vtrip_sel[22]
port 484 nsew signal input
rlabel metal2 s 41713 369817 42193 369873 6 mprj_io_in[22]
port 485 nsew signal output
rlabel metal2 s 41713 355097 42193 355153 6 mprj_io_in_3v3[22]
port 486 nsew signal output
rlabel metal2 s 41713 323933 42193 323989 6 mprj_gpio_analog[16]
port 487 nsew signal bidirectional
rlabel metal2 s 41713 322093 42193 322149 6 mprj_gpio_noesd[16]
port 488 nsew signal bidirectional
rlabel metal5 s 6598 313620 19088 326160 6 mprj_io[34]
port 489 nsew signal bidirectional
rlabel metal2 s 41713 321541 42193 321597 6 mprj_io_analog_en[23]
port 490 nsew signal input
rlabel metal2 s 41713 320253 42193 320309 6 mprj_io_analog_pol[23]
port 491 nsew signal input
rlabel metal2 s 41713 317217 42193 317273 6 mprj_io_analog_sel[23]
port 492 nsew signal input
rlabel metal2 s 41713 320897 42193 320953 6 mprj_io_dm[69]
port 493 nsew signal input
rlabel metal2 s 41713 322737 42193 322793 6 mprj_io_dm[70]
port 494 nsew signal input
rlabel metal2 s 41713 316573 42193 316629 6 mprj_io_dm[71]
port 495 nsew signal input
rlabel metal2 s 41713 315929 42193 315985 6 mprj_io_holdover[23]
port 496 nsew signal input
rlabel metal2 s 41713 312893 42193 312949 6 mprj_io_ib_mode_sel[23]
port 497 nsew signal input
rlabel metal2 s 41713 319701 42193 319757 6 mprj_io_inp_dis[23]
port 498 nsew signal input
rlabel metal2 s 41713 312249 42193 312305 6 mprj_io_oeb[23]
port 499 nsew signal input
rlabel metal2 s 41713 315377 42193 315433 6 mprj_io_out[23]
port 500 nsew signal input
rlabel metal2 s 41713 324577 42193 324633 6 mprj_io_slow_sel[23]
port 501 nsew signal input
rlabel metal2 s 41713 313537 42193 313593 6 mprj_io_vtrip_sel[23]
port 502 nsew signal input
rlabel metal2 s 41713 326417 42193 326473 6 mprj_io_in[23]
port 503 nsew signal output
rlabel metal2 s 41713 311697 42193 311753 6 mprj_io_in_3v3[23]
port 504 nsew signal output
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145103 40000 145131 40174 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145103 40174 145144 40202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527455 41713 527511 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 523131 41713 523187 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472655 41713 472711 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468331 41713 468387 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472636 41806 472711 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468312 41806 468387 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417855 41713 417911 41820 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413531 41713 413587 41820 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527468 42193 527496 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 523144 42193 523172 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527456 44134 527508 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 523132 44134 523184 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527468 44198 527496 46854 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472636 42193 472664 44270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468312 42193 468340 44270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417855 41820 417924 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413531 41820 413600 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 363055 41713 363111 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 358731 41713 358787 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308255 41713 308311 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303931 41713 303987 41806 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308232 41806 308311 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303908 41806 303987 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199655 41713 199711 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 195331 41713 195387 42193 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417896 42193 417924 44270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413572 42193 413600 44270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 363064 42193 363092 44270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 358740 42193 358768 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308232 42193 308260 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303908 42193 303936 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199672 42193 199700 44118 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199672 44118 199884 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 195348 42193 195376 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145116 40202 145144 44134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199660 44134 199884 44146 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199856 44146 199884 44202 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199660 44146 199712 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 195336 44134 195388 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 145104 44134 145156 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 143632 44134 143684 44198 6 porb_h
port 505 nsew signal input
rlabel metal2 s 358728 44202 358780 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 308220 44202 308272 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 303896 44202 303948 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 199844 44202 199896 44266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 472624 44270 472676 44334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 468300 44270 468352 44334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 417884 44270 417936 44334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 413560 44270 413612 44334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 363052 44270 363104 44334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 143644 44198 143672 45562 6 porb_h
port 505 nsew signal input
rlabel metal2 s 143632 45562 143684 45626 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42340 45562 42392 45626 6 porb_h
port 505 nsew signal input
rlabel metal2 s 527456 46854 527508 46918 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 46922 673696 46986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 107275 675340 107306 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673656 46986 673684 107306 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 107331 675887 107358 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 107306 675352 107358 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 107358 675887 107370 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673644 107306 673696 107370 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 107370 675887 107386 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 107386 675887 107387 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 111655 675887 111669 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 107386 675340 111669 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 111669 675887 111697 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 111697 675887 111711 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 111711 675432 111794 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 111794 675444 111858 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 111794 673880 111858 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 151662 675340 151710 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673840 111858 673868 151710 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 151731 675887 151745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 151710 675352 151745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 151745 675887 151773 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 151773 675887 151787 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 151773 675352 151774 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 151710 673880 151774 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 156055 675887 156060 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 156060 675887 156111 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 156111 675432 156182 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 151774 675340 156182 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 156182 675432 156210 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 156210 675432 156266 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 156266 675444 156330 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 156266 673788 156330 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 156330 673776 195774 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 45626 42380 184503 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 184489 42193 184503 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 184503 42380 184531 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 184531 42288 188958 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 184531 42193 184545 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 188813 42193 188869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 188869 41920 188958 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 188958 42380 188986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 195774 675444 195838 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 195774 673788 195838 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 195838 675432 195931 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 195931 675887 195945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 195945 675887 195973 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 195973 675887 195987 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 195973 675340 199702 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 199702 675432 199730 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 199730 675432 200255 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 200255 675887 200311 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 200311 675432 200398 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 200398 675444 200462 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 200398 673788 200462 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 200462 673776 239634 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 188986 42380 226306 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 226306 42380 226334 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 226334 42288 227854 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 227689 42193 227745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 227745 41828 227746 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 227746 41828 227854 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 227854 42288 227882 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 227882 42288 232478 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 232013 42193 232069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 232069 41828 232478 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 232478 42380 232506 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 239634 675444 239698 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 239634 673788 239698 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 239698 675432 240131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 240131 675887 240145 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 240145 675887 240173 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 240173 675887 240187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 240173 675340 243902 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 243902 675432 243930 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 243930 675432 244455 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 244455 675887 244511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 244511 675432 244598 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 244598 675444 244662 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 244598 673788 244662 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 244662 673776 284038 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 232506 42380 264946 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 264946 42380 264974 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 264974 42288 270903 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 270889 42193 270903 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 270903 42288 270931 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 270931 42288 275318 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 270931 42193 270945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 275213 42193 275269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 275269 41828 275318 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 275318 42380 275346 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 275346 42380 283902 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42340 283902 42392 283966 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 284038 675444 284102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 284038 673788 284102 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 284102 675432 284531 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42340 284106 42392 284170 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 284531 675887 284587 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 284587 675432 285110 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 285110 675432 285138 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 288855 675887 288869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 285138 675340 288869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 288869 675887 288897 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 288897 675887 288911 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 288911 675432 289274 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 289274 675444 289338 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 289274 673788 289338 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 289338 673776 328238 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 284170 42380 312870 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42340 312870 42392 312934 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42248 313074 42300 313138 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 313138 42288 313942 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 313942 42288 313970 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 313970 42288 318294 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 313970 41920 314078 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 314078 41920 314089 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 314089 42193 314145 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 318294 42380 318322 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 328238 675444 328302 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 328238 673788 328302 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 328302 675432 328630 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 328630 675432 328658 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 328658 675432 328731 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 328731 675887 328780 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 328780 675887 328787 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 333055 675887 333069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 328658 675340 333066 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 333066 675352 333069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 333069 675887 333097 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 333097 675887 333111 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 333097 675352 333130 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673552 333066 673604 333130 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 333130 675340 333180 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673564 333130 673592 372778 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 318322 42380 357503 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 318322 41920 318413 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 318413 42193 318469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 357489 42193 357503 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 357503 42380 357531 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 357531 42288 361546 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 357531 42193 357545 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 361546 42380 361574 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 372778 675444 372830 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 372830 675444 372842 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673552 372778 673604 372842 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 372842 675432 372858 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 372858 675432 372931 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 372931 675887 372980 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 372980 675887 372987 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 377255 675887 377269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 372858 675340 377269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 377269 675887 377297 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 377297 675887 377311 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673564 372842 673592 380866 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 361574 42380 380866 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 361574 41828 361813 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 361813 42193 361869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673472 380866 673592 380894 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 380866 42380 380894 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673472 380894 673500 546994 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 380894 42288 400710 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 400689 42193 400710 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 400710 42288 400738 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 400738 42288 405470 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 400738 42193 400745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 405013 42193 405069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 405069 41828 405470 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 405470 42380 405498 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 405498 42380 419506 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 419506 42380 419534 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 419534 42288 528414 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 528414 42288 528442 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 528442 42288 532827 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 528442 41920 528489 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 528489 42193 528545 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 532813 42193 532827 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 532827 42380 532855 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 546994 675444 547058 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 546994 675260 547058 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673460 546994 673512 547058 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 547058 675432 547131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 547131 675887 547159 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 547159 675887 547187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 551455 675887 551469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 547058 675248 551469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 551469 675887 551482 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 551482 675887 551497 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 551497 675887 551511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 551497 675260 551546 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 551482 673788 551546 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 551546 675248 551580 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 551546 673776 590786 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 532855 42380 571703 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 532855 42193 532869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 571689 42193 571703 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 571703 42380 571731 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 571731 42288 576506 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 571731 42193 571745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 576013 42193 576069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 576069 41828 576506 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42432 576506 42484 576570 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42248 576506 42300 576570 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41788 576506 41840 576570 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 590786 675444 590850 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 590786 675260 590850 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 590786 673788 590850 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 590850 675432 591331 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 591331 675887 591359 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 591359 675887 591387 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 595655 675887 595683 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 595683 675887 595711 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 595711 675432 596090 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 590850 675248 596090 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 596090 675444 596154 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 596090 675260 596154 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 596090 673788 596154 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 635731 675887 635732 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 635732 675887 635787 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 596154 673776 635734 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42444 576570 42472 604426 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 604426 42472 604454 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 604454 42380 614774 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 614774 42380 614802 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 614802 42288 619126 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 614802 41828 614889 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 614889 42193 614945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 619126 42380 619154 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 635787 675432 635854 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 635734 675352 635798 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 635734 673788 635798 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 635798 675340 635854 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 635854 675432 635882 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 640055 675887 640070 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 635882 675340 640070 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 640070 675887 640086 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 640086 675887 640098 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 640098 675887 640111 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 640098 675352 640150 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 640086 673880 640150 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 640150 675340 640181 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 679931 675887 679932 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 679932 675887 679987 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 679987 675432 680070 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673840 640150 673868 680070 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 619154 42380 651346 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 619154 41920 619213 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 619213 42193 619269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 651346 42380 651374 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 651374 42288 658103 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 658089 42193 658103 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 658103 42288 658131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 658131 42288 662510 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 658131 42193 658145 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 662413 42193 662469 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 662469 41920 662510 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 662510 42380 662538 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 680070 675444 680134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673828 680070 673880 680134 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 680134 675432 680326 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 680326 675432 680354 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 684255 675887 684270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 680354 675340 684270 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 684270 675887 684286 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 684286 675887 684298 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 684298 675887 684311 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675300 684298 675352 684350 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673460 684286 673512 684350 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 684350 675340 684381 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673472 684350 673500 723998 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 662538 42380 689986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 689986 42380 690014 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 690014 42288 701406 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 701406 42288 701434 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 701434 42288 705827 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 701434 41920 701489 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 701489 42193 701545 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 705813 42193 705827 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 705827 42380 705855 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 723998 675444 724062 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673460 723998 673512 724062 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 724062 675432 724131 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 724131 675887 724187 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 724187 675432 724662 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 724662 675432 724690 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 728455 675887 728470 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 724690 675340 728470 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 728470 675887 728498 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 728498 675887 728511 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 728511 675432 728554 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 728554 675444 728618 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 728554 673788 728618 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 768531 675887 768559 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 768559 675887 768587 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 768587 675432 769082 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 728618 673776 769082 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42352 705855 42380 728626 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 705855 42193 705869 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 728626 42380 728654 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 728654 42288 744703 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 744689 42193 744703 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 744703 42288 744731 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 744731 42288 749550 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 744731 42193 744745 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 749006 41828 749013 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 749013 42193 749069 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 749069 41828 749550 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41800 749550 42472 749578 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 769082 675444 769146 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 769082 675260 769146 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 769082 673788 769146 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 772855 675887 772883 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 772883 675887 772911 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 772911 675432 773298 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675220 769146 675248 773298 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 773298 675444 773362 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675208 773298 675260 773362 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 773298 673788 773362 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673748 773362 673776 855374 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42444 749578 42472 787986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 787889 42193 787945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 787955 42288 787986 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42432 787986 42484 788050 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42248 787986 42300 788038 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 787945 41920 788038 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 788038 42300 788050 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41892 788050 42288 788066 6 porb_h
port 505 nsew signal input
rlabel metal2 s 42260 788066 42288 792254 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 792213 42193 792254 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41713 792254 42288 792269 6 porb_h
port 505 nsew signal input
rlabel metal2 s 41722 792269 42288 792282 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675392 855374 675444 855438 6 porb_h
port 505 nsew signal input
rlabel metal2 s 673736 855374 673788 855438 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 855438 675432 855931 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675404 855931 675887 855945 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 855945 675887 855973 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 855973 675887 855987 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 855973 675340 860254 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 860254 675418 860255 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675312 860255 675887 860282 6 porb_h
port 505 nsew signal input
rlabel metal2 s 675407 860282 675887 860311 6 porb_h
port 505 nsew signal input
rlabel via1 s 527456 44140 527508 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 523132 44140 523184 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 199660 44140 199712 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 195336 44140 195388 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 145104 44140 145156 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 143632 44140 143684 44192 6 porb_h
port 505 nsew signal input
rlabel via1 s 472624 44276 472676 44328 6 porb_h
port 505 nsew signal input
rlabel via1 s 468300 44276 468352 44328 6 porb_h
port 505 nsew signal input
rlabel via1 s 417884 44276 417936 44328 6 porb_h
port 505 nsew signal input
rlabel via1 s 413560 44276 413612 44328 6 porb_h
port 505 nsew signal input
rlabel via1 s 363052 44276 363104 44328 6 porb_h
port 505 nsew signal input
rlabel via1 s 358728 44208 358780 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 308220 44208 308272 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 303896 44208 303948 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 199844 44208 199896 44260 6 porb_h
port 505 nsew signal input
rlabel via1 s 143632 45568 143684 45620 6 porb_h
port 505 nsew signal input
rlabel via1 s 42340 45568 42392 45620 6 porb_h
port 505 nsew signal input
rlabel via1 s 527456 46860 527508 46912 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 46928 673696 46980 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 107312 675352 107364 6 porb_h
port 505 nsew signal input
rlabel via1 s 673644 107312 673696 107364 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 111800 675444 111852 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 111800 673880 111852 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 151716 675352 151768 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 151716 673880 151768 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 156272 675444 156324 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 156272 673788 156324 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 195780 675444 195832 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 195780 673788 195832 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 200404 675444 200456 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 200404 673788 200456 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 239640 675444 239692 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 239640 673788 239692 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 244604 675444 244656 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 244604 673788 244656 6 porb_h
port 505 nsew signal input
rlabel via1 s 42340 283908 42392 283960 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 284044 675444 284096 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 284044 673788 284096 6 porb_h
port 505 nsew signal input
rlabel via1 s 42340 284112 42392 284164 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 289280 675444 289332 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 289280 673788 289332 6 porb_h
port 505 nsew signal input
rlabel via1 s 42340 312876 42392 312928 6 porb_h
port 505 nsew signal input
rlabel via1 s 42248 313080 42300 313132 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 328244 675444 328296 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 328244 673788 328296 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 333072 675352 333124 6 porb_h
port 505 nsew signal input
rlabel via1 s 673552 333072 673604 333124 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 372784 675444 372836 6 porb_h
port 505 nsew signal input
rlabel via1 s 673552 372784 673604 372836 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 547000 675444 547052 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 547000 675260 547052 6 porb_h
port 505 nsew signal input
rlabel via1 s 673460 547000 673512 547052 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 551488 675260 551540 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 551488 673788 551540 6 porb_h
port 505 nsew signal input
rlabel via1 s 42432 576512 42484 576564 6 porb_h
port 505 nsew signal input
rlabel via1 s 42248 576512 42300 576564 6 porb_h
port 505 nsew signal input
rlabel via1 s 41788 576512 41840 576564 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 590792 675444 590844 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 590792 675260 590844 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 590792 673788 590844 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 596096 675444 596148 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 596096 675260 596148 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 596096 673788 596148 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 635740 675352 635792 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 635740 673788 635792 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 640092 675352 640144 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 640092 673880 640144 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 680076 675444 680128 6 porb_h
port 505 nsew signal input
rlabel via1 s 673828 680076 673880 680128 6 porb_h
port 505 nsew signal input
rlabel via1 s 675300 684292 675352 684344 6 porb_h
port 505 nsew signal input
rlabel via1 s 673460 684292 673512 684344 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 724004 675444 724056 6 porb_h
port 505 nsew signal input
rlabel via1 s 673460 724004 673512 724056 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 728560 675444 728612 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 728560 673788 728612 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 769088 675444 769140 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 769088 675260 769140 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 769088 673788 769140 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 773304 675444 773356 6 porb_h
port 505 nsew signal input
rlabel via1 s 675208 773304 675260 773356 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 773304 673788 773356 6 porb_h
port 505 nsew signal input
rlabel via1 s 42432 787992 42484 788044 6 porb_h
port 505 nsew signal input
rlabel via1 s 42248 787992 42300 788044 6 porb_h
port 505 nsew signal input
rlabel via1 s 675392 855380 675444 855432 6 porb_h
port 505 nsew signal input
rlabel via1 s 673736 855380 673788 855432 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527450 44140 527514 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523126 44140 523190 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523126 44152 527514 44180 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527450 44180 527514 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523126 44180 523190 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 199654 44140 199718 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 195330 44140 195394 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 145098 44140 145162 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143626 44140 143690 44152 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143626 44152 199718 44180 6 porb_h
port 505 nsew signal input
rlabel metal1 s 199654 44180 199718 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 195330 44180 195394 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 145098 44180 145162 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143626 44180 143690 44192 6 porb_h
port 505 nsew signal input
rlabel metal1 s 523144 44192 523172 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 358722 44208 358786 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 308214 44208 308278 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303890 44208 303954 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 199838 44208 199902 44220 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303890 44220 361574 44248 6 porb_h
port 505 nsew signal input
rlabel metal1 s 472618 44276 472682 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 468294 44276 468358 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 417878 44276 417942 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 413554 44276 413618 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 363046 44276 363110 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 361546 44248 361574 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 358722 44248 358786 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 308214 44248 308278 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303890 44248 303954 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 199838 44220 303614 44248 6 porb_h
port 505 nsew signal input
rlabel metal1 s 361546 44288 523172 44316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303908 44260 303936 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303586 44248 303614 44288 6 porb_h
port 505 nsew signal input
rlabel metal1 s 199838 44248 199902 44260 6 porb_h
port 505 nsew signal input
rlabel metal1 s 303586 44288 303936 44316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 472618 44316 472682 44328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 468294 44316 468358 44328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 417878 44316 417942 44328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 413554 44316 413618 44328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 363046 44316 363110 44328 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143626 45568 143690 45580 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42334 45568 42398 45580 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42334 45580 143690 45608 6 porb_h
port 505 nsew signal input
rlabel metal1 s 143626 45608 143690 45620 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42334 45608 42398 45620 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527450 46860 527514 46912 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 46928 673702 46940 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527468 46912 527496 46940 6 porb_h
port 505 nsew signal input
rlabel metal1 s 527468 46940 673702 46968 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 46968 673702 46980 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 107312 675358 107324 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 107312 673702 107324 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 107324 675358 107352 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 107352 675358 107364 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673638 107352 673702 107364 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 111800 675450 111812 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 111800 673886 111812 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 111812 675450 111840 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 111840 675450 111852 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 111840 673886 111852 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 151716 675358 151728 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 151716 673886 151728 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 151728 675358 151756 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 151756 675358 151768 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 151756 673886 151768 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 156272 675450 156284 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 156272 673794 156284 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 156284 675450 156312 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 156312 675450 156324 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 156312 673794 156324 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 195780 675450 195792 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 195780 673794 195792 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 195792 675450 195820 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 195820 675450 195832 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 195820 673794 195832 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 200404 675450 200416 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 200404 673794 200416 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 200416 675450 200444 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 200444 675450 200456 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 200444 673794 200456 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 239640 675450 239652 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 239640 673794 239652 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 239652 675450 239680 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 239680 675450 239692 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 239680 673794 239692 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 244604 675450 244616 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 244604 673794 244616 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 244616 675450 244644 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 244644 675450 244656 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 244644 673794 244656 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42334 283908 42398 283960 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 284044 675450 284056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 284044 673794 284056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 284056 675450 284084 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 284084 675450 284096 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 284084 673794 284096 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42352 283960 42380 284112 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42334 284112 42398 284164 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 289280 675450 289292 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 289280 673794 289292 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 289292 675450 289320 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 289320 675450 289332 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 289320 673794 289332 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42334 312876 42398 312928 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42352 312928 42380 313092 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 313080 42306 313092 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 313092 42380 313120 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 313120 42306 313132 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 328244 675450 328256 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 328244 673794 328256 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 328256 675450 328284 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 328284 675450 328296 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 328284 673794 328296 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 333072 675358 333084 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673546 333072 673610 333084 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673546 333084 675358 333112 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 333112 675358 333124 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673546 333112 673610 333124 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 372784 675450 372796 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673546 372784 673610 372796 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673546 372796 675450 372824 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 372824 675450 372836 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673546 372824 673610 372836 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 547000 675450 547012 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 547000 675266 547012 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 547000 673518 547012 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 547012 675450 547040 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 547040 675450 547052 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 547040 675266 547052 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 547040 673518 547052 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 551488 675266 551500 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 551488 673794 551500 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 551500 675266 551528 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 551528 675266 551540 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 551528 673794 551540 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 576512 42490 576524 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 576512 42306 576524 6 porb_h
port 505 nsew signal input
rlabel metal1 s 41782 576512 41846 576524 6 porb_h
port 505 nsew signal input
rlabel metal1 s 41782 576524 42490 576552 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 576552 42490 576564 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 576552 42306 576564 6 porb_h
port 505 nsew signal input
rlabel metal1 s 41782 576552 41846 576564 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 590792 675450 590804 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 590792 675266 590804 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 590792 673794 590804 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 590804 675450 590832 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 590832 675450 590844 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 590832 675266 590844 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 590832 673794 590844 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 596096 675450 596108 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 596096 675266 596108 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 596096 673794 596108 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 596108 675450 596136 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 596136 675450 596148 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 596136 675266 596148 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 596136 673794 596148 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 635740 675358 635752 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 635740 673794 635752 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 635752 675358 635780 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 635780 675358 635792 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 635780 673794 635792 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 640092 675358 640104 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 640092 673886 640104 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 640104 675358 640132 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 640132 675358 640144 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 640132 673886 640144 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 680076 675450 680088 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 680076 673886 680088 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 680088 675450 680116 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 680116 675450 680128 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673822 680116 673886 680128 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 684292 675358 684304 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 684292 673518 684304 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 684304 675358 684332 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675294 684332 675358 684344 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 684332 673518 684344 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 724004 675450 724016 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 724004 673518 724016 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 724016 675450 724044 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 724044 675450 724056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673454 724044 673518 724056 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 728560 675450 728572 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 728560 673794 728572 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 728572 675450 728600 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 728600 675450 728612 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 728600 673794 728612 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 769088 675450 769100 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 769088 675266 769100 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 769088 673794 769100 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 769100 675450 769128 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 769128 675450 769140 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 769128 675266 769140 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 769128 673794 769140 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 773304 675450 773316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 773304 675266 773316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 773304 673794 773316 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 773316 675450 773344 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 773344 675450 773356 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675202 773344 675266 773356 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 773344 673794 773356 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 787992 42490 788004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 787992 42306 788004 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 788004 42490 788032 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42426 788032 42490 788044 6 porb_h
port 505 nsew signal input
rlabel metal1 s 42242 788032 42306 788044 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 855380 675450 855392 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 855380 673794 855392 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 855392 675450 855420 6 porb_h
port 505 nsew signal input
rlabel metal1 s 675386 855420 675450 855432 6 porb_h
port 505 nsew signal input
rlabel metal1 s 673730 855420 673794 855432 6 porb_h
port 505 nsew signal input
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 506 nsew signal input
rlabel metal3 s 141820 37046 141966 37818 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 37818 141966 37911 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141873 37911 141966 37971 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 37911 141820 37971 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 37971 141873 38031 6 resetb_core_h
port 507 nsew signal output
rlabel metal3 s 141667 38031 141813 40000 6 resetb_core_h
port 507 nsew signal output
rlabel metal4 s 93607 36323 132793 37013 6 vdda
port 508 nsew signal bidirectional
rlabel metal4 s 93546 28653 192982 28719 6 vssa
port 509 nsew signal bidirectional
rlabel metal4 s 93546 30753 132854 30762 6 vssd
port 510 nsew signal bidirectional
rlabel metal4 s 93546 30762 132869 31674 6 vssd
port 510 nsew signal bidirectional
rlabel metal4 s 93546 31674 132854 31683 6 vssd
port 510 nsew signal bidirectional
rlabel metal3 s 631944 997600 636944 1014070 6 mprj_analog[1]
port 511 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030789 6 mprj_io[15]
port 512 nsew signal bidirectional
rlabel metal3 s 530744 997600 535744 1014070 6 mprj_analog[2]
port 513 nsew signal bidirectional
rlabel metal5 s 527210 1018624 539378 1030789 6 mprj_io[16]
port 514 nsew signal bidirectional
rlabel metal3 s 479144 997600 484144 1014070 6 mprj_analog[3]
port 515 nsew signal bidirectional
rlabel metal5 s 475610 1018624 487778 1030789 6 mprj_io[17]
port 516 nsew signal bidirectional
rlabel metal3 s 429744 997600 434744 1014070 6 mprj_analog[4]
port 517 nsew signal bidirectional
rlabel metal5 s 426210 1018624 438378 1030789 6 mprj_io[18]
port 518 nsew signal bidirectional
rlabel metal3 s 677600 934600 680737 948922 6 mprj_analog[0]
port 519 nsew signal bidirectional
rlabel metal2 s 677600 944142 682732 948922 6 mprj_clamp_high[0]
port 520 nsew signal input
rlabel metal2 s 677600 954121 678011 958901 6 mprj_clamp_low[0]
port 521 nsew signal input
rlabel metal5 s 698624 945422 710789 957590 6 mprj_io[14]
port 522 nsew signal bidirectional
rlabel metal5 s 697980 893466 711433 904346 6 vccd1_pad
port 523 nsew signal bidirectional
rlabel metal5 s 698624 805222 710789 817390 6 vdda1_pad
port 524 nsew signal bidirectional
rlabel metal5 s 698624 496422 710789 508590 6 vdda1_pad2
port 525 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1_pad
port 526 nsew signal bidirectional
rlabel metal5 s 698624 409822 710789 421990 6 vssa1_pad2
port 527 nsew signal bidirectional
rlabel metal4 s 679377 423146 680307 451854 6 vccd1
port 528 nsew signal bidirectional
rlabel metal4 s 680587 423207 681277 451793 6 vdda1
port 529 nsew signal bidirectional
rlabel metal4 s 688881 423146 688947 544782 6 vssa1
port 530 nsew signal bidirectional
rlabel metal3 s 678000 461700 685920 466500 6 vssd1
port 531 nsew signal bidirectional
rlabel metal5 s 697980 453666 711433 464546 6 vssd1_pad
port 532 nsew signal bidirectional
rlabel metal3 s 175944 997600 180944 1014070 6 mprj_analog[7]
port 533 nsew signal bidirectional
rlabel metal5 s 172410 1018624 184578 1030789 6 mprj_io[21]
port 534 nsew signal bidirectional
rlabel metal3 s 127944 997600 132944 1014070 6 mprj_analog[8]
port 535 nsew signal bidirectional
rlabel metal5 s 124410 1018624 136578 1030789 6 mprj_io[22]
port 536 nsew signal bidirectional
rlabel metal3 s 79944 997600 84944 1014070 6 mprj_analog[9]
port 537 nsew signal bidirectional
rlabel metal5 s 76410 1018624 88578 1030789 6 mprj_io[23]
port 538 nsew signal bidirectional
rlabel metal3 s 23530 960144 40000 965144 6 mprj_analog[10]
port 539 nsew signal bidirectional
rlabel metal5 s 6811 956610 18976 968778 6 mprj_io[24]
port 540 nsew signal bidirectional
rlabel metal3 s 290878 997600 305200 1000737 6 mprj_analog[5]
port 541 nsew signal bidirectional
rlabel metal2 s 290878 997600 295658 1002732 6 mprj_clamp_high[1]
port 542 nsew signal input
rlabel metal2 s 280899 997600 285679 998011 6 mprj_clamp_low[1]
port 543 nsew signal input
rlabel metal5 s 282210 1018624 294378 1030789 6 mprj_io[19]
port 544 nsew signal bidirectional
rlabel metal3 s 239478 997600 253800 1000737 6 mprj_analog[6]
port 545 nsew signal bidirectional
rlabel metal2 s 239478 997600 244258 1002732 6 mprj_clamp_high[2]
port 546 nsew signal input
rlabel metal2 s 229499 997600 234279 998011 6 mprj_clamp_low[2]
port 547 nsew signal input
rlabel metal5 s 230810 1018624 242978 1030789 6 mprj_io[20]
port 548 nsew signal bidirectional
rlabel metal5 s 6167 915054 19620 925934 6 vccd2_pad
port 549 nsew signal bidirectional
rlabel metal5 s 6811 484810 18976 496978 6 vdda2_pad
port 550 nsew signal bidirectional
rlabel metal5 s 6811 829810 18976 841978 6 vssa2_pad
port 551 nsew signal bidirectional
rlabel metal4 s 38503 455946 39593 483654 6 vccd
port 552 nsew signal bidirectional
rlabel metal4 s 37293 455946 38223 483654 6 vccd2
port 553 nsew signal bidirectional
rlabel metal4 s 36323 456007 37013 483593 6 vdda2
port 554 nsew signal bidirectional
rlabel metal4 s 32933 455946 33623 483654 6 vddio
port 555 nsew signal bidirectional
rlabel metal4 s 28653 407418 28719 526322 6 vssa2
port 556 nsew signal bidirectional
rlabel metal3 s 31680 441300 39600 446100 6 vssd2
port 557 nsew signal bidirectional
rlabel metal5 s 6167 443254 19620 454134 6 vssd2_pad
port 558 nsew signal bidirectional
rlabel metal4 s 0 455946 4843 456200 6 vssio
port 559 nsew signal bidirectional
rlabel metal4 s 7 456200 4843 456493 6 vssio
port 559 nsew signal bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 717600 1037600
string LEFview TRUE
string GDS_FILE /project/openlane/chip_io_alt/runs/chip_io_alt/results/magic/chip_io_alt.gds
string GDS_END 36733536
string GDS_START 36371924
<< end >>

