VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io
  CLASS BLOCK ;
  FOREIGN chip_io ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 938.200 32.990 1000.800 95.440 ;
    END
  END clock
  PIN clock_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.635 208.565 936.915 210.965 ;
    END
  END clock_core
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.215 208.565 970.495 210.965 ;
    END
  END por
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1755.200 32.990 1817.800 95.440 ;
    END
  END flash_clk
  PIN flash_clk_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.835 208.565 1809.115 210.965 ;
    END
  END flash_clk_core
  PIN flash_clk_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.215 208.565 1787.495 210.965 ;
    END
  END flash_clk_ieb_core
  PIN flash_clk_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.475 208.565 1824.755 210.965 ;
    END
  END flash_clk_oeb_core
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1481.200 32.990 1543.800 95.440 ;
    END
  END flash_csb
  PIN flash_csb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.835 208.565 1535.115 210.965 ;
    END
  END flash_csb_core
  PIN flash_csb_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.215 208.565 1513.495 210.965 ;
    END
  END flash_csb_ieb_core
  PIN flash_csb_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.475 208.565 1550.755 210.965 ;
    END
  END flash_csb_oeb_core
  PIN flash_io0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2029.200 32.990 2091.800 95.440 ;
    END
  END flash_io0
  PIN flash_io0_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.635 208.565 2027.915 210.965 ;
    END
  END flash_io0_di_core
  PIN flash_io0_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.835 208.565 2083.115 210.965 ;
    END
  END flash_io0_do_core
  PIN flash_io0_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2046.610 209.000 2046.930 209.060 ;
        RECT 2061.790 209.000 2062.110 209.060 ;
        RECT 2076.050 209.000 2076.370 209.060 ;
        RECT 2046.610 208.860 2076.370 209.000 ;
        RECT 2046.610 208.800 2046.930 208.860 ;
        RECT 2061.790 208.800 2062.110 208.860 ;
        RECT 2076.050 208.800 2076.370 208.860 ;
      LAYER via ;
        RECT 2046.640 208.800 2046.900 209.060 ;
        RECT 2061.820 208.800 2062.080 209.060 ;
        RECT 2076.080 208.800 2076.340 209.060 ;
      LAYER met2 ;
        RECT 2046.035 209.170 2046.315 210.965 ;
        RECT 2061.215 209.170 2061.495 210.965 ;
        RECT 2076.855 209.170 2077.135 210.965 ;
        RECT 2046.035 209.090 2046.840 209.170 ;
        RECT 2061.215 209.090 2062.020 209.170 ;
        RECT 2076.140 209.090 2077.135 209.170 ;
        RECT 2046.035 209.030 2046.900 209.090 ;
        RECT 2046.035 208.565 2046.315 209.030 ;
        RECT 2046.640 208.770 2046.900 209.030 ;
        RECT 2061.215 209.030 2062.080 209.090 ;
        RECT 2061.215 208.565 2061.495 209.030 ;
        RECT 2061.820 208.770 2062.080 209.030 ;
        RECT 2076.080 209.030 2077.135 209.090 ;
        RECT 2076.080 208.770 2076.340 209.030 ;
        RECT 2076.855 208.565 2077.135 209.030 ;
    END
  END flash_io0_ieb_core
  PIN flash_io0_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2055.350 221.240 2055.670 221.300 ;
        RECT 2098.590 221.240 2098.910 221.300 ;
        RECT 2055.350 221.100 2098.910 221.240 ;
        RECT 2055.350 221.040 2055.670 221.100 ;
        RECT 2098.590 221.040 2098.910 221.100 ;
      LAYER via ;
        RECT 2055.380 221.040 2055.640 221.300 ;
        RECT 2098.620 221.040 2098.880 221.300 ;
      LAYER met2 ;
        RECT 2055.380 221.010 2055.640 221.330 ;
        RECT 2098.620 221.010 2098.880 221.330 ;
        RECT 2055.440 210.965 2055.580 221.010 ;
        RECT 2098.680 210.965 2098.820 221.010 ;
        RECT 2055.235 209.100 2055.580 210.965 ;
        RECT 2098.475 209.100 2098.820 210.965 ;
        RECT 2055.235 208.565 2055.515 209.100 ;
        RECT 2098.475 208.565 2098.755 209.100 ;
    END
  END flash_io0_oeb_core
  PIN flash_io1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2303.200 32.990 2365.800 95.440 ;
    END
  END flash_io1
  PIN flash_io1_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.635 208.565 2301.915 210.965 ;
    END
  END flash_io1_di_core
  PIN flash_io1_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.835 208.565 2357.115 210.965 ;
    END
  END flash_io1_do_core
  PIN flash_io1_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2320.770 209.340 2321.090 209.400 ;
        RECT 2335.950 209.340 2336.270 209.400 ;
        RECT 2350.210 209.340 2350.530 209.400 ;
        RECT 2320.770 209.200 2350.530 209.340 ;
        RECT 2320.770 209.140 2321.090 209.200 ;
        RECT 2335.950 209.140 2336.270 209.200 ;
        RECT 2350.210 209.140 2350.530 209.200 ;
      LAYER via ;
        RECT 2320.800 209.140 2321.060 209.400 ;
        RECT 2335.980 209.140 2336.240 209.400 ;
        RECT 2350.240 209.140 2350.500 209.400 ;
      LAYER met2 ;
        RECT 2320.035 209.170 2320.315 210.965 ;
        RECT 2320.800 209.170 2321.060 209.430 ;
        RECT 2320.035 209.110 2321.060 209.170 ;
        RECT 2335.215 209.170 2335.495 210.965 ;
        RECT 2335.980 209.170 2336.240 209.430 ;
        RECT 2335.215 209.110 2336.240 209.170 ;
        RECT 2350.240 209.170 2350.500 209.430 ;
        RECT 2350.855 209.170 2351.135 210.965 ;
        RECT 2350.240 209.110 2351.135 209.170 ;
        RECT 2320.035 209.030 2321.000 209.110 ;
        RECT 2335.215 209.030 2336.180 209.110 ;
        RECT 2350.300 209.030 2351.135 209.110 ;
        RECT 2320.035 208.565 2320.315 209.030 ;
        RECT 2335.215 208.565 2335.495 209.030 ;
        RECT 2350.855 208.565 2351.135 209.030 ;
    END
  END flash_io1_ieb_core
  PIN flash_io1_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.070 221.155 2329.350 221.525 ;
        RECT 2372.310 221.155 2372.590 221.525 ;
        RECT 2329.140 210.965 2329.280 221.155 ;
        RECT 2372.380 210.965 2372.520 221.155 ;
        RECT 2329.140 209.030 2329.515 210.965 ;
        RECT 2372.380 209.030 2372.755 210.965 ;
        RECT 2329.235 208.565 2329.515 209.030 ;
        RECT 2372.475 208.565 2372.755 209.030 ;
      LAYER via2 ;
        RECT 2329.070 221.200 2329.350 221.480 ;
        RECT 2372.310 221.200 2372.590 221.480 ;
      LAYER met3 ;
        RECT 2329.045 221.490 2329.375 221.505 ;
        RECT 2372.285 221.490 2372.615 221.505 ;
        RECT 2329.045 221.190 2372.615 221.490 ;
        RECT 2329.045 221.175 2329.375 221.190 ;
        RECT 2372.285 221.175 2372.615 221.190 ;
    END
  END flash_io1_oeb_core
  PIN gpio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2577.200 32.990 2639.800 95.440 ;
    END
  END gpio
  PIN gpio_in_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.635 208.565 2575.915 210.965 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.215 208.565 2609.495 210.965 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.235 208.565 2603.515 210.965 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.030 221.155 2594.310 221.525 ;
        RECT 2624.850 221.155 2625.130 221.525 ;
        RECT 2594.100 210.965 2594.240 221.155 ;
        RECT 2624.920 210.965 2625.060 221.155 ;
        RECT 2594.035 208.565 2594.315 210.965 ;
        RECT 2624.855 208.565 2625.135 210.965 ;
      LAYER via2 ;
        RECT 2594.030 221.200 2594.310 221.480 ;
        RECT 2624.850 221.200 2625.130 221.480 ;
      LAYER met3 ;
        RECT 2594.005 221.490 2594.335 221.505 ;
        RECT 2624.825 221.490 2625.155 221.505 ;
        RECT 2594.005 221.190 2625.155 221.490 ;
        RECT 2594.005 221.175 2594.335 221.190 ;
        RECT 2624.825 221.175 2625.155 221.190 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.835 208.565 2631.115 210.965 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.475 208.565 2646.755 210.965 ;
    END
  END gpio_outenb_core
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 186.465 202.730 191.115 341.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 30.835 350.270 98.100 404.670 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 186.465 413.730 191.115 552.270 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 186.565 202.730 191.015 341.270 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 186.565 413.730 191.015 552.270 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 191.100 340.500 198.000 364.500 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1987.270 4954.040 1987.590 4954.100 ;
        RECT 1988.190 4954.040 1988.510 4954.100 ;
        RECT 2433.010 4954.040 2433.330 4954.100 ;
        RECT 2690.150 4954.040 2690.470 4954.100 ;
        RECT 3198.910 4954.040 3199.230 4954.100 ;
        RECT 1987.270 4953.900 3199.230 4954.040 ;
        RECT 1987.270 4953.840 1987.590 4953.900 ;
        RECT 1988.190 4953.840 1988.510 4953.900 ;
        RECT 2433.010 4953.840 2433.330 4953.900 ;
        RECT 2690.150 4953.840 2690.470 4953.900 ;
        RECT 3198.910 4953.840 3199.230 4953.900 ;
        RECT 449.950 4953.700 450.270 4953.760 ;
        RECT 707.090 4953.700 707.410 4953.760 ;
        RECT 964.230 4953.700 964.550 4953.760 ;
        RECT 449.950 4953.560 964.550 4953.700 ;
        RECT 449.950 4953.500 450.270 4953.560 ;
        RECT 707.090 4953.500 707.410 4953.560 ;
        RECT 964.230 4953.500 964.550 4953.560 ;
        RECT 974.810 4953.700 975.130 4953.760 ;
        RECT 1220.910 4953.700 1221.230 4953.760 ;
        RECT 1478.970 4953.700 1479.290 4953.760 ;
        RECT 974.810 4953.560 1479.290 4953.700 ;
        RECT 974.810 4953.500 975.130 4953.560 ;
        RECT 1220.910 4953.500 1221.230 4953.560 ;
        RECT 1478.970 4953.500 1479.290 4953.560 ;
        RECT 1478.970 4952.680 1479.290 4952.740 ;
        RECT 1987.270 4952.680 1987.590 4952.740 ;
        RECT 1478.970 4952.540 1987.590 4952.680 ;
        RECT 1478.970 4952.480 1479.290 4952.540 ;
        RECT 1987.270 4952.480 1987.590 4952.540 ;
        RECT 964.230 4952.340 964.550 4952.400 ;
        RECT 974.810 4952.340 975.130 4952.400 ;
        RECT 964.230 4952.200 975.130 4952.340 ;
        RECT 964.230 4952.140 964.550 4952.200 ;
        RECT 974.810 4952.140 975.130 4952.200 ;
        RECT 3198.910 4950.980 3199.230 4951.040 ;
        RECT 3368.190 4950.980 3368.510 4951.040 ;
        RECT 3198.910 4950.840 3368.510 4950.980 ;
        RECT 3198.910 4950.780 3199.230 4950.840 ;
        RECT 3368.190 4950.780 3368.510 4950.840 ;
        RECT 449.490 4950.440 449.810 4950.700 ;
        RECT 212.590 4950.300 212.910 4950.360 ;
        RECT 449.580 4950.300 449.720 4950.440 ;
        RECT 212.590 4950.160 449.720 4950.300 ;
        RECT 212.590 4950.100 212.910 4950.160 ;
        RECT 208.910 4842.520 209.230 4842.580 ;
        RECT 212.590 4842.520 212.910 4842.580 ;
        RECT 208.910 4842.380 212.910 4842.520 ;
        RECT 208.910 4842.320 209.230 4842.380 ;
        RECT 212.590 4842.320 212.910 4842.380 ;
        RECT 3368.190 4766.700 3368.510 4766.760 ;
        RECT 3376.930 4766.700 3377.250 4766.760 ;
        RECT 3368.190 4766.560 3377.250 4766.700 ;
        RECT 3368.190 4766.500 3368.510 4766.560 ;
        RECT 3376.930 4766.500 3377.250 4766.560 ;
        RECT 3368.190 4322.320 3368.510 4322.380 ;
        RECT 3376.930 4322.320 3377.250 4322.380 ;
        RECT 3368.190 4322.180 3377.250 4322.320 ;
        RECT 3368.190 4322.120 3368.510 4322.180 ;
        RECT 3376.930 4322.120 3377.250 4322.180 ;
        RECT 208.910 3988.780 209.230 3988.840 ;
        RECT 212.590 3988.780 212.910 3988.840 ;
        RECT 213.510 3988.780 213.830 3988.840 ;
        RECT 208.910 3988.640 213.830 3988.780 ;
        RECT 208.910 3988.580 209.230 3988.640 ;
        RECT 212.590 3988.580 212.910 3988.640 ;
        RECT 213.510 3988.580 213.830 3988.640 ;
        RECT 3367.270 3874.540 3367.590 3874.600 ;
        RECT 3368.190 3874.540 3368.510 3874.600 ;
        RECT 3376.930 3874.540 3377.250 3874.600 ;
        RECT 3367.270 3874.400 3377.250 3874.540 ;
        RECT 3367.270 3874.340 3367.590 3874.400 ;
        RECT 3368.190 3874.340 3368.510 3874.400 ;
        RECT 3376.930 3874.340 3377.250 3874.400 ;
        RECT 212.130 3836.800 212.450 3836.860 ;
        RECT 213.510 3836.800 213.830 3836.860 ;
        RECT 212.130 3836.660 213.830 3836.800 ;
        RECT 212.130 3836.600 212.450 3836.660 ;
        RECT 213.510 3836.600 213.830 3836.660 ;
        RECT 208.910 3772.540 209.230 3772.600 ;
        RECT 212.130 3772.540 212.450 3772.600 ;
        RECT 208.910 3772.400 212.450 3772.540 ;
        RECT 208.910 3772.340 209.230 3772.400 ;
        RECT 212.130 3772.340 212.450 3772.400 ;
        RECT 3367.270 3650.820 3367.590 3650.880 ;
        RECT 3376.930 3650.820 3377.250 3650.880 ;
        RECT 3367.270 3650.680 3377.250 3650.820 ;
        RECT 3367.270 3650.620 3367.590 3650.680 ;
        RECT 3376.930 3650.620 3377.250 3650.680 ;
        RECT 208.910 3556.640 209.230 3556.700 ;
        RECT 212.130 3556.640 212.450 3556.700 ;
        RECT 213.510 3556.640 213.830 3556.700 ;
        RECT 208.910 3556.500 213.830 3556.640 ;
        RECT 208.910 3556.440 209.230 3556.500 ;
        RECT 212.130 3556.440 212.450 3556.500 ;
        RECT 213.510 3556.440 213.830 3556.500 ;
        RECT 3367.270 3426.080 3367.590 3426.140 ;
        RECT 3376.930 3426.080 3377.250 3426.140 ;
        RECT 3367.270 3425.940 3377.250 3426.080 ;
        RECT 3367.270 3425.880 3367.590 3425.940 ;
        RECT 3376.930 3425.880 3377.250 3425.940 ;
        RECT 208.910 3345.500 209.230 3345.560 ;
        RECT 212.590 3345.500 212.910 3345.560 ;
        RECT 208.910 3345.360 212.910 3345.500 ;
        RECT 208.910 3345.300 209.230 3345.360 ;
        RECT 212.590 3345.300 212.910 3345.360 ;
        RECT 3367.270 3198.620 3367.590 3198.680 ;
        RECT 3369.570 3198.620 3369.890 3198.680 ;
        RECT 3376.930 3198.620 3377.250 3198.680 ;
        RECT 3367.270 3198.480 3377.250 3198.620 ;
        RECT 3367.270 3198.420 3367.590 3198.480 ;
        RECT 3369.570 3198.420 3369.890 3198.480 ;
        RECT 3376.930 3198.420 3377.250 3198.480 ;
        RECT 212.590 3160.000 212.910 3160.260 ;
        RECT 212.680 3159.520 212.820 3160.000 ;
        RECT 213.970 3159.520 214.290 3159.580 ;
        RECT 212.680 3159.380 214.290 3159.520 ;
        RECT 213.970 3159.320 214.290 3159.380 ;
        RECT 208.910 3124.840 209.230 3124.900 ;
        RECT 213.970 3124.840 214.290 3124.900 ;
        RECT 208.910 3124.700 214.290 3124.840 ;
        RECT 208.910 3124.640 209.230 3124.700 ;
        RECT 213.970 3124.640 214.290 3124.700 ;
        RECT 213.970 3064.120 214.290 3064.380 ;
        RECT 213.050 3063.980 213.370 3064.040 ;
        RECT 214.060 3063.980 214.200 3064.120 ;
        RECT 213.050 3063.840 214.200 3063.980 ;
        RECT 213.050 3063.780 213.370 3063.840 ;
        RECT 213.050 3063.300 213.370 3063.360 ;
        RECT 213.970 3063.300 214.290 3063.360 ;
        RECT 213.050 3063.160 214.290 3063.300 ;
        RECT 213.050 3063.100 213.370 3063.160 ;
        RECT 213.970 3063.100 214.290 3063.160 ;
        RECT 3368.190 2974.560 3368.510 2974.620 ;
        RECT 3369.570 2974.560 3369.890 2974.620 ;
        RECT 3376.930 2974.560 3377.250 2974.620 ;
        RECT 3368.190 2974.420 3377.250 2974.560 ;
        RECT 3368.190 2974.360 3368.510 2974.420 ;
        RECT 3369.570 2974.360 3369.890 2974.420 ;
        RECT 3376.930 2974.360 3377.250 2974.420 ;
        RECT 208.910 2913.360 209.230 2913.420 ;
        RECT 213.970 2913.360 214.290 2913.420 ;
        RECT 208.910 2913.220 214.290 2913.360 ;
        RECT 208.910 2913.160 209.230 2913.220 ;
        RECT 213.970 2913.160 214.290 2913.220 ;
        RECT 211.670 2870.520 211.990 2870.580 ;
        RECT 213.970 2870.520 214.290 2870.580 ;
        RECT 211.670 2870.380 214.290 2870.520 ;
        RECT 211.670 2870.320 211.990 2870.380 ;
        RECT 213.970 2870.320 214.290 2870.380 ;
        RECT 3368.190 2752.540 3368.510 2752.600 ;
        RECT 3376.930 2752.540 3377.250 2752.600 ;
        RECT 3368.190 2752.400 3377.250 2752.540 ;
        RECT 3368.190 2752.340 3368.510 2752.400 ;
        RECT 3376.930 2752.340 3377.250 2752.400 ;
        RECT 208.910 2697.460 209.230 2697.520 ;
        RECT 212.590 2697.460 212.910 2697.520 ;
        RECT 208.910 2697.320 212.910 2697.460 ;
        RECT 208.910 2697.260 209.230 2697.320 ;
        RECT 212.590 2697.260 212.910 2697.320 ;
        RECT 208.910 2056.220 209.230 2056.280 ;
        RECT 212.590 2056.220 212.910 2056.280 ;
        RECT 208.910 2056.080 212.910 2056.220 ;
        RECT 208.910 2056.020 209.230 2056.080 ;
        RECT 212.590 2056.020 212.910 2056.080 ;
        RECT 213.050 1931.780 213.370 1931.840 ;
        RECT 214.430 1931.780 214.750 1931.840 ;
        RECT 213.050 1931.640 214.750 1931.780 ;
        RECT 213.050 1931.580 213.370 1931.640 ;
        RECT 214.430 1931.580 214.750 1931.640 ;
        RECT 3368.650 1861.740 3368.970 1861.800 ;
        RECT 3376.930 1861.740 3377.250 1861.800 ;
        RECT 3368.650 1861.600 3377.250 1861.740 ;
        RECT 3368.650 1861.540 3368.970 1861.600 ;
        RECT 3376.930 1861.540 3377.250 1861.600 ;
        RECT 208.910 1843.380 209.230 1843.440 ;
        RECT 214.430 1843.380 214.750 1843.440 ;
        RECT 208.910 1843.240 214.750 1843.380 ;
        RECT 208.910 1843.180 209.230 1843.240 ;
        RECT 214.430 1843.180 214.750 1843.240 ;
        RECT 3368.650 1640.400 3368.970 1640.460 ;
        RECT 3376.930 1640.400 3377.250 1640.460 ;
        RECT 3368.650 1640.260 3377.250 1640.400 ;
        RECT 3368.650 1640.200 3368.970 1640.260 ;
        RECT 3376.930 1640.200 3377.250 1640.260 ;
        RECT 208.910 1627.480 209.230 1627.540 ;
        RECT 212.130 1627.480 212.450 1627.540 ;
        RECT 213.510 1627.480 213.830 1627.540 ;
        RECT 208.910 1627.340 213.830 1627.480 ;
        RECT 208.910 1627.280 209.230 1627.340 ;
        RECT 212.130 1627.280 212.450 1627.340 ;
        RECT 213.510 1627.280 213.830 1627.340 ;
        RECT 212.130 1614.560 212.450 1614.620 ;
        RECT 212.130 1614.420 213.740 1614.560 ;
        RECT 212.130 1614.360 212.450 1614.420 ;
        RECT 213.600 1614.280 213.740 1614.420 ;
        RECT 213.510 1614.020 213.830 1614.280 ;
        RECT 211.670 1571.040 211.990 1571.100 ;
        RECT 213.510 1571.040 213.830 1571.100 ;
        RECT 211.670 1570.900 213.830 1571.040 ;
        RECT 211.670 1570.840 211.990 1570.900 ;
        RECT 213.510 1570.840 213.830 1570.900 ;
        RECT 208.910 1411.580 209.230 1411.640 ;
        RECT 212.590 1411.580 212.910 1411.640 ;
        RECT 208.910 1411.440 212.910 1411.580 ;
        RECT 208.910 1411.380 209.230 1411.440 ;
        RECT 212.590 1411.380 212.910 1411.440 ;
        RECT 3368.650 1410.560 3368.970 1410.620 ;
        RECT 3376.930 1410.560 3377.250 1410.620 ;
        RECT 3368.650 1410.420 3377.250 1410.560 ;
        RECT 3368.650 1410.360 3368.970 1410.420 ;
        RECT 3376.930 1410.360 3377.250 1410.420 ;
        RECT 211.670 1227.980 211.990 1228.040 ;
        RECT 214.430 1227.980 214.750 1228.040 ;
        RECT 211.670 1227.840 214.750 1227.980 ;
        RECT 211.670 1227.780 211.990 1227.840 ;
        RECT 214.430 1227.780 214.750 1227.840 ;
        RECT 208.910 1190.580 209.230 1190.640 ;
        RECT 213.050 1190.580 213.370 1190.640 ;
        RECT 214.430 1190.580 214.750 1190.640 ;
        RECT 208.910 1190.440 214.750 1190.580 ;
        RECT 208.910 1190.380 209.230 1190.440 ;
        RECT 213.050 1190.380 213.370 1190.440 ;
        RECT 214.430 1190.380 214.750 1190.440 ;
        RECT 3369.570 1188.540 3369.890 1188.600 ;
        RECT 3376.930 1188.540 3377.250 1188.600 ;
        RECT 3369.570 1188.400 3377.250 1188.540 ;
        RECT 3369.570 1188.340 3369.890 1188.400 ;
        RECT 3376.930 1188.340 3377.250 1188.400 ;
        RECT 3369.570 1186.840 3369.890 1186.900 ;
        RECT 3370.490 1186.840 3370.810 1186.900 ;
        RECT 3369.570 1186.700 3370.810 1186.840 ;
        RECT 3369.570 1186.640 3369.890 1186.700 ;
        RECT 3370.490 1186.640 3370.810 1186.700 ;
        RECT 211.670 1164.400 211.990 1164.460 ;
        RECT 213.050 1164.400 213.370 1164.460 ;
        RECT 211.670 1164.260 213.370 1164.400 ;
        RECT 211.670 1164.200 211.990 1164.260 ;
        RECT 213.050 1164.200 213.370 1164.260 ;
        RECT 3370.490 1158.960 3370.810 1159.020 ;
        RECT 3371.410 1158.960 3371.730 1159.020 ;
        RECT 3370.490 1158.820 3371.730 1158.960 ;
        RECT 3370.490 1158.760 3370.810 1158.820 ;
        RECT 3371.410 1158.760 3371.730 1158.820 ;
        RECT 3370.030 1062.740 3370.350 1062.800 ;
        RECT 3371.410 1062.740 3371.730 1062.800 ;
        RECT 3370.030 1062.600 3371.730 1062.740 ;
        RECT 3370.030 1062.540 3370.350 1062.600 ;
        RECT 3371.410 1062.540 3371.730 1062.600 ;
        RECT 211.670 1042.000 211.990 1042.060 ;
        RECT 214.430 1042.000 214.750 1042.060 ;
        RECT 211.670 1041.860 214.750 1042.000 ;
        RECT 211.670 1041.800 211.990 1041.860 ;
        RECT 214.430 1041.800 214.750 1041.860 ;
        RECT 3370.030 993.720 3370.350 993.780 ;
        RECT 3376.010 993.720 3376.330 993.780 ;
        RECT 3370.030 993.580 3376.330 993.720 ;
        RECT 3370.030 993.520 3370.350 993.580 ;
        RECT 3376.010 993.520 3376.330 993.580 ;
        RECT 208.910 974.680 209.230 974.740 ;
        RECT 212.130 974.680 212.450 974.740 ;
        RECT 214.430 974.680 214.750 974.740 ;
        RECT 208.910 974.540 214.750 974.680 ;
        RECT 208.910 974.480 209.230 974.540 ;
        RECT 212.130 974.480 212.450 974.540 ;
        RECT 214.430 974.480 214.750 974.540 ;
        RECT 3373.710 960.740 3374.030 960.800 ;
        RECT 3376.010 960.740 3376.330 960.800 ;
        RECT 3376.930 960.740 3377.250 960.800 ;
        RECT 3373.710 960.600 3377.250 960.740 ;
        RECT 3373.710 960.540 3374.030 960.600 ;
        RECT 3376.010 960.540 3376.330 960.600 ;
        RECT 3376.930 960.540 3377.250 960.600 ;
        RECT 212.130 926.740 212.450 926.800 ;
        RECT 213.510 926.740 213.830 926.800 ;
        RECT 212.130 926.600 213.830 926.740 ;
        RECT 212.130 926.540 212.450 926.600 ;
        RECT 213.510 926.540 213.830 926.600 ;
        RECT 3369.110 869.620 3369.430 869.680 ;
        RECT 3373.710 869.620 3374.030 869.680 ;
        RECT 3369.110 869.480 3374.030 869.620 ;
        RECT 3369.110 869.420 3369.430 869.480 ;
        RECT 3373.710 869.420 3374.030 869.480 ;
        RECT 212.590 745.520 212.910 745.580 ;
        RECT 213.510 745.520 213.830 745.580 ;
        RECT 212.590 745.380 213.830 745.520 ;
        RECT 212.590 745.320 212.910 745.380 ;
        RECT 213.510 745.320 213.830 745.380 ;
        RECT 3368.190 735.660 3368.510 735.720 ;
        RECT 3375.090 735.660 3375.410 735.720 ;
        RECT 3376.930 735.660 3377.250 735.720 ;
        RECT 3368.190 735.520 3377.250 735.660 ;
        RECT 3368.190 735.460 3368.510 735.520 ;
        RECT 3375.090 735.460 3375.410 735.520 ;
        RECT 3376.930 735.460 3377.250 735.520 ;
        RECT 3370.030 703.360 3370.350 703.420 ;
        RECT 3375.090 703.360 3375.410 703.420 ;
        RECT 3370.030 703.220 3375.410 703.360 ;
        RECT 3370.030 703.160 3370.350 703.220 ;
        RECT 3375.090 703.160 3375.410 703.220 ;
        RECT 3369.110 579.940 3369.430 580.000 ;
        RECT 3370.030 579.940 3370.350 580.000 ;
        RECT 3369.110 579.800 3370.350 579.940 ;
        RECT 3369.110 579.740 3369.430 579.800 ;
        RECT 3370.030 579.740 3370.350 579.800 ;
        RECT 3369.110 579.260 3369.430 579.320 ;
        RECT 3375.090 579.260 3375.410 579.320 ;
        RECT 3369.110 579.120 3375.410 579.260 ;
        RECT 3369.110 579.060 3369.430 579.120 ;
        RECT 3375.090 579.060 3375.410 579.120 ;
        RECT 212.590 552.400 212.910 552.460 ;
        RECT 213.510 552.400 213.830 552.460 ;
        RECT 212.590 552.260 213.830 552.400 ;
        RECT 212.590 552.200 212.910 552.260 ;
        RECT 213.510 552.200 213.830 552.260 ;
        RECT 3368.190 511.600 3368.510 511.660 ;
        RECT 3375.090 511.600 3375.410 511.660 ;
        RECT 3376.930 511.600 3377.250 511.660 ;
        RECT 3368.190 511.460 3377.250 511.600 ;
        RECT 3368.190 511.400 3368.510 511.460 ;
        RECT 3375.090 511.400 3375.410 511.460 ;
        RECT 3376.930 511.400 3377.250 511.460 ;
        RECT 213.510 228.040 213.830 228.100 ;
        RECT 717.670 228.040 717.990 228.100 ;
        RECT 213.510 227.900 717.990 228.040 ;
        RECT 213.510 227.840 213.830 227.900 ;
        RECT 717.670 227.840 717.990 227.900 ;
        RECT 2581.590 227.700 2581.910 227.760 ;
        RECT 3368.190 227.700 3368.510 227.760 ;
        RECT 2581.590 227.560 3368.510 227.700 ;
        RECT 2581.590 227.500 2581.910 227.560 ;
        RECT 3368.190 227.500 3368.510 227.560 ;
        RECT 2033.730 223.620 2034.050 223.680 ;
        RECT 2125.270 223.620 2125.590 223.680 ;
        RECT 2220.950 223.620 2221.270 223.680 ;
        RECT 2033.730 223.480 2056.500 223.620 ;
        RECT 2033.730 223.420 2034.050 223.480 ;
        RECT 2056.360 222.940 2056.500 223.480 ;
        RECT 2125.270 223.480 2221.270 223.620 ;
        RECT 2125.270 223.420 2125.590 223.480 ;
        RECT 2220.950 223.420 2221.270 223.480 ;
        RECT 2415.070 223.280 2415.390 223.340 ;
        RECT 2366.400 223.140 2415.390 223.280 ;
        RECT 2125.270 222.940 2125.590 223.000 ;
        RECT 2307.430 222.940 2307.750 223.000 ;
        RECT 2345.610 222.940 2345.930 223.000 ;
        RECT 2056.360 222.800 2125.590 222.940 ;
        RECT 2125.270 222.740 2125.590 222.800 ;
        RECT 2249.100 222.800 2345.930 222.940 ;
        RECT 1771.990 222.600 1772.310 222.660 ;
        RECT 1802.810 222.600 1803.130 222.660 ;
        RECT 1771.990 222.460 1803.130 222.600 ;
        RECT 1771.990 222.400 1772.310 222.460 ;
        RECT 1802.810 222.400 1803.130 222.460 ;
        RECT 1998.310 222.600 1998.630 222.660 ;
        RECT 2033.730 222.600 2034.050 222.660 ;
        RECT 1998.310 222.460 2034.050 222.600 ;
        RECT 1998.310 222.400 1998.630 222.460 ;
        RECT 2033.730 222.400 2034.050 222.460 ;
        RECT 2221.410 222.600 2221.730 222.660 ;
        RECT 2249.100 222.600 2249.240 222.800 ;
        RECT 2307.430 222.740 2307.750 222.800 ;
        RECT 2345.610 222.740 2345.930 222.800 ;
        RECT 2346.070 222.940 2346.390 223.000 ;
        RECT 2366.400 222.940 2366.540 223.140 ;
        RECT 2415.070 223.080 2415.390 223.140 ;
        RECT 2346.070 222.800 2366.540 222.940 ;
        RECT 2511.300 222.800 2511.900 222.940 ;
        RECT 2346.070 222.740 2346.390 222.800 ;
        RECT 2511.300 222.660 2511.440 222.800 ;
        RECT 2221.410 222.460 2249.240 222.600 ;
        RECT 2221.410 222.400 2221.730 222.460 ;
        RECT 2511.210 222.400 2511.530 222.660 ;
        RECT 2511.760 222.600 2511.900 222.800 ;
        RECT 2581.590 222.600 2581.910 222.660 ;
        RECT 2511.760 222.460 2581.910 222.600 ;
        RECT 2581.590 222.400 2581.910 222.460 ;
        RECT 942.610 221.580 942.930 221.640 ;
        RECT 964.230 221.580 964.550 221.640 ;
        RECT 1007.470 221.580 1007.790 221.640 ;
        RECT 1485.410 221.580 1485.730 221.640 ;
        RECT 1497.830 221.580 1498.150 221.640 ;
        RECT 1528.650 221.580 1528.970 221.640 ;
        RECT 1759.570 221.580 1759.890 221.640 ;
        RECT 1771.990 221.580 1772.310 221.640 ;
        RECT 942.610 221.440 1772.310 221.580 ;
        RECT 942.610 221.380 942.930 221.440 ;
        RECT 964.230 221.380 964.550 221.440 ;
        RECT 1007.470 221.380 1007.790 221.440 ;
        RECT 1485.410 221.380 1485.730 221.440 ;
        RECT 1497.830 221.380 1498.150 221.440 ;
        RECT 1528.650 221.380 1528.970 221.440 ;
        RECT 1759.570 221.380 1759.890 221.440 ;
        RECT 1771.990 221.380 1772.310 221.440 ;
        RECT 1802.810 221.580 1803.130 221.640 ;
        RECT 1998.310 221.580 1998.630 221.640 ;
        RECT 1802.810 221.440 1998.630 221.580 ;
        RECT 1802.810 221.380 1803.130 221.440 ;
        RECT 1998.310 221.380 1998.630 221.440 ;
        RECT 938.470 209.680 938.790 209.740 ;
        RECT 942.150 209.680 942.470 209.740 ;
        RECT 938.470 209.540 942.470 209.680 ;
        RECT 938.470 209.480 938.790 209.540 ;
        RECT 942.150 209.480 942.470 209.540 ;
        RECT 748.030 209.000 748.350 209.060 ;
        RECT 938.470 209.000 938.790 209.060 ;
        RECT 748.030 208.860 938.790 209.000 ;
        RECT 748.030 208.800 748.350 208.860 ;
        RECT 938.470 208.800 938.790 208.860 ;
      LAYER via ;
        RECT 1987.300 4953.840 1987.560 4954.100 ;
        RECT 1988.220 4953.840 1988.480 4954.100 ;
        RECT 2433.040 4953.840 2433.300 4954.100 ;
        RECT 2690.180 4953.840 2690.440 4954.100 ;
        RECT 3198.940 4953.840 3199.200 4954.100 ;
        RECT 449.980 4953.500 450.240 4953.760 ;
        RECT 707.120 4953.500 707.380 4953.760 ;
        RECT 964.260 4953.500 964.520 4953.760 ;
        RECT 974.840 4953.500 975.100 4953.760 ;
        RECT 1220.940 4953.500 1221.200 4953.760 ;
        RECT 1479.000 4953.500 1479.260 4953.760 ;
        RECT 1479.000 4952.480 1479.260 4952.740 ;
        RECT 1987.300 4952.480 1987.560 4952.740 ;
        RECT 964.260 4952.140 964.520 4952.400 ;
        RECT 974.840 4952.140 975.100 4952.400 ;
        RECT 3198.940 4950.780 3199.200 4951.040 ;
        RECT 3368.220 4950.780 3368.480 4951.040 ;
        RECT 449.520 4950.440 449.780 4950.700 ;
        RECT 212.620 4950.100 212.880 4950.360 ;
        RECT 208.940 4842.320 209.200 4842.580 ;
        RECT 212.620 4842.320 212.880 4842.580 ;
        RECT 3368.220 4766.500 3368.480 4766.760 ;
        RECT 3376.960 4766.500 3377.220 4766.760 ;
        RECT 3368.220 4322.120 3368.480 4322.380 ;
        RECT 3376.960 4322.120 3377.220 4322.380 ;
        RECT 208.940 3988.580 209.200 3988.840 ;
        RECT 212.620 3988.580 212.880 3988.840 ;
        RECT 213.540 3988.580 213.800 3988.840 ;
        RECT 3367.300 3874.340 3367.560 3874.600 ;
        RECT 3368.220 3874.340 3368.480 3874.600 ;
        RECT 3376.960 3874.340 3377.220 3874.600 ;
        RECT 212.160 3836.600 212.420 3836.860 ;
        RECT 213.540 3836.600 213.800 3836.860 ;
        RECT 208.940 3772.340 209.200 3772.600 ;
        RECT 212.160 3772.340 212.420 3772.600 ;
        RECT 3367.300 3650.620 3367.560 3650.880 ;
        RECT 3376.960 3650.620 3377.220 3650.880 ;
        RECT 208.940 3556.440 209.200 3556.700 ;
        RECT 212.160 3556.440 212.420 3556.700 ;
        RECT 213.540 3556.440 213.800 3556.700 ;
        RECT 3367.300 3425.880 3367.560 3426.140 ;
        RECT 3376.960 3425.880 3377.220 3426.140 ;
        RECT 208.940 3345.300 209.200 3345.560 ;
        RECT 212.620 3345.300 212.880 3345.560 ;
        RECT 3367.300 3198.420 3367.560 3198.680 ;
        RECT 3369.600 3198.420 3369.860 3198.680 ;
        RECT 3376.960 3198.420 3377.220 3198.680 ;
        RECT 212.620 3160.000 212.880 3160.260 ;
        RECT 214.000 3159.320 214.260 3159.580 ;
        RECT 208.940 3124.640 209.200 3124.900 ;
        RECT 214.000 3124.640 214.260 3124.900 ;
        RECT 214.000 3064.120 214.260 3064.380 ;
        RECT 213.080 3063.780 213.340 3064.040 ;
        RECT 213.080 3063.100 213.340 3063.360 ;
        RECT 214.000 3063.100 214.260 3063.360 ;
        RECT 3368.220 2974.360 3368.480 2974.620 ;
        RECT 3369.600 2974.360 3369.860 2974.620 ;
        RECT 3376.960 2974.360 3377.220 2974.620 ;
        RECT 208.940 2913.160 209.200 2913.420 ;
        RECT 214.000 2913.160 214.260 2913.420 ;
        RECT 211.700 2870.320 211.960 2870.580 ;
        RECT 214.000 2870.320 214.260 2870.580 ;
        RECT 3368.220 2752.340 3368.480 2752.600 ;
        RECT 3376.960 2752.340 3377.220 2752.600 ;
        RECT 208.940 2697.260 209.200 2697.520 ;
        RECT 212.620 2697.260 212.880 2697.520 ;
        RECT 208.940 2056.020 209.200 2056.280 ;
        RECT 212.620 2056.020 212.880 2056.280 ;
        RECT 213.080 1931.580 213.340 1931.840 ;
        RECT 214.460 1931.580 214.720 1931.840 ;
        RECT 3368.680 1861.540 3368.940 1861.800 ;
        RECT 3376.960 1861.540 3377.220 1861.800 ;
        RECT 208.940 1843.180 209.200 1843.440 ;
        RECT 214.460 1843.180 214.720 1843.440 ;
        RECT 3368.680 1640.200 3368.940 1640.460 ;
        RECT 3376.960 1640.200 3377.220 1640.460 ;
        RECT 208.940 1627.280 209.200 1627.540 ;
        RECT 212.160 1627.280 212.420 1627.540 ;
        RECT 213.540 1627.280 213.800 1627.540 ;
        RECT 212.160 1614.360 212.420 1614.620 ;
        RECT 213.540 1614.020 213.800 1614.280 ;
        RECT 211.700 1570.840 211.960 1571.100 ;
        RECT 213.540 1570.840 213.800 1571.100 ;
        RECT 208.940 1411.380 209.200 1411.640 ;
        RECT 212.620 1411.380 212.880 1411.640 ;
        RECT 3368.680 1410.360 3368.940 1410.620 ;
        RECT 3376.960 1410.360 3377.220 1410.620 ;
        RECT 211.700 1227.780 211.960 1228.040 ;
        RECT 214.460 1227.780 214.720 1228.040 ;
        RECT 208.940 1190.380 209.200 1190.640 ;
        RECT 213.080 1190.380 213.340 1190.640 ;
        RECT 214.460 1190.380 214.720 1190.640 ;
        RECT 3369.600 1188.340 3369.860 1188.600 ;
        RECT 3376.960 1188.340 3377.220 1188.600 ;
        RECT 3369.600 1186.640 3369.860 1186.900 ;
        RECT 3370.520 1186.640 3370.780 1186.900 ;
        RECT 211.700 1164.200 211.960 1164.460 ;
        RECT 213.080 1164.200 213.340 1164.460 ;
        RECT 3370.520 1158.760 3370.780 1159.020 ;
        RECT 3371.440 1158.760 3371.700 1159.020 ;
        RECT 3370.060 1062.540 3370.320 1062.800 ;
        RECT 3371.440 1062.540 3371.700 1062.800 ;
        RECT 211.700 1041.800 211.960 1042.060 ;
        RECT 214.460 1041.800 214.720 1042.060 ;
        RECT 3370.060 993.520 3370.320 993.780 ;
        RECT 3376.040 993.520 3376.300 993.780 ;
        RECT 208.940 974.480 209.200 974.740 ;
        RECT 212.160 974.480 212.420 974.740 ;
        RECT 214.460 974.480 214.720 974.740 ;
        RECT 3373.740 960.540 3374.000 960.800 ;
        RECT 3376.040 960.540 3376.300 960.800 ;
        RECT 3376.960 960.540 3377.220 960.800 ;
        RECT 212.160 926.540 212.420 926.800 ;
        RECT 213.540 926.540 213.800 926.800 ;
        RECT 3369.140 869.420 3369.400 869.680 ;
        RECT 3373.740 869.420 3374.000 869.680 ;
        RECT 212.620 745.320 212.880 745.580 ;
        RECT 213.540 745.320 213.800 745.580 ;
        RECT 3368.220 735.460 3368.480 735.720 ;
        RECT 3375.120 735.460 3375.380 735.720 ;
        RECT 3376.960 735.460 3377.220 735.720 ;
        RECT 3370.060 703.160 3370.320 703.420 ;
        RECT 3375.120 703.160 3375.380 703.420 ;
        RECT 3369.140 579.740 3369.400 580.000 ;
        RECT 3370.060 579.740 3370.320 580.000 ;
        RECT 3369.140 579.060 3369.400 579.320 ;
        RECT 3375.120 579.060 3375.380 579.320 ;
        RECT 212.620 552.200 212.880 552.460 ;
        RECT 213.540 552.200 213.800 552.460 ;
        RECT 3368.220 511.400 3368.480 511.660 ;
        RECT 3375.120 511.400 3375.380 511.660 ;
        RECT 3376.960 511.400 3377.220 511.660 ;
        RECT 213.540 227.840 213.800 228.100 ;
        RECT 717.700 227.840 717.960 228.100 ;
        RECT 2581.620 227.500 2581.880 227.760 ;
        RECT 3368.220 227.500 3368.480 227.760 ;
        RECT 2033.760 223.420 2034.020 223.680 ;
        RECT 2125.300 223.420 2125.560 223.680 ;
        RECT 2220.980 223.420 2221.240 223.680 ;
        RECT 2125.300 222.740 2125.560 223.000 ;
        RECT 1772.020 222.400 1772.280 222.660 ;
        RECT 1802.840 222.400 1803.100 222.660 ;
        RECT 1998.340 222.400 1998.600 222.660 ;
        RECT 2033.760 222.400 2034.020 222.660 ;
        RECT 2221.440 222.400 2221.700 222.660 ;
        RECT 2307.460 222.740 2307.720 223.000 ;
        RECT 2345.640 222.740 2345.900 223.000 ;
        RECT 2346.100 222.740 2346.360 223.000 ;
        RECT 2415.100 223.080 2415.360 223.340 ;
        RECT 2511.240 222.400 2511.500 222.660 ;
        RECT 2581.620 222.400 2581.880 222.660 ;
        RECT 942.640 221.380 942.900 221.640 ;
        RECT 964.260 221.380 964.520 221.640 ;
        RECT 1007.500 221.380 1007.760 221.640 ;
        RECT 1485.440 221.380 1485.700 221.640 ;
        RECT 1497.860 221.380 1498.120 221.640 ;
        RECT 1528.680 221.380 1528.940 221.640 ;
        RECT 1759.600 221.380 1759.860 221.640 ;
        RECT 1772.020 221.380 1772.280 221.640 ;
        RECT 1802.840 221.380 1803.100 221.640 ;
        RECT 1998.340 221.380 1998.600 221.640 ;
        RECT 938.500 209.480 938.760 209.740 ;
        RECT 942.180 209.480 942.440 209.740 ;
        RECT 748.060 208.800 748.320 209.060 ;
        RECT 938.500 208.800 938.760 209.060 ;
      LAYER met2 ;
        RECT 450.105 4977.260 450.385 4979.435 ;
        RECT 450.040 4977.035 450.385 4977.260 ;
        RECT 707.105 4977.035 707.385 4979.435 ;
        RECT 964.105 4977.330 964.385 4979.435 ;
        RECT 1221.105 4977.330 1221.385 4979.435 ;
        RECT 964.105 4977.035 964.460 4977.330 ;
        RECT 450.040 4953.790 450.180 4977.035 ;
        RECT 707.180 4953.790 707.320 4977.035 ;
        RECT 964.320 4953.790 964.460 4977.035 ;
        RECT 1221.000 4977.035 1221.385 4977.330 ;
        RECT 1479.105 4977.260 1479.385 4979.435 ;
        RECT 1479.060 4977.035 1479.385 4977.260 ;
        RECT 1988.105 4977.260 1988.385 4979.435 ;
        RECT 2433.105 4977.260 2433.385 4979.435 ;
        RECT 1988.105 4977.035 1988.420 4977.260 ;
        RECT 1221.000 4953.790 1221.140 4977.035 ;
        RECT 1479.060 4953.790 1479.200 4977.035 ;
        RECT 1988.280 4954.130 1988.420 4977.035 ;
        RECT 2433.100 4977.035 2433.385 4977.260 ;
        RECT 2690.105 4977.035 2690.385 4979.435 ;
        RECT 3199.105 4977.330 3199.385 4979.435 ;
        RECT 3199.000 4977.035 3199.385 4977.330 ;
        RECT 2433.100 4954.130 2433.240 4977.035 ;
        RECT 2690.240 4954.130 2690.380 4977.035 ;
        RECT 3199.000 4954.130 3199.140 4977.035 ;
        RECT 1987.300 4953.810 1987.560 4954.130 ;
        RECT 1988.220 4953.810 1988.480 4954.130 ;
        RECT 2433.040 4953.810 2433.300 4954.130 ;
        RECT 2690.180 4953.810 2690.440 4954.130 ;
        RECT 3198.940 4953.810 3199.200 4954.130 ;
        RECT 449.980 4953.470 450.240 4953.790 ;
        RECT 707.120 4953.470 707.380 4953.790 ;
        RECT 964.260 4953.470 964.520 4953.790 ;
        RECT 974.840 4953.470 975.100 4953.790 ;
        RECT 1220.940 4953.470 1221.200 4953.790 ;
        RECT 1479.000 4953.470 1479.260 4953.790 ;
        RECT 450.040 4950.810 450.180 4953.470 ;
        RECT 964.320 4952.430 964.460 4953.470 ;
        RECT 974.900 4952.430 975.040 4953.470 ;
        RECT 1479.060 4952.770 1479.200 4953.470 ;
        RECT 1987.360 4952.770 1987.500 4953.810 ;
        RECT 1479.000 4952.450 1479.260 4952.770 ;
        RECT 1987.300 4952.450 1987.560 4952.770 ;
        RECT 964.260 4952.110 964.520 4952.430 ;
        RECT 974.840 4952.110 975.100 4952.430 ;
        RECT 3199.000 4951.070 3199.140 4953.810 ;
        RECT 449.580 4950.730 450.180 4950.810 ;
        RECT 3198.940 4950.750 3199.200 4951.070 ;
        RECT 3368.220 4950.750 3368.480 4951.070 ;
        RECT 449.520 4950.670 450.180 4950.730 ;
        RECT 449.520 4950.410 449.780 4950.670 ;
        RECT 212.620 4950.070 212.880 4950.390 ;
        RECT 212.680 4842.610 212.820 4950.070 ;
        RECT 208.940 4842.290 209.200 4842.610 ;
        RECT 212.620 4842.290 212.880 4842.610 ;
        RECT 209.000 4840.385 209.140 4842.290 ;
        RECT 208.565 4840.105 210.965 4840.385 ;
        RECT 208.565 3991.105 210.965 3991.385 ;
        RECT 209.000 3988.870 209.140 3991.105 ;
        RECT 212.680 3988.870 212.820 4842.290 ;
        RECT 3368.280 4766.790 3368.420 4950.750 ;
        RECT 3377.035 4768.755 3379.435 4768.895 ;
        RECT 3377.020 4768.615 3379.435 4768.755 ;
        RECT 3377.020 4766.790 3377.160 4768.615 ;
        RECT 3368.220 4766.470 3368.480 4766.790 ;
        RECT 3376.960 4766.470 3377.220 4766.790 ;
        RECT 3368.280 4322.410 3368.420 4766.470 ;
        RECT 3377.035 4322.755 3379.435 4322.895 ;
        RECT 3377.020 4322.615 3379.435 4322.755 ;
        RECT 3377.020 4322.410 3377.160 4322.615 ;
        RECT 3368.220 4322.090 3368.480 4322.410 ;
        RECT 3376.960 4322.090 3377.220 4322.410 ;
        RECT 208.940 3988.550 209.200 3988.870 ;
        RECT 212.620 3988.550 212.880 3988.870 ;
        RECT 213.540 3988.550 213.800 3988.870 ;
        RECT 213.600 3836.890 213.740 3988.550 ;
        RECT 3368.280 3874.630 3368.420 4322.090 ;
        RECT 3377.035 3876.755 3379.435 3876.895 ;
        RECT 3377.020 3876.615 3379.435 3876.755 ;
        RECT 3377.020 3874.630 3377.160 3876.615 ;
        RECT 3367.300 3874.310 3367.560 3874.630 ;
        RECT 3368.220 3874.310 3368.480 3874.630 ;
        RECT 3376.960 3874.310 3377.220 3874.630 ;
        RECT 212.160 3836.570 212.420 3836.890 ;
        RECT 213.540 3836.570 213.800 3836.890 ;
        RECT 208.565 3775.105 210.965 3775.385 ;
        RECT 209.000 3772.630 209.140 3775.105 ;
        RECT 212.220 3772.630 212.360 3836.570 ;
        RECT 208.940 3772.310 209.200 3772.630 ;
        RECT 212.160 3772.310 212.420 3772.630 ;
        RECT 208.565 3559.105 210.965 3559.385 ;
        RECT 209.000 3556.730 209.140 3559.105 ;
        RECT 212.220 3556.730 212.360 3772.310 ;
        RECT 3367.360 3650.910 3367.500 3874.310 ;
        RECT 3377.035 3651.755 3379.435 3651.895 ;
        RECT 3377.020 3651.615 3379.435 3651.755 ;
        RECT 3377.020 3650.910 3377.160 3651.615 ;
        RECT 3367.300 3650.590 3367.560 3650.910 ;
        RECT 3376.960 3650.590 3377.220 3650.910 ;
        RECT 208.940 3556.410 209.200 3556.730 ;
        RECT 212.160 3556.410 212.420 3556.730 ;
        RECT 213.540 3556.410 213.800 3556.730 ;
        RECT 213.600 3392.250 213.740 3556.410 ;
        RECT 3367.360 3426.170 3367.500 3650.590 ;
        RECT 3377.035 3426.860 3379.435 3426.895 ;
        RECT 3377.020 3426.615 3379.435 3426.860 ;
        RECT 3377.020 3426.170 3377.160 3426.615 ;
        RECT 3367.300 3425.850 3367.560 3426.170 ;
        RECT 3376.960 3425.850 3377.220 3426.170 ;
        RECT 213.140 3392.110 213.740 3392.250 ;
        RECT 213.140 3360.970 213.280 3392.110 ;
        RECT 212.680 3360.830 213.280 3360.970 ;
        RECT 212.680 3345.590 212.820 3360.830 ;
        RECT 208.940 3345.270 209.200 3345.590 ;
        RECT 212.620 3345.270 212.880 3345.590 ;
        RECT 209.000 3343.385 209.140 3345.270 ;
        RECT 208.565 3343.105 210.965 3343.385 ;
        RECT 212.680 3160.290 212.820 3345.270 ;
        RECT 3367.360 3198.710 3367.500 3425.850 ;
        RECT 3377.035 3200.755 3379.435 3200.895 ;
        RECT 3377.020 3200.615 3379.435 3200.755 ;
        RECT 3377.020 3198.710 3377.160 3200.615 ;
        RECT 3367.300 3198.390 3367.560 3198.710 ;
        RECT 3369.600 3198.390 3369.860 3198.710 ;
        RECT 3376.960 3198.390 3377.220 3198.710 ;
        RECT 212.620 3159.970 212.880 3160.290 ;
        RECT 214.000 3159.290 214.260 3159.610 ;
        RECT 208.565 3127.105 210.965 3127.385 ;
        RECT 209.000 3124.930 209.140 3127.105 ;
        RECT 214.060 3124.930 214.200 3159.290 ;
        RECT 208.940 3124.610 209.200 3124.930 ;
        RECT 214.000 3124.610 214.260 3124.930 ;
        RECT 214.060 3064.410 214.200 3124.610 ;
        RECT 214.000 3064.090 214.260 3064.410 ;
        RECT 213.080 3063.750 213.340 3064.070 ;
        RECT 213.140 3063.390 213.280 3063.750 ;
        RECT 213.080 3063.070 213.340 3063.390 ;
        RECT 214.000 3063.070 214.260 3063.390 ;
        RECT 214.060 2913.450 214.200 3063.070 ;
        RECT 3369.660 2974.650 3369.800 3198.390 ;
        RECT 3377.035 2975.755 3379.435 2975.895 ;
        RECT 3377.020 2975.615 3379.435 2975.755 ;
        RECT 3377.020 2974.650 3377.160 2975.615 ;
        RECT 3368.220 2974.330 3368.480 2974.650 ;
        RECT 3369.600 2974.330 3369.860 2974.650 ;
        RECT 3376.960 2974.330 3377.220 2974.650 ;
        RECT 208.940 2913.130 209.200 2913.450 ;
        RECT 214.000 2913.130 214.260 2913.450 ;
        RECT 209.000 2911.385 209.140 2913.130 ;
        RECT 208.565 2911.105 210.965 2911.385 ;
        RECT 214.060 2870.610 214.200 2913.130 ;
        RECT 211.700 2870.290 211.960 2870.610 ;
        RECT 214.000 2870.290 214.260 2870.610 ;
        RECT 211.760 2702.730 211.900 2870.290 ;
        RECT 3368.280 2752.630 3368.420 2974.330 ;
        RECT 3368.220 2752.310 3368.480 2752.630 ;
        RECT 3376.960 2752.310 3377.220 2752.630 ;
        RECT 3377.020 2749.895 3377.160 2752.310 ;
        RECT 3377.020 2749.755 3379.435 2749.895 ;
        RECT 3377.035 2749.615 3379.435 2749.755 ;
        RECT 211.760 2702.590 212.820 2702.730 ;
        RECT 212.680 2697.550 212.820 2702.590 ;
        RECT 208.940 2697.230 209.200 2697.550 ;
        RECT 212.620 2697.230 212.880 2697.550 ;
        RECT 209.000 2695.385 209.140 2697.230 ;
        RECT 208.565 2695.105 210.965 2695.385 ;
        RECT 208.565 2057.105 210.965 2057.385 ;
        RECT 209.000 2056.310 209.140 2057.105 ;
        RECT 212.680 2056.310 212.820 2697.230 ;
        RECT 208.940 2055.990 209.200 2056.310 ;
        RECT 212.620 2055.990 212.880 2056.310 ;
        RECT 212.680 1959.490 212.820 2055.990 ;
        RECT 212.680 1959.350 213.280 1959.490 ;
        RECT 213.140 1931.870 213.280 1959.350 ;
        RECT 213.080 1931.550 213.340 1931.870 ;
        RECT 214.460 1931.550 214.720 1931.870 ;
        RECT 214.520 1843.470 214.660 1931.550 ;
        RECT 3377.035 1863.755 3379.435 1863.895 ;
        RECT 3377.020 1863.615 3379.435 1863.755 ;
        RECT 3377.020 1861.830 3377.160 1863.615 ;
        RECT 3368.680 1861.510 3368.940 1861.830 ;
        RECT 3376.960 1861.510 3377.220 1861.830 ;
        RECT 208.940 1843.150 209.200 1843.470 ;
        RECT 214.460 1843.150 214.720 1843.470 ;
        RECT 209.000 1841.385 209.140 1843.150 ;
        RECT 208.565 1841.105 210.965 1841.385 ;
        RECT 214.520 1838.620 214.660 1843.150 ;
        RECT 214.060 1838.480 214.660 1838.620 ;
        RECT 214.060 1711.290 214.200 1838.480 ;
        RECT 213.600 1711.150 214.200 1711.290 ;
        RECT 213.600 1627.570 213.740 1711.150 ;
        RECT 3368.740 1640.490 3368.880 1861.510 ;
        RECT 3368.680 1640.170 3368.940 1640.490 ;
        RECT 3376.960 1640.170 3377.220 1640.490 ;
        RECT 208.940 1627.250 209.200 1627.570 ;
        RECT 212.160 1627.250 212.420 1627.570 ;
        RECT 213.540 1627.250 213.800 1627.570 ;
        RECT 209.000 1625.385 209.140 1627.250 ;
        RECT 208.565 1625.105 210.965 1625.385 ;
        RECT 212.220 1614.650 212.360 1627.250 ;
        RECT 212.160 1614.330 212.420 1614.650 ;
        RECT 213.540 1613.990 213.800 1614.310 ;
        RECT 213.600 1571.130 213.740 1613.990 ;
        RECT 211.700 1570.810 211.960 1571.130 ;
        RECT 213.540 1570.810 213.800 1571.130 ;
        RECT 211.760 1418.515 211.900 1570.810 ;
        RECT 211.760 1418.375 212.820 1418.515 ;
        RECT 212.680 1411.670 212.820 1418.375 ;
        RECT 208.940 1411.350 209.200 1411.670 ;
        RECT 212.620 1411.350 212.880 1411.670 ;
        RECT 209.000 1409.385 209.140 1411.350 ;
        RECT 208.565 1409.105 210.965 1409.385 ;
        RECT 212.680 1380.130 212.820 1411.350 ;
        RECT 3368.740 1410.650 3368.880 1640.170 ;
        RECT 3377.020 1637.895 3377.160 1640.170 ;
        RECT 3377.020 1637.780 3379.435 1637.895 ;
        RECT 3377.035 1637.615 3379.435 1637.780 ;
        RECT 3377.035 1412.700 3379.435 1412.895 ;
        RECT 3377.020 1412.615 3379.435 1412.700 ;
        RECT 3377.020 1410.650 3377.160 1412.615 ;
        RECT 3368.680 1410.330 3368.940 1410.650 ;
        RECT 3376.960 1410.330 3377.220 1410.650 ;
        RECT 211.760 1379.990 212.820 1380.130 ;
        RECT 211.760 1228.070 211.900 1379.990 ;
        RECT 211.700 1227.750 211.960 1228.070 ;
        RECT 214.460 1227.750 214.720 1228.070 ;
        RECT 208.565 1193.105 210.965 1193.385 ;
        RECT 209.000 1190.670 209.140 1193.105 ;
        RECT 214.520 1190.670 214.660 1227.750 ;
        RECT 3368.740 1220.330 3368.880 1410.330 ;
        RECT 3368.740 1220.190 3369.800 1220.330 ;
        RECT 208.940 1190.350 209.200 1190.670 ;
        RECT 213.080 1190.350 213.340 1190.670 ;
        RECT 214.460 1190.350 214.720 1190.670 ;
        RECT 213.140 1164.490 213.280 1190.350 ;
        RECT 3369.660 1188.630 3369.800 1220.190 ;
        RECT 3369.600 1188.310 3369.860 1188.630 ;
        RECT 3376.960 1188.310 3377.220 1188.630 ;
        RECT 3369.660 1186.930 3369.800 1188.310 ;
        RECT 3377.020 1187.895 3377.160 1188.310 ;
        RECT 3377.020 1187.620 3379.435 1187.895 ;
        RECT 3377.035 1187.615 3379.435 1187.620 ;
        RECT 3369.600 1186.610 3369.860 1186.930 ;
        RECT 3370.520 1186.610 3370.780 1186.930 ;
        RECT 211.700 1164.170 211.960 1164.490 ;
        RECT 213.080 1164.170 213.340 1164.490 ;
        RECT 211.760 1042.090 211.900 1164.170 ;
        RECT 3370.580 1159.050 3370.720 1186.610 ;
        RECT 3370.520 1158.730 3370.780 1159.050 ;
        RECT 3371.440 1158.730 3371.700 1159.050 ;
        RECT 3371.500 1062.830 3371.640 1158.730 ;
        RECT 3370.060 1062.510 3370.320 1062.830 ;
        RECT 3371.440 1062.510 3371.700 1062.830 ;
        RECT 211.700 1041.770 211.960 1042.090 ;
        RECT 214.460 1041.770 214.720 1042.090 ;
        RECT 208.565 977.105 210.965 977.385 ;
        RECT 209.000 974.770 209.140 977.105 ;
        RECT 214.520 974.770 214.660 1041.770 ;
        RECT 3370.120 993.810 3370.260 1062.510 ;
        RECT 3370.060 993.490 3370.320 993.810 ;
        RECT 3376.040 993.490 3376.300 993.810 ;
        RECT 208.940 974.450 209.200 974.770 ;
        RECT 212.160 974.450 212.420 974.770 ;
        RECT 214.460 974.450 214.720 974.770 ;
        RECT 212.220 926.830 212.360 974.450 ;
        RECT 3376.100 960.830 3376.240 993.490 ;
        RECT 3377.035 961.860 3379.435 961.895 ;
        RECT 3377.020 961.615 3379.435 961.860 ;
        RECT 3377.020 960.830 3377.160 961.615 ;
        RECT 3373.740 960.510 3374.000 960.830 ;
        RECT 3376.040 960.510 3376.300 960.830 ;
        RECT 3376.960 960.510 3377.220 960.830 ;
        RECT 212.160 926.510 212.420 926.830 ;
        RECT 213.540 926.510 213.800 926.830 ;
        RECT 213.600 745.610 213.740 926.510 ;
        RECT 3373.800 869.710 3373.940 960.510 ;
        RECT 3369.140 869.390 3369.400 869.710 ;
        RECT 3373.740 869.390 3374.000 869.710 ;
        RECT 3369.200 773.005 3369.340 869.390 ;
        RECT 3368.210 772.635 3368.490 773.005 ;
        RECT 3369.130 772.635 3369.410 773.005 ;
        RECT 212.620 745.290 212.880 745.610 ;
        RECT 213.540 745.290 213.800 745.610 ;
        RECT 212.680 648.450 212.820 745.290 ;
        RECT 3368.280 735.750 3368.420 772.635 ;
        RECT 3377.035 736.780 3379.435 736.895 ;
        RECT 3377.020 736.615 3379.435 736.780 ;
        RECT 3377.020 735.750 3377.160 736.615 ;
        RECT 3368.220 735.430 3368.480 735.750 ;
        RECT 3375.120 735.430 3375.380 735.750 ;
        RECT 3376.960 735.430 3377.220 735.750 ;
        RECT 3375.180 703.450 3375.320 735.430 ;
        RECT 3370.060 703.130 3370.320 703.450 ;
        RECT 3375.120 703.130 3375.380 703.450 ;
        RECT 212.680 648.310 213.740 648.450 ;
        RECT 213.600 552.490 213.740 648.310 ;
        RECT 3370.120 580.030 3370.260 703.130 ;
        RECT 3369.140 579.710 3369.400 580.030 ;
        RECT 3370.060 579.710 3370.320 580.030 ;
        RECT 3369.200 579.350 3369.340 579.710 ;
        RECT 3369.140 579.030 3369.400 579.350 ;
        RECT 3375.120 579.030 3375.380 579.350 ;
        RECT 212.620 552.170 212.880 552.490 ;
        RECT 213.540 552.170 213.800 552.490 ;
        RECT 212.680 455.330 212.820 552.170 ;
        RECT 3375.180 511.690 3375.320 579.030 ;
        RECT 3368.220 511.370 3368.480 511.690 ;
        RECT 3375.120 511.370 3375.380 511.690 ;
        RECT 3376.960 511.370 3377.220 511.690 ;
        RECT 212.680 455.190 213.740 455.330 ;
        RECT 213.600 403.085 213.740 455.190 ;
        RECT 207.090 402.715 207.370 403.085 ;
        RECT 213.530 402.715 213.810 403.085 ;
        RECT 207.160 391.525 207.300 402.715 ;
        RECT 207.090 391.155 207.370 391.525 ;
        RECT 213.600 228.130 213.740 402.715 ;
        RECT 213.540 227.810 213.800 228.130 ;
        RECT 717.700 227.810 717.960 228.130 ;
        RECT 717.760 202.485 717.900 227.810 ;
        RECT 3368.280 227.790 3368.420 511.370 ;
        RECT 3377.020 510.895 3377.160 511.370 ;
        RECT 3377.020 510.755 3379.435 510.895 ;
        RECT 3377.035 510.615 3379.435 510.755 ;
        RECT 2581.620 227.470 2581.880 227.790 ;
        RECT 3368.220 227.470 3368.480 227.790 ;
        RECT 2033.760 223.390 2034.020 223.710 ;
        RECT 2125.300 223.390 2125.560 223.710 ;
        RECT 2220.980 223.390 2221.240 223.710 ;
        RECT 2033.820 222.690 2033.960 223.390 ;
        RECT 2125.360 223.030 2125.500 223.390 ;
        RECT 2125.300 222.710 2125.560 223.030 ;
        RECT 1772.020 222.370 1772.280 222.690 ;
        RECT 1802.840 222.370 1803.100 222.690 ;
        RECT 1998.340 222.370 1998.600 222.690 ;
        RECT 2033.760 222.370 2034.020 222.690 ;
        RECT 1772.080 221.670 1772.220 222.370 ;
        RECT 1802.900 221.670 1803.040 222.370 ;
        RECT 1998.400 221.670 1998.540 222.370 ;
        RECT 942.640 221.350 942.900 221.670 ;
        RECT 964.260 221.350 964.520 221.670 ;
        RECT 1007.500 221.350 1007.760 221.670 ;
        RECT 1485.440 221.350 1485.700 221.670 ;
        RECT 1497.860 221.350 1498.120 221.670 ;
        RECT 1528.680 221.350 1528.940 221.670 ;
        RECT 1759.600 221.350 1759.860 221.670 ;
        RECT 1772.020 221.350 1772.280 221.670 ;
        RECT 1802.840 221.350 1803.100 221.670 ;
        RECT 1998.340 221.350 1998.600 221.670 ;
        RECT 942.700 210.965 942.840 221.350 ;
        RECT 964.320 210.965 964.460 221.350 ;
        RECT 1007.560 210.965 1007.700 221.350 ;
        RECT 1485.500 210.965 1485.640 221.350 ;
        RECT 1497.920 210.965 1498.060 221.350 ;
        RECT 1528.740 210.965 1528.880 221.350 ;
        RECT 1759.660 210.965 1759.800 221.350 ;
        RECT 1772.080 210.965 1772.220 221.350 ;
        RECT 1802.900 210.965 1803.040 221.350 ;
        RECT 2033.820 210.965 2033.960 222.370 ;
        RECT 2221.040 222.090 2221.180 223.390 ;
        RECT 2415.090 223.195 2415.370 223.565 ;
        RECT 2510.310 223.195 2510.590 223.565 ;
        RECT 2415.100 223.050 2415.360 223.195 ;
        RECT 2307.460 222.710 2307.720 223.030 ;
        RECT 2345.640 222.770 2345.900 223.030 ;
        RECT 2346.100 222.770 2346.360 223.030 ;
        RECT 2345.640 222.710 2346.360 222.770 ;
        RECT 2221.440 222.370 2221.700 222.690 ;
        RECT 2221.500 222.090 2221.640 222.370 ;
        RECT 2221.040 221.950 2221.640 222.090 ;
        RECT 942.615 209.850 942.895 210.965 ;
        RECT 942.240 209.770 942.895 209.850 ;
        RECT 938.500 209.450 938.760 209.770 ;
        RECT 942.180 209.710 942.895 209.770 ;
        RECT 942.180 209.450 942.440 209.710 ;
        RECT 938.560 209.090 938.700 209.450 ;
        RECT 748.060 208.770 748.320 209.090 ;
        RECT 938.500 208.770 938.760 209.090 ;
        RECT 717.690 202.115 717.970 202.485 ;
        RECT 748.120 201.805 748.260 208.770 ;
        RECT 942.615 208.565 942.895 209.710 ;
        RECT 964.235 208.565 964.515 210.965 ;
        RECT 1007.475 208.565 1007.755 210.965 ;
        RECT 1485.500 209.030 1485.895 210.965 ;
        RECT 1497.920 209.030 1498.315 210.965 ;
        RECT 1528.740 209.030 1529.135 210.965 ;
        RECT 1485.615 208.565 1485.895 209.030 ;
        RECT 1498.035 208.565 1498.315 209.030 ;
        RECT 1528.855 208.565 1529.135 209.030 ;
        RECT 1759.615 208.565 1759.895 210.965 ;
        RECT 1772.035 208.565 1772.315 210.965 ;
        RECT 1802.855 208.565 1803.135 210.965 ;
        RECT 2033.615 209.100 2033.960 210.965 ;
        RECT 2307.520 210.965 2307.660 222.710 ;
        RECT 2345.700 222.630 2346.300 222.710 ;
        RECT 2510.380 222.090 2510.520 223.195 ;
        RECT 2581.680 222.690 2581.820 227.470 ;
        RECT 2511.240 222.370 2511.500 222.690 ;
        RECT 2581.620 222.370 2581.880 222.690 ;
        RECT 2511.300 222.090 2511.440 222.370 ;
        RECT 2510.380 221.950 2511.440 222.090 ;
        RECT 2581.680 210.965 2581.820 222.370 ;
        RECT 2033.615 208.565 2033.895 209.100 ;
        RECT 2307.520 209.030 2307.895 210.965 ;
        RECT 2307.615 208.565 2307.895 209.030 ;
        RECT 2581.615 208.565 2581.895 210.965 ;
        RECT 748.050 201.435 748.330 201.805 ;
      LAYER via2 ;
        RECT 3368.210 772.680 3368.490 772.960 ;
        RECT 3369.130 772.680 3369.410 772.960 ;
        RECT 207.090 402.760 207.370 403.040 ;
        RECT 213.530 402.760 213.810 403.040 ;
        RECT 207.090 391.200 207.370 391.480 ;
        RECT 2415.090 223.240 2415.370 223.520 ;
        RECT 2510.310 223.240 2510.590 223.520 ;
        RECT 717.690 202.160 717.970 202.440 ;
        RECT 748.050 201.480 748.330 201.760 ;
      LAYER met3 ;
        RECT 3368.185 772.970 3368.515 772.985 ;
        RECT 3369.105 772.970 3369.435 772.985 ;
        RECT 3368.185 772.670 3369.435 772.970 ;
        RECT 3368.185 772.655 3368.515 772.670 ;
        RECT 3369.105 772.655 3369.435 772.670 ;
        RECT 191.100 391.490 198.000 414.700 ;
        RECT 207.065 403.050 207.395 403.065 ;
        RECT 213.505 403.050 213.835 403.065 ;
        RECT 207.065 402.750 213.835 403.050 ;
        RECT 207.065 402.735 207.395 402.750 ;
        RECT 213.505 402.735 213.835 402.750 ;
        RECT 207.065 391.490 207.395 391.505 ;
        RECT 191.100 391.190 207.395 391.490 ;
        RECT 191.100 390.755 198.000 391.190 ;
        RECT 207.065 391.175 207.395 391.190 ;
        RECT 2415.065 223.530 2415.395 223.545 ;
        RECT 2510.285 223.530 2510.615 223.545 ;
        RECT 2415.065 223.230 2510.615 223.530 ;
        RECT 2415.065 223.215 2415.395 223.230 ;
        RECT 2510.285 223.215 2510.615 223.230 ;
        RECT 717.665 202.450 717.995 202.465 ;
        RECT 717.665 202.150 729.250 202.450 ;
        RECT 717.665 202.135 717.995 202.150 ;
        RECT 728.950 201.770 729.250 202.150 ;
        RECT 748.025 201.770 748.355 201.785 ;
        RECT 728.950 201.470 748.355 201.770 ;
        RECT 729.190 200.070 729.490 201.470 ;
        RECT 748.025 201.455 748.355 201.470 ;
        RECT 729.100 200.000 729.490 200.070 ;
        RECT 729.080 184.215 729.600 200.000 ;
        RECT 729.080 184.005 729.810 184.215 ;
        RECT 729.080 183.705 729.670 184.005 ;
        RECT 729.810 183.705 730.260 184.005 ;
        RECT 729.080 183.555 730.260 183.705 ;
        RECT 729.080 183.415 729.670 183.555 ;
    END
  END vccd
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3188.035 181.615 3385.255 185.065 ;
    END
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.880 ;
    END
  END vdda
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2919.035 181.615 3114.965 185.065 ;
    END
  END vdda
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3188.035 181.715 3385.255 184.965 ;
    END
  END vdda
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2919.035 181.715 3114.965 184.965 ;
    END
  END vdda
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3164.605 185.040 3188.505 200.000 ;
    END
  END vdda
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3114.710 185.040 3138.610 200.000 ;
    END
  END vdda
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.000 549.000 129.965 552.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 34.055 558.050 94.880 618.890 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 175.565 413.730 180.215 552.270 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.000 624.730 129.965 627.000 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 175.565 624.730 180.215 909.270 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 175.665 413.730 180.115 552.270 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 105.015 549.000 129.965 552.270 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 175.665 624.730 180.115 909.270 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 105.015 624.730 129.965 627.000 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 211.210 607.480 211.530 607.540 ;
        RECT 223.630 607.480 223.950 607.540 ;
        RECT 211.210 607.340 223.950 607.480 ;
        RECT 211.210 607.280 211.530 607.340 ;
        RECT 223.630 607.280 223.950 607.340 ;
        RECT 214.890 579.600 215.210 579.660 ;
        RECT 223.630 579.600 223.950 579.660 ;
        RECT 214.890 579.460 223.950 579.600 ;
        RECT 214.890 579.400 215.210 579.460 ;
        RECT 223.630 579.400 223.950 579.460 ;
        RECT 223.170 414.160 223.490 414.420 ;
        RECT 223.260 414.020 223.400 414.160 ;
        RECT 224.090 414.020 224.410 414.080 ;
        RECT 223.260 413.880 224.410 414.020 ;
        RECT 224.090 413.820 224.410 413.880 ;
        RECT 224.550 227.700 224.870 227.760 ;
        RECT 979.870 227.700 980.190 227.760 ;
        RECT 224.550 227.560 980.190 227.700 ;
        RECT 224.550 227.500 224.870 227.560 ;
        RECT 979.870 227.500 980.190 227.560 ;
        RECT 2028.210 223.960 2028.530 224.020 ;
        RECT 2056.270 223.960 2056.590 224.020 ;
        RECT 2028.210 223.820 2056.590 223.960 ;
        RECT 2028.210 223.760 2028.530 223.820 ;
        RECT 2056.270 223.760 2056.590 223.820 ;
        RECT 1796.830 223.620 1797.150 223.680 ;
        RECT 1711.360 223.480 1797.150 223.620 ;
        RECT 979.870 222.260 980.190 222.320 ;
        RECT 1522.670 222.260 1522.990 222.320 ;
        RECT 1711.360 222.260 1711.500 223.480 ;
        RECT 1796.830 223.420 1797.150 223.480 ;
        RECT 1803.270 222.600 1803.590 222.660 ;
        RECT 1932.070 222.600 1932.390 222.660 ;
        RECT 1803.270 222.460 1932.390 222.600 ;
        RECT 1803.270 222.400 1803.590 222.460 ;
        RECT 1932.070 222.400 1932.390 222.460 ;
        RECT 2056.270 222.600 2056.590 222.660 ;
        RECT 2056.270 222.460 2071.220 222.600 ;
        RECT 2056.270 222.400 2056.590 222.460 ;
        RECT 2071.080 222.320 2071.220 222.460 ;
        RECT 979.870 222.120 1711.500 222.260 ;
        RECT 2070.990 222.260 2071.310 222.320 ;
        RECT 2099.050 222.260 2099.370 222.320 ;
        RECT 2070.990 222.120 2099.370 222.260 ;
        RECT 979.870 222.060 980.190 222.120 ;
        RECT 1522.670 222.060 1522.990 222.120 ;
        RECT 2070.990 222.060 2071.310 222.120 ;
        RECT 2099.050 222.060 2099.370 222.120 ;
        RECT 1796.830 221.920 1797.150 221.980 ;
        RECT 1803.270 221.920 1803.590 221.980 ;
        RECT 1796.830 221.780 1803.590 221.920 ;
        RECT 1796.830 221.720 1797.150 221.780 ;
        RECT 1803.270 221.720 1803.590 221.780 ;
        RECT 2099.050 221.240 2099.370 221.300 ;
        RECT 2344.690 221.240 2345.010 221.300 ;
        RECT 2618.850 221.240 2619.170 221.300 ;
        RECT 2099.050 221.100 2619.170 221.240 ;
        RECT 2099.050 221.040 2099.370 221.100 ;
        RECT 2344.690 221.040 2345.010 221.100 ;
        RECT 2618.850 221.040 2619.170 221.100 ;
      LAYER via ;
        RECT 211.240 607.280 211.500 607.540 ;
        RECT 223.660 607.280 223.920 607.540 ;
        RECT 214.920 579.400 215.180 579.660 ;
        RECT 223.660 579.400 223.920 579.660 ;
        RECT 223.200 414.160 223.460 414.420 ;
        RECT 224.120 413.820 224.380 414.080 ;
        RECT 224.580 227.500 224.840 227.760 ;
        RECT 979.900 227.500 980.160 227.760 ;
        RECT 2028.240 223.760 2028.500 224.020 ;
        RECT 2056.300 223.760 2056.560 224.020 ;
        RECT 979.900 222.060 980.160 222.320 ;
        RECT 1522.700 222.060 1522.960 222.320 ;
        RECT 1796.860 223.420 1797.120 223.680 ;
        RECT 1803.300 222.400 1803.560 222.660 ;
        RECT 1932.100 222.400 1932.360 222.660 ;
        RECT 2056.300 222.400 2056.560 222.660 ;
        RECT 2071.020 222.060 2071.280 222.320 ;
        RECT 2099.080 222.060 2099.340 222.320 ;
        RECT 1796.860 221.720 1797.120 221.980 ;
        RECT 1803.300 221.720 1803.560 221.980 ;
        RECT 2099.080 221.040 2099.340 221.300 ;
        RECT 2344.720 221.040 2344.980 221.300 ;
        RECT 2618.880 221.040 2619.140 221.300 ;
      LAYER met2 ;
        RECT 211.230 4350.115 211.510 4350.485 ;
        RECT 211.300 607.570 211.440 4350.115 ;
        RECT 211.240 607.250 211.500 607.570 ;
        RECT 223.660 607.250 223.920 607.570 ;
        RECT 223.720 579.690 223.860 607.250 ;
        RECT 214.920 579.370 215.180 579.690 ;
        RECT 223.660 579.370 223.920 579.690 ;
        RECT 214.980 552.005 215.120 579.370 ;
        RECT 214.910 551.635 215.190 552.005 ;
        RECT 214.980 483.325 215.120 551.635 ;
        RECT 214.910 482.955 215.190 483.325 ;
        RECT 223.190 482.955 223.470 483.325 ;
        RECT 223.260 414.450 223.400 482.955 ;
        RECT 223.200 414.130 223.460 414.450 ;
        RECT 224.120 413.790 224.380 414.110 ;
        RECT 224.180 413.170 224.320 413.790 ;
        RECT 224.180 413.030 224.780 413.170 ;
        RECT 224.640 227.790 224.780 413.030 ;
        RECT 224.580 227.470 224.840 227.790 ;
        RECT 979.900 227.470 980.160 227.790 ;
        RECT 979.960 222.350 980.100 227.470 ;
        RECT 2028.240 223.730 2028.500 224.050 ;
        RECT 2056.300 223.730 2056.560 224.050 ;
        RECT 1796.860 223.390 1797.120 223.710 ;
        RECT 979.900 222.030 980.160 222.350 ;
        RECT 1522.700 222.030 1522.960 222.350 ;
        RECT 979.960 210.965 980.100 222.030 ;
        RECT 1522.760 210.965 1522.900 222.030 ;
        RECT 1796.920 222.010 1797.060 223.390 ;
        RECT 2028.300 222.885 2028.440 223.730 ;
        RECT 1803.300 222.370 1803.560 222.690 ;
        RECT 1932.090 222.515 1932.370 222.885 ;
        RECT 2028.230 222.515 2028.510 222.885 ;
        RECT 2056.360 222.690 2056.500 223.730 ;
        RECT 1932.100 222.370 1932.360 222.515 ;
        RECT 2056.300 222.370 2056.560 222.690 ;
        RECT 1803.360 222.010 1803.500 222.370 ;
        RECT 2071.020 222.030 2071.280 222.350 ;
        RECT 2099.080 222.030 2099.340 222.350 ;
        RECT 1796.860 221.690 1797.120 222.010 ;
        RECT 1803.300 221.690 1803.560 222.010 ;
        RECT 1796.920 210.965 1797.060 221.690 ;
        RECT 2071.080 210.965 2071.220 222.030 ;
        RECT 2099.140 221.330 2099.280 222.030 ;
        RECT 2099.080 221.010 2099.340 221.330 ;
        RECT 2344.720 221.010 2344.980 221.330 ;
        RECT 2618.880 221.010 2619.140 221.330 ;
        RECT 979.875 208.565 980.155 210.965 ;
        RECT 1522.760 209.030 1523.155 210.965 ;
        RECT 1522.875 208.565 1523.155 209.030 ;
        RECT 1796.875 208.565 1797.155 210.965 ;
        RECT 2070.875 209.100 2071.220 210.965 ;
        RECT 2344.780 210.965 2344.920 221.010 ;
        RECT 2618.940 210.965 2619.080 221.010 ;
        RECT 2070.875 208.565 2071.155 209.100 ;
        RECT 2344.780 209.030 2345.155 210.965 ;
        RECT 2344.875 208.565 2345.155 209.030 ;
        RECT 2618.875 208.565 2619.155 210.965 ;
      LAYER via2 ;
        RECT 211.230 4350.160 211.510 4350.440 ;
        RECT 214.910 551.680 215.190 551.960 ;
        RECT 214.910 483.000 215.190 483.280 ;
        RECT 223.190 483.000 223.470 483.280 ;
        RECT 1932.090 222.560 1932.370 222.840 ;
        RECT 2028.230 222.560 2028.510 222.840 ;
      LAYER met3 ;
        RECT 180.200 4350.450 200.000 4373.395 ;
        RECT 211.205 4350.450 211.535 4350.465 ;
        RECT 180.200 4350.150 211.535 4350.450 ;
        RECT 180.200 4349.495 200.000 4350.150 ;
        RECT 211.205 4350.135 211.535 4350.150 ;
        RECT 180.200 551.970 200.000 575.395 ;
        RECT 214.885 551.970 215.215 551.985 ;
        RECT 180.200 551.670 215.215 551.970 ;
        RECT 180.200 551.495 200.000 551.670 ;
        RECT 214.885 551.655 215.215 551.670 ;
        RECT 214.885 483.290 215.215 483.305 ;
        RECT 223.165 483.290 223.495 483.305 ;
        RECT 214.885 482.990 223.495 483.290 ;
        RECT 214.885 482.975 215.215 482.990 ;
        RECT 223.165 482.975 223.495 482.990 ;
        RECT 1932.065 222.850 1932.395 222.865 ;
        RECT 2028.205 222.850 2028.535 222.865 ;
        RECT 1932.065 222.550 2028.535 222.850 ;
        RECT 1932.065 222.535 1932.395 222.550 ;
        RECT 2028.205 222.535 2028.535 222.550 ;
    END
  END vddio
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 180.200 601.390 200.000 625.290 ;
    END
  END vddio
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 159.815 664.270 163.265 ;
    END
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.880 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 143.265 964.910 143.595 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 147.175 469.000 148.355 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 151.935 964.910 152.265 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 198.665 159.815 395.270 163.265 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 180.425 151.935 395.270 152.265 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 176.825 143.265 395.270 143.595 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 394.000 147.175 395.270 148.355 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 469.000 163.160 663.000 163.165 ;
        RECT 467.730 159.915 664.270 163.160 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 467.730 143.265 664.270 152.265 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 198.665 163.160 394.000 163.165 ;
        RECT 198.665 159.915 395.270 163.160 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 176.845 143.265 395.270 152.265 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 394.710 163.240 418.610 200.000 ;
    END
  END vssa
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 994.590 209.680 994.910 209.740 ;
        RECT 1537.390 209.680 1537.710 209.740 ;
        RECT 994.590 209.540 1537.710 209.680 ;
        RECT 994.590 209.480 994.910 209.540 ;
        RECT 994.130 209.000 994.450 209.060 ;
        RECT 993.760 208.860 994.450 209.000 ;
        RECT 841.410 208.660 841.730 208.720 ;
        RECT 800.100 208.520 841.730 208.660 ;
        RECT 800.100 208.320 800.240 208.520 ;
        RECT 841.410 208.460 841.730 208.520 ;
        RECT 772.500 208.180 800.240 208.320 ;
        RECT 468.810 207.980 469.130 208.040 ;
        RECT 607.730 207.980 608.050 208.040 ;
        RECT 704.330 207.980 704.650 208.040 ;
        RECT 772.500 207.980 772.640 208.180 ;
        RECT 468.810 207.840 510.900 207.980 ;
        RECT 468.810 207.780 469.130 207.840 ;
        RECT 510.760 207.640 510.900 207.840 ;
        RECT 607.730 207.840 676.500 207.980 ;
        RECT 607.730 207.780 608.050 207.840 ;
        RECT 606.350 207.640 606.670 207.700 ;
        RECT 510.760 207.500 606.670 207.640 ;
        RECT 676.360 207.640 676.500 207.840 ;
        RECT 704.330 207.840 772.640 207.980 ;
        RECT 704.330 207.780 704.650 207.840 ;
        RECT 703.410 207.640 703.730 207.700 ;
        RECT 676.360 207.500 703.730 207.640 ;
        RECT 606.350 207.440 606.670 207.500 ;
        RECT 703.410 207.440 703.730 207.500 ;
        RECT 841.410 207.640 841.730 207.700 ;
        RECT 993.760 207.640 993.900 208.860 ;
        RECT 994.130 208.800 994.450 208.860 ;
        RECT 1537.020 208.660 1537.160 209.540 ;
        RECT 1537.390 209.480 1537.710 209.540 ;
        RECT 1812.470 209.680 1812.790 209.740 ;
        RECT 1835.470 209.680 1835.790 209.740 ;
        RECT 1812.470 209.540 1835.790 209.680 ;
        RECT 1812.470 209.480 1812.790 209.540 ;
        RECT 1835.470 209.480 1835.790 209.540 ;
        RECT 2085.250 209.000 2085.570 209.060 ;
        RECT 2359.410 209.000 2359.730 209.060 ;
        RECT 2085.250 208.860 2086.400 209.000 ;
        RECT 2085.250 208.800 2085.570 208.860 ;
        RECT 1537.020 208.520 1545.900 208.660 ;
        RECT 1545.760 208.320 1545.900 208.520 ;
        RECT 1572.810 208.320 1573.130 208.380 ;
        RECT 1545.760 208.180 1573.130 208.320 ;
        RECT 1572.810 208.120 1573.130 208.180 ;
        RECT 1573.270 208.320 1573.590 208.380 ;
        RECT 1931.610 208.320 1931.930 208.380 ;
        RECT 2086.260 208.320 2086.400 208.860 ;
        RECT 2359.410 208.860 2360.560 209.000 ;
        RECT 2359.410 208.800 2359.730 208.860 ;
        RECT 2360.420 208.320 2360.560 208.860 ;
        RECT 2633.570 208.800 2633.890 209.060 ;
        RECT 1573.270 208.180 1642.040 208.320 ;
        RECT 1573.270 208.120 1573.590 208.180 ;
        RECT 1641.900 207.980 1642.040 208.180 ;
        RECT 1931.610 208.180 1959.440 208.320 ;
        RECT 1931.610 208.120 1931.930 208.180 ;
        RECT 1748.070 207.980 1748.390 208.040 ;
        RECT 1641.900 207.840 1669.640 207.980 ;
        RECT 841.410 207.500 993.900 207.640 ;
        RECT 1669.500 207.640 1669.640 207.840 ;
        RECT 1669.960 207.840 1748.390 207.980 ;
        RECT 1669.960 207.640 1670.100 207.840 ;
        RECT 1748.070 207.780 1748.390 207.840 ;
        RECT 1669.500 207.500 1670.100 207.640 ;
        RECT 841.410 207.440 841.730 207.500 ;
        RECT 1959.300 207.300 1959.440 208.180 ;
        RECT 2086.260 208.180 2152.640 208.320 ;
        RECT 2086.260 207.300 2086.400 208.180 ;
        RECT 2152.500 207.640 2152.640 208.180 ;
        RECT 2360.420 208.180 2442.440 208.320 ;
        RECT 2360.420 207.640 2360.560 208.180 ;
        RECT 2442.300 207.980 2442.440 208.180 ;
        RECT 2539.270 207.980 2539.590 208.040 ;
        RECT 2442.300 207.840 2511.900 207.980 ;
        RECT 2152.500 207.500 2360.560 207.640 ;
        RECT 2511.760 207.640 2511.900 207.840 ;
        RECT 2539.270 207.840 2608.040 207.980 ;
        RECT 2539.270 207.780 2539.590 207.840 ;
        RECT 2538.810 207.640 2539.130 207.700 ;
        RECT 2511.760 207.500 2539.130 207.640 ;
        RECT 2607.900 207.640 2608.040 207.840 ;
        RECT 2633.660 207.640 2633.800 208.800 ;
        RECT 2607.900 207.500 2633.800 207.640 ;
        RECT 2538.810 207.440 2539.130 207.500 ;
        RECT 1959.300 207.160 2086.400 207.300 ;
      LAYER via ;
        RECT 994.620 209.480 994.880 209.740 ;
        RECT 841.440 208.460 841.700 208.720 ;
        RECT 468.840 207.780 469.100 208.040 ;
        RECT 607.760 207.780 608.020 208.040 ;
        RECT 606.380 207.440 606.640 207.700 ;
        RECT 704.360 207.780 704.620 208.040 ;
        RECT 703.440 207.440 703.700 207.700 ;
        RECT 841.440 207.440 841.700 207.700 ;
        RECT 994.160 208.800 994.420 209.060 ;
        RECT 1537.420 209.480 1537.680 209.740 ;
        RECT 1812.500 209.480 1812.760 209.740 ;
        RECT 1835.500 209.480 1835.760 209.740 ;
        RECT 2085.280 208.800 2085.540 209.060 ;
        RECT 1572.840 208.120 1573.100 208.380 ;
        RECT 1573.300 208.120 1573.560 208.380 ;
        RECT 1931.640 208.120 1931.900 208.380 ;
        RECT 2359.440 208.800 2359.700 209.060 ;
        RECT 2633.600 208.800 2633.860 209.060 ;
        RECT 1748.100 207.780 1748.360 208.040 ;
        RECT 2539.300 207.780 2539.560 208.040 ;
        RECT 2538.840 207.440 2539.100 207.700 ;
      LAYER met2 ;
        RECT 994.620 209.450 994.880 209.770 ;
        RECT 994.680 209.170 994.820 209.450 ;
        RECT 995.055 209.170 995.335 210.965 ;
        RECT 1537.420 209.450 1537.680 209.770 ;
        RECT 994.220 209.090 995.335 209.170 ;
        RECT 994.160 209.030 995.335 209.090 ;
        RECT 1537.480 209.170 1537.620 209.450 ;
        RECT 1538.055 209.170 1538.335 210.965 ;
        RECT 1812.055 209.680 1812.335 210.965 ;
        RECT 1812.500 209.680 1812.760 209.770 ;
        RECT 1812.055 209.540 1812.760 209.680 ;
        RECT 1835.490 209.595 1835.770 209.965 ;
        RECT 1930.710 209.595 1930.990 209.965 ;
        RECT 1812.055 209.285 1812.335 209.540 ;
        RECT 1812.500 209.450 1812.760 209.540 ;
        RECT 1835.500 209.450 1835.760 209.595 ;
        RECT 1537.480 209.030 1538.335 209.170 ;
        RECT 994.160 208.770 994.420 209.030 ;
        RECT 841.440 208.430 841.700 208.750 ;
        RECT 995.055 208.565 995.335 209.030 ;
        RECT 1538.055 208.565 1538.335 209.030 ;
        RECT 1748.090 208.915 1748.370 209.285 ;
        RECT 1812.030 208.915 1812.335 209.285 ;
        RECT 468.840 207.750 469.100 208.070 ;
        RECT 607.760 207.810 608.020 208.070 ;
        RECT 704.360 207.810 704.620 208.070 ;
        RECT 606.440 207.750 608.020 207.810 ;
        RECT 703.500 207.750 704.620 207.810 ;
        RECT 468.900 201.125 469.040 207.750 ;
        RECT 606.440 207.730 607.960 207.750 ;
        RECT 703.500 207.730 704.560 207.750 ;
        RECT 841.500 207.730 841.640 208.430 ;
        RECT 1572.900 208.410 1573.500 208.490 ;
        RECT 1572.840 208.350 1573.560 208.410 ;
        RECT 1572.840 208.090 1573.100 208.350 ;
        RECT 1573.300 208.090 1573.560 208.350 ;
        RECT 1748.160 208.070 1748.300 208.915 ;
        RECT 1812.055 208.565 1812.335 208.915 ;
        RECT 1748.100 207.750 1748.360 208.070 ;
        RECT 1930.780 207.810 1930.920 209.595 ;
        RECT 2086.055 209.170 2086.335 210.965 ;
        RECT 2360.055 209.170 2360.335 210.965 ;
        RECT 2634.055 209.170 2634.335 210.965 ;
        RECT 2085.340 209.090 2086.335 209.170 ;
        RECT 2359.500 209.090 2360.335 209.170 ;
        RECT 2633.660 209.090 2634.335 209.170 ;
        RECT 2085.280 209.030 2086.335 209.090 ;
        RECT 2085.280 208.770 2085.540 209.030 ;
        RECT 2086.055 208.565 2086.335 209.030 ;
        RECT 2359.440 209.030 2360.335 209.090 ;
        RECT 2359.440 208.770 2359.700 209.030 ;
        RECT 2360.055 208.565 2360.335 209.030 ;
        RECT 2633.600 209.030 2634.335 209.090 ;
        RECT 2633.600 208.770 2633.860 209.030 ;
        RECT 2634.055 208.565 2634.335 209.030 ;
        RECT 1931.640 208.090 1931.900 208.410 ;
        RECT 1931.700 207.810 1931.840 208.090 ;
        RECT 2539.300 207.810 2539.560 208.070 ;
        RECT 606.380 207.670 607.960 207.730 ;
        RECT 703.440 207.670 704.560 207.730 ;
        RECT 606.380 207.410 606.640 207.670 ;
        RECT 703.440 207.410 703.700 207.670 ;
        RECT 841.440 207.410 841.700 207.730 ;
        RECT 1930.780 207.670 1931.840 207.810 ;
        RECT 2538.900 207.750 2539.560 207.810 ;
        RECT 2538.900 207.730 2539.500 207.750 ;
        RECT 2538.840 207.670 2539.500 207.730 ;
        RECT 2538.840 207.410 2539.100 207.670 ;
        RECT 468.830 200.755 469.110 201.125 ;
      LAYER via2 ;
        RECT 1835.490 209.640 1835.770 209.920 ;
        RECT 1930.710 209.640 1930.990 209.920 ;
        RECT 1748.090 208.960 1748.370 209.240 ;
        RECT 1812.030 208.960 1812.310 209.240 ;
        RECT 468.830 200.800 469.110 201.080 ;
      LAYER met3 ;
        RECT 1835.465 209.930 1835.795 209.945 ;
        RECT 1930.685 209.930 1931.015 209.945 ;
        RECT 1835.465 209.630 1931.015 209.930 ;
        RECT 1835.465 209.615 1835.795 209.630 ;
        RECT 1930.685 209.615 1931.015 209.630 ;
        RECT 1748.065 209.250 1748.395 209.265 ;
        RECT 1812.005 209.250 1812.335 209.265 ;
        RECT 1748.065 208.950 1812.335 209.250 ;
        RECT 1748.065 208.935 1748.395 208.950 ;
        RECT 1812.005 208.935 1812.335 208.950 ;
        RECT 468.805 201.090 469.135 201.105 ;
        RECT 455.710 200.790 469.135 201.090 ;
        RECT 455.710 200.000 456.010 200.790 ;
        RECT 468.805 200.775 469.135 200.790 ;
        RECT 444.605 167.485 468.505 200.000 ;
    END
  END vssa
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1279.730 153.765 1476.270 158.415 ;
    END
    PORT
      LAYER met5 ;
        RECT 1216.330 30.835 1270.730 98.100 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1010.730 153.765 1207.270 158.415 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1279.730 153.865 1476.270 158.315 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1010.730 153.865 1207.270 158.315 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1256.500 158.400 1280.500 198.000 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1004.250 221.920 1004.570 221.980 ;
        RECT 1206.650 221.920 1206.970 221.980 ;
        RECT 1255.410 221.920 1255.730 221.980 ;
        RECT 1004.250 221.780 1255.730 221.920 ;
        RECT 1004.250 221.720 1004.570 221.780 ;
        RECT 1206.650 221.720 1206.970 221.780 ;
        RECT 1255.410 221.720 1255.730 221.780 ;
        RECT 1531.870 221.920 1532.190 221.980 ;
        RECT 1547.050 221.920 1547.370 221.980 ;
        RECT 1762.790 221.920 1763.110 221.980 ;
        RECT 1777.050 221.920 1777.370 221.980 ;
        RECT 1531.870 221.780 1777.370 221.920 ;
        RECT 1531.870 221.720 1532.190 221.780 ;
        RECT 1547.050 221.720 1547.370 221.780 ;
        RECT 1762.790 221.720 1763.110 221.780 ;
        RECT 1777.050 221.720 1777.370 221.780 ;
        RECT 1821.210 221.920 1821.530 221.980 ;
        RECT 2036.950 221.920 2037.270 221.980 ;
        RECT 2052.130 221.920 2052.450 221.980 ;
        RECT 1821.210 221.780 2052.450 221.920 ;
        RECT 1821.210 221.720 1821.530 221.780 ;
        RECT 2036.950 221.720 2037.270 221.780 ;
        RECT 2052.130 221.720 2052.450 221.780 ;
        RECT 2095.370 221.920 2095.690 221.980 ;
        RECT 2310.650 221.920 2310.970 221.980 ;
        RECT 2325.830 221.920 2326.150 221.980 ;
        RECT 2095.370 221.780 2326.150 221.920 ;
        RECT 2095.370 221.720 2095.690 221.780 ;
        RECT 2310.650 221.720 2310.970 221.780 ;
        RECT 2325.830 221.720 2326.150 221.780 ;
        RECT 2369.070 221.920 2369.390 221.980 ;
        RECT 2584.810 221.920 2585.130 221.980 ;
        RECT 2599.990 221.920 2600.310 221.980 ;
        RECT 2369.070 221.780 2600.310 221.920 ;
        RECT 2369.070 221.720 2369.390 221.780 ;
        RECT 2584.810 221.720 2585.130 221.780 ;
        RECT 2599.990 221.720 2600.310 221.780 ;
        RECT 1777.970 221.240 1778.290 221.300 ;
        RECT 1799.590 221.240 1799.910 221.300 ;
        RECT 1777.970 221.100 1799.910 221.240 ;
        RECT 1777.970 221.040 1778.290 221.100 ;
        RECT 1799.590 221.040 1799.910 221.100 ;
        RECT 1255.410 210.360 1255.730 210.420 ;
        RECT 1276.110 210.360 1276.430 210.420 ;
        RECT 1255.410 210.220 1276.430 210.360 ;
        RECT 1255.410 210.160 1255.730 210.220 ;
        RECT 1276.110 210.160 1276.430 210.220 ;
        RECT 992.290 209.340 992.610 209.400 ;
        RECT 1000.570 209.340 1000.890 209.400 ;
        RECT 992.290 209.200 1000.890 209.340 ;
        RECT 992.290 209.140 992.610 209.200 ;
        RECT 1000.570 209.140 1000.890 209.200 ;
        RECT 1276.110 209.340 1276.430 209.400 ;
        RECT 1488.170 209.340 1488.490 209.400 ;
        RECT 1503.350 209.340 1503.670 209.400 ;
        RECT 1276.110 209.200 1503.670 209.340 ;
        RECT 1276.110 209.140 1276.430 209.200 ;
        RECT 1488.170 209.140 1488.490 209.200 ;
        RECT 1503.350 209.140 1503.670 209.200 ;
        RECT 1800.050 209.340 1800.370 209.400 ;
        RECT 1805.570 209.340 1805.890 209.400 ;
        RECT 1817.530 209.340 1817.850 209.400 ;
        RECT 1800.050 209.200 1817.850 209.340 ;
        RECT 1800.050 209.140 1800.370 209.200 ;
        RECT 1805.570 209.140 1805.890 209.200 ;
        RECT 1817.530 209.140 1817.850 209.200 ;
        RECT 2052.590 209.340 2052.910 209.400 ;
        RECT 2059.030 209.340 2059.350 209.400 ;
        RECT 2074.210 209.340 2074.530 209.400 ;
        RECT 2080.650 209.340 2080.970 209.400 ;
        RECT 2092.610 209.340 2092.930 209.400 ;
        RECT 2354.810 209.340 2355.130 209.400 ;
        RECT 2365.390 209.340 2365.710 209.400 ;
        RECT 2052.590 209.200 2092.930 209.340 ;
        RECT 2052.590 209.140 2052.910 209.200 ;
        RECT 2059.030 209.140 2059.350 209.200 ;
        RECT 2074.210 209.140 2074.530 209.200 ;
        RECT 2080.650 209.140 2080.970 209.200 ;
        RECT 2092.610 209.140 2092.930 209.200 ;
        RECT 2350.760 209.200 2365.710 209.340 ;
        RECT 946.290 209.000 946.610 209.060 ;
        RECT 955.490 209.000 955.810 209.060 ;
        RECT 961.470 209.000 961.790 209.060 ;
        RECT 967.910 209.000 968.230 209.060 ;
        RECT 982.170 209.000 982.490 209.060 ;
        RECT 946.290 208.860 982.490 209.000 ;
        RECT 946.290 208.800 946.610 208.860 ;
        RECT 955.490 208.800 955.810 208.860 ;
        RECT 961.470 208.800 961.790 208.860 ;
        RECT 967.910 208.800 968.230 208.860 ;
        RECT 982.170 208.800 982.490 208.860 ;
        RECT 1511.170 209.000 1511.490 209.060 ;
        RECT 1524.970 209.000 1525.290 209.060 ;
        RECT 1531.410 209.000 1531.730 209.060 ;
        RECT 1511.170 208.860 1531.730 209.000 ;
        RECT 1511.170 208.800 1511.490 208.860 ;
        RECT 1524.970 208.800 1525.290 208.860 ;
        RECT 1531.410 208.800 1531.730 208.860 ;
        RECT 2326.750 209.000 2327.070 209.060 ;
        RECT 2331.810 209.000 2332.130 209.060 ;
        RECT 2348.370 209.000 2348.690 209.060 ;
        RECT 2350.760 209.000 2350.900 209.200 ;
        RECT 2354.810 209.140 2355.130 209.200 ;
        RECT 2365.390 209.140 2365.710 209.200 ;
        RECT 2600.450 209.340 2600.770 209.400 ;
        RECT 2605.970 209.340 2606.290 209.400 ;
        RECT 2621.150 209.340 2621.470 209.400 ;
        RECT 2627.590 209.340 2627.910 209.400 ;
        RECT 2639.550 209.340 2639.870 209.400 ;
        RECT 2600.450 209.200 2639.870 209.340 ;
        RECT 2600.450 209.140 2600.770 209.200 ;
        RECT 2605.970 209.140 2606.290 209.200 ;
        RECT 2621.150 209.140 2621.470 209.200 ;
        RECT 2627.590 209.140 2627.910 209.200 ;
        RECT 2639.550 209.140 2639.870 209.200 ;
        RECT 2326.750 208.860 2350.900 209.000 ;
        RECT 2326.750 208.800 2327.070 208.860 ;
        RECT 2331.810 208.800 2332.130 208.860 ;
        RECT 2348.370 208.800 2348.690 208.860 ;
      LAYER via ;
        RECT 1004.280 221.720 1004.540 221.980 ;
        RECT 1206.680 221.720 1206.940 221.980 ;
        RECT 1255.440 221.720 1255.700 221.980 ;
        RECT 1531.900 221.720 1532.160 221.980 ;
        RECT 1547.080 221.720 1547.340 221.980 ;
        RECT 1762.820 221.720 1763.080 221.980 ;
        RECT 1777.080 221.720 1777.340 221.980 ;
        RECT 1821.240 221.720 1821.500 221.980 ;
        RECT 2036.980 221.720 2037.240 221.980 ;
        RECT 2052.160 221.720 2052.420 221.980 ;
        RECT 2095.400 221.720 2095.660 221.980 ;
        RECT 2310.680 221.720 2310.940 221.980 ;
        RECT 2325.860 221.720 2326.120 221.980 ;
        RECT 2369.100 221.720 2369.360 221.980 ;
        RECT 2584.840 221.720 2585.100 221.980 ;
        RECT 2600.020 221.720 2600.280 221.980 ;
        RECT 1778.000 221.040 1778.260 221.300 ;
        RECT 1799.620 221.040 1799.880 221.300 ;
        RECT 1255.440 210.160 1255.700 210.420 ;
        RECT 1276.140 210.160 1276.400 210.420 ;
        RECT 992.320 209.140 992.580 209.400 ;
        RECT 1000.600 209.140 1000.860 209.400 ;
        RECT 1276.140 209.140 1276.400 209.400 ;
        RECT 1488.200 209.140 1488.460 209.400 ;
        RECT 1503.380 209.140 1503.640 209.400 ;
        RECT 1800.080 209.140 1800.340 209.400 ;
        RECT 1805.600 209.140 1805.860 209.400 ;
        RECT 1817.560 209.140 1817.820 209.400 ;
        RECT 2052.620 209.140 2052.880 209.400 ;
        RECT 2059.060 209.140 2059.320 209.400 ;
        RECT 2074.240 209.140 2074.500 209.400 ;
        RECT 2080.680 209.140 2080.940 209.400 ;
        RECT 2092.640 209.140 2092.900 209.400 ;
        RECT 946.320 208.800 946.580 209.060 ;
        RECT 955.520 208.800 955.780 209.060 ;
        RECT 961.500 208.800 961.760 209.060 ;
        RECT 967.940 208.800 968.200 209.060 ;
        RECT 982.200 208.800 982.460 209.060 ;
        RECT 1511.200 208.800 1511.460 209.060 ;
        RECT 1525.000 208.800 1525.260 209.060 ;
        RECT 1531.440 208.800 1531.700 209.060 ;
        RECT 2326.780 208.800 2327.040 209.060 ;
        RECT 2331.840 208.800 2332.100 209.060 ;
        RECT 2348.400 208.800 2348.660 209.060 ;
        RECT 2354.840 209.140 2355.100 209.400 ;
        RECT 2365.420 209.140 2365.680 209.400 ;
        RECT 2600.480 209.140 2600.740 209.400 ;
        RECT 2606.000 209.140 2606.260 209.400 ;
        RECT 2621.180 209.140 2621.440 209.400 ;
        RECT 2627.620 209.140 2627.880 209.400 ;
        RECT 2639.580 209.140 2639.840 209.400 ;
      LAYER met2 ;
        RECT 1004.280 221.690 1004.540 222.010 ;
        RECT 1206.680 221.690 1206.940 222.010 ;
        RECT 1255.440 221.690 1255.700 222.010 ;
        RECT 1531.900 221.690 1532.160 222.010 ;
        RECT 1547.080 221.690 1547.340 222.010 ;
        RECT 1762.820 221.690 1763.080 222.010 ;
        RECT 1777.080 221.690 1777.340 222.010 ;
        RECT 1821.240 221.690 1821.500 222.010 ;
        RECT 2036.980 221.690 2037.240 222.010 ;
        RECT 2052.160 221.690 2052.420 222.010 ;
        RECT 2095.400 221.690 2095.660 222.010 ;
        RECT 2310.680 221.690 2310.940 222.010 ;
        RECT 2325.860 221.690 2326.120 222.010 ;
        RECT 2369.100 221.690 2369.360 222.010 ;
        RECT 2584.840 221.690 2585.100 222.010 ;
        RECT 2600.020 221.690 2600.280 222.010 ;
        RECT 1004.340 210.965 1004.480 221.690 ;
        RECT 945.835 209.170 946.115 210.965 ;
        RECT 955.035 209.170 955.315 210.965 ;
        RECT 961.015 209.170 961.295 210.965 ;
        RECT 967.455 209.170 967.735 210.965 ;
        RECT 982.635 209.170 982.915 210.965 ;
        RECT 985.855 209.170 986.135 210.965 ;
        RECT 989.075 209.170 989.355 210.965 ;
        RECT 991.835 209.170 992.115 210.965 ;
        RECT 992.320 209.170 992.580 209.430 ;
        RECT 945.835 209.090 946.520 209.170 ;
        RECT 955.035 209.090 955.720 209.170 ;
        RECT 961.015 209.090 961.700 209.170 ;
        RECT 967.455 209.090 968.140 209.170 ;
        RECT 982.260 209.110 992.580 209.170 ;
        RECT 1000.600 209.170 1000.860 209.430 ;
        RECT 1001.035 209.170 1001.315 210.965 ;
        RECT 1004.255 209.170 1004.535 210.965 ;
        RECT 1000.600 209.110 1004.535 209.170 ;
        RECT 982.260 209.090 992.520 209.110 ;
        RECT 945.835 209.030 946.580 209.090 ;
        RECT 945.835 208.565 946.115 209.030 ;
        RECT 946.320 208.770 946.580 209.030 ;
        RECT 955.035 209.030 955.780 209.090 ;
        RECT 955.035 208.565 955.315 209.030 ;
        RECT 955.520 208.770 955.780 209.030 ;
        RECT 961.015 209.030 961.760 209.090 ;
        RECT 961.015 208.565 961.295 209.030 ;
        RECT 961.500 208.770 961.760 209.030 ;
        RECT 967.455 209.030 968.200 209.090 ;
        RECT 967.455 208.565 967.735 209.030 ;
        RECT 967.940 208.770 968.200 209.030 ;
        RECT 982.200 209.030 992.520 209.090 ;
        RECT 1000.660 209.030 1004.535 209.110 ;
        RECT 982.200 208.770 982.460 209.030 ;
        RECT 982.635 208.565 982.915 209.030 ;
        RECT 985.855 208.565 986.135 209.030 ;
        RECT 989.075 208.565 989.355 209.030 ;
        RECT 991.835 208.565 992.115 209.030 ;
        RECT 1001.035 208.565 1001.315 209.030 ;
        RECT 1004.255 208.565 1004.535 209.030 ;
        RECT 1206.740 202.550 1206.880 221.690 ;
        RECT 1255.500 210.450 1255.640 221.690 ;
        RECT 1531.960 210.965 1532.100 221.690 ;
        RECT 1547.140 210.965 1547.280 221.690 ;
        RECT 1762.880 210.965 1763.020 221.690 ;
        RECT 1777.140 221.410 1777.280 221.690 ;
        RECT 1777.140 221.330 1778.200 221.410 ;
        RECT 1777.140 221.270 1778.260 221.330 ;
        RECT 1778.000 221.010 1778.260 221.270 ;
        RECT 1799.620 221.010 1799.880 221.330 ;
        RECT 1778.060 210.965 1778.200 221.010 ;
        RECT 1799.680 210.965 1799.820 221.010 ;
        RECT 1821.300 210.965 1821.440 221.690 ;
        RECT 2037.040 210.965 2037.180 221.690 ;
        RECT 2052.220 210.965 2052.360 221.690 ;
        RECT 2095.460 210.965 2095.600 221.690 ;
        RECT 1255.440 210.130 1255.700 210.450 ;
        RECT 1276.140 210.130 1276.400 210.450 ;
        RECT 1276.200 209.430 1276.340 210.130 ;
        RECT 1276.140 209.110 1276.400 209.430 ;
        RECT 1488.200 209.170 1488.460 209.430 ;
        RECT 1488.835 209.170 1489.115 210.965 ;
        RECT 1488.200 209.110 1489.115 209.170 ;
        RECT 1503.380 209.170 1503.640 209.430 ;
        RECT 1504.015 209.170 1504.295 210.965 ;
        RECT 1507.235 209.170 1507.515 210.965 ;
        RECT 1510.455 209.170 1510.735 210.965 ;
        RECT 1525.635 209.170 1525.915 210.965 ;
        RECT 1531.960 209.170 1532.355 210.965 ;
        RECT 1503.380 209.110 1511.400 209.170 ;
        RECT 1488.260 209.030 1489.115 209.110 ;
        RECT 1503.440 209.090 1511.400 209.110 ;
        RECT 1525.060 209.090 1525.915 209.170 ;
        RECT 1531.500 209.090 1532.355 209.170 ;
        RECT 1503.440 209.030 1511.460 209.090 ;
        RECT 1488.835 208.565 1489.115 209.030 ;
        RECT 1504.015 208.565 1504.295 209.030 ;
        RECT 1507.235 208.565 1507.515 209.030 ;
        RECT 1510.455 208.565 1510.735 209.030 ;
        RECT 1511.200 208.770 1511.460 209.030 ;
        RECT 1525.000 209.030 1525.915 209.090 ;
        RECT 1525.000 208.770 1525.260 209.030 ;
        RECT 1525.635 208.565 1525.915 209.030 ;
        RECT 1531.440 209.030 1532.355 209.090 ;
        RECT 1531.440 208.770 1531.700 209.030 ;
        RECT 1532.075 208.565 1532.355 209.030 ;
        RECT 1544.035 209.170 1544.315 210.965 ;
        RECT 1547.140 209.170 1547.535 210.965 ;
        RECT 1544.035 209.030 1547.535 209.170 ;
        RECT 1544.035 208.565 1544.315 209.030 ;
        RECT 1547.255 208.565 1547.535 209.030 ;
        RECT 1762.835 208.565 1763.115 210.965 ;
        RECT 1778.015 209.170 1778.295 210.965 ;
        RECT 1781.235 209.170 1781.515 210.965 ;
        RECT 1784.455 209.170 1784.735 210.965 ;
        RECT 1778.015 209.030 1784.735 209.170 ;
        RECT 1778.015 208.565 1778.295 209.030 ;
        RECT 1781.235 208.565 1781.515 209.030 ;
        RECT 1784.455 208.565 1784.735 209.030 ;
        RECT 1799.635 209.170 1799.915 210.965 ;
        RECT 1800.080 209.170 1800.340 209.430 ;
        RECT 1799.635 209.110 1800.340 209.170 ;
        RECT 1805.600 209.170 1805.860 209.430 ;
        RECT 1806.075 209.170 1806.355 210.965 ;
        RECT 1805.600 209.110 1806.355 209.170 ;
        RECT 1817.560 209.170 1817.820 209.430 ;
        RECT 1818.035 209.170 1818.315 210.965 ;
        RECT 1821.255 209.170 1821.535 210.965 ;
        RECT 1817.560 209.110 1821.535 209.170 ;
        RECT 1799.635 209.030 1800.280 209.110 ;
        RECT 1805.660 209.030 1806.355 209.110 ;
        RECT 1817.620 209.030 1821.535 209.110 ;
        RECT 1799.635 208.565 1799.915 209.030 ;
        RECT 1806.075 208.565 1806.355 209.030 ;
        RECT 1818.035 208.565 1818.315 209.030 ;
        RECT 1821.255 208.565 1821.535 209.030 ;
        RECT 2036.835 209.100 2037.180 210.965 ;
        RECT 2052.015 209.170 2052.360 210.965 ;
        RECT 2052.620 209.170 2052.880 209.430 ;
        RECT 2052.015 209.110 2052.880 209.170 ;
        RECT 2058.455 209.170 2058.735 210.965 ;
        RECT 2059.060 209.170 2059.320 209.430 ;
        RECT 2058.455 209.110 2059.320 209.170 ;
        RECT 2073.635 209.170 2073.915 210.965 ;
        RECT 2074.240 209.170 2074.500 209.430 ;
        RECT 2073.635 209.110 2074.500 209.170 ;
        RECT 2080.075 209.170 2080.355 210.965 ;
        RECT 2080.680 209.170 2080.940 209.430 ;
        RECT 2080.075 209.110 2080.940 209.170 ;
        RECT 2092.035 209.170 2092.315 210.965 ;
        RECT 2092.700 209.430 2092.840 209.585 ;
        RECT 2092.640 209.170 2092.900 209.430 ;
        RECT 2095.255 209.170 2095.600 210.965 ;
        RECT 2036.835 208.565 2037.115 209.100 ;
        RECT 2052.015 209.030 2052.820 209.110 ;
        RECT 2058.455 209.030 2059.260 209.110 ;
        RECT 2073.635 209.030 2074.440 209.110 ;
        RECT 2080.075 209.030 2080.880 209.110 ;
        RECT 2092.035 209.100 2095.600 209.170 ;
        RECT 2310.740 210.965 2310.880 221.690 ;
        RECT 2325.920 210.965 2326.060 221.690 ;
        RECT 2369.160 210.965 2369.300 221.690 ;
        RECT 2584.900 210.965 2585.040 221.690 ;
        RECT 2600.080 210.965 2600.220 221.690 ;
        RECT 2092.035 209.030 2095.535 209.100 ;
        RECT 2310.740 209.030 2311.115 210.965 ;
        RECT 2325.920 209.170 2326.295 210.965 ;
        RECT 2332.455 209.170 2332.735 210.965 ;
        RECT 2325.920 209.090 2326.980 209.170 ;
        RECT 2331.900 209.090 2332.735 209.170 ;
        RECT 2325.920 209.030 2327.040 209.090 ;
        RECT 2052.015 208.565 2052.295 209.030 ;
        RECT 2058.455 208.565 2058.735 209.030 ;
        RECT 2073.635 208.565 2073.915 209.030 ;
        RECT 2080.075 208.565 2080.355 209.030 ;
        RECT 2092.035 208.565 2092.315 209.030 ;
        RECT 2095.255 208.565 2095.535 209.030 ;
        RECT 2310.835 208.565 2311.115 209.030 ;
        RECT 2326.015 208.565 2326.295 209.030 ;
        RECT 2326.780 208.770 2327.040 209.030 ;
        RECT 2331.840 209.030 2332.735 209.090 ;
        RECT 2331.840 208.770 2332.100 209.030 ;
        RECT 2332.455 208.565 2332.735 209.030 ;
        RECT 2347.635 209.170 2347.915 210.965 ;
        RECT 2354.075 209.170 2354.355 210.965 ;
        RECT 2354.840 209.170 2355.100 209.430 ;
        RECT 2347.635 209.090 2348.600 209.170 ;
        RECT 2354.075 209.110 2355.100 209.170 ;
        RECT 2365.420 209.170 2365.680 209.430 ;
        RECT 2366.035 209.170 2366.315 210.965 ;
        RECT 2369.160 209.170 2369.535 210.965 ;
        RECT 2365.420 209.110 2369.535 209.170 ;
        RECT 2347.635 209.030 2348.660 209.090 ;
        RECT 2347.635 208.565 2347.915 209.030 ;
        RECT 2348.400 208.770 2348.660 209.030 ;
        RECT 2354.075 209.030 2355.040 209.110 ;
        RECT 2365.480 209.030 2369.535 209.110 ;
        RECT 2354.075 208.565 2354.355 209.030 ;
        RECT 2366.035 208.565 2366.315 209.030 ;
        RECT 2369.255 208.565 2369.535 209.030 ;
        RECT 2584.835 208.565 2585.115 210.965 ;
        RECT 2600.015 209.170 2600.295 210.965 ;
        RECT 2600.480 209.170 2600.740 209.430 ;
        RECT 2600.015 209.110 2600.740 209.170 ;
        RECT 2606.000 209.170 2606.260 209.430 ;
        RECT 2606.455 209.170 2606.735 210.965 ;
        RECT 2606.000 209.110 2606.735 209.170 ;
        RECT 2621.180 209.170 2621.440 209.430 ;
        RECT 2621.635 209.170 2621.915 210.965 ;
        RECT 2621.180 209.110 2621.915 209.170 ;
        RECT 2627.620 209.170 2627.880 209.430 ;
        RECT 2628.075 209.170 2628.355 210.965 ;
        RECT 2627.620 209.110 2628.355 209.170 ;
        RECT 2639.580 209.170 2639.840 209.430 ;
        RECT 2640.035 209.170 2640.315 210.965 ;
        RECT 2643.255 209.170 2643.535 210.965 ;
        RECT 2639.580 209.110 2643.535 209.170 ;
        RECT 2600.015 209.030 2600.680 209.110 ;
        RECT 2606.060 209.030 2606.735 209.110 ;
        RECT 2621.240 209.030 2621.915 209.110 ;
        RECT 2627.680 209.030 2628.355 209.110 ;
        RECT 2639.640 209.030 2643.535 209.110 ;
        RECT 2600.015 208.565 2600.295 209.030 ;
        RECT 2606.455 208.565 2606.735 209.030 ;
        RECT 2621.635 208.565 2621.915 209.030 ;
        RECT 2628.075 208.565 2628.355 209.030 ;
        RECT 2640.035 208.565 2640.315 209.030 ;
        RECT 2643.255 208.565 2643.535 209.030 ;
        RECT 1203.740 202.410 1206.880 202.550 ;
        RECT 1203.740 201.920 1203.880 202.410 ;
        RECT 1202.800 200.040 1204.750 201.920 ;
      LAYER via2 ;
        RECT 1203.660 200.840 1203.960 201.140 ;
      LAYER met3 ;
        RECT 1198.650 199.950 1200.570 201.890 ;
        RECT 1202.800 200.040 1204.750 201.920 ;
        RECT 1199.480 199.350 1199.780 199.950 ;
        RECT 1199.480 199.050 1206.730 199.350 ;
        RECT 1206.430 198.000 1206.730 199.050 ;
        RECT 1206.300 158.400 1230.245 198.000 ;
      LAYER via3 ;
        RECT 1199.470 200.730 1199.790 201.050 ;
        RECT 1203.635 200.815 1203.985 201.165 ;
      LAYER met4 ;
        RECT 1198.650 199.950 1200.570 201.890 ;
        RECT 1203.010 200.190 1204.610 201.790 ;
      LAYER via4 ;
        RECT 1198.830 200.090 1200.430 201.690 ;
      LAYER met5 ;
        RECT 1202.890 201.900 1204.730 201.910 ;
        RECT 1201.030 201.890 1204.730 201.900 ;
        RECT 1198.650 200.070 1204.730 201.890 ;
        RECT 1198.650 200.030 1204.330 200.070 ;
        RECT 1198.650 199.950 1200.570 200.030 ;
    END
  END vssd
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1488.730 5013.835 1668.270 5018.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2895.605 174.150 2919.505 200.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1725.530 4954.040 1725.850 4954.100 ;
        RECT 1862.610 4954.040 1862.930 4954.100 ;
        RECT 1725.530 4953.900 1862.930 4954.040 ;
        RECT 1725.530 4953.840 1725.850 4953.900 ;
        RECT 1862.610 4953.840 1862.930 4953.900 ;
        RECT 1863.070 4954.040 1863.390 4954.100 ;
        RECT 1863.070 4953.900 1918.040 4954.040 ;
        RECT 1863.070 4953.840 1863.390 4953.900 ;
        RECT 1168.470 4953.360 1168.790 4953.420 ;
        RECT 1426.530 4953.360 1426.850 4953.420 ;
        RECT 1710.810 4953.360 1711.130 4953.420 ;
        RECT 1725.070 4953.360 1725.390 4953.420 ;
        RECT 975.360 4953.220 1725.390 4953.360 ;
        RECT 1917.900 4953.360 1918.040 4953.900 ;
        RECT 2000.610 4953.700 2000.930 4953.760 ;
        RECT 2097.670 4953.700 2097.990 4953.760 ;
        RECT 2000.610 4953.560 2097.990 4953.700 ;
        RECT 2000.610 4953.500 2000.930 4953.560 ;
        RECT 2097.670 4953.500 2097.990 4953.560 ;
        RECT 2193.810 4953.700 2194.130 4953.760 ;
        RECT 2290.870 4953.700 2291.190 4953.760 ;
        RECT 2193.810 4953.560 2291.190 4953.700 ;
        RECT 2193.810 4953.500 2194.130 4953.560 ;
        RECT 2290.870 4953.500 2291.190 4953.560 ;
        RECT 2387.010 4953.700 2387.330 4953.760 ;
        RECT 2637.710 4953.700 2638.030 4953.760 ;
        RECT 3146.470 4953.700 3146.790 4953.760 ;
        RECT 3156.130 4953.700 3156.450 4953.760 ;
        RECT 2387.010 4953.560 3156.450 4953.700 ;
        RECT 2387.010 4953.500 2387.330 4953.560 ;
        RECT 2637.710 4953.500 2638.030 4953.560 ;
        RECT 3146.470 4953.500 3146.790 4953.560 ;
        RECT 3156.130 4953.500 3156.450 4953.560 ;
        RECT 1932.070 4953.360 1932.390 4953.420 ;
        RECT 1917.900 4953.220 1932.390 4953.360 ;
        RECT 606.350 4953.020 606.670 4953.080 ;
        RECT 510.300 4952.880 606.670 4953.020 ;
        RECT 510.300 4952.680 510.440 4952.880 ;
        RECT 606.350 4952.820 606.670 4952.880 ;
        RECT 482.700 4952.540 510.440 4952.680 ;
        RECT 482.700 4951.320 482.840 4952.540 ;
        RECT 800.930 4952.340 801.250 4952.400 ;
        RECT 800.930 4952.200 869.700 4952.340 ;
        RECT 800.930 4952.140 801.250 4952.200 ;
        RECT 869.560 4952.060 869.700 4952.200 ;
        RECT 869.470 4951.800 869.790 4952.060 ;
        RECT 912.250 4952.000 912.570 4952.060 ;
        RECT 975.360 4952.000 975.500 4953.220 ;
        RECT 1168.470 4953.160 1168.790 4953.220 ;
        RECT 1426.530 4953.160 1426.850 4953.220 ;
        RECT 1710.810 4953.160 1711.130 4953.220 ;
        RECT 1725.070 4953.160 1725.390 4953.220 ;
        RECT 1932.070 4953.160 1932.390 4953.220 ;
        RECT 2097.670 4952.680 2097.990 4952.740 ;
        RECT 2193.810 4952.680 2194.130 4952.740 ;
        RECT 2097.670 4952.540 2194.130 4952.680 ;
        RECT 2097.670 4952.480 2097.990 4952.540 ;
        RECT 2193.810 4952.480 2194.130 4952.540 ;
        RECT 2290.870 4952.680 2291.190 4952.740 ;
        RECT 2380.570 4952.680 2380.890 4952.740 ;
        RECT 2387.010 4952.680 2387.330 4952.740 ;
        RECT 2290.870 4952.540 2387.330 4952.680 ;
        RECT 2290.870 4952.480 2291.190 4952.540 ;
        RECT 2380.570 4952.480 2380.890 4952.540 ;
        RECT 2387.010 4952.480 2387.330 4952.540 ;
        RECT 1932.070 4952.340 1932.390 4952.400 ;
        RECT 1935.750 4952.340 1936.070 4952.400 ;
        RECT 2000.610 4952.340 2000.930 4952.400 ;
        RECT 1932.070 4952.200 2000.930 4952.340 ;
        RECT 1932.070 4952.140 1932.390 4952.200 ;
        RECT 1935.750 4952.140 1936.070 4952.200 ;
        RECT 2000.610 4952.140 2000.930 4952.200 ;
        RECT 912.250 4951.860 975.500 4952.000 ;
        RECT 912.250 4951.800 912.570 4951.860 ;
        RECT 703.410 4951.660 703.730 4951.720 ;
        RECT 800.010 4951.660 800.330 4951.720 ;
        RECT 676.360 4951.520 703.730 4951.660 ;
        RECT 421.980 4951.180 482.840 4951.320 ;
        RECT 655.110 4951.320 655.430 4951.380 ;
        RECT 676.360 4951.320 676.500 4951.520 ;
        RECT 703.410 4951.460 703.730 4951.520 ;
        RECT 772.500 4951.520 800.330 4951.660 ;
        RECT 655.110 4951.180 676.500 4951.320 ;
        RECT 703.870 4951.320 704.190 4951.380 ;
        RECT 772.500 4951.320 772.640 4951.520 ;
        RECT 800.010 4951.460 800.330 4951.520 ;
        RECT 703.870 4951.180 772.640 4951.320 ;
        RECT 869.470 4951.320 869.790 4951.380 ;
        RECT 912.340 4951.320 912.480 4951.800 ;
        RECT 869.470 4951.180 912.480 4951.320 ;
        RECT 211.670 4950.640 211.990 4950.700 ;
        RECT 397.510 4950.640 397.830 4950.700 ;
        RECT 421.980 4950.640 422.120 4951.180 ;
        RECT 655.110 4951.120 655.430 4951.180 ;
        RECT 703.870 4951.120 704.190 4951.180 ;
        RECT 869.470 4951.120 869.790 4951.180 ;
        RECT 211.670 4950.500 422.120 4950.640 ;
        RECT 3156.130 4950.640 3156.450 4950.700 ;
        RECT 3367.730 4950.640 3368.050 4950.700 ;
        RECT 3156.130 4950.500 3368.050 4950.640 ;
        RECT 211.670 4950.440 211.990 4950.500 ;
        RECT 397.510 4950.440 397.830 4950.500 ;
        RECT 3156.130 4950.440 3156.450 4950.500 ;
        RECT 3367.730 4950.440 3368.050 4950.500 ;
        RECT 3367.730 4823.820 3368.050 4823.880 ;
        RECT 3376.930 4823.820 3377.250 4823.880 ;
        RECT 3367.730 4823.680 3377.250 4823.820 ;
        RECT 3367.730 4823.620 3368.050 4823.680 ;
        RECT 3376.930 4823.620 3377.250 4823.680 ;
        RECT 208.910 4790.500 209.230 4790.560 ;
        RECT 211.670 4790.500 211.990 4790.560 ;
        RECT 208.910 4790.360 211.990 4790.500 ;
        RECT 208.910 4790.300 209.230 4790.360 ;
        RECT 211.670 4790.300 211.990 4790.360 ;
        RECT 3367.730 4372.640 3368.050 4372.700 ;
        RECT 3376.930 4372.640 3377.250 4372.700 ;
        RECT 3367.730 4372.500 3377.250 4372.640 ;
        RECT 3367.730 4372.440 3368.050 4372.500 ;
        RECT 3376.930 4372.440 3377.250 4372.500 ;
        RECT 208.910 3936.420 209.230 3936.480 ;
        RECT 213.050 3936.420 213.370 3936.480 ;
        RECT 208.910 3936.280 213.370 3936.420 ;
        RECT 208.910 3936.220 209.230 3936.280 ;
        RECT 213.050 3936.220 213.370 3936.280 ;
        RECT 3367.730 3932.000 3368.050 3932.060 ;
        RECT 3376.930 3932.000 3377.250 3932.060 ;
        RECT 3367.730 3931.860 3377.250 3932.000 ;
        RECT 3367.730 3931.800 3368.050 3931.860 ;
        RECT 3376.930 3931.800 3377.250 3931.860 ;
        RECT 208.910 3720.860 209.230 3720.920 ;
        RECT 211.670 3720.860 211.990 3720.920 ;
        RECT 213.050 3720.860 213.370 3720.920 ;
        RECT 208.910 3720.720 213.370 3720.860 ;
        RECT 208.910 3720.660 209.230 3720.720 ;
        RECT 211.670 3720.660 211.990 3720.720 ;
        RECT 213.050 3720.660 213.370 3720.720 ;
        RECT 3367.730 3703.520 3368.050 3703.580 ;
        RECT 3376.930 3703.520 3377.250 3703.580 ;
        RECT 3367.730 3703.380 3377.250 3703.520 ;
        RECT 3367.730 3703.320 3368.050 3703.380 ;
        RECT 3376.930 3703.320 3377.250 3703.380 ;
        RECT 211.670 3698.080 211.990 3698.140 ;
        RECT 213.050 3698.080 213.370 3698.140 ;
        RECT 211.670 3697.940 213.370 3698.080 ;
        RECT 211.670 3697.880 211.990 3697.940 ;
        RECT 213.050 3697.880 213.370 3697.940 ;
        RECT 208.910 3504.960 209.230 3505.020 ;
        RECT 213.050 3504.960 213.370 3505.020 ;
        RECT 208.910 3504.820 213.370 3504.960 ;
        RECT 208.910 3504.760 209.230 3504.820 ;
        RECT 213.050 3504.760 213.370 3504.820 ;
        RECT 3367.730 3476.740 3368.050 3476.800 ;
        RECT 3376.930 3476.740 3377.250 3476.800 ;
        RECT 3367.730 3476.600 3377.250 3476.740 ;
        RECT 3367.730 3476.540 3368.050 3476.600 ;
        RECT 3376.930 3476.540 3377.250 3476.600 ;
        RECT 213.050 3392.760 213.370 3392.820 ;
        RECT 214.890 3392.760 215.210 3392.820 ;
        RECT 213.050 3392.620 215.210 3392.760 ;
        RECT 213.050 3392.560 213.370 3392.620 ;
        RECT 214.890 3392.560 215.210 3392.620 ;
        RECT 212.130 3380.860 212.450 3380.920 ;
        RECT 214.890 3380.860 215.210 3380.920 ;
        RECT 212.130 3380.720 215.210 3380.860 ;
        RECT 212.130 3380.660 212.450 3380.720 ;
        RECT 214.890 3380.660 215.210 3380.720 ;
        RECT 208.910 3293.480 209.230 3293.540 ;
        RECT 212.130 3293.480 212.450 3293.540 ;
        RECT 213.510 3293.480 213.830 3293.540 ;
        RECT 208.910 3293.340 213.830 3293.480 ;
        RECT 208.910 3293.280 209.230 3293.340 ;
        RECT 212.130 3293.280 212.450 3293.340 ;
        RECT 213.510 3293.280 213.830 3293.340 ;
        RECT 3367.730 3255.740 3368.050 3255.800 ;
        RECT 3376.930 3255.740 3377.250 3255.800 ;
        RECT 3367.730 3255.600 3377.250 3255.740 ;
        RECT 3367.730 3255.540 3368.050 3255.600 ;
        RECT 3376.930 3255.540 3377.250 3255.600 ;
        RECT 213.510 3160.200 213.830 3160.260 ;
        RECT 214.890 3160.200 215.210 3160.260 ;
        RECT 213.510 3160.060 215.210 3160.200 ;
        RECT 213.510 3160.000 213.830 3160.060 ;
        RECT 214.890 3160.000 215.210 3160.060 ;
        RECT 208.910 3077.580 209.230 3077.640 ;
        RECT 214.890 3077.580 215.210 3077.640 ;
        RECT 208.910 3077.440 215.210 3077.580 ;
        RECT 208.910 3077.380 209.230 3077.440 ;
        RECT 214.890 3077.380 215.210 3077.440 ;
        RECT 3367.730 3031.000 3368.050 3031.060 ;
        RECT 3375.090 3031.000 3375.410 3031.060 ;
        RECT 3376.930 3031.000 3377.250 3031.060 ;
        RECT 3367.730 3030.860 3377.250 3031.000 ;
        RECT 3367.730 3030.800 3368.050 3030.860 ;
        RECT 3375.090 3030.800 3375.410 3030.860 ;
        RECT 3376.930 3030.800 3377.250 3030.860 ;
        RECT 3368.650 2973.880 3368.970 2973.940 ;
        RECT 3375.090 2973.880 3375.410 2973.940 ;
        RECT 3368.650 2973.740 3375.410 2973.880 ;
        RECT 3368.650 2973.680 3368.970 2973.740 ;
        RECT 3375.090 2973.680 3375.410 2973.740 ;
        RECT 3368.650 2877.320 3368.970 2877.380 ;
        RECT 3371.870 2877.320 3372.190 2877.380 ;
        RECT 3368.650 2877.180 3372.190 2877.320 ;
        RECT 3368.650 2877.120 3368.970 2877.180 ;
        RECT 3371.870 2877.120 3372.190 2877.180 ;
        RECT 208.910 2856.240 209.230 2856.300 ;
        RECT 213.970 2856.240 214.290 2856.300 ;
        RECT 208.910 2856.100 214.290 2856.240 ;
        RECT 208.910 2856.040 209.230 2856.100 ;
        RECT 213.970 2856.040 214.290 2856.100 ;
        RECT 3370.030 2799.800 3370.350 2799.860 ;
        RECT 3371.870 2799.800 3372.190 2799.860 ;
        RECT 3376.930 2799.800 3377.250 2799.860 ;
        RECT 3370.030 2799.660 3377.250 2799.800 ;
        RECT 3370.030 2799.600 3370.350 2799.660 ;
        RECT 3371.870 2799.600 3372.190 2799.660 ;
        RECT 3376.930 2799.600 3377.250 2799.660 ;
        RECT 213.050 2773.960 213.370 2774.020 ;
        RECT 213.970 2773.960 214.290 2774.020 ;
        RECT 213.050 2773.820 214.290 2773.960 ;
        RECT 213.050 2773.760 213.370 2773.820 ;
        RECT 213.970 2773.760 214.290 2773.820 ;
        RECT 208.910 2640.340 209.230 2640.400 ;
        RECT 213.050 2640.340 213.370 2640.400 ;
        RECT 208.910 2640.200 213.370 2640.340 ;
        RECT 208.910 2640.140 209.230 2640.200 ;
        RECT 213.050 2640.140 213.370 2640.200 ;
        RECT 3368.650 2511.820 3368.970 2511.880 ;
        RECT 3369.570 2511.820 3369.890 2511.880 ;
        RECT 3368.650 2511.680 3369.890 2511.820 ;
        RECT 3368.650 2511.620 3368.970 2511.680 ;
        RECT 3369.570 2511.620 3369.890 2511.680 ;
        RECT 3369.110 2346.580 3369.430 2346.640 ;
        RECT 3368.740 2346.440 3369.430 2346.580 ;
        RECT 3368.740 2345.960 3368.880 2346.440 ;
        RECT 3369.110 2346.380 3369.430 2346.440 ;
        RECT 3368.650 2345.700 3368.970 2345.960 ;
        RECT 3368.650 2318.360 3368.970 2318.420 ;
        RECT 3370.030 2318.360 3370.350 2318.420 ;
        RECT 3368.650 2318.220 3370.350 2318.360 ;
        RECT 3368.650 2318.160 3368.970 2318.220 ;
        RECT 3370.030 2318.160 3370.350 2318.220 ;
        RECT 213.050 2221.800 213.370 2221.860 ;
        RECT 213.970 2221.800 214.290 2221.860 ;
        RECT 213.050 2221.660 214.290 2221.800 ;
        RECT 213.050 2221.600 213.370 2221.660 ;
        RECT 213.970 2221.600 214.290 2221.660 ;
        RECT 3368.650 2221.800 3368.970 2221.860 ;
        RECT 3370.030 2221.800 3370.350 2221.860 ;
        RECT 3368.650 2221.660 3370.350 2221.800 ;
        RECT 3368.650 2221.600 3368.970 2221.660 ;
        RECT 3370.030 2221.600 3370.350 2221.660 ;
        RECT 213.510 2207.860 213.830 2207.920 ;
        RECT 213.970 2207.860 214.290 2207.920 ;
        RECT 213.510 2207.720 214.290 2207.860 ;
        RECT 213.510 2207.660 213.830 2207.720 ;
        RECT 213.970 2207.660 214.290 2207.720 ;
        RECT 213.050 2111.640 213.370 2111.700 ;
        RECT 213.510 2111.640 213.830 2111.700 ;
        RECT 213.050 2111.500 213.830 2111.640 ;
        RECT 213.050 2111.440 213.370 2111.500 ;
        RECT 213.510 2111.440 213.830 2111.500 ;
        RECT 3368.190 2103.820 3368.510 2103.880 ;
        RECT 3369.110 2103.820 3369.430 2103.880 ;
        RECT 3368.190 2103.680 3369.430 2103.820 ;
        RECT 3368.190 2103.620 3368.510 2103.680 ;
        RECT 3369.110 2103.620 3369.430 2103.680 ;
        RECT 213.050 2028.680 213.370 2028.740 ;
        RECT 214.430 2028.680 214.750 2028.740 ;
        RECT 213.050 2028.540 214.750 2028.680 ;
        RECT 213.050 2028.480 213.370 2028.540 ;
        RECT 214.430 2028.480 214.750 2028.540 ;
        RECT 3369.110 2007.940 3369.430 2008.000 ;
        RECT 3376.470 2007.940 3376.790 2008.000 ;
        RECT 3369.110 2007.800 3376.790 2007.940 ;
        RECT 3369.110 2007.740 3369.430 2007.800 ;
        RECT 3376.470 2007.740 3376.790 2007.800 ;
        RECT 208.910 2006.920 209.230 2006.980 ;
        RECT 214.430 2006.920 214.750 2006.980 ;
        RECT 208.910 2006.780 214.750 2006.920 ;
        RECT 208.910 2006.720 209.230 2006.780 ;
        RECT 214.430 2006.720 214.750 2006.780 ;
        RECT 3368.190 1916.140 3368.510 1916.200 ;
        RECT 3376.470 1916.140 3376.790 1916.200 ;
        RECT 3368.190 1916.000 3376.790 1916.140 ;
        RECT 3368.190 1915.940 3368.510 1916.000 ;
        RECT 3376.470 1915.940 3376.790 1916.000 ;
        RECT 213.970 1863.100 214.290 1863.160 ;
        RECT 214.890 1863.100 215.210 1863.160 ;
        RECT 213.970 1862.960 215.210 1863.100 ;
        RECT 213.970 1862.900 214.290 1862.960 ;
        RECT 214.890 1862.900 215.210 1862.960 ;
        RECT 212.590 1839.300 212.910 1839.360 ;
        RECT 213.970 1839.300 214.290 1839.360 ;
        RECT 212.590 1839.160 214.290 1839.300 ;
        RECT 212.590 1839.100 212.910 1839.160 ;
        RECT 213.970 1839.100 214.290 1839.160 ;
        RECT 208.910 1791.360 209.230 1791.420 ;
        RECT 212.590 1791.360 212.910 1791.420 ;
        RECT 208.910 1791.220 212.910 1791.360 ;
        RECT 208.910 1791.160 209.230 1791.220 ;
        RECT 212.590 1791.160 212.910 1791.220 ;
        RECT 3368.190 1687.660 3368.510 1687.720 ;
        RECT 3376.930 1687.660 3377.250 1687.720 ;
        RECT 3368.190 1687.520 3377.250 1687.660 ;
        RECT 3368.190 1687.460 3368.510 1687.520 ;
        RECT 3376.930 1687.460 3377.250 1687.520 ;
        RECT 208.910 1570.360 209.230 1570.420 ;
        RECT 212.590 1570.360 212.910 1570.420 ;
        RECT 213.510 1570.360 213.830 1570.420 ;
        RECT 208.910 1570.220 213.830 1570.360 ;
        RECT 208.910 1570.160 209.230 1570.220 ;
        RECT 212.590 1570.160 212.910 1570.220 ;
        RECT 213.510 1570.160 213.830 1570.220 ;
        RECT 3368.190 1468.020 3368.510 1468.080 ;
        RECT 3369.570 1468.020 3369.890 1468.080 ;
        RECT 3376.930 1468.020 3377.250 1468.080 ;
        RECT 3368.190 1467.880 3377.250 1468.020 ;
        RECT 3368.190 1467.820 3368.510 1467.880 ;
        RECT 3369.570 1467.820 3369.890 1467.880 ;
        RECT 3376.930 1467.820 3377.250 1467.880 ;
        RECT 208.910 1359.560 209.230 1359.620 ;
        RECT 213.510 1359.560 213.830 1359.620 ;
        RECT 208.910 1359.420 213.830 1359.560 ;
        RECT 208.910 1359.360 209.230 1359.420 ;
        RECT 213.510 1359.360 213.830 1359.420 ;
        RECT 3368.190 1237.500 3368.510 1237.560 ;
        RECT 3369.570 1237.500 3369.890 1237.560 ;
        RECT 3376.930 1237.500 3377.250 1237.560 ;
        RECT 3368.190 1237.360 3377.250 1237.500 ;
        RECT 3368.190 1237.300 3368.510 1237.360 ;
        RECT 3369.570 1237.300 3369.890 1237.360 ;
        RECT 3376.930 1237.300 3377.250 1237.360 ;
        RECT 208.910 1143.320 209.230 1143.380 ;
        RECT 213.510 1143.320 213.830 1143.380 ;
        RECT 208.910 1143.180 213.830 1143.320 ;
        RECT 208.910 1143.120 209.230 1143.180 ;
        RECT 213.510 1143.120 213.830 1143.180 ;
        RECT 3368.190 1016.840 3368.510 1016.900 ;
        RECT 3376.930 1016.840 3377.250 1016.900 ;
        RECT 3368.190 1016.700 3377.250 1016.840 ;
        RECT 3368.190 1016.640 3368.510 1016.700 ;
        RECT 3376.930 1016.640 3377.250 1016.700 ;
        RECT 208.910 927.420 209.230 927.480 ;
        RECT 211.670 927.420 211.990 927.480 ;
        RECT 213.510 927.420 213.830 927.480 ;
        RECT 208.910 927.280 213.830 927.420 ;
        RECT 208.910 927.220 209.230 927.280 ;
        RECT 211.670 927.220 211.990 927.280 ;
        RECT 213.510 927.220 213.830 927.280 ;
        RECT 3367.270 786.660 3367.590 786.720 ;
        RECT 3376.930 786.660 3377.250 786.720 ;
        RECT 3367.270 786.520 3377.250 786.660 ;
        RECT 3367.270 786.460 3367.590 786.520 ;
        RECT 3376.930 786.460 3377.250 786.520 ;
        RECT 3367.270 560.560 3367.590 560.620 ;
        RECT 3376.930 560.560 3377.250 560.620 ;
        RECT 3367.270 560.420 3377.250 560.560 ;
        RECT 3367.270 560.360 3367.590 560.420 ;
        RECT 3376.930 560.360 3377.250 560.420 ;
        RECT 211.670 228.720 211.990 228.780 ;
        RECT 704.790 228.720 705.110 228.780 ;
        RECT 211.670 228.580 705.110 228.720 ;
        RECT 211.670 228.520 211.990 228.580 ;
        RECT 704.790 228.520 705.110 228.580 ;
        RECT 2883.810 213.760 2884.130 213.820 ;
        RECT 3367.270 213.760 3367.590 213.820 ;
        RECT 2883.810 213.620 3367.590 213.760 ;
        RECT 2883.810 213.560 2884.130 213.620 ;
        RECT 3367.270 213.560 3367.590 213.620 ;
        RECT 731.470 210.020 731.790 210.080 ;
        RECT 2845.630 210.020 2845.950 210.080 ;
        RECT 2883.810 210.020 2884.130 210.080 ;
        RECT 731.470 209.880 2884.130 210.020 ;
        RECT 731.470 209.820 731.790 209.880 ;
        RECT 2845.630 209.820 2845.950 209.880 ;
        RECT 2883.810 209.820 2884.130 209.880 ;
        RECT 723.190 203.900 723.510 203.960 ;
        RECT 731.470 203.900 731.790 203.960 ;
        RECT 723.190 203.760 731.790 203.900 ;
        RECT 723.190 203.700 723.510 203.760 ;
        RECT 731.470 203.700 731.790 203.760 ;
        RECT 704.950 200.500 705.270 200.560 ;
        RECT 715.370 200.500 715.690 200.560 ;
        RECT 723.190 200.500 723.510 200.560 ;
        RECT 704.950 200.360 723.510 200.500 ;
        RECT 704.950 200.300 705.270 200.360 ;
        RECT 712.930 200.000 713.070 200.360 ;
        RECT 715.370 200.300 715.690 200.360 ;
        RECT 723.190 200.300 723.510 200.360 ;
        RECT 712.865 190.025 713.095 200.000 ;
      LAYER via ;
        RECT 1725.560 4953.840 1725.820 4954.100 ;
        RECT 1862.640 4953.840 1862.900 4954.100 ;
        RECT 1863.100 4953.840 1863.360 4954.100 ;
        RECT 606.380 4952.820 606.640 4953.080 ;
        RECT 800.960 4952.140 801.220 4952.400 ;
        RECT 869.500 4951.800 869.760 4952.060 ;
        RECT 912.280 4951.800 912.540 4952.060 ;
        RECT 1168.500 4953.160 1168.760 4953.420 ;
        RECT 1426.560 4953.160 1426.820 4953.420 ;
        RECT 1710.840 4953.160 1711.100 4953.420 ;
        RECT 1725.100 4953.160 1725.360 4953.420 ;
        RECT 2000.640 4953.500 2000.900 4953.760 ;
        RECT 2097.700 4953.500 2097.960 4953.760 ;
        RECT 2193.840 4953.500 2194.100 4953.760 ;
        RECT 2290.900 4953.500 2291.160 4953.760 ;
        RECT 2387.040 4953.500 2387.300 4953.760 ;
        RECT 2637.740 4953.500 2638.000 4953.760 ;
        RECT 3146.500 4953.500 3146.760 4953.760 ;
        RECT 3156.160 4953.500 3156.420 4953.760 ;
        RECT 1932.100 4953.160 1932.360 4953.420 ;
        RECT 2097.700 4952.480 2097.960 4952.740 ;
        RECT 2193.840 4952.480 2194.100 4952.740 ;
        RECT 2290.900 4952.480 2291.160 4952.740 ;
        RECT 2380.600 4952.480 2380.860 4952.740 ;
        RECT 2387.040 4952.480 2387.300 4952.740 ;
        RECT 1932.100 4952.140 1932.360 4952.400 ;
        RECT 1935.780 4952.140 1936.040 4952.400 ;
        RECT 2000.640 4952.140 2000.900 4952.400 ;
        RECT 211.700 4950.440 211.960 4950.700 ;
        RECT 397.540 4950.440 397.800 4950.700 ;
        RECT 655.140 4951.120 655.400 4951.380 ;
        RECT 703.440 4951.460 703.700 4951.720 ;
        RECT 703.900 4951.120 704.160 4951.380 ;
        RECT 800.040 4951.460 800.300 4951.720 ;
        RECT 869.500 4951.120 869.760 4951.380 ;
        RECT 3156.160 4950.440 3156.420 4950.700 ;
        RECT 3367.760 4950.440 3368.020 4950.700 ;
        RECT 3367.760 4823.620 3368.020 4823.880 ;
        RECT 3376.960 4823.620 3377.220 4823.880 ;
        RECT 208.940 4790.300 209.200 4790.560 ;
        RECT 211.700 4790.300 211.960 4790.560 ;
        RECT 3367.760 4372.440 3368.020 4372.700 ;
        RECT 3376.960 4372.440 3377.220 4372.700 ;
        RECT 208.940 3936.220 209.200 3936.480 ;
        RECT 213.080 3936.220 213.340 3936.480 ;
        RECT 3367.760 3931.800 3368.020 3932.060 ;
        RECT 3376.960 3931.800 3377.220 3932.060 ;
        RECT 208.940 3720.660 209.200 3720.920 ;
        RECT 211.700 3720.660 211.960 3720.920 ;
        RECT 213.080 3720.660 213.340 3720.920 ;
        RECT 3367.760 3703.320 3368.020 3703.580 ;
        RECT 3376.960 3703.320 3377.220 3703.580 ;
        RECT 211.700 3697.880 211.960 3698.140 ;
        RECT 213.080 3697.880 213.340 3698.140 ;
        RECT 208.940 3504.760 209.200 3505.020 ;
        RECT 213.080 3504.760 213.340 3505.020 ;
        RECT 3367.760 3476.540 3368.020 3476.800 ;
        RECT 3376.960 3476.540 3377.220 3476.800 ;
        RECT 213.080 3392.560 213.340 3392.820 ;
        RECT 214.920 3392.560 215.180 3392.820 ;
        RECT 212.160 3380.660 212.420 3380.920 ;
        RECT 214.920 3380.660 215.180 3380.920 ;
        RECT 208.940 3293.280 209.200 3293.540 ;
        RECT 212.160 3293.280 212.420 3293.540 ;
        RECT 213.540 3293.280 213.800 3293.540 ;
        RECT 3367.760 3255.540 3368.020 3255.800 ;
        RECT 3376.960 3255.540 3377.220 3255.800 ;
        RECT 213.540 3160.000 213.800 3160.260 ;
        RECT 214.920 3160.000 215.180 3160.260 ;
        RECT 208.940 3077.380 209.200 3077.640 ;
        RECT 214.920 3077.380 215.180 3077.640 ;
        RECT 3367.760 3030.800 3368.020 3031.060 ;
        RECT 3375.120 3030.800 3375.380 3031.060 ;
        RECT 3376.960 3030.800 3377.220 3031.060 ;
        RECT 3368.680 2973.680 3368.940 2973.940 ;
        RECT 3375.120 2973.680 3375.380 2973.940 ;
        RECT 3368.680 2877.120 3368.940 2877.380 ;
        RECT 3371.900 2877.120 3372.160 2877.380 ;
        RECT 208.940 2856.040 209.200 2856.300 ;
        RECT 214.000 2856.040 214.260 2856.300 ;
        RECT 3370.060 2799.600 3370.320 2799.860 ;
        RECT 3371.900 2799.600 3372.160 2799.860 ;
        RECT 3376.960 2799.600 3377.220 2799.860 ;
        RECT 213.080 2773.760 213.340 2774.020 ;
        RECT 214.000 2773.760 214.260 2774.020 ;
        RECT 208.940 2640.140 209.200 2640.400 ;
        RECT 213.080 2640.140 213.340 2640.400 ;
        RECT 3368.680 2511.620 3368.940 2511.880 ;
        RECT 3369.600 2511.620 3369.860 2511.880 ;
        RECT 3369.140 2346.380 3369.400 2346.640 ;
        RECT 3368.680 2345.700 3368.940 2345.960 ;
        RECT 3368.680 2318.160 3368.940 2318.420 ;
        RECT 3370.060 2318.160 3370.320 2318.420 ;
        RECT 213.080 2221.600 213.340 2221.860 ;
        RECT 214.000 2221.600 214.260 2221.860 ;
        RECT 3368.680 2221.600 3368.940 2221.860 ;
        RECT 3370.060 2221.600 3370.320 2221.860 ;
        RECT 213.540 2207.660 213.800 2207.920 ;
        RECT 214.000 2207.660 214.260 2207.920 ;
        RECT 213.080 2111.440 213.340 2111.700 ;
        RECT 213.540 2111.440 213.800 2111.700 ;
        RECT 3368.220 2103.620 3368.480 2103.880 ;
        RECT 3369.140 2103.620 3369.400 2103.880 ;
        RECT 213.080 2028.480 213.340 2028.740 ;
        RECT 214.460 2028.480 214.720 2028.740 ;
        RECT 3369.140 2007.740 3369.400 2008.000 ;
        RECT 3376.500 2007.740 3376.760 2008.000 ;
        RECT 208.940 2006.720 209.200 2006.980 ;
        RECT 214.460 2006.720 214.720 2006.980 ;
        RECT 3368.220 1915.940 3368.480 1916.200 ;
        RECT 3376.500 1915.940 3376.760 1916.200 ;
        RECT 214.000 1862.900 214.260 1863.160 ;
        RECT 214.920 1862.900 215.180 1863.160 ;
        RECT 212.620 1839.100 212.880 1839.360 ;
        RECT 214.000 1839.100 214.260 1839.360 ;
        RECT 208.940 1791.160 209.200 1791.420 ;
        RECT 212.620 1791.160 212.880 1791.420 ;
        RECT 3368.220 1687.460 3368.480 1687.720 ;
        RECT 3376.960 1687.460 3377.220 1687.720 ;
        RECT 208.940 1570.160 209.200 1570.420 ;
        RECT 212.620 1570.160 212.880 1570.420 ;
        RECT 213.540 1570.160 213.800 1570.420 ;
        RECT 3368.220 1467.820 3368.480 1468.080 ;
        RECT 3369.600 1467.820 3369.860 1468.080 ;
        RECT 3376.960 1467.820 3377.220 1468.080 ;
        RECT 208.940 1359.360 209.200 1359.620 ;
        RECT 213.540 1359.360 213.800 1359.620 ;
        RECT 3368.220 1237.300 3368.480 1237.560 ;
        RECT 3369.600 1237.300 3369.860 1237.560 ;
        RECT 3376.960 1237.300 3377.220 1237.560 ;
        RECT 208.940 1143.120 209.200 1143.380 ;
        RECT 213.540 1143.120 213.800 1143.380 ;
        RECT 3368.220 1016.640 3368.480 1016.900 ;
        RECT 3376.960 1016.640 3377.220 1016.900 ;
        RECT 208.940 927.220 209.200 927.480 ;
        RECT 211.700 927.220 211.960 927.480 ;
        RECT 213.540 927.220 213.800 927.480 ;
        RECT 3367.300 786.460 3367.560 786.720 ;
        RECT 3376.960 786.460 3377.220 786.720 ;
        RECT 3367.300 560.360 3367.560 560.620 ;
        RECT 3376.960 560.360 3377.220 560.620 ;
        RECT 211.700 228.520 211.960 228.780 ;
        RECT 704.820 228.520 705.080 228.780 ;
        RECT 2883.840 213.560 2884.100 213.820 ;
        RECT 3367.300 213.560 3367.560 213.820 ;
        RECT 731.500 209.820 731.760 210.080 ;
        RECT 2845.660 209.820 2845.920 210.080 ;
        RECT 2883.840 209.820 2884.100 210.080 ;
        RECT 723.220 203.700 723.480 203.960 ;
        RECT 731.500 203.700 731.760 203.960 ;
        RECT 704.980 200.300 705.240 200.560 ;
        RECT 715.400 200.300 715.660 200.560 ;
        RECT 723.220 200.300 723.480 200.560 ;
      LAYER met2 ;
        RECT 1710.820 4987.025 1711.120 4987.415 ;
        RECT 397.665 4977.260 397.945 4979.435 ;
        RECT 397.600 4977.035 397.945 4977.260 ;
        RECT 654.665 4977.330 654.945 4979.435 ;
        RECT 911.665 4977.330 911.945 4979.435 ;
        RECT 1168.665 4977.330 1168.945 4979.435 ;
        RECT 654.665 4977.190 655.340 4977.330 ;
        RECT 654.665 4977.035 654.945 4977.190 ;
        RECT 397.600 4950.730 397.740 4977.035 ;
        RECT 606.380 4952.790 606.640 4953.110 ;
        RECT 606.440 4952.285 606.580 4952.790 ;
        RECT 655.200 4952.285 655.340 4977.190 ;
        RECT 911.665 4977.190 912.480 4977.330 ;
        RECT 911.665 4977.035 911.945 4977.190 ;
        RECT 606.370 4951.915 606.650 4952.285 ;
        RECT 655.130 4951.915 655.410 4952.285 ;
        RECT 800.960 4952.170 801.220 4952.430 ;
        RECT 800.100 4952.110 801.220 4952.170 ;
        RECT 800.100 4952.030 801.160 4952.110 ;
        RECT 912.340 4952.090 912.480 4977.190 ;
        RECT 1168.560 4977.035 1168.945 4977.330 ;
        RECT 1426.665 4977.260 1426.945 4979.435 ;
        RECT 1426.620 4977.035 1426.945 4977.260 ;
        RECT 1168.560 4953.450 1168.700 4977.035 ;
        RECT 1426.620 4953.450 1426.760 4977.035 ;
        RECT 1710.900 4953.450 1711.040 4987.025 ;
        RECT 1935.665 4977.260 1935.945 4979.435 ;
        RECT 2380.665 4977.260 2380.945 4979.435 ;
        RECT 1935.665 4977.035 1935.980 4977.260 ;
        RECT 1862.700 4954.130 1863.300 4954.210 ;
        RECT 1725.560 4953.810 1725.820 4954.130 ;
        RECT 1862.640 4954.070 1863.360 4954.130 ;
        RECT 1862.640 4953.810 1862.900 4954.070 ;
        RECT 1863.100 4953.810 1863.360 4954.070 ;
        RECT 1168.500 4953.130 1168.760 4953.450 ;
        RECT 1426.560 4953.130 1426.820 4953.450 ;
        RECT 1710.840 4953.130 1711.100 4953.450 ;
        RECT 1725.100 4953.360 1725.360 4953.450 ;
        RECT 1725.620 4953.360 1725.760 4953.810 ;
        RECT 1725.100 4953.220 1725.760 4953.360 ;
        RECT 1725.100 4953.130 1725.360 4953.220 ;
        RECT 1932.100 4953.130 1932.360 4953.450 ;
        RECT 1932.160 4952.430 1932.300 4953.130 ;
        RECT 1935.840 4952.430 1935.980 4977.035 ;
        RECT 2380.660 4977.035 2380.945 4977.260 ;
        RECT 2637.665 4977.035 2637.945 4979.435 ;
        RECT 3146.665 4977.330 3146.945 4979.435 ;
        RECT 3146.560 4977.035 3146.945 4977.330 ;
        RECT 2000.640 4953.470 2000.900 4953.790 ;
        RECT 2097.700 4953.470 2097.960 4953.790 ;
        RECT 2193.840 4953.470 2194.100 4953.790 ;
        RECT 2290.900 4953.470 2291.160 4953.790 ;
        RECT 2000.700 4952.430 2000.840 4953.470 ;
        RECT 2097.760 4952.770 2097.900 4953.470 ;
        RECT 2193.900 4952.770 2194.040 4953.470 ;
        RECT 2290.960 4952.770 2291.100 4953.470 ;
        RECT 2380.660 4952.770 2380.800 4977.035 ;
        RECT 2637.800 4953.790 2637.940 4977.035 ;
        RECT 3146.560 4953.790 3146.700 4977.035 ;
        RECT 2387.040 4953.470 2387.300 4953.790 ;
        RECT 2637.740 4953.470 2638.000 4953.790 ;
        RECT 3146.500 4953.470 3146.760 4953.790 ;
        RECT 3156.160 4953.470 3156.420 4953.790 ;
        RECT 2387.100 4952.770 2387.240 4953.470 ;
        RECT 2097.700 4952.450 2097.960 4952.770 ;
        RECT 2193.840 4952.450 2194.100 4952.770 ;
        RECT 2290.900 4952.450 2291.160 4952.770 ;
        RECT 2380.600 4952.450 2380.860 4952.770 ;
        RECT 2387.040 4952.450 2387.300 4952.770 ;
        RECT 1932.100 4952.110 1932.360 4952.430 ;
        RECT 1935.780 4952.110 1936.040 4952.430 ;
        RECT 2000.640 4952.110 2000.900 4952.430 ;
        RECT 655.200 4951.410 655.340 4951.915 ;
        RECT 800.100 4951.750 800.240 4952.030 ;
        RECT 869.500 4951.770 869.760 4952.090 ;
        RECT 912.280 4951.770 912.540 4952.090 ;
        RECT 703.440 4951.490 703.700 4951.750 ;
        RECT 703.440 4951.430 704.100 4951.490 ;
        RECT 800.040 4951.430 800.300 4951.750 ;
        RECT 703.500 4951.410 704.100 4951.430 ;
        RECT 869.560 4951.410 869.700 4951.770 ;
        RECT 655.140 4951.090 655.400 4951.410 ;
        RECT 703.500 4951.350 704.160 4951.410 ;
        RECT 703.900 4951.090 704.160 4951.350 ;
        RECT 869.500 4951.090 869.760 4951.410 ;
        RECT 3156.220 4950.730 3156.360 4953.470 ;
        RECT 211.700 4950.410 211.960 4950.730 ;
        RECT 397.540 4950.410 397.800 4950.730 ;
        RECT 3156.160 4950.410 3156.420 4950.730 ;
        RECT 3367.760 4950.410 3368.020 4950.730 ;
        RECT 211.760 4790.590 211.900 4950.410 ;
        RECT 3367.820 4823.910 3367.960 4950.410 ;
        RECT 3367.760 4823.590 3368.020 4823.910 ;
        RECT 3376.960 4823.590 3377.220 4823.910 ;
        RECT 208.940 4790.270 209.200 4790.590 ;
        RECT 211.700 4790.270 211.960 4790.590 ;
        RECT 209.000 4787.945 209.140 4790.270 ;
        RECT 208.565 4787.665 210.965 4787.945 ;
        RECT 3367.820 4372.730 3367.960 4823.590 ;
        RECT 3377.020 4821.335 3377.160 4823.590 ;
        RECT 3377.020 4821.195 3379.435 4821.335 ;
        RECT 3377.035 4821.055 3379.435 4821.195 ;
        RECT 3377.035 4375.195 3379.435 4375.335 ;
        RECT 3377.020 4375.055 3379.435 4375.195 ;
        RECT 3377.020 4372.730 3377.160 4375.055 ;
        RECT 3367.760 4372.410 3368.020 4372.730 ;
        RECT 3376.960 4372.410 3377.220 4372.730 ;
        RECT 208.565 3938.665 210.965 3938.945 ;
        RECT 209.000 3936.510 209.140 3938.665 ;
        RECT 208.940 3936.190 209.200 3936.510 ;
        RECT 213.080 3936.190 213.340 3936.510 ;
        RECT 208.565 3722.665 210.965 3722.945 ;
        RECT 209.000 3720.950 209.140 3722.665 ;
        RECT 213.140 3720.950 213.280 3936.190 ;
        RECT 3367.820 3932.090 3367.960 4372.410 ;
        RECT 3367.760 3931.770 3368.020 3932.090 ;
        RECT 3376.960 3931.770 3377.220 3932.090 ;
        RECT 208.940 3720.630 209.200 3720.950 ;
        RECT 211.700 3720.630 211.960 3720.950 ;
        RECT 213.080 3720.630 213.340 3720.950 ;
        RECT 211.760 3698.170 211.900 3720.630 ;
        RECT 3367.820 3703.610 3367.960 3931.770 ;
        RECT 3377.020 3929.335 3377.160 3931.770 ;
        RECT 3377.020 3929.195 3379.435 3929.335 ;
        RECT 3377.035 3929.055 3379.435 3929.195 ;
        RECT 3377.035 3704.300 3379.435 3704.335 ;
        RECT 3377.020 3704.055 3379.435 3704.300 ;
        RECT 3377.020 3703.610 3377.160 3704.055 ;
        RECT 3367.760 3703.290 3368.020 3703.610 ;
        RECT 3376.960 3703.290 3377.220 3703.610 ;
        RECT 211.700 3697.850 211.960 3698.170 ;
        RECT 213.080 3697.850 213.340 3698.170 ;
        RECT 208.565 3506.665 210.965 3506.945 ;
        RECT 209.000 3505.050 209.140 3506.665 ;
        RECT 213.140 3505.050 213.280 3697.850 ;
        RECT 208.940 3504.730 209.200 3505.050 ;
        RECT 213.080 3504.730 213.340 3505.050 ;
        RECT 213.140 3392.850 213.280 3504.730 ;
        RECT 3367.820 3476.830 3367.960 3703.290 ;
        RECT 3377.035 3479.220 3379.435 3479.335 ;
        RECT 3377.020 3479.055 3379.435 3479.220 ;
        RECT 3377.020 3476.830 3377.160 3479.055 ;
        RECT 3367.760 3476.510 3368.020 3476.830 ;
        RECT 3376.960 3476.510 3377.220 3476.830 ;
        RECT 213.080 3392.530 213.340 3392.850 ;
        RECT 214.920 3392.530 215.180 3392.850 ;
        RECT 214.980 3380.950 215.120 3392.530 ;
        RECT 212.160 3380.630 212.420 3380.950 ;
        RECT 214.920 3380.630 215.180 3380.950 ;
        RECT 212.220 3293.570 212.360 3380.630 ;
        RECT 208.940 3293.250 209.200 3293.570 ;
        RECT 212.160 3293.250 212.420 3293.570 ;
        RECT 213.540 3293.250 213.800 3293.570 ;
        RECT 209.000 3290.945 209.140 3293.250 ;
        RECT 208.565 3290.665 210.965 3290.945 ;
        RECT 213.600 3160.290 213.740 3293.250 ;
        RECT 3367.820 3255.830 3367.960 3476.510 ;
        RECT 3367.760 3255.510 3368.020 3255.830 ;
        RECT 3376.960 3255.510 3377.220 3255.830 ;
        RECT 213.540 3159.970 213.800 3160.290 ;
        RECT 214.920 3159.970 215.180 3160.290 ;
        RECT 214.980 3077.670 215.120 3159.970 ;
        RECT 208.940 3077.350 209.200 3077.670 ;
        RECT 214.920 3077.350 215.180 3077.670 ;
        RECT 209.000 3074.945 209.140 3077.350 ;
        RECT 208.565 3074.665 210.965 3074.945 ;
        RECT 214.980 3063.810 215.120 3077.350 ;
        RECT 213.600 3063.670 215.120 3063.810 ;
        RECT 208.565 2858.665 210.965 2858.945 ;
        RECT 209.000 2856.330 209.140 2858.665 ;
        RECT 213.600 2856.410 213.740 3063.670 ;
        RECT 3367.820 3031.090 3367.960 3255.510 ;
        RECT 3377.020 3253.335 3377.160 3255.510 ;
        RECT 3377.020 3253.195 3379.435 3253.335 ;
        RECT 3377.035 3253.055 3379.435 3253.195 ;
        RECT 3367.760 3030.770 3368.020 3031.090 ;
        RECT 3375.120 3030.770 3375.380 3031.090 ;
        RECT 3376.960 3030.770 3377.220 3031.090 ;
        RECT 3375.180 2973.970 3375.320 3030.770 ;
        RECT 3377.020 3028.335 3377.160 3030.770 ;
        RECT 3377.020 3028.195 3379.435 3028.335 ;
        RECT 3377.035 3028.055 3379.435 3028.195 ;
        RECT 3368.680 2973.650 3368.940 2973.970 ;
        RECT 3375.120 2973.650 3375.380 2973.970 ;
        RECT 3368.740 2877.410 3368.880 2973.650 ;
        RECT 3368.680 2877.090 3368.940 2877.410 ;
        RECT 3371.900 2877.090 3372.160 2877.410 ;
        RECT 213.600 2856.330 214.200 2856.410 ;
        RECT 208.940 2856.010 209.200 2856.330 ;
        RECT 213.600 2856.270 214.260 2856.330 ;
        RECT 214.000 2856.010 214.260 2856.270 ;
        RECT 214.060 2774.050 214.200 2856.010 ;
        RECT 3371.960 2799.890 3372.100 2877.090 ;
        RECT 3377.035 2802.195 3379.435 2802.335 ;
        RECT 3377.020 2802.055 3379.435 2802.195 ;
        RECT 3377.020 2799.890 3377.160 2802.055 ;
        RECT 3370.060 2799.570 3370.320 2799.890 ;
        RECT 3371.900 2799.570 3372.160 2799.890 ;
        RECT 3376.960 2799.570 3377.220 2799.890 ;
        RECT 213.080 2773.730 213.340 2774.050 ;
        RECT 214.000 2773.730 214.260 2774.050 ;
        RECT 208.565 2642.665 210.965 2642.945 ;
        RECT 209.000 2640.430 209.140 2642.665 ;
        RECT 213.140 2640.430 213.280 2773.730 ;
        RECT 208.940 2640.110 209.200 2640.430 ;
        RECT 213.080 2640.110 213.340 2640.430 ;
        RECT 213.140 2221.890 213.280 2640.110 ;
        RECT 3370.120 2608.325 3370.260 2799.570 ;
        RECT 3368.670 2607.955 3368.950 2608.325 ;
        RECT 3370.050 2607.955 3370.330 2608.325 ;
        RECT 3368.740 2511.910 3368.880 2607.955 ;
        RECT 3368.680 2511.590 3368.940 2511.910 ;
        RECT 3369.600 2511.590 3369.860 2511.910 ;
        RECT 3369.660 2442.290 3369.800 2511.590 ;
        RECT 3369.200 2442.150 3369.800 2442.290 ;
        RECT 3369.200 2346.670 3369.340 2442.150 ;
        RECT 3369.140 2346.350 3369.400 2346.670 ;
        RECT 3368.680 2345.670 3368.940 2345.990 ;
        RECT 3368.740 2318.450 3368.880 2345.670 ;
        RECT 3368.680 2318.130 3368.940 2318.450 ;
        RECT 3370.060 2318.130 3370.320 2318.450 ;
        RECT 3370.120 2221.890 3370.260 2318.130 ;
        RECT 213.080 2221.570 213.340 2221.890 ;
        RECT 214.000 2221.570 214.260 2221.890 ;
        RECT 3368.680 2221.570 3368.940 2221.890 ;
        RECT 3370.060 2221.570 3370.320 2221.890 ;
        RECT 214.060 2207.950 214.200 2221.570 ;
        RECT 213.540 2207.630 213.800 2207.950 ;
        RECT 214.000 2207.630 214.260 2207.950 ;
        RECT 213.600 2111.730 213.740 2207.630 ;
        RECT 213.080 2111.410 213.340 2111.730 ;
        RECT 213.540 2111.410 213.800 2111.730 ;
        RECT 213.140 2028.770 213.280 2111.410 ;
        RECT 3368.740 2105.010 3368.880 2221.570 ;
        RECT 3368.280 2104.870 3368.880 2105.010 ;
        RECT 3368.280 2103.910 3368.420 2104.870 ;
        RECT 3368.220 2103.590 3368.480 2103.910 ;
        RECT 3369.140 2103.590 3369.400 2103.910 ;
        RECT 213.080 2028.450 213.340 2028.770 ;
        RECT 214.460 2028.450 214.720 2028.770 ;
        RECT 214.520 2007.010 214.660 2028.450 ;
        RECT 3369.200 2008.030 3369.340 2103.590 ;
        RECT 3369.140 2007.710 3369.400 2008.030 ;
        RECT 3376.500 2007.710 3376.760 2008.030 ;
        RECT 208.940 2006.690 209.200 2007.010 ;
        RECT 214.460 2006.690 214.720 2007.010 ;
        RECT 209.000 2004.945 209.140 2006.690 ;
        RECT 214.520 2006.410 214.660 2006.690 ;
        RECT 214.520 2006.270 215.120 2006.410 ;
        RECT 208.565 2004.665 210.965 2004.945 ;
        RECT 214.980 1863.190 215.120 2006.270 ;
        RECT 3376.560 1916.265 3376.700 2007.710 ;
        RECT 3377.035 1916.265 3379.435 1916.335 ;
        RECT 3376.560 1916.230 3379.435 1916.265 ;
        RECT 3368.220 1915.910 3368.480 1916.230 ;
        RECT 3376.500 1916.125 3379.435 1916.230 ;
        RECT 3376.500 1915.910 3376.760 1916.125 ;
        RECT 3377.035 1916.055 3379.435 1916.125 ;
        RECT 214.000 1862.870 214.260 1863.190 ;
        RECT 214.920 1862.870 215.180 1863.190 ;
        RECT 214.060 1839.390 214.200 1862.870 ;
        RECT 212.620 1839.070 212.880 1839.390 ;
        RECT 214.000 1839.070 214.260 1839.390 ;
        RECT 212.680 1791.450 212.820 1839.070 ;
        RECT 208.940 1791.130 209.200 1791.450 ;
        RECT 212.620 1791.130 212.880 1791.450 ;
        RECT 209.000 1788.945 209.140 1791.130 ;
        RECT 208.565 1788.665 210.965 1788.945 ;
        RECT 208.565 1572.665 210.965 1572.945 ;
        RECT 209.000 1570.450 209.140 1572.665 ;
        RECT 212.680 1570.450 212.820 1791.130 ;
        RECT 3368.280 1687.750 3368.420 1915.910 ;
        RECT 3376.560 1915.710 3376.700 1915.910 ;
        RECT 3377.035 1690.140 3379.435 1690.335 ;
        RECT 3377.020 1690.055 3379.435 1690.140 ;
        RECT 3377.020 1687.750 3377.160 1690.055 ;
        RECT 3368.220 1687.430 3368.480 1687.750 ;
        RECT 3376.960 1687.430 3377.220 1687.750 ;
        RECT 208.940 1570.130 209.200 1570.450 ;
        RECT 212.620 1570.130 212.880 1570.450 ;
        RECT 213.540 1570.130 213.800 1570.450 ;
        RECT 213.600 1359.650 213.740 1570.130 ;
        RECT 3368.280 1468.110 3368.420 1687.430 ;
        RECT 3368.220 1467.790 3368.480 1468.110 ;
        RECT 3369.600 1467.790 3369.860 1468.110 ;
        RECT 3376.960 1467.790 3377.220 1468.110 ;
        RECT 208.940 1359.330 209.200 1359.650 ;
        RECT 213.540 1359.330 213.800 1359.650 ;
        RECT 209.000 1356.945 209.140 1359.330 ;
        RECT 208.565 1356.665 210.965 1356.945 ;
        RECT 213.600 1143.410 213.740 1359.330 ;
        RECT 3369.660 1237.590 3369.800 1467.790 ;
        RECT 3377.020 1465.335 3377.160 1467.790 ;
        RECT 3377.020 1465.060 3379.435 1465.335 ;
        RECT 3377.035 1465.055 3379.435 1465.060 ;
        RECT 3377.035 1240.195 3379.435 1240.335 ;
        RECT 3377.020 1240.055 3379.435 1240.195 ;
        RECT 3377.020 1237.590 3377.160 1240.055 ;
        RECT 3368.220 1237.270 3368.480 1237.590 ;
        RECT 3369.600 1237.270 3369.860 1237.590 ;
        RECT 3376.960 1237.270 3377.220 1237.590 ;
        RECT 208.940 1143.090 209.200 1143.410 ;
        RECT 213.540 1143.090 213.800 1143.410 ;
        RECT 209.000 1140.945 209.140 1143.090 ;
        RECT 208.565 1140.665 210.965 1140.945 ;
        RECT 213.600 927.510 213.740 1143.090 ;
        RECT 3368.280 1016.930 3368.420 1237.270 ;
        RECT 3368.220 1016.610 3368.480 1016.930 ;
        RECT 3376.960 1016.610 3377.220 1016.930 ;
        RECT 3368.280 1016.330 3368.420 1016.610 ;
        RECT 3367.360 1016.190 3368.420 1016.330 ;
        RECT 208.940 927.190 209.200 927.510 ;
        RECT 211.700 927.190 211.960 927.510 ;
        RECT 213.540 927.190 213.800 927.510 ;
        RECT 209.000 924.945 209.140 927.190 ;
        RECT 208.565 924.665 210.965 924.945 ;
        RECT 211.760 228.810 211.900 927.190 ;
        RECT 3367.360 786.750 3367.500 1016.190 ;
        RECT 3377.020 1014.335 3377.160 1016.610 ;
        RECT 3377.020 1014.220 3379.435 1014.335 ;
        RECT 3377.035 1014.055 3379.435 1014.220 ;
        RECT 3377.035 789.140 3379.435 789.335 ;
        RECT 3377.020 789.055 3379.435 789.140 ;
        RECT 3377.020 786.750 3377.160 789.055 ;
        RECT 3367.300 786.430 3367.560 786.750 ;
        RECT 3376.960 786.430 3377.220 786.750 ;
        RECT 3367.360 560.650 3367.500 786.430 ;
        RECT 3377.035 563.195 3379.435 563.335 ;
        RECT 3377.020 563.055 3379.435 563.195 ;
        RECT 3377.020 560.650 3377.160 563.055 ;
        RECT 3367.300 560.330 3367.560 560.650 ;
        RECT 3376.960 560.330 3377.220 560.650 ;
        RECT 211.700 228.490 211.960 228.810 ;
        RECT 704.820 228.490 705.080 228.810 ;
        RECT 704.880 201.010 705.020 228.490 ;
        RECT 3367.360 213.850 3367.500 560.330 ;
        RECT 2883.840 213.530 2884.100 213.850 ;
        RECT 3367.300 213.530 3367.560 213.850 ;
        RECT 2883.900 210.110 2884.040 213.530 ;
        RECT 731.500 209.790 731.760 210.110 ;
        RECT 2845.660 209.790 2845.920 210.110 ;
        RECT 2883.840 209.790 2884.100 210.110 ;
        RECT 731.560 203.990 731.700 209.790 ;
        RECT 723.220 203.670 723.480 203.990 ;
        RECT 731.500 203.670 731.760 203.990 ;
        RECT 704.880 200.870 705.180 201.010 ;
        RECT 705.040 200.590 705.180 200.870 ;
        RECT 715.390 200.755 715.670 201.125 ;
        RECT 715.460 200.590 715.600 200.755 ;
        RECT 723.280 200.590 723.420 203.670 ;
        RECT 2845.720 201.125 2845.860 209.790 ;
        RECT 2845.650 200.755 2845.930 201.125 ;
        RECT 704.980 200.270 705.240 200.590 ;
        RECT 715.400 200.270 715.660 200.590 ;
        RECT 723.220 200.270 723.480 200.590 ;
        RECT 705.040 200.000 705.180 200.270 ;
        RECT 715.460 200.000 715.600 200.270 ;
        RECT 723.280 200.000 723.420 200.270 ;
        RECT 704.980 199.360 705.240 200.000 ;
        RECT 715.340 195.755 715.640 200.000 ;
        RECT 722.865 199.015 723.445 200.000 ;
        RECT 722.755 196.425 727.320 196.565 ;
        RECT 722.755 196.355 727.650 196.425 ;
        RECT 722.755 196.305 727.180 196.355 ;
        RECT 722.755 196.205 723.115 196.305 ;
        RECT 723.125 196.205 723.225 196.305 ;
        RECT 727.070 196.235 727.305 196.305 ;
        RECT 727.320 196.235 727.650 196.355 ;
        RECT 722.485 196.165 722.755 196.205 ;
        RECT 722.855 196.165 723.125 196.205 ;
        RECT 722.485 196.025 723.125 196.165 ;
        RECT 727.070 196.095 727.650 196.235 ;
        RECT 727.070 196.070 727.305 196.095 ;
        RECT 722.485 195.935 722.755 196.025 ;
        RECT 722.855 195.935 723.125 196.025 ;
        RECT 715.340 195.740 715.940 195.755 ;
        RECT 715.055 195.455 715.940 195.740 ;
        RECT 722.115 195.565 722.855 195.935 ;
        RECT 722.005 195.455 722.485 195.565 ;
        RECT 708.880 195.315 722.485 195.455 ;
        RECT 708.880 195.245 709.235 195.315 ;
        RECT 715.340 195.245 715.640 195.315 ;
        RECT 722.115 195.245 722.485 195.315 ;
        RECT 708.880 195.195 722.485 195.245 ;
        RECT 708.880 195.100 709.235 195.195 ;
        RECT 709.250 195.100 709.345 195.195 ;
        RECT 708.550 195.055 708.880 195.100 ;
        RECT 708.920 195.055 709.250 195.100 ;
        RECT 708.550 194.845 709.250 195.055 ;
        RECT 708.550 194.770 708.880 194.845 ;
        RECT 708.920 194.770 709.250 194.845 ;
        RECT 708.420 194.640 708.550 194.770 ;
        RECT 708.680 194.640 708.920 194.770 ;
        RECT 708.420 194.530 708.920 194.640 ;
        RECT 708.420 189.025 708.680 194.530 ;
        RECT 708.230 188.915 708.680 189.025 ;
        RECT 708.230 188.835 708.420 188.915 ;
        RECT 708.600 188.835 708.680 188.915 ;
        RECT 707.970 188.465 708.600 188.835 ;
        RECT 707.970 184.355 708.230 188.465 ;
        RECT 707.635 184.105 708.230 184.355 ;
        RECT 707.635 184.020 707.970 184.105 ;
        RECT 708.005 184.020 708.230 184.105 ;
        RECT 707.375 183.650 708.005 184.020 ;
        RECT 707.375 179.505 707.635 183.650 ;
      LAYER via2 ;
        RECT 1710.820 4987.070 1711.120 4987.370 ;
        RECT 606.370 4951.960 606.650 4952.240 ;
        RECT 655.130 4951.960 655.410 4952.240 ;
        RECT 3368.670 2608.000 3368.950 2608.280 ;
        RECT 3370.050 2608.000 3370.330 2608.280 ;
        RECT 715.390 200.800 715.670 201.080 ;
        RECT 2845.650 200.800 2845.930 201.080 ;
      LAYER met3 ;
        RECT 1717.390 4988.000 1741.290 5013.850 ;
        RECT 1710.795 4987.390 1711.145 4987.395 ;
        RECT 1717.950 4987.390 1718.250 4988.000 ;
        RECT 1710.795 4987.090 1718.250 4987.390 ;
        RECT 1710.795 4987.045 1711.145 4987.090 ;
        RECT 606.345 4952.250 606.675 4952.265 ;
        RECT 655.105 4952.250 655.435 4952.265 ;
        RECT 606.345 4951.950 655.435 4952.250 ;
        RECT 606.345 4951.935 606.675 4951.950 ;
        RECT 655.105 4951.935 655.435 4951.950 ;
        RECT 3368.645 2608.290 3368.975 2608.305 ;
        RECT 3370.025 2608.290 3370.355 2608.305 ;
        RECT 3368.645 2607.990 3370.355 2608.290 ;
        RECT 3368.645 2607.975 3368.975 2607.990 ;
        RECT 3370.025 2607.975 3370.355 2607.990 ;
        RECT 715.365 201.090 715.695 201.105 ;
        RECT 2845.625 201.090 2845.955 201.105 ;
        RECT 715.365 200.790 717.290 201.090 ;
        RECT 715.365 200.775 715.695 200.790 ;
        RECT 716.990 200.000 717.290 200.790 ;
        RECT 2845.625 200.775 2846.170 201.090 ;
        RECT 2845.870 200.000 2846.170 200.775 ;
        RECT 716.775 193.330 717.925 200.000 ;
        RECT 715.310 192.100 717.925 193.330 ;
        RECT 715.310 191.865 716.775 192.100 ;
        RECT 716.940 191.865 717.925 192.100 ;
        RECT 716.660 191.585 716.940 191.865 ;
        RECT 2845.710 174.150 2869.610 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 1674.050 5093.120 1734.890 5153.945 ;
    END
  END vssio
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1667.000 5163.785 1668.270 5188.000 ;
    END
  END vssio
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1740.730 5163.785 1742.000 5188.000 ;
    END
  END vssio
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1740.730 5013.835 1920.270 5018.485 ;
    END
  END vssio
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1488.730 5013.935 1668.270 5018.385 ;
    END
  END vssio
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1740.730 5013.935 1920.270 5018.385 ;
    END
  END vssio
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1667.495 4988.000 1691.395 5013.850 ;
    END
  END vssio
  PIN mprj_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 506.200 3555.010 568.800 ;
    END
  END mprj_io[0]
  PIN mprj_io_analog_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 529.015 3379.435 529.295 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_pol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 535.455 3379.435 535.735 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 550.635 3379.435 550.915 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_dm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 532.235 3379.435 532.515 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 523.035 3379.435 523.315 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 553.855 3379.435 554.135 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_enh[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 544.655 3379.435 544.935 ;
    END
  END mprj_io_enh[0]
  PIN mprj_io_hldh_n[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 547.875 3379.435 548.155 ;
    END
  END mprj_io_hldh_n[0]
  PIN mprj_io_holdover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 557.075 3379.435 557.355 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 572.255 3379.435 572.535 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 538.215 3379.435 538.495 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 575.475 3379.435 575.755 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 559.835 3379.435 560.115 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_slow_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 513.835 3379.435 514.115 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 569.035 3379.435 569.315 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 504.635 3379.435 504.915 ;
    END
  END mprj_io_in[0]
  PIN mprj_analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3433.055 3379.435 3433.335 ;
    END
  END mprj_analog_io[3]
  PIN mprj_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3422.200 3555.010 3484.800 ;
    END
  END mprj_io[10]
  PIN mprj_io_analog_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3445.015 3379.435 3445.295 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_pol[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3451.455 3379.435 3451.735 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3466.635 3379.435 3466.915 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_dm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3448.235 3379.435 3448.515 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3439.035 3379.435 3439.315 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3469.855 3379.435 3470.135 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_enh[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3460.655 3379.435 3460.935 ;
    END
  END mprj_io_enh[10]
  PIN mprj_io_hldh_n[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3463.875 3379.435 3464.155 ;
    END
  END mprj_io_hldh_n[10]
  PIN mprj_io_holdover[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3473.075 3379.435 3473.355 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3488.255 3379.435 3488.535 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_inp_dis[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3454.215 3379.435 3454.495 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3491.475 3379.435 3491.755 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3475.835 3379.435 3476.115 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_slow_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3429.835 3379.435 3430.115 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3485.035 3379.435 3485.315 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3420.635 3379.435 3420.915 ;
    END
  END mprj_io_in[10]
  PIN mprj_analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3658.055 3379.435 3658.335 ;
    END
  END mprj_analog_io[4]
  PIN mprj_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3647.200 3555.010 3709.800 ;
    END
  END mprj_io[11]
  PIN mprj_io_analog_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3670.015 3379.435 3670.295 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_pol[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3676.455 3379.435 3676.735 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3691.635 3379.435 3691.915 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_dm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3673.235 3379.435 3673.515 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3664.035 3379.435 3664.315 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3694.855 3379.435 3695.135 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_enh[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3685.655 3379.435 3685.935 ;
    END
  END mprj_io_enh[11]
  PIN mprj_io_hldh_n[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3688.875 3379.435 3689.155 ;
    END
  END mprj_io_hldh_n[11]
  PIN mprj_io_holdover[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3698.075 3379.435 3698.355 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3713.255 3379.435 3713.535 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_inp_dis[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3679.215 3379.435 3679.495 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3716.475 3379.435 3716.755 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3700.835 3379.435 3701.115 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_slow_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3654.835 3379.435 3655.115 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3710.035 3379.435 3710.315 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3645.635 3379.435 3645.915 ;
    END
  END mprj_io_in[11]
  PIN mprj_analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3883.055 3379.435 3883.335 ;
    END
  END mprj_analog_io[5]
  PIN mprj_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3872.200 3555.010 3934.800 ;
    END
  END mprj_io[12]
  PIN mprj_io_analog_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3895.015 3379.435 3895.295 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_pol[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3901.455 3379.435 3901.735 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3916.635 3379.435 3916.915 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_dm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3898.235 3379.435 3898.515 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3889.035 3379.435 3889.315 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3919.855 3379.435 3920.135 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_enh[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3910.655 3379.435 3910.935 ;
    END
  END mprj_io_enh[12]
  PIN mprj_io_hldh_n[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3913.875 3379.435 3914.155 ;
    END
  END mprj_io_hldh_n[12]
  PIN mprj_io_holdover[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3923.075 3379.435 3923.355 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3938.255 3379.435 3938.535 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_inp_dis[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3904.215 3379.435 3904.495 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3941.475 3379.435 3941.755 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3925.835 3379.435 3926.115 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_slow_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3879.835 3379.435 3880.115 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3935.035 3379.435 3935.315 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3870.635 3379.435 3870.915 ;
    END
  END mprj_io_in[12]
  PIN mprj_analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4329.055 3379.435 4329.335 ;
    END
  END mprj_analog_io[6]
  PIN mprj_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4318.200 3555.010 4380.800 ;
    END
  END mprj_io[13]
  PIN mprj_io_analog_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4341.015 3379.435 4341.295 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_pol[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4347.455 3379.435 4347.735 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4362.635 3379.435 4362.915 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_dm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4344.235 3379.435 4344.515 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4335.035 3379.435 4335.315 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4365.855 3379.435 4366.135 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_enh[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4356.655 3379.435 4356.935 ;
    END
  END mprj_io_enh[13]
  PIN mprj_io_hldh_n[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4359.875 3379.435 4360.155 ;
    END
  END mprj_io_hldh_n[13]
  PIN mprj_io_holdover[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4369.075 3379.435 4369.355 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4384.255 3379.435 4384.535 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_inp_dis[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4350.215 3379.435 4350.495 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4387.475 3379.435 4387.755 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4371.835 3379.435 4372.115 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_slow_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4325.835 3379.435 4326.115 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4381.035 3379.435 4381.315 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4316.635 3379.435 4316.915 ;
    END
  END mprj_io_in[13]
  PIN mprj_analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4775.055 3379.435 4775.335 ;
    END
  END mprj_analog_io[7]
  PIN mprj_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4764.200 3555.010 4826.800 ;
    END
  END mprj_io[14]
  PIN mprj_io_analog_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4787.015 3379.435 4787.295 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_pol[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4793.455 3379.435 4793.735 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4808.635 3379.435 4808.915 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_dm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4790.235 3379.435 4790.515 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4781.035 3379.435 4781.315 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4811.855 3379.435 4812.135 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_enh[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4802.655 3379.435 4802.935 ;
    END
  END mprj_io_enh[14]
  PIN mprj_io_hldh_n[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4805.875 3379.435 4806.155 ;
    END
  END mprj_io_hldh_n[14]
  PIN mprj_io_holdover[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4815.075 3379.435 4815.355 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4830.255 3379.435 4830.535 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_inp_dis[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4796.215 3379.435 4796.495 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4833.475 3379.435 4833.755 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4817.835 3379.435 4818.115 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_slow_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4771.835 3379.435 4772.115 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4827.035 3379.435 4827.315 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4762.635 3379.435 4762.915 ;
    END
  END mprj_io_in[14]
  PIN mprj_analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3192.665 4977.035 3192.945 4979.435 ;
    END
  END mprj_analog_io[8]
  PIN mprj_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3141.200 5092.560 3203.800 5155.010 ;
    END
  END mprj_io[15]
  PIN mprj_io_analog_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3180.705 4977.035 3180.985 4979.435 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_pol[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3174.265 4977.035 3174.545 4979.435 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3159.085 4977.035 3159.365 4979.435 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_dm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3177.485 4977.035 3177.765 4979.435 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3186.685 4977.035 3186.965 4979.435 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3155.865 4977.035 3156.145 4979.435 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_enh[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3165.065 4977.035 3165.345 4979.435 ;
    END
  END mprj_io_enh[15]
  PIN mprj_io_hldh_n[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3161.845 4977.035 3162.125 4979.435 ;
    END
  END mprj_io_hldh_n[15]
  PIN mprj_io_holdover[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3152.645 4977.035 3152.925 4979.435 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3137.465 4977.035 3137.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_inp_dis[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3171.505 4977.035 3171.785 4979.435 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3134.245 4977.035 3134.525 4979.435 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3149.885 4977.035 3150.165 4979.435 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_slow_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3195.885 4977.035 3196.165 4979.435 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3140.685 4977.035 3140.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3205.085 4977.035 3205.365 4979.435 ;
    END
  END mprj_io_in[15]
  PIN mprj_analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2683.665 4977.035 2683.945 4979.435 ;
    END
  END mprj_analog_io[9]
  PIN mprj_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2632.200 5092.560 2694.800 5155.010 ;
    END
  END mprj_io[16]
  PIN mprj_io_analog_en[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.705 4977.035 2671.985 4979.435 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_pol[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.265 4977.035 2665.545 4979.435 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.085 4977.035 2650.365 4979.435 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_dm[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.485 4977.035 2668.765 4979.435 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2677.685 4977.035 2677.965 4979.435 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.865 4977.035 2647.145 4979.435 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_enh[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.065 4977.035 2656.345 4979.435 ;
    END
  END mprj_io_enh[16]
  PIN mprj_io_hldh_n[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2652.845 4977.035 2653.125 4979.435 ;
    END
  END mprj_io_hldh_n[16]
  PIN mprj_io_holdover[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.645 4977.035 2643.925 4979.435 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2628.465 4977.035 2628.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_inp_dis[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.505 4977.035 2662.785 4979.435 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.245 4977.035 2625.525 4979.435 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2640.885 4977.035 2641.165 4979.435 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_slow_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2686.885 4977.035 2687.165 4979.435 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.685 4977.035 2631.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.085 4977.035 2696.365 4979.435 ;
    END
  END mprj_io_in[16]
  PIN mprj_analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2426.665 4977.035 2426.945 4979.435 ;
    END
  END mprj_analog_io[10]
  PIN mprj_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2375.200 5092.560 2437.800 5155.010 ;
    END
  END mprj_io[17]
  PIN mprj_io_analog_en[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.705 4977.035 2414.985 4979.435 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_pol[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.265 4977.035 2408.545 4979.435 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.085 4977.035 2393.365 4979.435 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_dm[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.485 4977.035 2411.765 4979.435 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.685 4977.035 2420.965 4979.435 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.865 4977.035 2390.145 4979.435 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_enh[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.065 4977.035 2399.345 4979.435 ;
    END
  END mprj_io_enh[17]
  PIN mprj_io_hldh_n[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.845 4977.035 2396.125 4979.435 ;
    END
  END mprj_io_hldh_n[17]
  PIN mprj_io_holdover[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.645 4977.035 2386.925 4979.435 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2371.465 4977.035 2371.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_inp_dis[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.505 4977.035 2405.785 4979.435 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.245 4977.035 2368.525 4979.435 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2383.885 4977.035 2384.165 4979.435 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_slow_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.885 4977.035 2430.165 4979.435 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.685 4977.035 2374.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.085 4977.035 2439.365 4979.435 ;
    END
  END mprj_io_in[17]
  PIN mprj_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 732.200 3555.010 794.800 ;
    END
  END mprj_io[1]
  PIN mprj_io_analog_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 755.015 3379.435 755.295 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_pol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 761.455 3379.435 761.735 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 776.635 3379.435 776.915 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_dm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 758.235 3379.435 758.515 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 749.035 3379.435 749.315 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 779.855 3379.435 780.135 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_enh[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 770.655 3379.435 770.935 ;
    END
  END mprj_io_enh[1]
  PIN mprj_io_hldh_n[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 773.875 3379.435 774.155 ;
    END
  END mprj_io_hldh_n[1]
  PIN mprj_io_holdover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 783.075 3379.435 783.355 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 798.255 3379.435 798.535 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 764.215 3379.435 764.495 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 801.475 3379.435 801.755 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 785.835 3379.435 786.115 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_slow_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 739.835 3379.435 740.115 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 795.035 3379.435 795.315 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 730.635 3379.435 730.915 ;
    END
  END mprj_io_in[1]
  PIN mprj_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 957.200 3555.010 1019.800 ;
    END
  END mprj_io[2]
  PIN mprj_io_analog_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 980.015 3379.435 980.295 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_pol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 986.455 3379.435 986.735 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1001.635 3379.435 1001.915 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_dm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 983.235 3379.435 983.515 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 974.035 3379.435 974.315 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1004.855 3379.435 1005.135 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_enh[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 995.655 3379.435 995.935 ;
    END
  END mprj_io_enh[2]
  PIN mprj_io_hldh_n[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 998.875 3379.435 999.155 ;
    END
  END mprj_io_hldh_n[2]
  PIN mprj_io_holdover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1008.075 3379.435 1008.355 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1023.255 3379.435 1023.535 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_inp_dis[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 989.215 3379.435 989.495 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1026.475 3379.435 1026.755 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1010.835 3379.435 1011.115 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_slow_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 964.835 3379.435 965.115 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1020.035 3379.435 1020.315 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 955.635 3379.435 955.915 ;
    END
  END mprj_io_in[2]
  PIN mprj_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1183.200 3555.010 1245.800 ;
    END
  END mprj_io[3]
  PIN mprj_io_analog_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1206.015 3379.435 1206.295 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_pol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1212.455 3379.435 1212.735 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1227.635 3379.435 1227.915 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_dm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1200.035 3379.435 1200.315 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1230.855 3379.435 1231.135 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1209.235 3379.435 1209.515 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_enh[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1221.655 3379.435 1221.935 ;
    END
  END mprj_io_enh[3]
  PIN mprj_io_hldh_n[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1224.875 3379.435 1225.155 ;
    END
  END mprj_io_hldh_n[3]
  PIN mprj_io_holdover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1234.075 3379.435 1234.355 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1249.255 3379.435 1249.535 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_inp_dis[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1215.215 3379.435 1215.495 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1252.475 3379.435 1252.755 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1236.835 3379.435 1237.115 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_slow_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1190.835 3379.435 1191.115 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1246.035 3379.435 1246.315 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1181.635 3379.435 1181.915 ;
    END
  END mprj_io_in[3]
  PIN mprj_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1408.200 3555.010 1470.800 ;
    END
  END mprj_io[4]
  PIN mprj_io_analog_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1431.015 3379.435 1431.295 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_pol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1437.455 3379.435 1437.735 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1452.635 3379.435 1452.915 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_dm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1434.235 3379.435 1434.515 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1425.035 3379.435 1425.315 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1455.855 3379.435 1456.135 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_enh[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1446.655 3379.435 1446.935 ;
    END
  END mprj_io_enh[4]
  PIN mprj_io_hldh_n[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1449.875 3379.435 1450.155 ;
    END
  END mprj_io_hldh_n[4]
  PIN mprj_io_holdover[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1459.075 3379.435 1459.355 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1474.255 3379.435 1474.535 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_inp_dis[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1440.215 3379.435 1440.495 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1477.475 3379.435 1477.755 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1461.835 3379.435 1462.115 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_slow_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1415.835 3379.435 1416.115 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1471.035 3379.435 1471.315 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1406.635 3379.435 1406.915 ;
    END
  END mprj_io_in[4]
  PIN mprj_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1633.200 3555.010 1695.800 ;
    END
  END mprj_io[5]
  PIN mprj_io_analog_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1656.015 3379.435 1656.295 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_pol[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1662.455 3379.435 1662.735 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1677.635 3379.435 1677.915 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_dm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1659.235 3379.435 1659.515 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1650.035 3379.435 1650.315 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1680.855 3379.435 1681.135 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_enh[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1671.655 3379.435 1671.935 ;
    END
  END mprj_io_enh[5]
  PIN mprj_io_hldh_n[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1674.875 3379.435 1675.155 ;
    END
  END mprj_io_hldh_n[5]
  PIN mprj_io_holdover[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1684.075 3379.435 1684.355 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1699.255 3379.435 1699.535 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_inp_dis[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1665.215 3379.435 1665.495 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1702.475 3379.435 1702.755 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1686.835 3379.435 1687.115 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_slow_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1640.835 3379.435 1641.115 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1696.035 3379.435 1696.315 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1631.635 3379.435 1631.915 ;
    END
  END mprj_io_in[5]
  PIN mprj_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1859.200 3555.010 1921.800 ;
    END
  END mprj_io[6]
  PIN mprj_io_analog_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1882.015 3379.435 1882.295 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_pol[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1888.455 3379.435 1888.735 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1903.635 3379.435 1903.915 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_dm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1885.235 3379.435 1885.515 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1876.035 3379.435 1876.315 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1906.855 3379.435 1907.135 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_enh[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1897.655 3379.435 1897.935 ;
    END
  END mprj_io_enh[6]
  PIN mprj_io_hldh_n[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1900.875 3379.435 1901.155 ;
    END
  END mprj_io_hldh_n[6]
  PIN mprj_io_holdover[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1910.075 3379.435 1910.355 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1925.255 3379.435 1925.535 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_inp_dis[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1891.215 3379.435 1891.495 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1928.475 3379.435 1928.755 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1912.835 3379.435 1913.115 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_slow_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1866.835 3379.435 1867.115 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1922.035 3379.435 1922.315 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1857.635 3379.435 1857.915 ;
    END
  END mprj_io_in[6]
  PIN mprj_analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2756.055 3379.435 2756.335 ;
    END
  END mprj_analog_io[0]
  PIN mprj_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2745.200 3555.010 2807.800 ;
    END
  END mprj_io[7]
  PIN mprj_io_analog_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2768.015 3379.435 2768.295 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_pol[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2774.455 3379.435 2774.735 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2789.635 3379.435 2789.915 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_dm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2771.235 3379.435 2771.515 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2762.035 3379.435 2762.315 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2792.855 3379.435 2793.135 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_enh[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2783.655 3379.435 2783.935 ;
    END
  END mprj_io_enh[7]
  PIN mprj_io_hldh_n[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2786.875 3379.435 2787.155 ;
    END
  END mprj_io_hldh_n[7]
  PIN mprj_io_holdover[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2796.075 3379.435 2796.355 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2811.255 3379.435 2811.535 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_inp_dis[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2777.215 3379.435 2777.495 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2814.475 3379.435 2814.755 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2798.835 3379.435 2799.115 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_slow_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2752.835 3379.435 2753.115 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2808.035 3379.435 2808.315 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2743.635 3379.435 2743.915 ;
    END
  END mprj_io_in[7]
  PIN mprj_analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2982.055 3379.435 2982.335 ;
    END
  END mprj_analog_io[1]
  PIN mprj_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2971.200 3555.010 3033.800 ;
    END
  END mprj_io[8]
  PIN mprj_io_analog_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2994.015 3379.435 2994.295 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_pol[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3000.455 3379.435 3000.735 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3015.635 3379.435 3015.915 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_dm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2997.235 3379.435 2997.515 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2988.035 3379.435 2988.315 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3018.855 3379.435 3019.135 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_enh[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3009.655 3379.435 3009.935 ;
    END
  END mprj_io_enh[8]
  PIN mprj_io_hldh_n[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3012.875 3379.435 3013.155 ;
    END
  END mprj_io_hldh_n[8]
  PIN mprj_io_holdover[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3022.075 3379.435 3022.355 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3037.255 3379.435 3037.535 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_inp_dis[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3003.215 3379.435 3003.495 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3040.475 3379.435 3040.755 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3024.835 3379.435 3025.115 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_slow_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2978.835 3379.435 2979.115 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3034.035 3379.435 3034.315 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2969.635 3379.435 2969.915 ;
    END
  END mprj_io_in[8]
  PIN mprj_analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3207.055 3379.435 3207.335 ;
    END
  END mprj_analog_io[2]
  PIN mprj_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3196.200 3555.010 3258.800 ;
    END
  END mprj_io[9]
  PIN mprj_io_analog_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3219.015 3379.435 3219.295 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3225.455 3379.435 3225.735 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3240.635 3379.435 3240.915 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3222.235 3379.435 3222.515 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3213.035 3379.435 3213.315 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3243.855 3379.435 3244.135 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_enh[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3234.655 3379.435 3234.935 ;
    END
  END mprj_io_enh[9]
  PIN mprj_io_hldh_n[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3237.875 3379.435 3238.155 ;
    END
  END mprj_io_hldh_n[9]
  PIN mprj_io_holdover[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3247.075 3379.435 3247.355 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3262.255 3379.435 3262.535 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_inp_dis[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3228.215 3379.435 3228.495 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3265.475 3379.435 3265.755 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3249.835 3379.435 3250.115 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3203.835 3379.435 3204.115 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3259.035 3379.435 3259.315 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN mprj_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3194.635 3379.435 3194.915 ;
    END
  END mprj_io_in[9]
  PIN mprj_analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.665 4977.035 1981.945 4979.435 ;
    END
  END mprj_analog_io[11]
  PIN mprj_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1930.200 5092.560 1992.800 5155.010 ;
    END
  END mprj_io[18]
  PIN mprj_io_analog_en[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.705 4977.035 1969.985 4979.435 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_pol[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.265 4977.035 1963.545 4979.435 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.085 4977.035 1948.365 4979.435 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_dm[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.485 4977.035 1966.765 4979.435 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.685 4977.035 1975.965 4979.435 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.865 4977.035 1945.145 4979.435 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_enh[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.065 4977.035 1954.345 4979.435 ;
    END
  END mprj_io_enh[18]
  PIN mprj_io_hldh_n[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.845 4977.035 1951.125 4979.435 ;
    END
  END mprj_io_hldh_n[18]
  PIN mprj_io_holdover[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.645 4977.035 1941.925 4979.435 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.465 4977.035 1926.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_inp_dis[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1960.505 4977.035 1960.785 4979.435 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.245 4977.035 1923.525 4979.435 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.885 4977.035 1939.165 4979.435 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_slow_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.885 4977.035 1985.165 4979.435 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.685 4977.035 1929.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.085 4977.035 1994.365 4979.435 ;
    END
  END mprj_io_in[18]
  PIN mprj_analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3336.665 210.965 3336.945 ;
    END
  END mprj_analog_io[21]
  PIN mprj_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3285.200 95.440 3347.800 ;
    END
  END mprj_io[28]
  PIN mprj_io_analog_en[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3324.705 210.965 3324.985 ;
    END
  END mprj_io_analog_en[28]
  PIN mprj_io_analog_pol[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3318.265 210.965 3318.545 ;
    END
  END mprj_io_analog_pol[28]
  PIN mprj_io_analog_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3303.085 210.965 3303.365 ;
    END
  END mprj_io_analog_sel[28]
  PIN mprj_io_dm[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3321.485 210.965 3321.765 ;
    END
  END mprj_io_dm[84]
  PIN mprj_io_dm[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3330.685 210.965 3330.965 ;
    END
  END mprj_io_dm[85]
  PIN mprj_io_dm[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3299.865 210.965 3300.145 ;
    END
  END mprj_io_dm[86]
  PIN mprj_io_enh[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3309.065 210.965 3309.345 ;
    END
  END mprj_io_enh[28]
  PIN mprj_io_hldh_n[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3305.845 210.965 3306.125 ;
    END
  END mprj_io_hldh_n[28]
  PIN mprj_io_holdover[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3296.645 210.965 3296.925 ;
    END
  END mprj_io_holdover[28]
  PIN mprj_io_ib_mode_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3281.465 210.965 3281.745 ;
    END
  END mprj_io_ib_mode_sel[28]
  PIN mprj_io_inp_dis[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3315.505 210.965 3315.785 ;
    END
  END mprj_io_inp_dis[28]
  PIN mprj_io_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3278.245 210.965 3278.525 ;
    END
  END mprj_io_oeb[28]
  PIN mprj_io_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3293.885 210.965 3294.165 ;
    END
  END mprj_io_out[28]
  PIN mprj_io_slow_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3339.885 210.965 3340.165 ;
    END
  END mprj_io_slow_sel[28]
  PIN mprj_io_vtrip_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3284.685 210.965 3284.965 ;
    END
  END mprj_io_vtrip_sel[28]
  PIN mprj_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3349.085 210.965 3349.365 ;
    END
  END mprj_io_in[28]
  PIN mprj_analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3120.665 210.965 3120.945 ;
    END
  END mprj_analog_io[22]
  PIN mprj_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3069.200 95.440 3131.800 ;
    END
  END mprj_io[29]
  PIN mprj_io_analog_en[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3108.705 210.965 3108.985 ;
    END
  END mprj_io_analog_en[29]
  PIN mprj_io_analog_pol[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3102.265 210.965 3102.545 ;
    END
  END mprj_io_analog_pol[29]
  PIN mprj_io_analog_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3087.085 210.965 3087.365 ;
    END
  END mprj_io_analog_sel[29]
  PIN mprj_io_dm[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3105.485 210.965 3105.765 ;
    END
  END mprj_io_dm[87]
  PIN mprj_io_dm[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3114.685 210.965 3114.965 ;
    END
  END mprj_io_dm[88]
  PIN mprj_io_dm[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3083.865 210.965 3084.145 ;
    END
  END mprj_io_dm[89]
  PIN mprj_io_enh[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3093.065 210.965 3093.345 ;
    END
  END mprj_io_enh[29]
  PIN mprj_io_hldh_n[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3089.845 210.965 3090.125 ;
    END
  END mprj_io_hldh_n[29]
  PIN mprj_io_holdover[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3080.645 210.965 3080.925 ;
    END
  END mprj_io_holdover[29]
  PIN mprj_io_ib_mode_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3065.465 210.965 3065.745 ;
    END
  END mprj_io_ib_mode_sel[29]
  PIN mprj_io_inp_dis[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3099.505 210.965 3099.785 ;
    END
  END mprj_io_inp_dis[29]
  PIN mprj_io_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3062.245 210.965 3062.525 ;
    END
  END mprj_io_oeb[29]
  PIN mprj_io_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3077.885 210.965 3078.165 ;
    END
  END mprj_io_out[29]
  PIN mprj_io_slow_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3123.885 210.965 3124.165 ;
    END
  END mprj_io_slow_sel[29]
  PIN mprj_io_vtrip_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3068.685 210.965 3068.965 ;
    END
  END mprj_io_vtrip_sel[29]
  PIN mprj_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3133.085 210.965 3133.365 ;
    END
  END mprj_io_in[29]
  PIN mprj_analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2904.665 210.965 2904.945 ;
    END
  END mprj_analog_io[23]
  PIN mprj_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2853.200 95.440 2915.800 ;
    END
  END mprj_io[30]
  PIN mprj_io_analog_en[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2892.705 210.965 2892.985 ;
    END
  END mprj_io_analog_en[30]
  PIN mprj_io_analog_pol[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2886.265 210.965 2886.545 ;
    END
  END mprj_io_analog_pol[30]
  PIN mprj_io_analog_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2871.085 210.965 2871.365 ;
    END
  END mprj_io_analog_sel[30]
  PIN mprj_io_dm[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2889.485 210.965 2889.765 ;
    END
  END mprj_io_dm[90]
  PIN mprj_io_dm[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2898.685 210.965 2898.965 ;
    END
  END mprj_io_dm[91]
  PIN mprj_io_dm[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2867.865 210.965 2868.145 ;
    END
  END mprj_io_dm[92]
  PIN mprj_io_enh[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2877.065 210.965 2877.345 ;
    END
  END mprj_io_enh[30]
  PIN mprj_io_hldh_n[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2873.845 210.965 2874.125 ;
    END
  END mprj_io_hldh_n[30]
  PIN mprj_io_holdover[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2864.645 210.965 2864.925 ;
    END
  END mprj_io_holdover[30]
  PIN mprj_io_ib_mode_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2849.465 210.965 2849.745 ;
    END
  END mprj_io_ib_mode_sel[30]
  PIN mprj_io_inp_dis[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2883.505 210.965 2883.785 ;
    END
  END mprj_io_inp_dis[30]
  PIN mprj_io_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2846.245 210.965 2846.525 ;
    END
  END mprj_io_oeb[30]
  PIN mprj_io_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2861.885 210.965 2862.165 ;
    END
  END mprj_io_out[30]
  PIN mprj_io_slow_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2907.885 210.965 2908.165 ;
    END
  END mprj_io_slow_sel[30]
  PIN mprj_io_vtrip_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2852.685 210.965 2852.965 ;
    END
  END mprj_io_vtrip_sel[30]
  PIN mprj_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2917.085 210.965 2917.365 ;
    END
  END mprj_io_in[30]
  PIN mprj_analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2688.665 210.965 2688.945 ;
    END
  END mprj_analog_io[24]
  PIN mprj_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2637.200 95.440 2699.800 ;
    END
  END mprj_io[31]
  PIN mprj_io_analog_en[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2676.705 210.965 2676.985 ;
    END
  END mprj_io_analog_en[31]
  PIN mprj_io_analog_pol[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2670.265 210.965 2670.545 ;
    END
  END mprj_io_analog_pol[31]
  PIN mprj_io_analog_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2655.085 210.965 2655.365 ;
    END
  END mprj_io_analog_sel[31]
  PIN mprj_io_dm[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2673.485 210.965 2673.765 ;
    END
  END mprj_io_dm[93]
  PIN mprj_io_dm[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2682.685 210.965 2682.965 ;
    END
  END mprj_io_dm[94]
  PIN mprj_io_dm[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2651.865 210.965 2652.145 ;
    END
  END mprj_io_dm[95]
  PIN mprj_io_enh[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2661.065 210.965 2661.345 ;
    END
  END mprj_io_enh[31]
  PIN mprj_io_hldh_n[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2657.845 210.965 2658.125 ;
    END
  END mprj_io_hldh_n[31]
  PIN mprj_io_holdover[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2648.645 210.965 2648.925 ;
    END
  END mprj_io_holdover[31]
  PIN mprj_io_ib_mode_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.465 210.965 2633.745 ;
    END
  END mprj_io_ib_mode_sel[31]
  PIN mprj_io_inp_dis[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2667.505 210.965 2667.785 ;
    END
  END mprj_io_inp_dis[31]
  PIN mprj_io_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2630.245 210.965 2630.525 ;
    END
  END mprj_io_oeb[31]
  PIN mprj_io_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2645.885 210.965 2646.165 ;
    END
  END mprj_io_out[31]
  PIN mprj_io_slow_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2691.885 210.965 2692.165 ;
    END
  END mprj_io_slow_sel[31]
  PIN mprj_io_vtrip_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2636.685 210.965 2636.965 ;
    END
  END mprj_io_vtrip_sel[31]
  PIN mprj_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2701.085 210.965 2701.365 ;
    END
  END mprj_io_in[31]
  PIN mprj_analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2050.665 210.965 2050.945 ;
    END
  END mprj_analog_io[25]
  PIN mprj_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1999.200 95.440 2061.800 ;
    END
  END mprj_io[32]
  PIN mprj_io_analog_en[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2038.705 210.965 2038.985 ;
    END
  END mprj_io_analog_en[32]
  PIN mprj_io_analog_pol[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2032.265 210.965 2032.545 ;
    END
  END mprj_io_analog_pol[32]
  PIN mprj_io_analog_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2017.085 210.965 2017.365 ;
    END
  END mprj_io_analog_sel[32]
  PIN mprj_io_dm[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2035.485 210.965 2035.765 ;
    END
  END mprj_io_dm[96]
  PIN mprj_io_dm[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2044.685 210.965 2044.965 ;
    END
  END mprj_io_dm[97]
  PIN mprj_io_dm[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2013.865 210.965 2014.145 ;
    END
  END mprj_io_dm[98]
  PIN mprj_io_enh[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2023.065 210.965 2023.345 ;
    END
  END mprj_io_enh[32]
  PIN mprj_io_hldh_n[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2019.845 210.965 2020.125 ;
    END
  END mprj_io_hldh_n[32]
  PIN mprj_io_holdover[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2010.645 210.965 2010.925 ;
    END
  END mprj_io_holdover[32]
  PIN mprj_io_ib_mode_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1995.465 210.965 1995.745 ;
    END
  END mprj_io_ib_mode_sel[32]
  PIN mprj_io_inp_dis[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2029.505 210.965 2029.785 ;
    END
  END mprj_io_inp_dis[32]
  PIN mprj_io_oeb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1992.245 210.965 1992.525 ;
    END
  END mprj_io_oeb[32]
  PIN mprj_io_out[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2007.885 210.965 2008.165 ;
    END
  END mprj_io_out[32]
  PIN mprj_io_slow_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2053.885 210.965 2054.165 ;
    END
  END mprj_io_slow_sel[32]
  PIN mprj_io_vtrip_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1998.685 210.965 1998.965 ;
    END
  END mprj_io_vtrip_sel[32]
  PIN mprj_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2063.085 210.965 2063.365 ;
    END
  END mprj_io_in[32]
  PIN mprj_analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1834.665 210.965 1834.945 ;
    END
  END mprj_analog_io[26]
  PIN mprj_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1783.200 95.440 1845.800 ;
    END
  END mprj_io[33]
  PIN mprj_io_analog_en[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1822.705 210.965 1822.985 ;
    END
  END mprj_io_analog_en[33]
  PIN mprj_io_analog_pol[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1816.265 210.965 1816.545 ;
    END
  END mprj_io_analog_pol[33]
  PIN mprj_io_analog_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1801.085 210.965 1801.365 ;
    END
  END mprj_io_analog_sel[33]
  PIN mprj_io_dm[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1828.685 210.965 1828.965 ;
    END
  END mprj_io_dm[100]
  PIN mprj_io_dm[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1797.865 210.965 1798.145 ;
    END
  END mprj_io_dm[101]
  PIN mprj_io_dm[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1819.485 210.965 1819.765 ;
    END
  END mprj_io_dm[99]
  PIN mprj_io_enh[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1807.065 210.965 1807.345 ;
    END
  END mprj_io_enh[33]
  PIN mprj_io_hldh_n[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1803.845 210.965 1804.125 ;
    END
  END mprj_io_hldh_n[33]
  PIN mprj_io_holdover[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1794.645 210.965 1794.925 ;
    END
  END mprj_io_holdover[33]
  PIN mprj_io_ib_mode_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1779.465 210.965 1779.745 ;
    END
  END mprj_io_ib_mode_sel[33]
  PIN mprj_io_inp_dis[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1813.505 210.965 1813.785 ;
    END
  END mprj_io_inp_dis[33]
  PIN mprj_io_oeb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1776.245 210.965 1776.525 ;
    END
  END mprj_io_oeb[33]
  PIN mprj_io_out[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1791.885 210.965 1792.165 ;
    END
  END mprj_io_out[33]
  PIN mprj_io_slow_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1837.885 210.965 1838.165 ;
    END
  END mprj_io_slow_sel[33]
  PIN mprj_io_vtrip_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1782.685 210.965 1782.965 ;
    END
  END mprj_io_vtrip_sel[33]
  PIN mprj_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1847.085 210.965 1847.365 ;
    END
  END mprj_io_in[33]
  PIN mprj_analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1618.665 210.965 1618.945 ;
    END
  END mprj_analog_io[27]
  PIN mprj_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1567.200 95.440 1629.800 ;
    END
  END mprj_io[34]
  PIN mprj_io_analog_en[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1606.705 210.965 1606.985 ;
    END
  END mprj_io_analog_en[34]
  PIN mprj_io_analog_pol[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1600.265 210.965 1600.545 ;
    END
  END mprj_io_analog_pol[34]
  PIN mprj_io_analog_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1585.085 210.965 1585.365 ;
    END
  END mprj_io_analog_sel[34]
  PIN mprj_io_dm[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1603.485 210.965 1603.765 ;
    END
  END mprj_io_dm[102]
  PIN mprj_io_dm[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1612.685 210.965 1612.965 ;
    END
  END mprj_io_dm[103]
  PIN mprj_io_dm[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1581.865 210.965 1582.145 ;
    END
  END mprj_io_dm[104]
  PIN mprj_io_enh[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1591.065 210.965 1591.345 ;
    END
  END mprj_io_enh[34]
  PIN mprj_io_hldh_n[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1587.845 210.965 1588.125 ;
    END
  END mprj_io_hldh_n[34]
  PIN mprj_io_holdover[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1578.645 210.965 1578.925 ;
    END
  END mprj_io_holdover[34]
  PIN mprj_io_ib_mode_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1563.465 210.965 1563.745 ;
    END
  END mprj_io_ib_mode_sel[34]
  PIN mprj_io_inp_dis[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1597.505 210.965 1597.785 ;
    END
  END mprj_io_inp_dis[34]
  PIN mprj_io_oeb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1560.245 210.965 1560.525 ;
    END
  END mprj_io_oeb[34]
  PIN mprj_io_out[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1575.885 210.965 1576.165 ;
    END
  END mprj_io_out[34]
  PIN mprj_io_slow_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1621.885 210.965 1622.165 ;
    END
  END mprj_io_slow_sel[34]
  PIN mprj_io_vtrip_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1566.685 210.965 1566.965 ;
    END
  END mprj_io_vtrip_sel[34]
  PIN mprj_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1631.085 210.965 1631.365 ;
    END
  END mprj_io_in[34]
  PIN mprj_analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1402.665 210.965 1402.945 ;
    END
  END mprj_analog_io[28]
  PIN mprj_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1351.200 95.440 1413.800 ;
    END
  END mprj_io[35]
  PIN mprj_io_analog_en[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1390.705 210.965 1390.985 ;
    END
  END mprj_io_analog_en[35]
  PIN mprj_io_analog_pol[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1384.265 210.965 1384.545 ;
    END
  END mprj_io_analog_pol[35]
  PIN mprj_io_analog_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1369.085 210.965 1369.365 ;
    END
  END mprj_io_analog_sel[35]
  PIN mprj_io_dm[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1387.485 210.965 1387.765 ;
    END
  END mprj_io_dm[105]
  PIN mprj_io_dm[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1396.685 210.965 1396.965 ;
    END
  END mprj_io_dm[106]
  PIN mprj_io_dm[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1365.865 210.965 1366.145 ;
    END
  END mprj_io_dm[107]
  PIN mprj_io_enh[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1375.065 210.965 1375.345 ;
    END
  END mprj_io_enh[35]
  PIN mprj_io_hldh_n[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1371.845 210.965 1372.125 ;
    END
  END mprj_io_hldh_n[35]
  PIN mprj_io_holdover[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1362.645 210.965 1362.925 ;
    END
  END mprj_io_holdover[35]
  PIN mprj_io_ib_mode_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1347.465 210.965 1347.745 ;
    END
  END mprj_io_ib_mode_sel[35]
  PIN mprj_io_inp_dis[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1381.505 210.965 1381.785 ;
    END
  END mprj_io_inp_dis[35]
  PIN mprj_io_oeb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1344.245 210.965 1344.525 ;
    END
  END mprj_io_oeb[35]
  PIN mprj_io_out[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1359.885 210.965 1360.165 ;
    END
  END mprj_io_out[35]
  PIN mprj_io_slow_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1405.885 210.965 1406.165 ;
    END
  END mprj_io_slow_sel[35]
  PIN mprj_io_vtrip_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1350.685 210.965 1350.965 ;
    END
  END mprj_io_vtrip_sel[35]
  PIN mprj_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1415.085 210.965 1415.365 ;
    END
  END mprj_io_in[35]
  PIN mprj_analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1186.665 210.965 1186.945 ;
    END
  END mprj_analog_io[29]
  PIN mprj_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1135.200 95.440 1197.800 ;
    END
  END mprj_io[36]
  PIN mprj_io_analog_en[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1174.705 210.965 1174.985 ;
    END
  END mprj_io_analog_en[36]
  PIN mprj_io_analog_pol[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1168.265 210.965 1168.545 ;
    END
  END mprj_io_analog_pol[36]
  PIN mprj_io_analog_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1153.085 210.965 1153.365 ;
    END
  END mprj_io_analog_sel[36]
  PIN mprj_io_dm[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1171.485 210.965 1171.765 ;
    END
  END mprj_io_dm[108]
  PIN mprj_io_dm[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1180.685 210.965 1180.965 ;
    END
  END mprj_io_dm[109]
  PIN mprj_io_dm[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1149.865 210.965 1150.145 ;
    END
  END mprj_io_dm[110]
  PIN mprj_io_enh[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1159.065 210.965 1159.345 ;
    END
  END mprj_io_enh[36]
  PIN mprj_io_hldh_n[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1155.845 210.965 1156.125 ;
    END
  END mprj_io_hldh_n[36]
  PIN mprj_io_holdover[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1146.645 210.965 1146.925 ;
    END
  END mprj_io_holdover[36]
  PIN mprj_io_ib_mode_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1131.465 210.965 1131.745 ;
    END
  END mprj_io_ib_mode_sel[36]
  PIN mprj_io_inp_dis[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1165.505 210.965 1165.785 ;
    END
  END mprj_io_inp_dis[36]
  PIN mprj_io_oeb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1128.245 210.965 1128.525 ;
    END
  END mprj_io_oeb[36]
  PIN mprj_io_out[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1143.885 210.965 1144.165 ;
    END
  END mprj_io_out[36]
  PIN mprj_io_slow_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1189.885 210.965 1190.165 ;
    END
  END mprj_io_slow_sel[36]
  PIN mprj_io_vtrip_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1134.685 210.965 1134.965 ;
    END
  END mprj_io_vtrip_sel[36]
  PIN mprj_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1199.085 210.965 1199.365 ;
    END
  END mprj_io_in[36]
  PIN mprj_analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 970.665 210.965 970.945 ;
    END
  END mprj_analog_io[30]
  PIN mprj_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 919.200 95.440 981.800 ;
    END
  END mprj_io[37]
  PIN mprj_io_analog_en[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 958.705 210.965 958.985 ;
    END
  END mprj_io_analog_en[37]
  PIN mprj_io_analog_pol[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 952.265 210.965 952.545 ;
    END
  END mprj_io_analog_pol[37]
  PIN mprj_io_analog_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 937.085 210.965 937.365 ;
    END
  END mprj_io_analog_sel[37]
  PIN mprj_io_dm[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 955.485 210.965 955.765 ;
    END
  END mprj_io_dm[111]
  PIN mprj_io_dm[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 964.685 210.965 964.965 ;
    END
  END mprj_io_dm[112]
  PIN mprj_io_dm[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 933.865 210.965 934.145 ;
    END
  END mprj_io_dm[113]
  PIN mprj_io_enh[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 943.065 210.965 943.345 ;
    END
  END mprj_io_enh[37]
  PIN mprj_io_hldh_n[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 939.845 210.965 940.125 ;
    END
  END mprj_io_hldh_n[37]
  PIN mprj_io_holdover[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 930.645 210.965 930.925 ;
    END
  END mprj_io_holdover[37]
  PIN mprj_io_ib_mode_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 915.465 210.965 915.745 ;
    END
  END mprj_io_ib_mode_sel[37]
  PIN mprj_io_inp_dis[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 949.505 210.965 949.785 ;
    END
  END mprj_io_inp_dis[37]
  PIN mprj_io_oeb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 912.245 210.965 912.525 ;
    END
  END mprj_io_oeb[37]
  PIN mprj_io_out[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 927.885 210.965 928.165 ;
    END
  END mprj_io_out[37]
  PIN mprj_io_slow_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 973.885 210.965 974.165 ;
    END
  END mprj_io_slow_sel[37]
  PIN mprj_io_vtrip_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 918.685 210.965 918.965 ;
    END
  END mprj_io_vtrip_sel[37]
  PIN mprj_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 983.085 210.965 983.365 ;
    END
  END mprj_io_in[37]
  PIN mprj_analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.665 4977.035 1472.945 4979.435 ;
    END
  END mprj_analog_io[12]
  PIN mprj_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1421.200 5092.560 1483.800 5155.010 ;
    END
  END mprj_io[19]
  PIN mprj_io_analog_en[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.705 4977.035 1460.985 4979.435 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_pol[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.265 4977.035 1454.545 4979.435 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.085 4977.035 1439.365 4979.435 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_dm[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.485 4977.035 1457.765 4979.435 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.685 4977.035 1466.965 4979.435 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.865 4977.035 1436.145 4979.435 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_enh[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.065 4977.035 1445.345 4979.435 ;
    END
  END mprj_io_enh[19]
  PIN mprj_io_hldh_n[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.845 4977.035 1442.125 4979.435 ;
    END
  END mprj_io_hldh_n[19]
  PIN mprj_io_holdover[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.645 4977.035 1432.925 4979.435 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.465 4977.035 1417.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_inp_dis[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.505 4977.035 1451.785 4979.435 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.245 4977.035 1414.525 4979.435 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.885 4977.035 1430.165 4979.435 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_slow_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.885 4977.035 1476.165 4979.435 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.685 4977.035 1420.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.085 4977.035 1485.365 4979.435 ;
    END
  END mprj_io_in[19]
  PIN mprj_analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.665 4977.035 1214.945 4979.435 ;
    END
  END mprj_analog_io[13]
  PIN mprj_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1163.200 5092.560 1225.800 5155.010 ;
    END
  END mprj_io[20]
  PIN mprj_io_analog_en[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.705 4977.035 1202.985 4979.435 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_pol[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.265 4977.035 1196.545 4979.435 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.085 4977.035 1181.365 4979.435 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_dm[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.485 4977.035 1199.765 4979.435 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.685 4977.035 1208.965 4979.435 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.865 4977.035 1178.145 4979.435 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_enh[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.065 4977.035 1187.345 4979.435 ;
    END
  END mprj_io_enh[20]
  PIN mprj_io_hldh_n[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.845 4977.035 1184.125 4979.435 ;
    END
  END mprj_io_hldh_n[20]
  PIN mprj_io_holdover[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.645 4977.035 1174.925 4979.435 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.465 4977.035 1159.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_inp_dis[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.505 4977.035 1193.785 4979.435 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.245 4977.035 1156.525 4979.435 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.885 4977.035 1172.165 4979.435 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_slow_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.885 4977.035 1218.165 4979.435 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.685 4977.035 1162.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.085 4977.035 1227.365 4979.435 ;
    END
  END mprj_io_in[20]
  PIN mprj_analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.665 4977.035 957.945 4979.435 ;
    END
  END mprj_analog_io[14]
  PIN mprj_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 906.200 5092.560 968.800 5155.010 ;
    END
  END mprj_io[21]
  PIN mprj_io_analog_en[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.705 4977.035 945.985 4979.435 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_pol[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.265 4977.035 939.545 4979.435 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.085 4977.035 924.365 4979.435 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_dm[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.485 4977.035 942.765 4979.435 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.685 4977.035 951.965 4979.435 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.865 4977.035 921.145 4979.435 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_enh[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.065 4977.035 930.345 4979.435 ;
    END
  END mprj_io_enh[21]
  PIN mprj_io_hldh_n[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.845 4977.035 927.125 4979.435 ;
    END
  END mprj_io_hldh_n[21]
  PIN mprj_io_holdover[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.645 4977.035 917.925 4979.435 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.465 4977.035 902.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_inp_dis[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.505 4977.035 936.785 4979.435 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.245 4977.035 899.525 4979.435 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.885 4977.035 915.165 4979.435 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_slow_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.885 4977.035 961.165 4979.435 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.685 4977.035 905.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.085 4977.035 970.365 4979.435 ;
    END
  END mprj_io_in[21]
  PIN mprj_analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.665 4977.035 700.945 4979.435 ;
    END
  END mprj_analog_io[15]
  PIN mprj_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 649.200 5092.560 711.800 5155.010 ;
    END
  END mprj_io[22]
  PIN mprj_io_analog_en[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.705 4977.035 688.985 4979.435 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_pol[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.265 4977.035 682.545 4979.435 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.085 4977.035 667.365 4979.435 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_dm[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.485 4977.035 685.765 4979.435 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.685 4977.035 694.965 4979.435 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.865 4977.035 664.145 4979.435 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_enh[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.065 4977.035 673.345 4979.435 ;
    END
  END mprj_io_enh[22]
  PIN mprj_io_hldh_n[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.845 4977.035 670.125 4979.435 ;
    END
  END mprj_io_hldh_n[22]
  PIN mprj_io_holdover[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.645 4977.035 660.925 4979.435 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.465 4977.035 645.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_inp_dis[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.505 4977.035 679.785 4979.435 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.245 4977.035 642.525 4979.435 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.885 4977.035 658.165 4979.435 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_slow_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.885 4977.035 704.165 4979.435 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.685 4977.035 648.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.085 4977.035 713.365 4979.435 ;
    END
  END mprj_io_in[22]
  PIN mprj_analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.665 4977.035 443.945 4979.435 ;
    END
  END mprj_analog_io[16]
  PIN mprj_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 392.200 5092.560 454.800 5155.010 ;
    END
  END mprj_io[23]
  PIN mprj_io_analog_en[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.705 4977.035 431.985 4979.435 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_pol[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.265 4977.035 425.545 4979.435 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.085 4977.035 410.365 4979.435 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_dm[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.485 4977.035 428.765 4979.435 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.685 4977.035 437.965 4979.435 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.865 4977.035 407.145 4979.435 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_enh[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.065 4977.035 416.345 4979.435 ;
    END
  END mprj_io_enh[23]
  PIN mprj_io_hldh_n[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.845 4977.035 413.125 4979.435 ;
    END
  END mprj_io_hldh_n[23]
  PIN mprj_io_holdover[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.645 4977.035 403.925 4979.435 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.465 4977.035 388.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_inp_dis[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.505 4977.035 422.785 4979.435 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.245 4977.035 385.525 4979.435 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.885 4977.035 401.165 4979.435 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_slow_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.885 4977.035 447.165 4979.435 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.685 4977.035 391.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.085 4977.035 456.365 4979.435 ;
    END
  END mprj_io_in[23]
  PIN mprj_analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4833.665 210.965 4833.945 ;
    END
  END mprj_analog_io[17]
  PIN mprj_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 4782.200 95.440 4844.800 ;
    END
  END mprj_io[24]
  PIN mprj_io_analog_en[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4821.705 210.965 4821.985 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_pol[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4815.265 210.965 4815.545 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4800.085 210.965 4800.365 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_dm[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4818.485 210.965 4818.765 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4827.685 210.965 4827.965 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4796.865 210.965 4797.145 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_enh[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4806.065 210.965 4806.345 ;
    END
  END mprj_io_enh[24]
  PIN mprj_io_hldh_n[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4802.845 210.965 4803.125 ;
    END
  END mprj_io_hldh_n[24]
  PIN mprj_io_holdover[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4793.645 210.965 4793.925 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4778.465 210.965 4778.745 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_inp_dis[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4812.505 210.965 4812.785 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4775.245 210.965 4775.525 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4790.885 210.965 4791.165 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_slow_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4836.885 210.965 4837.165 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4781.685 210.965 4781.965 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4846.085 210.965 4846.365 ;
    END
  END mprj_io_in[24]
  PIN mprj_analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3984.665 210.965 3984.945 ;
    END
  END mprj_analog_io[18]
  PIN mprj_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3933.200 95.440 3995.800 ;
    END
  END mprj_io[25]
  PIN mprj_io_analog_en[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3972.705 210.965 3972.985 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_pol[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3966.265 210.965 3966.545 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3951.085 210.965 3951.365 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_dm[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3969.485 210.965 3969.765 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3978.685 210.965 3978.965 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3947.865 210.965 3948.145 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_enh[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3957.065 210.965 3957.345 ;
    END
  END mprj_io_enh[25]
  PIN mprj_io_hldh_n[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3953.845 210.965 3954.125 ;
    END
  END mprj_io_hldh_n[25]
  PIN mprj_io_holdover[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3944.645 210.965 3944.925 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3929.465 210.965 3929.745 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_inp_dis[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3963.505 210.965 3963.785 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3926.245 210.965 3926.525 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3941.885 210.965 3942.165 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_slow_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3987.885 210.965 3988.165 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3932.685 210.965 3932.965 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3997.085 210.965 3997.365 ;
    END
  END mprj_io_in[25]
  PIN mprj_analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3768.665 210.965 3768.945 ;
    END
  END mprj_analog_io[19]
  PIN mprj_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3717.200 95.440 3779.800 ;
    END
  END mprj_io[26]
  PIN mprj_io_analog_en[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3756.705 210.965 3756.985 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_pol[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3750.265 210.965 3750.545 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3735.085 210.965 3735.365 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_dm[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3753.485 210.965 3753.765 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3762.685 210.965 3762.965 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3731.865 210.965 3732.145 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_enh[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3741.065 210.965 3741.345 ;
    END
  END mprj_io_enh[26]
  PIN mprj_io_hldh_n[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3737.845 210.965 3738.125 ;
    END
  END mprj_io_hldh_n[26]
  PIN mprj_io_holdover[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3728.645 210.965 3728.925 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3713.465 210.965 3713.745 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_inp_dis[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3747.505 210.965 3747.785 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3710.245 210.965 3710.525 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3725.885 210.965 3726.165 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_slow_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3771.885 210.965 3772.165 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3716.685 210.965 3716.965 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3781.085 210.965 3781.365 ;
    END
  END mprj_io_in[26]
  PIN mprj_analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3552.665 210.965 3552.945 ;
    END
  END mprj_analog_io[20]
  PIN mprj_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3501.200 95.440 3563.800 ;
    END
  END mprj_io[27]
  PIN mprj_io_analog_en[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3540.705 210.965 3540.985 ;
    END
  END mprj_io_analog_en[27]
  PIN mprj_io_analog_pol[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3534.265 210.965 3534.545 ;
    END
  END mprj_io_analog_pol[27]
  PIN mprj_io_analog_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3519.085 210.965 3519.365 ;
    END
  END mprj_io_analog_sel[27]
  PIN mprj_io_dm[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3537.485 210.965 3537.765 ;
    END
  END mprj_io_dm[81]
  PIN mprj_io_dm[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3546.685 210.965 3546.965 ;
    END
  END mprj_io_dm[82]
  PIN mprj_io_dm[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3515.865 210.965 3516.145 ;
    END
  END mprj_io_dm[83]
  PIN mprj_io_enh[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3525.065 210.965 3525.345 ;
    END
  END mprj_io_enh[27]
  PIN mprj_io_hldh_n[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3521.845 210.965 3522.125 ;
    END
  END mprj_io_hldh_n[27]
  PIN mprj_io_holdover[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3512.645 210.965 3512.925 ;
    END
  END mprj_io_holdover[27]
  PIN mprj_io_ib_mode_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3497.465 210.965 3497.745 ;
    END
  END mprj_io_ib_mode_sel[27]
  PIN mprj_io_inp_dis[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3531.505 210.965 3531.785 ;
    END
  END mprj_io_inp_dis[27]
  PIN mprj_io_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3494.245 210.965 3494.525 ;
    END
  END mprj_io_oeb[27]
  PIN mprj_io_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3509.885 210.965 3510.165 ;
    END
  END mprj_io_out[27]
  PIN mprj_io_slow_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3555.885 210.965 3556.165 ;
    END
  END mprj_io_slow_sel[27]
  PIN mprj_io_vtrip_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3500.685 210.965 3500.965 ;
    END
  END mprj_io_vtrip_sel[27]
  PIN mprj_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3565.085 210.965 3565.365 ;
    END
  END mprj_io_in[27]
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.290 4954.040 394.610 4954.100 ;
        RECT 651.430 4954.040 651.750 4954.100 ;
        RECT 1165.250 4954.040 1165.570 4954.100 ;
        RECT 1423.310 4954.040 1423.630 4954.100 ;
        RECT 1434.810 4954.040 1435.130 4954.100 ;
        RECT 394.290 4953.900 651.750 4954.040 ;
        RECT 394.290 4953.840 394.610 4953.900 ;
        RECT 651.430 4953.840 651.750 4953.900 ;
        RECT 973.520 4953.900 1435.130 4954.040 ;
        RECT 651.430 4953.360 651.750 4953.420 ;
        RECT 908.570 4953.360 908.890 4953.420 ;
        RECT 973.520 4953.360 973.660 4953.900 ;
        RECT 1165.250 4953.840 1165.570 4953.900 ;
        RECT 1423.310 4953.840 1423.630 4953.900 ;
        RECT 1434.810 4953.840 1435.130 4953.900 ;
        RECT 651.430 4953.220 973.660 4953.360 ;
        RECT 1932.530 4953.360 1932.850 4953.420 ;
        RECT 2377.350 4953.360 2377.670 4953.420 ;
        RECT 2634.490 4953.360 2634.810 4953.420 ;
        RECT 3132.670 4953.360 3132.990 4953.420 ;
        RECT 1932.530 4953.220 3132.990 4953.360 ;
        RECT 651.430 4953.160 651.750 4953.220 ;
        RECT 908.570 4953.160 908.890 4953.220 ;
        RECT 1932.530 4953.160 1932.850 4953.220 ;
        RECT 2377.350 4953.160 2377.670 4953.220 ;
        RECT 2634.490 4953.160 2634.810 4953.220 ;
        RECT 3132.670 4953.160 3132.990 4953.220 ;
        RECT 1434.810 4953.020 1435.130 4953.080 ;
        RECT 1932.620 4953.020 1932.760 4953.160 ;
        RECT 1434.810 4952.880 1932.760 4953.020 ;
        RECT 1434.810 4952.820 1435.130 4952.880 ;
        RECT 211.210 4950.980 211.530 4951.040 ;
        RECT 394.290 4950.980 394.610 4951.040 ;
        RECT 211.210 4950.840 394.610 4950.980 ;
        RECT 211.210 4950.780 211.530 4950.840 ;
        RECT 394.290 4950.780 394.610 4950.840 ;
        RECT 3132.670 4950.440 3132.990 4950.700 ;
        RECT 3143.250 4950.440 3143.570 4950.700 ;
        RECT 3132.760 4950.300 3132.900 4950.440 ;
        RECT 3143.340 4950.300 3143.480 4950.440 ;
        RECT 3367.270 4950.300 3367.590 4950.360 ;
        RECT 3132.760 4950.160 3367.590 4950.300 ;
        RECT 3367.270 4950.100 3367.590 4950.160 ;
        RECT 3367.270 4826.540 3367.590 4826.600 ;
        RECT 3376.930 4826.540 3377.250 4826.600 ;
        RECT 3367.270 4826.400 3377.250 4826.540 ;
        RECT 3367.270 4826.340 3367.590 4826.400 ;
        RECT 3376.930 4826.340 3377.250 4826.400 ;
        RECT 211.210 4788.600 211.530 4788.860 ;
        RECT 211.300 4787.840 211.440 4788.600 ;
        RECT 211.210 4787.580 211.530 4787.840 ;
        RECT 3367.270 4376.040 3367.590 4376.100 ;
        RECT 3376.930 4376.040 3377.250 4376.100 ;
        RECT 3367.270 4375.900 3377.250 4376.040 ;
        RECT 3367.270 4375.840 3367.590 4375.900 ;
        RECT 3376.930 4375.840 3377.250 4375.900 ;
        RECT 208.910 3933.360 209.230 3933.420 ;
        RECT 212.590 3933.360 212.910 3933.420 ;
        RECT 208.910 3933.220 212.910 3933.360 ;
        RECT 208.910 3933.160 209.230 3933.220 ;
        RECT 212.590 3933.160 212.910 3933.220 ;
        RECT 3367.270 3933.020 3367.590 3933.080 ;
        RECT 3370.030 3933.020 3370.350 3933.080 ;
        RECT 3376.930 3933.020 3377.250 3933.080 ;
        RECT 3367.270 3932.880 3377.250 3933.020 ;
        RECT 3367.270 3932.820 3367.590 3932.880 ;
        RECT 3370.030 3932.820 3370.350 3932.880 ;
        RECT 3376.930 3932.820 3377.250 3932.880 ;
        RECT 3368.650 3864.000 3368.970 3864.060 ;
        RECT 3370.030 3864.000 3370.350 3864.060 ;
        RECT 3368.650 3863.860 3370.350 3864.000 ;
        RECT 3368.650 3863.800 3368.970 3863.860 ;
        RECT 3370.030 3863.800 3370.350 3863.860 ;
        RECT 212.590 3794.980 212.910 3795.040 ;
        RECT 213.970 3794.980 214.290 3795.040 ;
        RECT 212.590 3794.840 214.290 3794.980 ;
        RECT 212.590 3794.780 212.910 3794.840 ;
        RECT 213.970 3794.780 214.290 3794.840 ;
        RECT 3368.650 3767.780 3368.970 3767.840 ;
        RECT 3369.570 3767.780 3369.890 3767.840 ;
        RECT 3368.650 3767.640 3369.890 3767.780 ;
        RECT 3368.650 3767.580 3368.970 3767.640 ;
        RECT 3369.570 3767.580 3369.890 3767.640 ;
        RECT 212.590 3767.440 212.910 3767.500 ;
        RECT 213.970 3767.440 214.290 3767.500 ;
        RECT 212.590 3767.300 214.290 3767.440 ;
        RECT 212.590 3767.240 212.910 3767.300 ;
        RECT 213.970 3767.240 214.290 3767.300 ;
        RECT 208.910 3720.180 209.230 3720.240 ;
        RECT 212.590 3720.180 212.910 3720.240 ;
        RECT 214.890 3720.180 215.210 3720.240 ;
        RECT 208.910 3720.040 215.210 3720.180 ;
        RECT 208.910 3719.980 209.230 3720.040 ;
        RECT 212.590 3719.980 212.910 3720.040 ;
        RECT 214.890 3719.980 215.210 3720.040 ;
        RECT 3368.190 3709.980 3368.510 3710.040 ;
        RECT 3369.570 3709.980 3369.890 3710.040 ;
        RECT 3368.190 3709.840 3377.160 3709.980 ;
        RECT 3368.190 3709.780 3368.510 3709.840 ;
        RECT 3369.570 3709.780 3369.890 3709.840 ;
        RECT 3377.020 3709.700 3377.160 3709.840 ;
        RECT 3376.930 3709.440 3377.250 3709.700 ;
        RECT 3368.190 3698.900 3368.510 3699.160 ;
        RECT 3368.280 3698.480 3368.420 3698.900 ;
        RECT 3368.190 3698.220 3368.510 3698.480 ;
        RECT 212.590 3670.880 212.910 3670.940 ;
        RECT 214.890 3670.880 215.210 3670.940 ;
        RECT 212.590 3670.740 215.210 3670.880 ;
        RECT 212.590 3670.680 212.910 3670.740 ;
        RECT 214.890 3670.680 215.210 3670.740 ;
        RECT 212.590 3601.860 212.910 3601.920 ;
        RECT 214.430 3601.860 214.750 3601.920 ;
        RECT 212.590 3601.720 214.750 3601.860 ;
        RECT 212.590 3601.660 212.910 3601.720 ;
        RECT 214.430 3601.660 214.750 3601.720 ;
        RECT 3368.190 3505.300 3368.510 3505.360 ;
        RECT 3369.110 3505.300 3369.430 3505.360 ;
        RECT 3368.190 3505.160 3369.430 3505.300 ;
        RECT 3368.190 3505.100 3368.510 3505.160 ;
        RECT 3369.110 3505.100 3369.430 3505.160 ;
        RECT 208.910 3504.280 209.230 3504.340 ;
        RECT 214.430 3504.280 214.750 3504.340 ;
        RECT 208.910 3504.140 214.750 3504.280 ;
        RECT 208.910 3504.080 209.230 3504.140 ;
        RECT 214.430 3504.080 214.750 3504.140 ;
        RECT 3376.930 3479.600 3377.250 3479.860 ;
        RECT 3368.190 3479.460 3368.510 3479.520 ;
        RECT 3377.020 3479.460 3377.160 3479.600 ;
        RECT 3368.190 3479.320 3377.160 3479.460 ;
        RECT 3368.190 3479.260 3368.510 3479.320 ;
        RECT 212.130 3477.760 212.450 3477.820 ;
        RECT 214.430 3477.760 214.750 3477.820 ;
        RECT 212.130 3477.620 214.750 3477.760 ;
        RECT 212.130 3477.560 212.450 3477.620 ;
        RECT 214.430 3477.560 214.750 3477.620 ;
        RECT 212.130 3408.200 212.450 3408.460 ;
        RECT 212.220 3408.060 212.360 3408.200 ;
        RECT 213.970 3408.060 214.290 3408.120 ;
        RECT 212.220 3407.920 214.290 3408.060 ;
        RECT 213.970 3407.860 214.290 3407.920 ;
        RECT 208.910 3290.420 209.230 3290.480 ;
        RECT 213.970 3290.420 214.290 3290.480 ;
        RECT 208.910 3290.280 214.290 3290.420 ;
        RECT 208.910 3290.220 209.230 3290.280 ;
        RECT 213.970 3290.220 214.290 3290.280 ;
        RECT 3368.190 3258.800 3368.510 3258.860 ;
        RECT 3376.930 3258.800 3377.250 3258.860 ;
        RECT 3368.190 3258.660 3377.250 3258.800 ;
        RECT 3368.190 3258.600 3368.510 3258.660 ;
        RECT 3376.930 3258.600 3377.250 3258.660 ;
        RECT 212.130 3257.100 212.450 3257.160 ;
        RECT 213.970 3257.100 214.290 3257.160 ;
        RECT 212.130 3256.960 214.290 3257.100 ;
        RECT 212.130 3256.900 212.450 3256.960 ;
        RECT 213.970 3256.900 214.290 3256.960 ;
        RECT 208.910 3074.180 209.230 3074.240 ;
        RECT 212.590 3074.180 212.910 3074.240 ;
        RECT 208.910 3074.040 212.910 3074.180 ;
        RECT 208.910 3073.980 209.230 3074.040 ;
        RECT 212.590 3073.980 212.910 3074.040 ;
        RECT 3368.190 3033.720 3368.510 3033.780 ;
        RECT 3376.930 3033.720 3377.250 3033.780 ;
        RECT 3368.190 3033.580 3377.250 3033.720 ;
        RECT 3368.190 3033.520 3368.510 3033.580 ;
        RECT 3376.930 3033.520 3377.250 3033.580 ;
        RECT 3367.730 2925.940 3368.050 2926.000 ;
        RECT 3369.110 2925.940 3369.430 2926.000 ;
        RECT 3367.730 2925.800 3369.430 2925.940 ;
        RECT 3367.730 2925.740 3368.050 2925.800 ;
        RECT 3369.110 2925.740 3369.430 2925.800 ;
        RECT 208.910 2853.520 209.230 2853.580 ;
        RECT 212.590 2853.520 212.910 2853.580 ;
        RECT 213.510 2853.520 213.830 2853.580 ;
        RECT 208.910 2853.380 213.830 2853.520 ;
        RECT 208.910 2853.320 209.230 2853.380 ;
        RECT 212.590 2853.320 212.910 2853.380 ;
        RECT 213.510 2853.320 213.830 2853.380 ;
        RECT 3367.730 2802.860 3368.050 2802.920 ;
        RECT 3369.110 2802.860 3369.430 2802.920 ;
        RECT 3376.930 2802.860 3377.250 2802.920 ;
        RECT 3367.730 2802.720 3377.250 2802.860 ;
        RECT 3367.730 2802.660 3368.050 2802.720 ;
        RECT 3369.110 2802.660 3369.430 2802.720 ;
        RECT 3376.930 2802.660 3377.250 2802.720 ;
        RECT 3367.730 2731.940 3368.050 2732.200 ;
        RECT 3367.820 2731.800 3367.960 2731.940 ;
        RECT 3369.110 2731.800 3369.430 2731.860 ;
        RECT 3367.820 2731.660 3369.430 2731.800 ;
        RECT 3369.110 2731.600 3369.430 2731.660 ;
        RECT 208.910 2637.620 209.230 2637.680 ;
        RECT 212.130 2637.620 212.450 2637.680 ;
        RECT 213.510 2637.620 213.830 2637.680 ;
        RECT 208.910 2637.480 213.830 2637.620 ;
        RECT 208.910 2637.420 209.230 2637.480 ;
        RECT 212.130 2637.420 212.450 2637.480 ;
        RECT 213.510 2637.420 213.830 2637.480 ;
        RECT 3367.730 2491.080 3368.050 2491.140 ;
        RECT 3369.110 2491.080 3369.430 2491.140 ;
        RECT 3367.730 2490.940 3369.430 2491.080 ;
        RECT 3367.730 2490.880 3368.050 2490.940 ;
        RECT 3369.110 2490.880 3369.430 2490.940 ;
        RECT 3367.730 2247.980 3368.050 2248.040 ;
        RECT 3369.110 2247.980 3369.430 2248.040 ;
        RECT 3367.730 2247.840 3369.430 2247.980 ;
        RECT 3367.730 2247.780 3368.050 2247.840 ;
        RECT 3369.110 2247.780 3369.430 2247.840 ;
        RECT 208.910 2004.200 209.230 2004.260 ;
        RECT 212.130 2004.200 212.450 2004.260 ;
        RECT 208.910 2004.060 212.450 2004.200 ;
        RECT 208.910 2004.000 209.230 2004.060 ;
        RECT 212.130 2004.000 212.450 2004.060 ;
        RECT 3368.650 1921.580 3368.970 1921.640 ;
        RECT 3376.930 1921.580 3377.250 1921.640 ;
        RECT 3368.650 1921.440 3377.250 1921.580 ;
        RECT 3368.650 1921.380 3368.970 1921.440 ;
        RECT 3376.930 1921.380 3377.250 1921.440 ;
        RECT 3367.730 1904.580 3368.050 1904.640 ;
        RECT 3368.650 1904.580 3368.970 1904.640 ;
        RECT 3367.730 1904.440 3368.970 1904.580 ;
        RECT 3367.730 1904.380 3368.050 1904.440 ;
        RECT 3368.650 1904.380 3368.970 1904.440 ;
        RECT 208.910 1788.300 209.230 1788.360 ;
        RECT 212.130 1788.300 212.450 1788.360 ;
        RECT 213.050 1788.300 213.370 1788.360 ;
        RECT 208.910 1788.160 213.370 1788.300 ;
        RECT 208.910 1788.100 209.230 1788.160 ;
        RECT 212.130 1788.100 212.450 1788.160 ;
        RECT 213.050 1788.100 213.370 1788.160 ;
        RECT 3367.730 1690.720 3368.050 1690.780 ;
        RECT 3376.930 1690.720 3377.250 1690.780 ;
        RECT 3367.730 1690.580 3377.250 1690.720 ;
        RECT 3367.730 1690.520 3368.050 1690.580 ;
        RECT 3376.930 1690.520 3377.250 1690.580 ;
        RECT 213.050 1614.020 213.370 1614.280 ;
        RECT 213.140 1613.880 213.280 1614.020 ;
        RECT 214.430 1613.880 214.750 1613.940 ;
        RECT 213.140 1613.740 214.750 1613.880 ;
        RECT 214.430 1613.680 214.750 1613.740 ;
        RECT 208.910 1567.440 209.230 1567.700 ;
        RECT 209.000 1567.300 209.140 1567.440 ;
        RECT 213.970 1567.300 214.290 1567.360 ;
        RECT 209.000 1567.160 214.290 1567.300 ;
        RECT 213.970 1567.100 214.290 1567.160 ;
        RECT 3367.730 1518.000 3368.050 1518.060 ;
        RECT 3376.470 1518.000 3376.790 1518.060 ;
        RECT 3367.730 1517.860 3376.790 1518.000 ;
        RECT 3367.730 1517.800 3368.050 1517.860 ;
        RECT 3376.470 1517.800 3376.790 1517.860 ;
        RECT 3368.190 1467.340 3368.510 1467.400 ;
        RECT 3376.470 1467.340 3376.790 1467.400 ;
        RECT 3368.190 1467.200 3376.790 1467.340 ;
        RECT 3368.190 1467.140 3368.510 1467.200 ;
        RECT 3376.470 1467.140 3376.790 1467.200 ;
        RECT 208.910 1356.160 209.230 1356.220 ;
        RECT 212.590 1356.160 212.910 1356.220 ;
        RECT 213.970 1356.160 214.290 1356.220 ;
        RECT 208.910 1356.020 214.290 1356.160 ;
        RECT 208.910 1355.960 209.230 1356.020 ;
        RECT 212.590 1355.960 212.910 1356.020 ;
        RECT 213.970 1355.960 214.290 1356.020 ;
        RECT 3367.270 1324.880 3367.590 1324.940 ;
        RECT 3368.190 1324.880 3368.510 1324.940 ;
        RECT 3367.270 1324.740 3368.510 1324.880 ;
        RECT 3367.270 1324.680 3367.590 1324.740 ;
        RECT 3368.190 1324.680 3368.510 1324.740 ;
        RECT 3367.270 1243.620 3367.590 1243.680 ;
        RECT 3376.470 1243.620 3376.790 1243.680 ;
        RECT 3367.270 1243.480 3376.790 1243.620 ;
        RECT 3367.270 1243.420 3367.590 1243.480 ;
        RECT 3376.470 1243.420 3376.790 1243.480 ;
        RECT 212.590 1227.640 212.910 1227.700 ;
        RECT 213.970 1227.640 214.290 1227.700 ;
        RECT 212.590 1227.500 214.290 1227.640 ;
        RECT 212.590 1227.440 212.910 1227.500 ;
        RECT 213.970 1227.440 214.290 1227.500 ;
        RECT 3369.110 1219.140 3369.430 1219.200 ;
        RECT 3376.470 1219.140 3376.790 1219.200 ;
        RECT 3369.110 1219.000 3376.790 1219.140 ;
        RECT 3369.110 1218.940 3369.430 1219.000 ;
        RECT 3376.470 1218.940 3376.790 1219.000 ;
        RECT 208.910 1140.260 209.230 1140.320 ;
        RECT 213.050 1140.260 213.370 1140.320 ;
        RECT 213.970 1140.260 214.290 1140.320 ;
        RECT 208.910 1140.120 214.290 1140.260 ;
        RECT 208.910 1140.060 209.230 1140.120 ;
        RECT 213.050 1140.060 213.370 1140.120 ;
        RECT 213.970 1140.060 214.290 1140.120 ;
        RECT 3369.110 1090.420 3369.430 1090.680 ;
        RECT 3369.200 1090.000 3369.340 1090.420 ;
        RECT 3369.110 1089.740 3369.430 1090.000 ;
        RECT 3368.650 1062.740 3368.970 1062.800 ;
        RECT 3369.110 1062.740 3369.430 1062.800 ;
        RECT 3368.650 1062.600 3369.430 1062.740 ;
        RECT 3368.650 1062.540 3368.970 1062.600 ;
        RECT 3369.110 1062.540 3369.430 1062.600 ;
        RECT 3368.650 1019.560 3368.970 1019.620 ;
        RECT 3376.930 1019.560 3377.250 1019.620 ;
        RECT 3368.650 1019.420 3377.250 1019.560 ;
        RECT 3368.650 1019.360 3368.970 1019.420 ;
        RECT 3376.930 1019.360 3377.250 1019.420 ;
        RECT 208.910 924.360 209.230 924.420 ;
        RECT 212.130 924.360 212.450 924.420 ;
        RECT 213.050 924.360 213.370 924.420 ;
        RECT 208.910 924.220 213.370 924.360 ;
        RECT 208.910 924.160 209.230 924.220 ;
        RECT 212.130 924.160 212.450 924.220 ;
        RECT 213.050 924.160 213.370 924.220 ;
        RECT 3367.730 791.760 3368.050 791.820 ;
        RECT 3376.930 791.760 3377.250 791.820 ;
        RECT 3367.730 791.620 3377.250 791.760 ;
        RECT 3367.730 791.560 3368.050 791.620 ;
        RECT 3376.930 791.560 3377.250 791.620 ;
        RECT 3367.730 563.960 3368.050 564.020 ;
        RECT 3376.930 563.960 3377.250 564.020 ;
        RECT 3367.730 563.820 3377.250 563.960 ;
        RECT 3367.730 563.760 3368.050 563.820 ;
        RECT 3376.930 563.760 3377.250 563.820 ;
        RECT 212.130 228.380 212.450 228.440 ;
        RECT 718.130 228.380 718.450 228.440 ;
        RECT 212.130 228.240 718.450 228.380 ;
        RECT 212.130 228.180 212.450 228.240 ;
        RECT 718.130 228.180 718.450 228.240 ;
        RECT 2637.250 228.040 2637.570 228.100 ;
        RECT 3367.730 228.040 3368.050 228.100 ;
        RECT 2637.250 227.900 3368.050 228.040 ;
        RECT 2637.250 227.840 2637.570 227.900 ;
        RECT 3367.730 227.840 3368.050 227.900 ;
        RECT 718.130 221.920 718.450 221.980 ;
        RECT 725.490 221.920 725.810 221.980 ;
        RECT 976.650 221.920 976.970 221.980 ;
        RECT 998.270 221.920 998.590 221.980 ;
        RECT 718.130 221.780 998.590 221.920 ;
        RECT 718.130 221.720 718.450 221.780 ;
        RECT 725.490 221.720 725.810 221.780 ;
        RECT 976.650 221.720 976.970 221.780 ;
        RECT 998.270 221.720 998.590 221.780 ;
        RECT 1793.610 221.580 1793.930 221.640 ;
        RECT 2067.770 221.580 2068.090 221.640 ;
        RECT 2089.390 221.580 2089.710 221.640 ;
        RECT 2341.470 221.580 2341.790 221.640 ;
        RECT 2363.090 221.580 2363.410 221.640 ;
        RECT 2615.630 221.580 2615.950 221.640 ;
        RECT 1777.600 221.440 1793.930 221.580 ;
        RECT 998.270 221.240 998.590 221.300 ;
        RECT 1519.450 221.240 1519.770 221.300 ;
        RECT 1541.070 221.240 1541.390 221.300 ;
        RECT 1777.600 221.240 1777.740 221.440 ;
        RECT 1793.610 221.380 1793.930 221.440 ;
        RECT 1998.860 221.440 2615.950 221.580 ;
        RECT 998.270 221.100 1777.740 221.240 ;
        RECT 1815.230 221.240 1815.550 221.300 ;
        RECT 1998.860 221.240 1999.000 221.440 ;
        RECT 2067.770 221.380 2068.090 221.440 ;
        RECT 2089.390 221.380 2089.710 221.440 ;
        RECT 2341.470 221.380 2341.790 221.440 ;
        RECT 2363.090 221.380 2363.410 221.440 ;
        RECT 2615.630 221.380 2615.950 221.440 ;
        RECT 1815.230 221.100 1999.000 221.240 ;
        RECT 998.270 221.040 998.590 221.100 ;
        RECT 1519.450 221.040 1519.770 221.100 ;
        RECT 1541.070 221.040 1541.390 221.100 ;
        RECT 1815.230 221.040 1815.550 221.100 ;
        RECT 1793.610 220.900 1793.930 220.960 ;
        RECT 1815.320 220.900 1815.460 221.040 ;
        RECT 1793.610 220.760 1815.460 220.900 ;
        RECT 2615.630 220.900 2615.950 220.960 ;
        RECT 2637.250 220.900 2637.570 220.960 ;
        RECT 2615.630 220.760 2637.570 220.900 ;
        RECT 1793.610 220.700 1793.930 220.760 ;
        RECT 2615.630 220.700 2615.950 220.760 ;
        RECT 2637.250 220.700 2637.570 220.760 ;
      LAYER via ;
        RECT 394.320 4953.840 394.580 4954.100 ;
        RECT 651.460 4953.840 651.720 4954.100 ;
        RECT 651.460 4953.160 651.720 4953.420 ;
        RECT 908.600 4953.160 908.860 4953.420 ;
        RECT 1165.280 4953.840 1165.540 4954.100 ;
        RECT 1423.340 4953.840 1423.600 4954.100 ;
        RECT 1434.840 4953.840 1435.100 4954.100 ;
        RECT 1932.560 4953.160 1932.820 4953.420 ;
        RECT 2377.380 4953.160 2377.640 4953.420 ;
        RECT 2634.520 4953.160 2634.780 4953.420 ;
        RECT 3132.700 4953.160 3132.960 4953.420 ;
        RECT 1434.840 4952.820 1435.100 4953.080 ;
        RECT 211.240 4950.780 211.500 4951.040 ;
        RECT 394.320 4950.780 394.580 4951.040 ;
        RECT 3132.700 4950.440 3132.960 4950.700 ;
        RECT 3143.280 4950.440 3143.540 4950.700 ;
        RECT 3367.300 4950.100 3367.560 4950.360 ;
        RECT 3367.300 4826.340 3367.560 4826.600 ;
        RECT 3376.960 4826.340 3377.220 4826.600 ;
        RECT 211.240 4788.600 211.500 4788.860 ;
        RECT 211.240 4787.580 211.500 4787.840 ;
        RECT 3367.300 4375.840 3367.560 4376.100 ;
        RECT 3376.960 4375.840 3377.220 4376.100 ;
        RECT 208.940 3933.160 209.200 3933.420 ;
        RECT 212.620 3933.160 212.880 3933.420 ;
        RECT 3367.300 3932.820 3367.560 3933.080 ;
        RECT 3370.060 3932.820 3370.320 3933.080 ;
        RECT 3376.960 3932.820 3377.220 3933.080 ;
        RECT 3368.680 3863.800 3368.940 3864.060 ;
        RECT 3370.060 3863.800 3370.320 3864.060 ;
        RECT 212.620 3794.780 212.880 3795.040 ;
        RECT 214.000 3794.780 214.260 3795.040 ;
        RECT 3368.680 3767.580 3368.940 3767.840 ;
        RECT 3369.600 3767.580 3369.860 3767.840 ;
        RECT 212.620 3767.240 212.880 3767.500 ;
        RECT 214.000 3767.240 214.260 3767.500 ;
        RECT 208.940 3719.980 209.200 3720.240 ;
        RECT 212.620 3719.980 212.880 3720.240 ;
        RECT 214.920 3719.980 215.180 3720.240 ;
        RECT 3368.220 3709.780 3368.480 3710.040 ;
        RECT 3369.600 3709.780 3369.860 3710.040 ;
        RECT 3376.960 3709.440 3377.220 3709.700 ;
        RECT 3368.220 3698.900 3368.480 3699.160 ;
        RECT 3368.220 3698.220 3368.480 3698.480 ;
        RECT 212.620 3670.680 212.880 3670.940 ;
        RECT 214.920 3670.680 215.180 3670.940 ;
        RECT 212.620 3601.660 212.880 3601.920 ;
        RECT 214.460 3601.660 214.720 3601.920 ;
        RECT 3368.220 3505.100 3368.480 3505.360 ;
        RECT 3369.140 3505.100 3369.400 3505.360 ;
        RECT 208.940 3504.080 209.200 3504.340 ;
        RECT 214.460 3504.080 214.720 3504.340 ;
        RECT 3376.960 3479.600 3377.220 3479.860 ;
        RECT 3368.220 3479.260 3368.480 3479.520 ;
        RECT 212.160 3477.560 212.420 3477.820 ;
        RECT 214.460 3477.560 214.720 3477.820 ;
        RECT 212.160 3408.200 212.420 3408.460 ;
        RECT 214.000 3407.860 214.260 3408.120 ;
        RECT 208.940 3290.220 209.200 3290.480 ;
        RECT 214.000 3290.220 214.260 3290.480 ;
        RECT 3368.220 3258.600 3368.480 3258.860 ;
        RECT 3376.960 3258.600 3377.220 3258.860 ;
        RECT 212.160 3256.900 212.420 3257.160 ;
        RECT 214.000 3256.900 214.260 3257.160 ;
        RECT 208.940 3073.980 209.200 3074.240 ;
        RECT 212.620 3073.980 212.880 3074.240 ;
        RECT 3368.220 3033.520 3368.480 3033.780 ;
        RECT 3376.960 3033.520 3377.220 3033.780 ;
        RECT 3367.760 2925.740 3368.020 2926.000 ;
        RECT 3369.140 2925.740 3369.400 2926.000 ;
        RECT 208.940 2853.320 209.200 2853.580 ;
        RECT 212.620 2853.320 212.880 2853.580 ;
        RECT 213.540 2853.320 213.800 2853.580 ;
        RECT 3367.760 2802.660 3368.020 2802.920 ;
        RECT 3369.140 2802.660 3369.400 2802.920 ;
        RECT 3376.960 2802.660 3377.220 2802.920 ;
        RECT 3367.760 2731.940 3368.020 2732.200 ;
        RECT 3369.140 2731.600 3369.400 2731.860 ;
        RECT 208.940 2637.420 209.200 2637.680 ;
        RECT 212.160 2637.420 212.420 2637.680 ;
        RECT 213.540 2637.420 213.800 2637.680 ;
        RECT 3367.760 2490.880 3368.020 2491.140 ;
        RECT 3369.140 2490.880 3369.400 2491.140 ;
        RECT 3367.760 2247.780 3368.020 2248.040 ;
        RECT 3369.140 2247.780 3369.400 2248.040 ;
        RECT 208.940 2004.000 209.200 2004.260 ;
        RECT 212.160 2004.000 212.420 2004.260 ;
        RECT 3368.680 1921.380 3368.940 1921.640 ;
        RECT 3376.960 1921.380 3377.220 1921.640 ;
        RECT 3367.760 1904.380 3368.020 1904.640 ;
        RECT 3368.680 1904.380 3368.940 1904.640 ;
        RECT 208.940 1788.100 209.200 1788.360 ;
        RECT 212.160 1788.100 212.420 1788.360 ;
        RECT 213.080 1788.100 213.340 1788.360 ;
        RECT 3367.760 1690.520 3368.020 1690.780 ;
        RECT 3376.960 1690.520 3377.220 1690.780 ;
        RECT 213.080 1614.020 213.340 1614.280 ;
        RECT 214.460 1613.680 214.720 1613.940 ;
        RECT 208.940 1567.440 209.200 1567.700 ;
        RECT 214.000 1567.100 214.260 1567.360 ;
        RECT 3367.760 1517.800 3368.020 1518.060 ;
        RECT 3376.500 1517.800 3376.760 1518.060 ;
        RECT 3368.220 1467.140 3368.480 1467.400 ;
        RECT 3376.500 1467.140 3376.760 1467.400 ;
        RECT 208.940 1355.960 209.200 1356.220 ;
        RECT 212.620 1355.960 212.880 1356.220 ;
        RECT 214.000 1355.960 214.260 1356.220 ;
        RECT 3367.300 1324.680 3367.560 1324.940 ;
        RECT 3368.220 1324.680 3368.480 1324.940 ;
        RECT 3367.300 1243.420 3367.560 1243.680 ;
        RECT 3376.500 1243.420 3376.760 1243.680 ;
        RECT 212.620 1227.440 212.880 1227.700 ;
        RECT 214.000 1227.440 214.260 1227.700 ;
        RECT 3369.140 1218.940 3369.400 1219.200 ;
        RECT 3376.500 1218.940 3376.760 1219.200 ;
        RECT 208.940 1140.060 209.200 1140.320 ;
        RECT 213.080 1140.060 213.340 1140.320 ;
        RECT 214.000 1140.060 214.260 1140.320 ;
        RECT 3369.140 1090.420 3369.400 1090.680 ;
        RECT 3369.140 1089.740 3369.400 1090.000 ;
        RECT 3368.680 1062.540 3368.940 1062.800 ;
        RECT 3369.140 1062.540 3369.400 1062.800 ;
        RECT 3368.680 1019.360 3368.940 1019.620 ;
        RECT 3376.960 1019.360 3377.220 1019.620 ;
        RECT 208.940 924.160 209.200 924.420 ;
        RECT 212.160 924.160 212.420 924.420 ;
        RECT 213.080 924.160 213.340 924.420 ;
        RECT 3367.760 791.560 3368.020 791.820 ;
        RECT 3376.960 791.560 3377.220 791.820 ;
        RECT 3367.760 563.760 3368.020 564.020 ;
        RECT 3376.960 563.760 3377.220 564.020 ;
        RECT 212.160 228.180 212.420 228.440 ;
        RECT 718.160 228.180 718.420 228.440 ;
        RECT 2637.280 227.840 2637.540 228.100 ;
        RECT 3367.760 227.840 3368.020 228.100 ;
        RECT 718.160 221.720 718.420 221.980 ;
        RECT 725.520 221.720 725.780 221.980 ;
        RECT 976.680 221.720 976.940 221.980 ;
        RECT 998.300 221.720 998.560 221.980 ;
        RECT 998.300 221.040 998.560 221.300 ;
        RECT 1519.480 221.040 1519.740 221.300 ;
        RECT 1541.100 221.040 1541.360 221.300 ;
        RECT 1793.640 221.380 1793.900 221.640 ;
        RECT 1815.260 221.040 1815.520 221.300 ;
        RECT 2067.800 221.380 2068.060 221.640 ;
        RECT 2089.420 221.380 2089.680 221.640 ;
        RECT 2341.500 221.380 2341.760 221.640 ;
        RECT 2363.120 221.380 2363.380 221.640 ;
        RECT 2615.660 221.380 2615.920 221.640 ;
        RECT 1793.640 220.700 1793.900 220.960 ;
        RECT 2615.660 220.700 2615.920 220.960 ;
        RECT 2637.280 220.700 2637.540 220.960 ;
      LAYER met2 ;
        RECT 394.445 4977.260 394.725 4979.435 ;
        RECT 394.380 4977.035 394.725 4977.260 ;
        RECT 651.445 4977.035 651.725 4979.435 ;
        RECT 908.445 4977.330 908.725 4979.435 ;
        RECT 1165.445 4977.330 1165.725 4979.435 ;
        RECT 908.445 4977.035 908.800 4977.330 ;
        RECT 394.380 4954.130 394.520 4977.035 ;
        RECT 651.520 4954.130 651.660 4977.035 ;
        RECT 394.320 4953.810 394.580 4954.130 ;
        RECT 651.460 4953.810 651.720 4954.130 ;
        RECT 394.380 4951.070 394.520 4953.810 ;
        RECT 651.520 4953.450 651.660 4953.810 ;
        RECT 908.660 4953.450 908.800 4977.035 ;
        RECT 1165.340 4977.035 1165.725 4977.330 ;
        RECT 1423.445 4977.260 1423.725 4979.435 ;
        RECT 1423.400 4977.035 1423.725 4977.260 ;
        RECT 1932.445 4977.260 1932.725 4979.435 ;
        RECT 2377.445 4977.260 2377.725 4979.435 ;
        RECT 1932.445 4977.035 1932.760 4977.260 ;
        RECT 1165.340 4954.130 1165.480 4977.035 ;
        RECT 1423.400 4954.130 1423.540 4977.035 ;
        RECT 1165.280 4953.810 1165.540 4954.130 ;
        RECT 1423.340 4953.810 1423.600 4954.130 ;
        RECT 1434.840 4953.810 1435.100 4954.130 ;
        RECT 651.460 4953.130 651.720 4953.450 ;
        RECT 908.600 4953.130 908.860 4953.450 ;
        RECT 1434.900 4953.110 1435.040 4953.810 ;
        RECT 1932.620 4953.450 1932.760 4977.035 ;
        RECT 2377.440 4977.035 2377.725 4977.260 ;
        RECT 2634.445 4977.035 2634.725 4979.435 ;
        RECT 3143.445 4977.330 3143.725 4979.435 ;
        RECT 3143.340 4977.035 3143.725 4977.330 ;
        RECT 2377.440 4953.450 2377.580 4977.035 ;
        RECT 2634.580 4953.450 2634.720 4977.035 ;
        RECT 1932.560 4953.130 1932.820 4953.450 ;
        RECT 2377.380 4953.130 2377.640 4953.450 ;
        RECT 2634.520 4953.130 2634.780 4953.450 ;
        RECT 3132.700 4953.130 3132.960 4953.450 ;
        RECT 1434.840 4952.790 1435.100 4953.110 ;
        RECT 211.240 4950.750 211.500 4951.070 ;
        RECT 394.320 4950.750 394.580 4951.070 ;
        RECT 211.300 4788.890 211.440 4950.750 ;
        RECT 3132.760 4950.730 3132.900 4953.130 ;
        RECT 3143.340 4950.730 3143.480 4977.035 ;
        RECT 3132.700 4950.410 3132.960 4950.730 ;
        RECT 3143.280 4950.410 3143.540 4950.730 ;
        RECT 3367.300 4950.070 3367.560 4950.390 ;
        RECT 3367.360 4826.630 3367.500 4950.070 ;
        RECT 3367.300 4826.310 3367.560 4826.630 ;
        RECT 3376.960 4826.310 3377.220 4826.630 ;
        RECT 211.240 4788.570 211.500 4788.890 ;
        RECT 211.240 4787.550 211.500 4787.870 ;
        RECT 208.565 4784.655 210.965 4784.725 ;
        RECT 211.300 4784.655 211.440 4787.550 ;
        RECT 208.565 4784.515 211.440 4784.655 ;
        RECT 208.565 4784.445 210.965 4784.515 ;
        RECT 3367.360 4376.130 3367.500 4826.310 ;
        RECT 3377.020 4824.555 3377.160 4826.310 ;
        RECT 3377.020 4824.415 3379.435 4824.555 ;
        RECT 3377.035 4824.275 3379.435 4824.415 ;
        RECT 3377.035 4378.415 3379.435 4378.555 ;
        RECT 3377.020 4378.275 3379.435 4378.415 ;
        RECT 3377.020 4376.130 3377.160 4378.275 ;
        RECT 3367.300 4375.810 3367.560 4376.130 ;
        RECT 3376.960 4375.810 3377.220 4376.130 ;
        RECT 208.565 3935.445 210.965 3935.725 ;
        RECT 209.000 3933.450 209.140 3935.445 ;
        RECT 208.940 3933.130 209.200 3933.450 ;
        RECT 212.620 3933.130 212.880 3933.450 ;
        RECT 212.680 3795.070 212.820 3933.130 ;
        RECT 3367.360 3933.110 3367.500 4375.810 ;
        RECT 3367.300 3932.790 3367.560 3933.110 ;
        RECT 3370.060 3932.790 3370.320 3933.110 ;
        RECT 3376.960 3932.790 3377.220 3933.110 ;
        RECT 3370.120 3864.090 3370.260 3932.790 ;
        RECT 3377.020 3932.555 3377.160 3932.790 ;
        RECT 3377.020 3932.415 3379.435 3932.555 ;
        RECT 3377.035 3932.275 3379.435 3932.415 ;
        RECT 3368.680 3863.770 3368.940 3864.090 ;
        RECT 3370.060 3863.770 3370.320 3864.090 ;
        RECT 212.620 3794.750 212.880 3795.070 ;
        RECT 214.000 3794.750 214.260 3795.070 ;
        RECT 214.060 3767.530 214.200 3794.750 ;
        RECT 3368.740 3767.870 3368.880 3863.770 ;
        RECT 3368.680 3767.550 3368.940 3767.870 ;
        RECT 3369.600 3767.550 3369.860 3767.870 ;
        RECT 212.620 3767.210 212.880 3767.530 ;
        RECT 214.000 3767.210 214.260 3767.530 ;
        RECT 212.680 3720.270 212.820 3767.210 ;
        RECT 208.940 3719.950 209.200 3720.270 ;
        RECT 212.620 3719.950 212.880 3720.270 ;
        RECT 214.920 3719.950 215.180 3720.270 ;
        RECT 209.000 3719.725 209.140 3719.950 ;
        RECT 208.565 3719.445 210.965 3719.725 ;
        RECT 214.980 3670.970 215.120 3719.950 ;
        RECT 3369.660 3710.070 3369.800 3767.550 ;
        RECT 3368.220 3709.750 3368.480 3710.070 ;
        RECT 3369.600 3709.750 3369.860 3710.070 ;
        RECT 3368.280 3699.190 3368.420 3709.750 ;
        RECT 3376.960 3709.410 3377.220 3709.730 ;
        RECT 3377.020 3707.555 3377.160 3709.410 ;
        RECT 3377.020 3707.415 3379.435 3707.555 ;
        RECT 3377.035 3707.275 3379.435 3707.415 ;
        RECT 3368.220 3698.870 3368.480 3699.190 ;
        RECT 3368.220 3698.190 3368.480 3698.510 ;
        RECT 212.620 3670.650 212.880 3670.970 ;
        RECT 214.920 3670.650 215.180 3670.970 ;
        RECT 212.680 3601.950 212.820 3670.650 ;
        RECT 212.620 3601.630 212.880 3601.950 ;
        RECT 214.460 3601.630 214.720 3601.950 ;
        RECT 3368.280 3601.690 3368.420 3698.190 ;
        RECT 214.520 3504.370 214.660 3601.630 ;
        RECT 3368.280 3601.550 3369.340 3601.690 ;
        RECT 3369.200 3505.390 3369.340 3601.550 ;
        RECT 3368.220 3505.070 3368.480 3505.390 ;
        RECT 3369.140 3505.070 3369.400 3505.390 ;
        RECT 208.940 3504.050 209.200 3504.370 ;
        RECT 214.460 3504.050 214.720 3504.370 ;
        RECT 209.000 3503.725 209.140 3504.050 ;
        RECT 208.565 3503.445 210.965 3503.725 ;
        RECT 214.520 3477.850 214.660 3504.050 ;
        RECT 3368.280 3479.550 3368.420 3505.070 ;
        RECT 3377.035 3482.415 3379.435 3482.555 ;
        RECT 3377.020 3482.275 3379.435 3482.415 ;
        RECT 3377.020 3479.890 3377.160 3482.275 ;
        RECT 3376.960 3479.570 3377.220 3479.890 ;
        RECT 3368.220 3479.230 3368.480 3479.550 ;
        RECT 212.160 3477.530 212.420 3477.850 ;
        RECT 214.460 3477.530 214.720 3477.850 ;
        RECT 212.220 3408.490 212.360 3477.530 ;
        RECT 212.160 3408.170 212.420 3408.490 ;
        RECT 214.000 3407.830 214.260 3408.150 ;
        RECT 214.060 3290.510 214.200 3407.830 ;
        RECT 208.940 3290.190 209.200 3290.510 ;
        RECT 214.000 3290.190 214.260 3290.510 ;
        RECT 209.000 3287.725 209.140 3290.190 ;
        RECT 208.565 3287.445 210.965 3287.725 ;
        RECT 214.060 3257.190 214.200 3290.190 ;
        RECT 3368.280 3258.890 3368.420 3479.230 ;
        RECT 3368.220 3258.570 3368.480 3258.890 ;
        RECT 3376.960 3258.570 3377.220 3258.890 ;
        RECT 212.160 3256.870 212.420 3257.190 ;
        RECT 214.000 3256.870 214.260 3257.190 ;
        RECT 212.220 3159.690 212.360 3256.870 ;
        RECT 212.220 3159.550 212.820 3159.690 ;
        RECT 212.680 3074.270 212.820 3159.550 ;
        RECT 208.940 3073.950 209.200 3074.270 ;
        RECT 212.620 3073.950 212.880 3074.270 ;
        RECT 209.000 3071.725 209.140 3073.950 ;
        RECT 208.565 3071.445 210.965 3071.725 ;
        RECT 208.565 2855.445 210.965 2855.725 ;
        RECT 209.000 2853.610 209.140 2855.445 ;
        RECT 212.680 2853.610 212.820 3073.950 ;
        RECT 3368.280 3033.810 3368.420 3258.570 ;
        RECT 3377.020 3256.555 3377.160 3258.570 ;
        RECT 3377.020 3256.415 3379.435 3256.555 ;
        RECT 3377.035 3256.275 3379.435 3256.415 ;
        RECT 3368.220 3033.490 3368.480 3033.810 ;
        RECT 3376.960 3033.490 3377.220 3033.810 ;
        RECT 3368.280 2975.410 3368.420 3033.490 ;
        RECT 3377.020 3031.555 3377.160 3033.490 ;
        RECT 3377.020 3031.415 3379.435 3031.555 ;
        RECT 3377.035 3031.275 3379.435 3031.415 ;
        RECT 3367.820 2975.270 3368.420 2975.410 ;
        RECT 3367.820 2926.030 3367.960 2975.270 ;
        RECT 3367.760 2925.710 3368.020 2926.030 ;
        RECT 3369.140 2925.710 3369.400 2926.030 ;
        RECT 208.940 2853.290 209.200 2853.610 ;
        RECT 212.620 2853.290 212.880 2853.610 ;
        RECT 213.540 2853.290 213.800 2853.610 ;
        RECT 208.565 2639.445 210.965 2639.725 ;
        RECT 209.000 2637.710 209.140 2639.445 ;
        RECT 213.600 2637.710 213.740 2853.290 ;
        RECT 3369.200 2802.950 3369.340 2925.710 ;
        RECT 3377.035 2805.340 3379.435 2805.555 ;
        RECT 3377.020 2805.275 3379.435 2805.340 ;
        RECT 3377.020 2802.950 3377.160 2805.275 ;
        RECT 3367.760 2802.630 3368.020 2802.950 ;
        RECT 3369.140 2802.630 3369.400 2802.950 ;
        RECT 3376.960 2802.630 3377.220 2802.950 ;
        RECT 3367.820 2732.230 3367.960 2802.630 ;
        RECT 3367.760 2731.910 3368.020 2732.230 ;
        RECT 3369.140 2731.570 3369.400 2731.890 ;
        RECT 208.940 2637.390 209.200 2637.710 ;
        RECT 212.160 2637.390 212.420 2637.710 ;
        RECT 213.540 2637.390 213.800 2637.710 ;
        RECT 212.220 2004.290 212.360 2637.390 ;
        RECT 3369.200 2491.170 3369.340 2731.570 ;
        RECT 3367.760 2490.850 3368.020 2491.170 ;
        RECT 3369.140 2490.850 3369.400 2491.170 ;
        RECT 3367.820 2248.070 3367.960 2490.850 ;
        RECT 3367.760 2247.750 3368.020 2248.070 ;
        RECT 3369.140 2247.750 3369.400 2248.070 ;
        RECT 3369.200 2104.330 3369.340 2247.750 ;
        RECT 3368.740 2104.190 3369.340 2104.330 ;
        RECT 208.940 2003.970 209.200 2004.290 ;
        RECT 212.160 2003.970 212.420 2004.290 ;
        RECT 209.000 2001.725 209.140 2003.970 ;
        RECT 208.565 2001.445 210.965 2001.725 ;
        RECT 212.220 1788.390 212.360 2003.970 ;
        RECT 3368.740 1921.670 3368.880 2104.190 ;
        RECT 3368.680 1921.350 3368.940 1921.670 ;
        RECT 3376.960 1921.350 3377.220 1921.670 ;
        RECT 3368.740 1904.670 3368.880 1921.350 ;
        RECT 3377.020 1919.555 3377.160 1921.350 ;
        RECT 3377.020 1919.300 3379.435 1919.555 ;
        RECT 3377.035 1919.275 3379.435 1919.300 ;
        RECT 3367.760 1904.350 3368.020 1904.670 ;
        RECT 3368.680 1904.350 3368.940 1904.670 ;
        RECT 208.940 1788.070 209.200 1788.390 ;
        RECT 212.160 1788.070 212.420 1788.390 ;
        RECT 213.080 1788.070 213.340 1788.390 ;
        RECT 209.000 1785.725 209.140 1788.070 ;
        RECT 208.565 1785.445 210.965 1785.725 ;
        RECT 213.140 1614.310 213.280 1788.070 ;
        RECT 3367.820 1690.810 3367.960 1904.350 ;
        RECT 3377.035 1693.540 3379.435 1693.555 ;
        RECT 3377.020 1693.275 3379.435 1693.540 ;
        RECT 3377.020 1690.810 3377.160 1693.275 ;
        RECT 3367.760 1690.490 3368.020 1690.810 ;
        RECT 3376.960 1690.490 3377.220 1690.810 ;
        RECT 213.080 1613.990 213.340 1614.310 ;
        RECT 214.460 1613.650 214.720 1613.970 ;
        RECT 208.565 1569.445 210.965 1569.725 ;
        RECT 209.000 1567.730 209.140 1569.445 ;
        RECT 208.940 1567.410 209.200 1567.730 ;
        RECT 214.000 1567.130 214.260 1567.390 ;
        RECT 214.520 1567.130 214.660 1613.650 ;
        RECT 214.000 1567.070 214.660 1567.130 ;
        RECT 214.060 1566.990 214.660 1567.070 ;
        RECT 214.060 1356.250 214.200 1566.990 ;
        RECT 3367.820 1518.090 3367.960 1690.490 ;
        RECT 3367.760 1517.770 3368.020 1518.090 ;
        RECT 3376.500 1517.770 3376.760 1518.090 ;
        RECT 3376.560 1468.530 3376.700 1517.770 ;
        RECT 3377.035 1468.530 3379.435 1468.555 ;
        RECT 3376.560 1468.390 3379.435 1468.530 ;
        RECT 3376.560 1467.430 3376.700 1468.390 ;
        RECT 3377.035 1468.275 3379.435 1468.390 ;
        RECT 3368.220 1467.110 3368.480 1467.430 ;
        RECT 3376.500 1467.110 3376.760 1467.430 ;
        RECT 208.940 1355.930 209.200 1356.250 ;
        RECT 212.620 1355.930 212.880 1356.250 ;
        RECT 214.000 1355.930 214.260 1356.250 ;
        RECT 209.000 1353.725 209.140 1355.930 ;
        RECT 208.565 1353.445 210.965 1353.725 ;
        RECT 212.680 1227.730 212.820 1355.930 ;
        RECT 3368.280 1324.970 3368.420 1467.110 ;
        RECT 3367.300 1324.650 3367.560 1324.970 ;
        RECT 3368.220 1324.650 3368.480 1324.970 ;
        RECT 3367.360 1243.710 3367.500 1324.650 ;
        RECT 3376.560 1243.710 3376.700 1243.865 ;
        RECT 3367.300 1243.390 3367.560 1243.710 ;
        RECT 3376.500 1243.450 3376.760 1243.710 ;
        RECT 3377.035 1243.450 3379.435 1243.555 ;
        RECT 3376.500 1243.390 3379.435 1243.450 ;
        RECT 3376.560 1243.310 3379.435 1243.390 ;
        RECT 212.620 1227.410 212.880 1227.730 ;
        RECT 214.000 1227.410 214.260 1227.730 ;
        RECT 214.060 1140.350 214.200 1227.410 ;
        RECT 3376.560 1219.230 3376.700 1243.310 ;
        RECT 3377.035 1243.275 3379.435 1243.310 ;
        RECT 3369.140 1218.910 3369.400 1219.230 ;
        RECT 3376.500 1218.910 3376.760 1219.230 ;
        RECT 208.940 1140.030 209.200 1140.350 ;
        RECT 213.080 1140.030 213.340 1140.350 ;
        RECT 214.000 1140.030 214.260 1140.350 ;
        RECT 209.000 1137.725 209.140 1140.030 ;
        RECT 208.565 1137.445 210.965 1137.725 ;
        RECT 213.140 924.450 213.280 1140.030 ;
        RECT 3369.200 1090.710 3369.340 1218.910 ;
        RECT 3369.140 1090.390 3369.400 1090.710 ;
        RECT 3369.140 1089.710 3369.400 1090.030 ;
        RECT 3369.200 1062.830 3369.340 1089.710 ;
        RECT 3368.680 1062.510 3368.940 1062.830 ;
        RECT 3369.140 1062.510 3369.400 1062.830 ;
        RECT 3368.740 1019.650 3368.880 1062.510 ;
        RECT 3368.680 1019.330 3368.940 1019.650 ;
        RECT 3376.960 1019.330 3377.220 1019.650 ;
        RECT 3368.740 1015.650 3368.880 1019.330 ;
        RECT 3377.020 1017.555 3377.160 1019.330 ;
        RECT 3377.020 1017.415 3379.435 1017.555 ;
        RECT 3377.035 1017.275 3379.435 1017.415 ;
        RECT 3367.820 1015.510 3368.880 1015.650 ;
        RECT 208.940 924.130 209.200 924.450 ;
        RECT 212.160 924.130 212.420 924.450 ;
        RECT 213.080 924.130 213.340 924.450 ;
        RECT 209.000 921.725 209.140 924.130 ;
        RECT 208.565 921.445 210.965 921.725 ;
        RECT 212.220 228.470 212.360 924.130 ;
        RECT 3367.820 791.850 3367.960 1015.510 ;
        RECT 3377.035 792.540 3379.435 792.555 ;
        RECT 3377.020 792.275 3379.435 792.540 ;
        RECT 3377.020 791.850 3377.160 792.275 ;
        RECT 3367.760 791.530 3368.020 791.850 ;
        RECT 3376.960 791.530 3377.220 791.850 ;
        RECT 3367.820 564.050 3367.960 791.530 ;
        RECT 3377.035 566.415 3379.435 566.555 ;
        RECT 3377.020 566.275 3379.435 566.415 ;
        RECT 3377.020 564.050 3377.160 566.275 ;
        RECT 3367.760 563.730 3368.020 564.050 ;
        RECT 3376.960 563.730 3377.220 564.050 ;
        RECT 212.160 228.150 212.420 228.470 ;
        RECT 718.160 228.150 718.420 228.470 ;
        RECT 718.220 222.010 718.360 228.150 ;
        RECT 3367.820 228.130 3367.960 563.730 ;
        RECT 2637.280 227.810 2637.540 228.130 ;
        RECT 3367.760 227.810 3368.020 228.130 ;
        RECT 718.160 221.690 718.420 222.010 ;
        RECT 725.520 221.690 725.780 222.010 ;
        RECT 976.680 221.690 976.940 222.010 ;
        RECT 998.300 221.690 998.560 222.010 ;
        RECT 725.580 201.010 725.720 221.690 ;
        RECT 976.740 210.965 976.880 221.690 ;
        RECT 998.360 221.330 998.500 221.690 ;
        RECT 1793.640 221.350 1793.900 221.670 ;
        RECT 2067.800 221.350 2068.060 221.670 ;
        RECT 2089.420 221.350 2089.680 221.670 ;
        RECT 2341.500 221.350 2341.760 221.670 ;
        RECT 2363.120 221.350 2363.380 221.670 ;
        RECT 2615.660 221.350 2615.920 221.670 ;
        RECT 998.300 221.010 998.560 221.330 ;
        RECT 1519.480 221.010 1519.740 221.330 ;
        RECT 1541.100 221.010 1541.360 221.330 ;
        RECT 998.360 210.965 998.500 221.010 ;
        RECT 1519.540 210.965 1519.680 221.010 ;
        RECT 1541.160 210.965 1541.300 221.010 ;
        RECT 1793.700 220.990 1793.840 221.350 ;
        RECT 1815.260 221.010 1815.520 221.330 ;
        RECT 1793.640 220.670 1793.900 220.990 ;
        RECT 1793.700 210.965 1793.840 220.670 ;
        RECT 1815.320 210.965 1815.460 221.010 ;
        RECT 2067.860 210.965 2068.000 221.350 ;
        RECT 2089.480 210.965 2089.620 221.350 ;
        RECT 976.655 208.565 976.935 210.965 ;
        RECT 998.275 208.565 998.555 210.965 ;
        RECT 1519.540 209.030 1519.935 210.965 ;
        RECT 1541.160 209.030 1541.555 210.965 ;
        RECT 1519.655 208.565 1519.935 209.030 ;
        RECT 1541.275 208.565 1541.555 209.030 ;
        RECT 1793.655 208.565 1793.935 210.965 ;
        RECT 1815.275 208.565 1815.555 210.965 ;
        RECT 2067.655 209.100 2068.000 210.965 ;
        RECT 2089.275 209.100 2089.620 210.965 ;
        RECT 2341.560 210.965 2341.700 221.350 ;
        RECT 2363.180 210.965 2363.320 221.350 ;
        RECT 2615.720 220.990 2615.860 221.350 ;
        RECT 2637.340 220.990 2637.480 227.810 ;
        RECT 2615.660 220.670 2615.920 220.990 ;
        RECT 2637.280 220.670 2637.540 220.990 ;
        RECT 2615.720 210.965 2615.860 220.670 ;
        RECT 2637.340 210.965 2637.480 220.670 ;
        RECT 2067.655 208.565 2067.935 209.100 ;
        RECT 2089.275 208.565 2089.555 209.100 ;
        RECT 2341.560 209.030 2341.935 210.965 ;
        RECT 2363.180 209.030 2363.555 210.965 ;
        RECT 2341.655 208.565 2341.935 209.030 ;
        RECT 2363.275 208.565 2363.555 209.030 ;
        RECT 2615.655 208.565 2615.935 210.965 ;
        RECT 2637.275 208.565 2637.555 210.965 ;
        RECT 725.515 200.870 725.720 201.010 ;
        RECT 725.515 200.000 725.655 200.870 ;
        RECT 725.455 198.530 725.715 200.000 ;
    END
  END porb_h
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.455 199.670 725.715 200.000 ;
    END
  END porb_h
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.750 91.545 ;
    END
  END resetb
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 708.335 190.155 709.065 200.000 ;
        RECT 708.335 189.855 709.365 190.155 ;
        RECT 708.335 189.555 709.100 189.855 ;
        RECT 709.365 189.555 709.830 189.855 ;
        RECT 708.335 189.090 709.830 189.555 ;
        RECT 709.100 185.230 709.830 189.090 ;
    END
  END resetb_core_h
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.335 199.670 709.065 200.000 ;
    END
  END resetb_core_h
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3396.885 4611.730 3401.535 4759.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 3489.900 4548.330 3557.165 4602.730 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3396.885 4390.730 3401.535 4539.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3396.985 4611.730 3401.435 4759.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3396.985 4390.730 3401.435 4539.270 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3390.000 4588.500 3396.900 4612.500 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3390.000 4538.300 3396.900 4562.245 ;
    END
  END vccd1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3402.935 4166.035 3406.385 4313.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 3493.120 4099.110 3553.945 4159.950 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3402.935 3945.035 3406.385 4092.965 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3403.035 4166.035 3406.285 4313.030 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3403.035 3945.035 3406.285 4092.965 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3388.000 4142.605 3402.960 4166.505 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 3376.470 4091.800 3376.790 4091.860 ;
        RECT 3387.510 4091.800 3387.830 4091.860 ;
        RECT 3376.470 4091.660 3387.830 4091.800 ;
        RECT 3376.470 4091.600 3376.790 4091.660 ;
        RECT 3387.510 4091.600 3387.830 4091.660 ;
        RECT 3376.470 3908.000 3376.790 3908.260 ;
        RECT 3376.560 3907.240 3376.700 3908.000 ;
        RECT 3376.470 3906.980 3376.790 3907.240 ;
        RECT 3376.010 3230.040 3376.330 3230.300 ;
        RECT 3376.100 3228.880 3376.240 3230.040 ;
        RECT 3376.470 3228.880 3376.790 3228.940 ;
        RECT 3376.100 3228.740 3376.790 3228.880 ;
        RECT 3376.470 3228.680 3376.790 3228.740 ;
        RECT 3376.470 2966.880 3376.790 2967.140 ;
        RECT 3376.560 2966.120 3376.700 2966.880 ;
        RECT 3376.470 2965.860 3376.790 2966.120 ;
        RECT 3376.470 2568.940 3376.790 2569.000 ;
        RECT 3388.430 2568.940 3388.750 2569.000 ;
        RECT 3376.470 2568.800 3388.750 2568.940 ;
        RECT 3376.470 2568.740 3376.790 2568.800 ;
        RECT 3388.430 2568.740 3388.750 2568.800 ;
      LAYER via ;
        RECT 3376.500 4091.600 3376.760 4091.860 ;
        RECT 3387.540 4091.600 3387.800 4091.860 ;
        RECT 3376.500 3908.000 3376.760 3908.260 ;
        RECT 3376.500 3906.980 3376.760 3907.240 ;
        RECT 3376.040 3230.040 3376.300 3230.300 ;
        RECT 3376.500 3228.680 3376.760 3228.940 ;
        RECT 3376.500 2966.880 3376.760 2967.140 ;
        RECT 3376.500 2965.860 3376.760 2966.120 ;
        RECT 3376.500 2568.740 3376.760 2569.000 ;
        RECT 3388.460 2568.740 3388.720 2569.000 ;
      LAYER met2 ;
        RECT 3376.500 4091.570 3376.760 4091.890 ;
        RECT 3387.530 4091.715 3387.810 4092.085 ;
        RECT 3387.540 4091.570 3387.800 4091.715 ;
        RECT 3376.560 3908.290 3376.700 4091.570 ;
        RECT 3376.500 3907.970 3376.760 3908.290 ;
        RECT 3376.500 3906.950 3376.760 3907.270 ;
        RECT 3376.560 3683.290 3376.700 3906.950 ;
        RECT 3376.100 3683.150 3376.700 3683.290 ;
        RECT 3376.100 3641.810 3376.240 3683.150 ;
        RECT 3376.100 3641.670 3376.700 3641.810 ;
        RECT 3376.560 3458.210 3376.700 3641.670 ;
        RECT 3376.100 3458.070 3376.700 3458.210 ;
        RECT 3376.100 3416.730 3376.240 3458.070 ;
        RECT 3376.100 3416.590 3376.700 3416.730 ;
        RECT 3376.560 3234.490 3376.700 3416.590 ;
        RECT 3376.100 3234.350 3376.700 3234.490 ;
        RECT 3376.100 3230.330 3376.240 3234.350 ;
        RECT 3376.040 3230.010 3376.300 3230.330 ;
        RECT 3376.500 3228.650 3376.760 3228.970 ;
        RECT 3376.560 2967.170 3376.700 3228.650 ;
        RECT 3376.500 2966.850 3376.760 2967.170 ;
        RECT 3376.500 2965.830 3376.760 2966.150 ;
        RECT 3376.560 2780.930 3376.700 2965.830 ;
        RECT 3376.100 2780.790 3376.700 2780.930 ;
        RECT 3376.100 2741.490 3376.240 2780.790 ;
        RECT 3376.100 2741.350 3376.700 2741.490 ;
        RECT 3376.560 2569.030 3376.700 2741.350 ;
        RECT 3376.500 2568.710 3376.760 2569.030 ;
        RECT 3388.460 2568.885 3388.720 2569.030 ;
        RECT 3388.450 2568.515 3388.730 2568.885 ;
      LAYER via2 ;
        RECT 3387.530 4091.760 3387.810 4092.040 ;
        RECT 3388.450 2568.560 3388.730 2568.840 ;
      LAYER met3 ;
        RECT 3388.000 4092.710 3402.960 4116.610 ;
        RECT 3387.505 4092.050 3387.835 4092.065 ;
        RECT 3388.670 4092.050 3388.970 4092.710 ;
        RECT 3387.505 4091.750 3388.970 4092.050 ;
        RECT 3387.505 4091.735 3387.835 4091.750 ;
        RECT 3388.000 2569.605 3402.960 2593.505 ;
        RECT 3388.670 2568.865 3388.970 2569.605 ;
        RECT 3388.425 2568.550 3388.970 2568.865 ;
        RECT 3388.425 2568.535 3388.755 2568.550 ;
        RECT 3388.000 2519.710 3402.960 2543.610 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2699.730 5024.735 2879.270 5028.185 ;
    END
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.945 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2668.090 5044.405 2879.270 5044.735 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2878.000 5039.645 2879.270 5040.825 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2668.090 5035.735 2879.270 5036.065 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2951.730 5024.735 3131.270 5028.185 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2951.730 5035.735 3132.610 5036.065 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2951.730 5044.405 3132.610 5044.735 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2951.730 5039.645 2953.000 5040.825 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2699.730 5024.840 2879.270 5028.085 ;
        RECT 2701.000 5024.835 2878.000 5024.840 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2699.730 5035.735 2879.270 5044.735 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2951.730 5024.840 3131.270 5028.085 ;
        RECT 2953.000 5024.835 3130.000 5024.840 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2951.730 5035.735 3131.270 5044.735 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2925.210 4961.180 2925.530 4961.240 ;
        RECT 3373.710 4961.180 3374.030 4961.240 ;
        RECT 2925.210 4961.040 3374.030 4961.180 ;
        RECT 2925.210 4960.980 2925.530 4961.040 ;
        RECT 3373.710 4960.980 3374.030 4961.040 ;
        RECT 3373.710 2139.180 3374.030 2139.240 ;
        RECT 3385.590 2139.180 3385.910 2139.240 ;
        RECT 3373.710 2139.040 3385.910 2139.180 ;
        RECT 3373.710 2138.980 3374.030 2139.040 ;
        RECT 3385.590 2138.980 3385.910 2139.040 ;
      LAYER via ;
        RECT 2925.240 4960.980 2925.500 4961.240 ;
        RECT 3373.740 4960.980 3374.000 4961.240 ;
        RECT 3373.740 2138.980 3374.000 2139.240 ;
        RECT 3385.620 2138.980 3385.880 2139.240 ;
      LAYER met2 ;
        RECT 2925.220 4986.895 2925.520 4987.285 ;
        RECT 2925.300 4961.270 2925.440 4986.895 ;
        RECT 2925.240 4960.950 2925.500 4961.270 ;
        RECT 3373.740 4960.950 3374.000 4961.270 ;
        RECT 3373.800 2139.270 3373.940 4960.950 ;
        RECT 3373.740 2138.950 3374.000 2139.270 ;
        RECT 3385.620 2139.180 3385.880 2139.270 ;
        RECT 3386.555 2139.180 3386.945 2139.260 ;
        RECT 3385.620 2139.040 3386.945 2139.180 ;
        RECT 3385.620 2138.950 3385.880 2139.040 ;
        RECT 3386.555 2138.960 3386.945 2139.040 ;
      LAYER via2 ;
        RECT 2925.220 4986.940 2925.520 4987.240 ;
        RECT 3386.600 2138.960 3386.900 2139.260 ;
      LAYER met3 ;
        RECT 2928.390 4988.000 2952.290 5024.760 ;
        RECT 2925.195 4987.230 2925.545 4987.265 ;
        RECT 2928.670 4987.230 2928.970 4988.000 ;
        RECT 2925.195 4986.930 2928.970 4987.230 ;
        RECT 2925.195 4986.915 2925.545 4986.930 ;
        RECT 3386.575 2139.260 3386.925 2139.285 ;
        RECT 3388.000 2139.260 3420.515 2152.505 ;
        RECT 3386.575 2138.960 3420.515 2139.260 ;
        RECT 3386.575 2138.935 3386.925 2138.960 ;
        RECT 3388.000 2128.605 3420.515 2138.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2878.495 4988.000 2902.395 5020.515 ;
    END
  END vssa1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3429.585 2372.730 3434.235 2520.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 3489.900 2309.330 3557.165 2363.730 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3429.585 2151.730 3434.235 2300.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3429.685 2372.730 3434.135 2520.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3429.685 2151.730 3434.135 2300.270 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3390.000 2349.500 3429.600 2373.500 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3390.000 2299.300 3429.600 2323.245 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 186.465 4422.730 191.115 4561.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 30.835 4570.270 98.100 4624.670 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 186.465 4633.730 191.115 4772.270 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 186.565 4422.730 191.015 4561.270 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 186.565 4633.730 191.015 4772.270 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 191.100 4560.500 198.000 4584.500 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 191.100 4610.755 198.000 4634.700 ;
    END
  END vccd2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 181.615 2278.035 185.065 2415.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 34.055 2422.050 94.880 2482.890 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 181.615 2489.035 185.065 2626.965 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 181.715 2278.035 184.965 2415.965 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 181.715 2489.035 184.965 2626.965 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 185.040 2415.495 200.000 2439.395 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 185.040 2465.390 200.000 2489.290 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 159.815 4000.730 163.265 4139.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 34.055 4145.050 94.880 4205.890 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.265 3969.090 143.595 4139.270 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.175 4138.000 148.355 4139.270 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.935 3969.090 152.265 4139.270 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 159.815 4211.730 163.265 4350.270 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.935 4211.730 152.265 4773.610 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.265 4211.730 143.595 4773.610 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.175 4211.730 148.355 4213.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 159.915 4138.000 163.160 4139.270 ;
        RECT 159.915 4002.000 163.165 4138.000 ;
        RECT 159.915 4000.730 163.160 4002.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 143.265 4000.730 152.265 4139.270 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 159.915 4349.000 163.160 4350.270 ;
        RECT 159.915 4213.000 163.165 4349.000 ;
        RECT 159.915 4211.730 163.160 4213.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 143.265 4211.730 152.265 4350.270 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 163.240 4188.390 200.000 4212.290 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 167.485 4138.495 200.000 4162.395 ;
    END
  END vssa2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 153.765 2066.730 158.415 2205.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 30.835 2214.270 98.100 2268.670 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 153.765 2277.730 158.415 2416.270 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 153.865 2066.730 158.315 2205.270 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 153.865 2277.730 158.315 2416.270 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.400 2204.500 198.000 2228.500 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.400 2254.755 198.000 2278.700 ;
    END
  END vssd2
  OBS
      LAYER nwell ;
        RECT 1678.860 4988.685 1737.965 4990.205 ;
        RECT 2889.860 4988.685 2948.965 4990.205 ;
        RECT 197.795 4360.860 199.315 4419.965 ;
      LAYER pwell ;
        RECT 176.080 4352.625 198.935 4360.155 ;
      LAYER nwell ;
        RECT 197.795 4149.860 199.315 4208.965 ;
      LAYER pwell ;
        RECT 3389.065 4155.845 3411.920 4163.375 ;
      LAYER nwell ;
        RECT 3388.685 4096.035 3390.205 4155.140 ;
      LAYER pwell ;
        RECT 3389.065 2582.845 3411.920 2590.375 ;
      LAYER nwell ;
        RECT 3388.685 2523.035 3390.205 2582.140 ;
        RECT 197.795 2426.860 199.315 2485.965 ;
      LAYER pwell ;
        RECT 176.080 2418.625 198.935 2426.155 ;
      LAYER nwell ;
        RECT 3388.685 2082.035 3390.205 2141.140 ;
        RECT 197.795 562.860 199.315 621.965 ;
      LAYER pwell ;
        RECT 176.080 554.625 198.935 562.155 ;
      LAYER nwell ;
        RECT 398.035 197.795 457.140 199.315 ;
        RECT 2849.035 197.795 2908.140 199.315 ;
        RECT 3118.035 197.795 3177.140 199.315 ;
      LAYER pwell ;
        RECT 3177.845 176.080 3185.375 198.935 ;
      LAYER li1 ;
        RECT 380.840 4988.230 461.160 5187.705 ;
        RECT 637.840 4988.230 718.160 5187.705 ;
        RECT 894.840 4988.230 975.160 5187.705 ;
        RECT 1151.840 4988.230 1232.160 5187.705 ;
        RECT 1409.840 4988.230 1490.160 5187.705 ;
        RECT 1668.070 4990.035 1739.775 5187.695 ;
        RECT 1679.065 4989.890 1680.045 4990.035 ;
        RECT 1736.760 4989.890 1737.650 4990.035 ;
        RECT 1679.065 4989.000 1737.650 4989.890 ;
        RECT 1918.840 4988.230 1999.160 5187.705 ;
        RECT 2363.840 4988.230 2444.160 5187.705 ;
        RECT 2620.840 4988.230 2701.160 5187.705 ;
        RECT 2879.070 4990.035 2950.775 5187.695 ;
        RECT 2890.065 4989.890 2891.045 4990.035 ;
        RECT 2947.760 4989.890 2948.650 4990.035 ;
        RECT 2890.065 4989.000 2948.650 4989.890 ;
        RECT 3129.840 4988.230 3210.160 5187.705 ;
        RECT 0.295 4770.840 199.770 4851.160 ;
        RECT 3388.230 4757.840 3587.705 4838.160 ;
        RECT 0.220 4560.240 196.980 4634.755 ;
        RECT 3391.020 4538.245 3587.780 4612.760 ;
        RECT 0.305 4419.680 197.965 4421.855 ;
        RECT 0.305 4418.730 199.030 4419.680 ;
        RECT 0.305 4362.045 197.965 4418.730 ;
        RECT 198.080 4362.045 199.030 4418.730 ;
        RECT 0.305 4361.035 199.030 4362.045 ;
        RECT 0.305 4360.155 197.965 4361.035 ;
        RECT 0.305 4349.610 198.935 4360.155 ;
        RECT 3388.230 4311.840 3587.705 4392.160 ;
        RECT 0.305 4208.650 197.965 4210.775 ;
        RECT 0.305 4207.760 199.000 4208.650 ;
        RECT 0.305 4151.045 197.965 4207.760 ;
        RECT 198.110 4151.045 199.000 4207.760 ;
        RECT 3389.065 4155.845 3587.695 4166.390 ;
        RECT 3390.035 4154.965 3587.695 4155.845 ;
        RECT 0.305 4150.065 199.000 4151.045 ;
        RECT 3388.970 4153.955 3587.695 4154.965 ;
        RECT 0.305 4139.070 197.965 4150.065 ;
        RECT 3388.970 4097.270 3389.920 4153.955 ;
        RECT 3390.035 4097.270 3587.695 4153.955 ;
        RECT 3388.970 4096.320 3587.695 4097.270 ;
        RECT 3390.035 4094.145 3587.695 4096.320 ;
        RECT 0.295 3921.840 199.770 4002.160 ;
        RECT 3388.230 3865.840 3587.705 3946.160 ;
        RECT 0.295 3705.840 199.770 3786.160 ;
        RECT 3388.230 3640.840 3587.705 3721.160 ;
        RECT 0.295 3489.840 199.770 3570.160 ;
        RECT 3388.230 3415.840 3587.705 3496.160 ;
        RECT 0.295 3273.840 199.770 3354.160 ;
        RECT 3388.230 3189.840 3587.705 3270.160 ;
        RECT 0.295 3057.840 199.770 3138.160 ;
        RECT 3388.230 2964.840 3587.705 3045.160 ;
        RECT 0.295 2841.840 199.770 2922.160 ;
        RECT 3388.230 2738.840 3587.705 2819.160 ;
        RECT 0.295 2625.840 199.770 2706.160 ;
        RECT 3389.065 2582.845 3587.695 2593.390 ;
        RECT 3390.035 2581.965 3587.695 2582.845 ;
        RECT 3388.970 2580.955 3587.695 2581.965 ;
        RECT 3388.970 2524.270 3389.920 2580.955 ;
        RECT 3390.035 2524.270 3587.695 2580.955 ;
        RECT 3388.970 2523.320 3587.695 2524.270 ;
        RECT 3390.035 2521.145 3587.695 2523.320 ;
        RECT 0.305 2485.680 197.965 2487.855 ;
        RECT 0.305 2484.730 199.030 2485.680 ;
        RECT 0.305 2428.045 197.965 2484.730 ;
        RECT 198.080 2428.045 199.030 2484.730 ;
        RECT 0.305 2427.035 199.030 2428.045 ;
        RECT 0.305 2426.155 197.965 2427.035 ;
        RECT 0.305 2415.610 198.935 2426.155 ;
        RECT 3391.020 2299.245 3587.780 2373.760 ;
        RECT 0.220 2204.240 196.980 2278.755 ;
        RECT 3390.035 2140.935 3587.695 2151.930 ;
        RECT 3389.000 2139.955 3587.695 2140.935 ;
        RECT 3389.000 2083.240 3389.890 2139.955 ;
        RECT 3390.035 2083.240 3587.695 2139.955 ;
        RECT 3389.000 2082.350 3587.695 2083.240 ;
        RECT 3390.035 2080.225 3587.695 2082.350 ;
        RECT 0.295 1987.840 199.770 2068.160 ;
        RECT 3388.230 1852.840 3587.705 1933.160 ;
        RECT 0.295 1771.840 199.770 1852.160 ;
        RECT 0.295 1555.840 199.770 1636.160 ;
        RECT 3388.230 1626.840 3587.705 1707.160 ;
        RECT 0.295 1339.840 199.770 1420.160 ;
        RECT 3388.230 1401.840 3587.705 1482.160 ;
        RECT 0.295 1123.840 199.770 1204.160 ;
        RECT 3388.230 1176.840 3587.705 1257.160 ;
        RECT 0.295 907.840 199.770 988.160 ;
        RECT 3388.230 950.840 3587.705 1031.160 ;
        RECT 3388.230 725.840 3587.705 806.160 ;
        RECT 0.305 621.680 197.965 623.855 ;
        RECT 0.305 620.730 199.030 621.680 ;
        RECT 0.305 564.045 197.965 620.730 ;
        RECT 198.080 564.045 199.030 620.730 ;
        RECT 0.305 563.035 199.030 564.045 ;
        RECT 0.305 562.155 197.965 563.035 ;
        RECT 0.305 551.610 198.935 562.155 ;
        RECT 3388.230 499.840 3587.705 580.160 ;
        RECT 0.220 340.240 196.980 414.755 ;
        RECT 398.350 198.110 456.935 199.000 ;
        RECT 398.350 197.965 399.240 198.110 ;
        RECT 455.955 197.965 456.935 198.110 ;
        RECT 396.225 0.305 467.930 197.965 ;
        RECT 663.000 0.780 738.000 199.815 ;
        RECT 931.840 0.295 1012.160 199.770 ;
        RECT 1206.245 0.220 1280.760 196.980 ;
        RECT 1474.840 0.295 1555.160 199.770 ;
        RECT 1748.840 0.295 1829.160 199.770 ;
        RECT 2022.840 0.295 2103.160 199.770 ;
        RECT 2296.840 0.295 2377.160 199.770 ;
        RECT 2570.840 0.295 2651.160 199.770 ;
        RECT 2849.350 198.110 2907.935 199.000 ;
        RECT 2849.350 197.965 2850.240 198.110 ;
        RECT 2906.955 197.965 2907.935 198.110 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.270 198.080 ;
        RECT 3175.955 197.965 3176.965 198.080 ;
        RECT 3177.845 197.965 3188.390 198.935 ;
        RECT 2847.225 0.305 2918.930 197.965 ;
        RECT 3116.145 0.305 3188.390 197.965 ;
      LAYER met1 ;
        RECT 380.855 4981.155 461.145 5188.000 ;
        RECT 637.855 4981.155 718.145 5188.000 ;
        RECT 894.855 4981.155 975.145 5188.000 ;
        RECT 1151.855 4981.155 1232.145 5188.000 ;
        RECT 1409.855 4981.155 1490.145 5188.000 ;
        RECT 1667.185 4990.035 1740.620 5187.725 ;
        RECT 1679.035 4989.920 1680.350 4990.035 ;
        POLYGON 1680.350 4990.035 1680.465 4989.920 1680.350 4989.920 ;
        POLYGON 1736.540 4990.035 1736.540 4989.920 1736.425 4989.920 ;
        RECT 1736.540 4989.920 1737.680 4990.035 ;
        RECT 1679.035 4988.970 1737.680 4989.920 ;
        RECT 1918.855 4981.155 1999.145 5188.000 ;
        RECT 2363.855 4981.155 2444.145 5188.000 ;
        RECT 2620.855 4981.155 2701.145 5188.000 ;
        RECT 2878.185 4990.035 2951.620 5187.725 ;
        RECT 2890.035 4989.920 2891.350 4990.035 ;
        POLYGON 2891.350 4990.035 2891.465 4989.920 2891.350 4989.920 ;
        POLYGON 2947.540 4990.035 2947.540 4989.920 2947.425 4989.920 ;
        RECT 2947.540 4989.920 2948.680 4990.035 ;
        RECT 2890.035 4988.970 2948.680 4989.920 ;
        RECT 3129.855 4981.155 3210.145 5188.000 ;
      LAYER met1 ;
        RECT 420.050 4978.180 420.370 4978.240 ;
        RECT 458.690 4978.180 459.010 4978.240 ;
        RECT 420.050 4978.040 459.010 4978.180 ;
        RECT 420.050 4977.980 420.370 4978.040 ;
        RECT 458.690 4977.980 459.010 4978.040 ;
        RECT 1191.010 4978.180 1191.330 4978.240 ;
        RECT 1229.650 4978.180 1229.970 4978.240 ;
        RECT 1191.010 4978.040 1229.970 4978.180 ;
        RECT 1191.010 4977.980 1191.330 4978.040 ;
        RECT 1229.650 4977.980 1229.970 4978.040 ;
        RECT 2659.790 4978.180 2660.110 4978.240 ;
        RECT 2698.430 4978.180 2698.750 4978.240 ;
        RECT 2659.790 4978.040 2698.750 4978.180 ;
        RECT 2659.790 4977.980 2660.110 4978.040 ;
        RECT 2698.430 4977.980 2698.750 4978.040 ;
        RECT 676.730 4977.500 677.050 4977.560 ;
        RECT 715.830 4977.500 716.150 4977.560 ;
        RECT 676.730 4977.360 716.150 4977.500 ;
        RECT 676.730 4977.300 677.050 4977.360 ;
        RECT 715.830 4977.300 716.150 4977.360 ;
        RECT 3169.010 4977.500 3169.330 4977.560 ;
        RECT 3207.650 4977.500 3207.970 4977.560 ;
        RECT 3169.010 4977.360 3207.970 4977.500 ;
        RECT 3169.010 4977.300 3169.330 4977.360 ;
        RECT 3207.650 4977.300 3207.970 4977.360 ;
        RECT 1448.150 4976.480 1448.470 4976.540 ;
        RECT 1488.170 4976.480 1488.490 4976.540 ;
        RECT 1448.150 4976.340 1488.490 4976.480 ;
        RECT 1448.150 4976.280 1448.470 4976.340 ;
        RECT 1488.170 4976.280 1488.490 4976.340 ;
        RECT 1957.370 4976.480 1957.690 4976.540 ;
        RECT 1997.390 4976.480 1997.710 4976.540 ;
        RECT 1957.370 4976.340 1997.710 4976.480 ;
        RECT 1957.370 4976.280 1957.690 4976.340 ;
        RECT 1997.390 4976.280 1997.710 4976.340 ;
        RECT 2402.190 4976.480 2402.510 4976.540 ;
        RECT 2442.210 4976.480 2442.530 4976.540 ;
        RECT 2402.190 4976.340 2442.530 4976.480 ;
        RECT 2402.190 4976.280 2402.510 4976.340 ;
        RECT 2442.210 4976.280 2442.530 4976.340 ;
        RECT 933.410 4953.020 933.730 4953.080 ;
        RECT 973.430 4953.020 973.750 4953.080 ;
        RECT 933.410 4952.880 973.750 4953.020 ;
        RECT 933.410 4952.820 933.730 4952.880 ;
        RECT 973.430 4952.820 973.750 4952.880 ;
      LAYER met1 ;
        RECT 0.000 4770.855 206.845 4851.145 ;
      LAYER met1 ;
        RECT 208.910 4846.940 209.230 4847.000 ;
        RECT 212.130 4846.940 212.450 4847.000 ;
        RECT 208.910 4846.800 212.450 4846.940 ;
        RECT 208.910 4846.740 209.230 4846.800 ;
        RECT 212.130 4846.740 212.450 4846.800 ;
        RECT 208.910 4812.260 209.230 4812.320 ;
        RECT 212.130 4812.260 212.450 4812.320 ;
        RECT 208.910 4812.120 212.450 4812.260 ;
        RECT 208.910 4812.060 209.230 4812.120 ;
        RECT 212.130 4812.060 212.450 4812.120 ;
      LAYER met1 ;
        RECT 3381.155 4757.855 3588.000 4838.145 ;
        RECT 159.640 4645.935 163.510 4646.195 ;
        RECT 159.640 4641.935 204.500 4645.935 ;
        POLYGON 204.500 4645.935 208.500 4641.935 204.500 4641.935 ;
        RECT 159.640 4636.200 208.500 4641.935 ;
        RECT 159.640 4635.245 163.510 4636.200 ;
        RECT 0.160 4616.565 197.965 4635.000 ;
        RECT 198.780 4616.565 208.500 4636.200 ;
        RECT 0.160 4580.495 208.500 4616.565 ;
        RECT 3390.035 4596.345 3587.840 4612.880 ;
        RECT 0.160 4576.655 198.000 4580.495 ;
        RECT 198.980 4578.655 208.500 4580.495 ;
        POLYGON 198.980 4578.655 200.980 4578.655 200.980 4576.655 ;
        RECT 200.980 4576.655 206.500 4578.655 ;
        POLYGON 206.500 4578.655 208.500 4578.655 206.500 4576.655 ;
        POLYGON 3381.500 4596.345 3381.500 4594.345 3379.500 4594.345 ;
        RECT 3381.500 4594.345 3387.020 4596.345 ;
        POLYGON 3387.020 4596.345 3389.020 4594.345 3387.020 4594.345 ;
        RECT 3379.500 4592.505 3389.020 4594.345 ;
        RECT 3390.000 4592.505 3587.840 4596.345 ;
        RECT 0.160 4560.120 197.965 4576.655 ;
        RECT 3379.500 4556.435 3587.840 4592.505 ;
        RECT 3379.500 4536.800 3389.220 4556.435 ;
        RECT 3390.035 4538.000 3587.840 4556.435 ;
        RECT 3424.490 4536.800 3428.360 4537.755 ;
        RECT 3379.500 4531.065 3428.360 4536.800 ;
        POLYGON 3379.500 4531.065 3383.500 4531.065 3383.500 4527.065 ;
        RECT 3383.500 4527.065 3428.360 4531.065 ;
        RECT 3424.490 4526.805 3428.360 4527.065 ;
        RECT 0.275 4419.680 197.965 4421.915 ;
        RECT 0.275 4418.540 199.030 4419.680 ;
        RECT 0.275 4362.350 197.965 4418.540 ;
        POLYGON 197.965 4418.540 198.080 4418.540 198.080 4418.425 ;
        POLYGON 198.080 4362.465 198.080 4362.350 197.965 4362.350 ;
        RECT 198.080 4362.350 199.030 4418.540 ;
        RECT 0.275 4361.035 199.030 4362.350 ;
        RECT 0.275 4357.855 197.965 4361.035 ;
        RECT 0.275 4352.625 198.870 4357.855 ;
        RECT 0.275 4349.185 197.965 4352.625 ;
      LAYER met1 ;
        RECT 3368.650 4350.880 3368.970 4350.940 ;
        RECT 3376.930 4350.880 3377.250 4350.940 ;
        RECT 3368.650 4350.740 3377.250 4350.880 ;
        RECT 3368.650 4350.680 3368.970 4350.740 ;
        RECT 3376.930 4350.680 3377.250 4350.740 ;
        RECT 3368.650 4316.200 3368.970 4316.260 ;
        RECT 3376.930 4316.200 3377.250 4316.260 ;
        RECT 3368.650 4316.060 3377.250 4316.200 ;
        RECT 3368.650 4316.000 3368.970 4316.060 ;
        RECT 3376.930 4316.000 3377.250 4316.060 ;
      LAYER met1 ;
        RECT 3381.155 4311.855 3588.000 4392.145 ;
        RECT 0.275 4208.680 197.965 4211.620 ;
        RECT 0.275 4207.540 199.030 4208.680 ;
        RECT 0.275 4151.350 197.965 4207.540 ;
        POLYGON 197.965 4207.540 198.080 4207.540 198.080 4207.425 ;
        POLYGON 198.080 4151.465 198.080 4151.350 197.965 4151.350 ;
        RECT 198.080 4151.350 199.030 4207.540 ;
        RECT 3390.035 4163.375 3587.725 4166.815 ;
        RECT 3389.130 4158.145 3587.725 4163.375 ;
        RECT 3390.035 4154.965 3587.725 4158.145 ;
        RECT 0.275 4150.035 199.030 4151.350 ;
        RECT 3388.970 4153.650 3587.725 4154.965 ;
        RECT 0.275 4138.185 197.965 4150.035 ;
        RECT 3388.970 4097.460 3389.920 4153.650 ;
        POLYGON 3389.920 4153.650 3390.035 4153.650 3389.920 4153.535 ;
        POLYGON 3389.920 4097.575 3390.035 4097.460 3389.920 4097.460 ;
        RECT 3390.035 4097.460 3587.725 4153.650 ;
        RECT 3388.970 4096.320 3587.725 4097.460 ;
        RECT 3390.035 4094.085 3587.725 4096.320 ;
        RECT 0.000 3921.855 206.845 4002.145 ;
      LAYER met1 ;
        RECT 208.910 3997.960 209.230 3998.020 ;
        RECT 211.670 3997.960 211.990 3998.020 ;
        RECT 208.910 3997.820 211.990 3997.960 ;
        RECT 208.910 3997.760 209.230 3997.820 ;
        RECT 211.670 3997.760 211.990 3997.820 ;
        RECT 208.910 3962.940 209.230 3963.000 ;
        RECT 211.670 3962.940 211.990 3963.000 ;
        RECT 208.910 3962.800 211.990 3962.940 ;
        RECT 208.910 3962.740 209.230 3962.800 ;
        RECT 211.670 3962.740 211.990 3962.800 ;
        RECT 3376.010 3870.120 3376.330 3870.180 ;
        RECT 3376.930 3870.120 3377.250 3870.180 ;
        RECT 3376.010 3869.980 3377.250 3870.120 ;
        RECT 3376.010 3869.920 3376.330 3869.980 ;
        RECT 3376.930 3869.920 3377.250 3869.980 ;
      LAYER met1 ;
        RECT 3381.155 3865.855 3588.000 3946.145 ;
        RECT 0.000 3705.855 206.845 3786.145 ;
      LAYER met1 ;
        RECT 208.910 3782.060 209.230 3782.120 ;
        RECT 211.670 3782.060 211.990 3782.120 ;
        RECT 208.910 3781.920 211.990 3782.060 ;
        RECT 208.910 3781.860 209.230 3781.920 ;
        RECT 211.670 3781.860 211.990 3781.920 ;
        RECT 208.910 3747.040 209.230 3747.100 ;
        RECT 211.670 3747.040 211.990 3747.100 ;
        RECT 208.910 3746.900 211.990 3747.040 ;
        RECT 208.910 3746.840 209.230 3746.900 ;
        RECT 211.670 3746.840 211.990 3746.900 ;
      LAYER met1 ;
        RECT 3381.155 3640.855 3588.000 3721.145 ;
        RECT 0.000 3489.855 206.845 3570.145 ;
      LAYER met1 ;
        RECT 208.910 3565.820 209.230 3565.880 ;
        RECT 211.670 3565.820 211.990 3565.880 ;
        RECT 208.910 3565.680 211.990 3565.820 ;
        RECT 208.910 3565.620 209.230 3565.680 ;
        RECT 211.670 3565.620 211.990 3565.680 ;
        RECT 208.910 3531.140 209.230 3531.200 ;
        RECT 211.670 3531.140 211.990 3531.200 ;
        RECT 208.910 3531.000 211.990 3531.140 ;
        RECT 208.910 3530.940 209.230 3531.000 ;
        RECT 211.670 3530.940 211.990 3531.000 ;
      LAYER met1 ;
        RECT 3381.155 3415.855 3588.000 3496.145 ;
        RECT 0.000 3273.855 206.845 3354.145 ;
      LAYER met1 ;
        RECT 208.910 3349.920 209.230 3349.980 ;
        RECT 211.670 3349.920 211.990 3349.980 ;
        RECT 208.910 3349.780 211.990 3349.920 ;
        RECT 208.910 3349.720 209.230 3349.780 ;
        RECT 211.670 3349.720 211.990 3349.780 ;
        RECT 208.910 3315.240 209.230 3315.300 ;
        RECT 211.670 3315.240 211.990 3315.300 ;
        RECT 208.910 3315.100 211.990 3315.240 ;
        RECT 208.910 3315.040 209.230 3315.100 ;
        RECT 211.670 3315.040 211.990 3315.100 ;
        RECT 3376.010 3194.200 3376.330 3194.260 ;
        RECT 3376.930 3194.200 3377.250 3194.260 ;
        RECT 3376.010 3194.060 3377.250 3194.200 ;
        RECT 3376.010 3194.000 3376.330 3194.060 ;
        RECT 3376.930 3194.000 3377.250 3194.060 ;
      LAYER met1 ;
        RECT 3381.155 3189.855 3588.000 3270.145 ;
        RECT 0.000 3057.855 206.845 3138.145 ;
      LAYER met1 ;
        RECT 208.910 3134.020 209.230 3134.080 ;
        RECT 211.670 3134.020 211.990 3134.080 ;
        RECT 208.910 3133.880 211.990 3134.020 ;
        RECT 208.910 3133.820 209.230 3133.880 ;
        RECT 211.670 3133.820 211.990 3133.880 ;
        RECT 208.910 3099.000 209.230 3099.060 ;
        RECT 211.670 3099.000 211.990 3099.060 ;
        RECT 208.910 3098.860 211.990 3099.000 ;
        RECT 208.910 3098.800 209.230 3098.860 ;
        RECT 211.670 3098.800 211.990 3098.860 ;
        RECT 3376.010 3004.140 3376.330 3004.200 ;
        RECT 3376.930 3004.140 3377.250 3004.200 ;
        RECT 3376.010 3004.000 3377.250 3004.140 ;
        RECT 3376.010 3003.940 3376.330 3004.000 ;
        RECT 3376.930 3003.940 3377.250 3004.000 ;
      LAYER met1 ;
        RECT 3381.155 2964.855 3588.000 3045.145 ;
        RECT 0.000 2841.855 206.845 2922.145 ;
      LAYER met1 ;
        RECT 208.910 2917.780 209.230 2917.840 ;
        RECT 211.670 2917.780 211.990 2917.840 ;
        RECT 208.910 2917.640 211.990 2917.780 ;
        RECT 208.910 2917.580 209.230 2917.640 ;
        RECT 211.670 2917.580 211.990 2917.640 ;
        RECT 208.910 2883.100 209.230 2883.160 ;
        RECT 211.670 2883.100 211.990 2883.160 ;
        RECT 208.910 2882.960 211.990 2883.100 ;
        RECT 208.910 2882.900 209.230 2882.960 ;
        RECT 211.670 2882.900 211.990 2882.960 ;
      LAYER met1 ;
        RECT 3381.155 2738.855 3588.000 2819.145 ;
        RECT 0.000 2625.855 206.845 2706.145 ;
      LAYER met1 ;
        RECT 208.910 2701.880 209.230 2701.940 ;
        RECT 211.670 2701.880 211.990 2701.940 ;
        RECT 208.910 2701.740 211.990 2701.880 ;
        RECT 208.910 2701.680 209.230 2701.740 ;
        RECT 211.670 2701.680 211.990 2701.740 ;
        RECT 208.910 2667.200 209.230 2667.260 ;
        RECT 211.670 2667.200 211.990 2667.260 ;
        RECT 208.910 2667.060 211.990 2667.200 ;
        RECT 208.910 2667.000 209.230 2667.060 ;
        RECT 211.670 2667.000 211.990 2667.060 ;
      LAYER met1 ;
        RECT 3390.035 2590.375 3587.725 2593.815 ;
        RECT 3389.130 2585.145 3587.725 2590.375 ;
        RECT 3390.035 2581.965 3587.725 2585.145 ;
        RECT 3388.970 2580.650 3587.725 2581.965 ;
        RECT 3388.970 2524.460 3389.920 2580.650 ;
        POLYGON 3389.920 2580.650 3390.035 2580.650 3389.920 2580.535 ;
        POLYGON 3389.920 2524.575 3390.035 2524.460 3389.920 2524.460 ;
        RECT 3390.035 2524.460 3587.725 2580.650 ;
        RECT 3388.970 2523.320 3587.725 2524.460 ;
        RECT 3390.035 2521.085 3587.725 2523.320 ;
        RECT 0.275 2485.680 197.965 2487.915 ;
        RECT 0.275 2484.540 199.030 2485.680 ;
        RECT 0.275 2428.350 197.965 2484.540 ;
        POLYGON 197.965 2484.540 198.080 2484.540 198.080 2484.425 ;
        POLYGON 198.080 2428.465 198.080 2428.350 197.965 2428.350 ;
        RECT 198.080 2428.350 199.030 2484.540 ;
        RECT 0.275 2427.035 199.030 2428.350 ;
        RECT 0.275 2423.855 197.965 2427.035 ;
        RECT 0.275 2418.625 198.870 2423.855 ;
        RECT 0.275 2415.185 197.965 2418.625 ;
        RECT 3390.035 2357.345 3587.840 2373.880 ;
        POLYGON 3381.500 2357.345 3381.500 2355.345 3379.500 2355.345 ;
        RECT 3381.500 2355.345 3387.020 2357.345 ;
        POLYGON 3387.020 2357.345 3389.020 2355.345 3387.020 2355.345 ;
        RECT 3379.500 2353.505 3389.020 2355.345 ;
        RECT 3390.000 2353.505 3587.840 2357.345 ;
        RECT 3379.500 2317.435 3587.840 2353.505 ;
        RECT 3379.500 2297.800 3389.220 2317.435 ;
        RECT 3390.035 2299.000 3587.840 2317.435 ;
        RECT 3424.490 2297.800 3428.360 2298.755 ;
        RECT 3379.500 2292.065 3428.360 2297.800 ;
        POLYGON 3379.500 2292.065 3381.370 2292.065 3381.370 2290.195 ;
        RECT 3381.370 2290.195 3428.360 2292.065 ;
        RECT 159.640 2289.935 163.510 2290.195 ;
        POLYGON 3381.370 2290.195 3381.630 2290.195 3381.630 2289.935 ;
        RECT 3381.630 2289.935 3428.360 2290.195 ;
        RECT 159.640 2285.935 204.500 2289.935 ;
        POLYGON 204.500 2289.935 208.500 2285.935 204.500 2285.935 ;
        POLYGON 3381.630 2289.935 3383.500 2289.935 3383.500 2288.065 ;
        RECT 3383.500 2288.065 3428.360 2289.935 ;
        RECT 3424.490 2287.805 3428.360 2288.065 ;
        RECT 159.640 2280.200 208.500 2285.935 ;
        RECT 159.640 2279.245 163.510 2280.200 ;
        RECT 0.160 2260.565 197.965 2279.000 ;
        RECT 198.780 2260.565 208.500 2280.200 ;
        RECT 0.160 2224.495 208.500 2260.565 ;
        RECT 0.160 2220.655 198.000 2224.495 ;
        RECT 198.980 2222.655 208.500 2224.495 ;
        POLYGON 198.980 2222.655 200.980 2222.655 200.980 2220.655 ;
        RECT 200.980 2220.655 206.500 2222.655 ;
        POLYGON 206.500 2222.655 208.500 2222.655 206.500 2220.655 ;
        RECT 0.160 2204.120 197.965 2220.655 ;
        RECT 3390.035 2140.965 3587.725 2152.815 ;
        RECT 3388.970 2139.650 3587.725 2140.965 ;
        RECT 3388.970 2083.460 3389.920 2139.650 ;
        POLYGON 3389.920 2139.650 3390.035 2139.650 3389.920 2139.535 ;
        POLYGON 3389.920 2083.575 3390.035 2083.460 3389.920 2083.460 ;
        RECT 3390.035 2083.460 3587.725 2139.650 ;
        RECT 3388.970 2082.320 3587.725 2083.460 ;
        RECT 3390.035 2079.380 3587.725 2082.320 ;
        RECT 0.000 1987.855 206.845 2068.145 ;
      LAYER met1 ;
        RECT 208.910 2064.040 209.230 2064.100 ;
        RECT 211.670 2064.040 211.990 2064.100 ;
        RECT 208.910 2063.900 211.990 2064.040 ;
        RECT 208.910 2063.840 209.230 2063.900 ;
        RECT 211.670 2063.840 211.990 2063.900 ;
        RECT 208.910 2029.020 209.230 2029.080 ;
        RECT 211.670 2029.020 211.990 2029.080 ;
        RECT 208.910 2028.880 211.990 2029.020 ;
        RECT 208.910 2028.820 209.230 2028.880 ;
        RECT 211.670 2028.820 211.990 2028.880 ;
      LAYER met1 ;
        RECT 3381.155 1852.855 3588.000 1933.145 ;
        RECT 0.000 1771.855 206.845 1852.145 ;
      LAYER met1 ;
        RECT 208.910 1847.800 209.230 1847.860 ;
        RECT 211.670 1847.800 211.990 1847.860 ;
        RECT 208.910 1847.660 211.990 1847.800 ;
        RECT 208.910 1847.600 209.230 1847.660 ;
        RECT 211.670 1847.600 211.990 1847.660 ;
        RECT 208.910 1813.120 209.230 1813.180 ;
        RECT 211.670 1813.120 211.990 1813.180 ;
        RECT 208.910 1812.980 211.990 1813.120 ;
        RECT 208.910 1812.920 209.230 1812.980 ;
        RECT 211.670 1812.920 211.990 1812.980 ;
      LAYER met1 ;
        RECT 0.000 1555.855 206.845 1636.145 ;
      LAYER met1 ;
        RECT 208.910 1631.900 209.230 1631.960 ;
        RECT 211.670 1631.900 211.990 1631.960 ;
        RECT 208.910 1631.760 211.990 1631.900 ;
        RECT 208.910 1631.700 209.230 1631.760 ;
        RECT 211.670 1631.700 211.990 1631.760 ;
      LAYER met1 ;
        RECT 3381.155 1626.855 3588.000 1707.145 ;
      LAYER met1 ;
        RECT 208.910 1597.220 209.230 1597.280 ;
        RECT 211.670 1597.220 211.990 1597.280 ;
        RECT 208.910 1597.080 211.990 1597.220 ;
        RECT 208.910 1597.020 209.230 1597.080 ;
        RECT 211.670 1597.020 211.990 1597.080 ;
      LAYER met1 ;
        RECT 0.000 1339.855 206.845 1420.145 ;
      LAYER met1 ;
        RECT 208.910 1416.000 209.230 1416.060 ;
        RECT 211.670 1416.000 211.990 1416.060 ;
        RECT 208.910 1415.860 211.990 1416.000 ;
        RECT 208.910 1415.800 209.230 1415.860 ;
        RECT 211.670 1415.800 211.990 1415.860 ;
      LAYER met1 ;
        RECT 3381.155 1401.855 3588.000 1482.145 ;
      LAYER met1 ;
        RECT 208.910 1380.980 209.230 1381.040 ;
        RECT 211.670 1380.980 211.990 1381.040 ;
        RECT 208.910 1380.840 211.990 1380.980 ;
        RECT 208.910 1380.780 209.230 1380.840 ;
        RECT 211.670 1380.780 211.990 1380.840 ;
      LAYER met1 ;
        RECT 0.000 1123.855 206.845 1204.145 ;
      LAYER met1 ;
        RECT 208.910 1199.760 209.230 1199.820 ;
        RECT 211.670 1199.760 211.990 1199.820 ;
        RECT 208.910 1199.620 211.990 1199.760 ;
        RECT 208.910 1199.560 209.230 1199.620 ;
        RECT 211.670 1199.560 211.990 1199.620 ;
      LAYER met1 ;
        RECT 3381.155 1176.855 3588.000 1257.145 ;
      LAYER met1 ;
        RECT 208.910 1165.080 209.230 1165.140 ;
        RECT 211.670 1165.080 211.990 1165.140 ;
        RECT 208.910 1164.940 211.990 1165.080 ;
        RECT 208.910 1164.880 209.230 1164.940 ;
        RECT 211.670 1164.880 211.990 1164.940 ;
      LAYER met1 ;
        RECT 0.000 907.855 206.845 988.145 ;
      LAYER met1 ;
        RECT 208.910 983.860 209.230 983.920 ;
        RECT 211.670 983.860 211.990 983.920 ;
        RECT 208.910 983.720 211.990 983.860 ;
        RECT 208.910 983.660 209.230 983.720 ;
        RECT 211.670 983.660 211.990 983.720 ;
      LAYER met1 ;
        RECT 3381.155 950.855 3588.000 1031.145 ;
      LAYER met1 ;
        RECT 208.910 949.180 209.230 949.240 ;
        RECT 211.670 949.180 211.990 949.240 ;
        RECT 208.910 949.040 211.990 949.180 ;
        RECT 208.910 948.980 209.230 949.040 ;
        RECT 211.670 948.980 211.990 949.040 ;
      LAYER met1 ;
        RECT 3381.155 725.855 3588.000 806.145 ;
        RECT 0.275 621.680 197.965 623.915 ;
        RECT 0.275 620.540 199.030 621.680 ;
        RECT 0.275 564.350 197.965 620.540 ;
        POLYGON 197.965 620.540 198.080 620.540 198.080 620.425 ;
        POLYGON 198.080 564.465 198.080 564.350 197.965 564.350 ;
        RECT 198.080 564.350 199.030 620.540 ;
        RECT 0.275 563.035 199.030 564.350 ;
        RECT 0.275 559.855 197.965 563.035 ;
        RECT 0.275 554.625 198.870 559.855 ;
        RECT 0.275 551.185 197.965 554.625 ;
        RECT 3381.155 499.855 3588.000 580.145 ;
        RECT 122.615 421.935 204.885 425.935 ;
        POLYGON 204.885 425.935 208.885 421.935 204.885 421.935 ;
        RECT 122.615 416.200 208.885 421.935 ;
        RECT 0.160 396.565 197.965 415.000 ;
        RECT 198.780 396.565 208.885 416.200 ;
        RECT 0.160 360.925 208.885 396.565 ;
        RECT 0.160 356.655 198.000 360.925 ;
        RECT 0.160 340.120 197.965 356.655 ;
      LAYER met1 ;
        RECT 933.410 221.240 933.730 221.300 ;
        RECT 973.430 221.240 973.750 221.300 ;
        RECT 933.410 221.100 973.750 221.240 ;
        RECT 933.410 221.040 933.730 221.100 ;
        RECT 973.430 221.040 973.750 221.100 ;
        RECT 1476.210 220.900 1476.530 220.960 ;
        RECT 1516.230 220.900 1516.550 220.960 ;
        RECT 1476.210 220.760 1516.550 220.900 ;
        RECT 1476.210 220.700 1476.530 220.760 ;
        RECT 1516.230 220.700 1516.550 220.760 ;
        RECT 1750.370 220.900 1750.690 220.960 ;
        RECT 1790.390 220.900 1790.710 220.960 ;
        RECT 1750.370 220.760 1790.710 220.900 ;
        RECT 1750.370 220.700 1750.690 220.760 ;
        RECT 1790.390 220.700 1790.710 220.760 ;
        RECT 2024.530 220.900 2024.850 220.960 ;
        RECT 2064.550 220.900 2064.870 220.960 ;
        RECT 2024.530 220.760 2064.870 220.900 ;
        RECT 2024.530 220.700 2024.850 220.760 ;
        RECT 2064.550 220.700 2064.870 220.760 ;
        RECT 2298.230 220.900 2298.550 220.960 ;
        RECT 2338.250 220.900 2338.570 220.960 ;
        RECT 2298.230 220.760 2338.570 220.900 ;
        RECT 2298.230 220.700 2298.550 220.760 ;
        RECT 2338.250 220.700 2338.570 220.760 ;
        RECT 2572.390 220.900 2572.710 220.960 ;
        RECT 2612.410 220.900 2612.730 220.960 ;
        RECT 2572.390 220.760 2612.730 220.900 ;
        RECT 2572.390 220.700 2572.710 220.760 ;
        RECT 2612.410 220.700 2612.730 220.760 ;
      LAYER met1 ;
        POLYGON 1199.065 208.885 1199.065 206.845 1197.025 206.845 ;
        RECT 1199.065 206.845 1260.075 208.885 ;
      LAYER met1 ;
        RECT 675.810 201.180 676.130 201.240 ;
        RECT 717.670 201.180 717.990 201.240 ;
        RECT 675.810 201.040 717.990 201.180 ;
        RECT 675.810 200.980 676.130 201.040 ;
        RECT 717.670 200.980 717.990 201.040 ;
      LAYER met1 ;
        RECT 663.000 199.390 704.700 199.815 ;
      LAYER met1 ;
        RECT 704.980 199.670 705.240 200.000 ;
      LAYER met1 ;
        RECT 705.520 199.390 706.565 199.815 ;
      LAYER met1 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met1 ;
        RECT 707.775 199.390 709.490 199.815 ;
      LAYER met1 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met1 ;
        RECT 710.700 199.390 712.585 199.815 ;
        RECT 398.320 198.080 456.965 199.030 ;
        RECT 398.320 197.965 399.460 198.080 ;
        POLYGON 399.460 198.080 399.575 198.080 399.460 197.965 ;
        POLYGON 455.535 198.080 455.650 198.080 455.650 197.965 ;
        RECT 455.650 197.965 456.965 198.080 ;
        RECT 395.380 0.275 468.815 197.965 ;
        RECT 663.000 189.745 712.585 199.390 ;
        RECT 713.375 199.390 715.060 199.815 ;
      LAYER met1 ;
        RECT 715.340 199.670 715.640 200.000 ;
      LAYER met1 ;
        RECT 715.920 199.390 722.585 199.815 ;
      LAYER met1 ;
        RECT 722.865 199.670 723.445 200.000 ;
      LAYER met1 ;
        RECT 723.725 199.390 725.175 199.815 ;
        RECT 725.995 199.390 738.000 199.815 ;
        RECT 713.375 189.745 738.000 199.390 ;
        RECT 663.000 0.790 738.000 189.745 ;
        RECT 931.855 0.000 1012.145 206.845 ;
        POLYGON 1197.025 206.845 1197.025 204.885 1195.065 204.885 ;
        RECT 1197.025 204.885 1260.075 206.845 ;
        RECT 1195.065 198.780 1260.075 204.885 ;
        RECT 1195.065 122.615 1204.800 198.780 ;
        RECT 1224.435 198.000 1260.075 198.780 ;
        RECT 1224.435 197.965 1264.345 198.000 ;
        RECT 1206.000 0.160 1280.880 197.965 ;
        RECT 1474.855 0.000 1555.145 206.845 ;
        RECT 1748.855 0.000 1829.145 206.845 ;
        RECT 2022.855 0.000 2103.145 206.845 ;
        RECT 2296.855 0.000 2377.145 206.845 ;
        RECT 2570.855 0.000 2651.145 206.845 ;
        RECT 2849.320 198.080 2907.965 199.030 ;
        RECT 2849.320 197.965 2850.460 198.080 ;
        POLYGON 2850.460 198.080 2850.575 198.080 2850.460 197.965 ;
        POLYGON 2906.535 198.080 2906.650 198.080 2906.650 197.965 ;
        RECT 2906.650 197.965 2907.965 198.080 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.460 198.080 ;
        POLYGON 3119.460 198.080 3119.575 198.080 3119.460 197.965 ;
        POLYGON 3175.535 198.080 3175.650 198.080 3175.650 197.965 ;
        RECT 3175.650 197.965 3176.965 198.080 ;
        RECT 3180.145 197.965 3185.375 198.870 ;
        RECT 2846.380 0.275 2919.815 197.965 ;
        RECT 3116.085 0.275 3188.815 197.965 ;
      LAYER via ;
        RECT 420.080 4977.980 420.340 4978.240 ;
        RECT 458.720 4977.980 458.980 4978.240 ;
        RECT 1191.040 4977.980 1191.300 4978.240 ;
        RECT 1229.680 4977.980 1229.940 4978.240 ;
        RECT 2659.820 4977.980 2660.080 4978.240 ;
        RECT 2698.460 4977.980 2698.720 4978.240 ;
        RECT 676.760 4977.300 677.020 4977.560 ;
        RECT 715.860 4977.300 716.120 4977.560 ;
        RECT 3169.040 4977.300 3169.300 4977.560 ;
        RECT 3207.680 4977.300 3207.940 4977.560 ;
        RECT 1448.180 4976.280 1448.440 4976.540 ;
        RECT 1488.200 4976.280 1488.460 4976.540 ;
        RECT 1957.400 4976.280 1957.660 4976.540 ;
        RECT 1997.420 4976.280 1997.680 4976.540 ;
        RECT 2402.220 4976.280 2402.480 4976.540 ;
        RECT 2442.240 4976.280 2442.500 4976.540 ;
        RECT 933.440 4952.820 933.700 4953.080 ;
        RECT 973.460 4952.820 973.720 4953.080 ;
        RECT 208.940 4846.740 209.200 4847.000 ;
        RECT 212.160 4846.740 212.420 4847.000 ;
        RECT 208.940 4812.060 209.200 4812.320 ;
        RECT 212.160 4812.060 212.420 4812.320 ;
        RECT 3368.680 4350.680 3368.940 4350.940 ;
        RECT 3376.960 4350.680 3377.220 4350.940 ;
        RECT 3368.680 4316.000 3368.940 4316.260 ;
        RECT 3376.960 4316.000 3377.220 4316.260 ;
        RECT 208.940 3997.760 209.200 3998.020 ;
        RECT 211.700 3997.760 211.960 3998.020 ;
        RECT 208.940 3962.740 209.200 3963.000 ;
        RECT 211.700 3962.740 211.960 3963.000 ;
        RECT 3376.040 3869.920 3376.300 3870.180 ;
        RECT 3376.960 3869.920 3377.220 3870.180 ;
        RECT 208.940 3781.860 209.200 3782.120 ;
        RECT 211.700 3781.860 211.960 3782.120 ;
        RECT 208.940 3746.840 209.200 3747.100 ;
        RECT 211.700 3746.840 211.960 3747.100 ;
        RECT 208.940 3565.620 209.200 3565.880 ;
        RECT 211.700 3565.620 211.960 3565.880 ;
        RECT 208.940 3530.940 209.200 3531.200 ;
        RECT 211.700 3530.940 211.960 3531.200 ;
        RECT 208.940 3349.720 209.200 3349.980 ;
        RECT 211.700 3349.720 211.960 3349.980 ;
        RECT 208.940 3315.040 209.200 3315.300 ;
        RECT 211.700 3315.040 211.960 3315.300 ;
        RECT 3376.040 3194.000 3376.300 3194.260 ;
        RECT 3376.960 3194.000 3377.220 3194.260 ;
        RECT 208.940 3133.820 209.200 3134.080 ;
        RECT 211.700 3133.820 211.960 3134.080 ;
        RECT 208.940 3098.800 209.200 3099.060 ;
        RECT 211.700 3098.800 211.960 3099.060 ;
        RECT 3376.040 3003.940 3376.300 3004.200 ;
        RECT 3376.960 3003.940 3377.220 3004.200 ;
        RECT 208.940 2917.580 209.200 2917.840 ;
        RECT 211.700 2917.580 211.960 2917.840 ;
        RECT 208.940 2882.900 209.200 2883.160 ;
        RECT 211.700 2882.900 211.960 2883.160 ;
        RECT 208.940 2701.680 209.200 2701.940 ;
        RECT 211.700 2701.680 211.960 2701.940 ;
        RECT 208.940 2667.000 209.200 2667.260 ;
        RECT 211.700 2667.000 211.960 2667.260 ;
        RECT 208.940 2063.840 209.200 2064.100 ;
        RECT 211.700 2063.840 211.960 2064.100 ;
        RECT 208.940 2028.820 209.200 2029.080 ;
        RECT 211.700 2028.820 211.960 2029.080 ;
        RECT 208.940 1847.600 209.200 1847.860 ;
        RECT 211.700 1847.600 211.960 1847.860 ;
        RECT 208.940 1812.920 209.200 1813.180 ;
        RECT 211.700 1812.920 211.960 1813.180 ;
        RECT 208.940 1631.700 209.200 1631.960 ;
        RECT 211.700 1631.700 211.960 1631.960 ;
        RECT 208.940 1597.020 209.200 1597.280 ;
        RECT 211.700 1597.020 211.960 1597.280 ;
        RECT 208.940 1415.800 209.200 1416.060 ;
        RECT 211.700 1415.800 211.960 1416.060 ;
        RECT 208.940 1380.780 209.200 1381.040 ;
        RECT 211.700 1380.780 211.960 1381.040 ;
        RECT 208.940 1199.560 209.200 1199.820 ;
        RECT 211.700 1199.560 211.960 1199.820 ;
        RECT 208.940 1164.880 209.200 1165.140 ;
        RECT 211.700 1164.880 211.960 1165.140 ;
        RECT 208.940 983.660 209.200 983.920 ;
        RECT 211.700 983.660 211.960 983.920 ;
        RECT 208.940 948.980 209.200 949.240 ;
        RECT 211.700 948.980 211.960 949.240 ;
        RECT 933.440 221.040 933.700 221.300 ;
        RECT 973.460 221.040 973.720 221.300 ;
        RECT 1476.240 220.700 1476.500 220.960 ;
        RECT 1516.260 220.700 1516.520 220.960 ;
        RECT 1750.400 220.700 1750.660 220.960 ;
        RECT 1790.420 220.700 1790.680 220.960 ;
        RECT 2024.560 220.700 2024.820 220.960 ;
        RECT 2064.580 220.700 2064.840 220.960 ;
        RECT 2298.260 220.700 2298.520 220.960 ;
        RECT 2338.280 220.700 2338.540 220.960 ;
        RECT 2572.420 220.700 2572.680 220.960 ;
        RECT 2612.440 220.700 2612.700 220.960 ;
        RECT 675.840 200.980 676.100 201.240 ;
        RECT 717.700 200.980 717.960 201.240 ;
      LAYER met2 ;
        RECT 381.210 4979.715 460.915 5188.000 ;
        RECT 381.210 4979.435 382.205 4979.715 ;
        RECT 383.045 4979.435 384.965 4979.715 ;
        RECT 385.805 4979.435 388.185 4979.715 ;
        RECT 389.025 4979.435 391.405 4979.715 ;
        RECT 392.245 4979.435 394.165 4979.715 ;
        RECT 395.005 4979.435 397.385 4979.715 ;
        RECT 398.225 4979.435 400.605 4979.715 ;
        RECT 401.445 4979.435 403.365 4979.715 ;
        RECT 404.205 4979.435 406.585 4979.715 ;
        RECT 407.425 4979.435 409.805 4979.715 ;
        RECT 410.645 4979.435 412.565 4979.715 ;
        RECT 413.405 4979.435 415.785 4979.715 ;
        RECT 416.625 4979.435 419.005 4979.715 ;
        RECT 419.845 4979.435 422.225 4979.715 ;
        RECT 423.065 4979.435 424.985 4979.715 ;
        RECT 425.825 4979.435 428.205 4979.715 ;
        RECT 429.045 4979.435 431.425 4979.715 ;
        RECT 432.265 4979.435 434.185 4979.715 ;
        RECT 435.025 4979.435 437.405 4979.715 ;
        RECT 438.245 4979.435 440.625 4979.715 ;
        RECT 441.465 4979.435 443.385 4979.715 ;
        RECT 444.225 4979.435 446.605 4979.715 ;
        RECT 447.445 4979.435 449.825 4979.715 ;
        RECT 450.665 4979.435 452.585 4979.715 ;
        RECT 453.425 4979.435 455.805 4979.715 ;
        RECT 456.645 4979.435 459.025 4979.715 ;
        RECT 459.865 4979.435 460.915 4979.715 ;
        RECT 638.210 4979.715 717.915 5188.000 ;
        RECT 638.210 4979.435 639.205 4979.715 ;
        RECT 640.045 4979.435 641.965 4979.715 ;
        RECT 642.805 4979.435 645.185 4979.715 ;
        RECT 646.025 4979.435 648.405 4979.715 ;
        RECT 649.245 4979.435 651.165 4979.715 ;
        RECT 652.005 4979.435 654.385 4979.715 ;
        RECT 655.225 4979.435 657.605 4979.715 ;
        RECT 658.445 4979.435 660.365 4979.715 ;
        RECT 661.205 4979.435 663.585 4979.715 ;
        RECT 664.425 4979.435 666.805 4979.715 ;
        RECT 667.645 4979.435 669.565 4979.715 ;
        RECT 670.405 4979.435 672.785 4979.715 ;
        RECT 673.625 4979.435 676.005 4979.715 ;
        RECT 676.845 4979.435 679.225 4979.715 ;
        RECT 680.065 4979.435 681.985 4979.715 ;
        RECT 682.825 4979.435 685.205 4979.715 ;
        RECT 686.045 4979.435 688.425 4979.715 ;
        RECT 689.265 4979.435 691.185 4979.715 ;
        RECT 692.025 4979.435 694.405 4979.715 ;
        RECT 695.245 4979.435 697.625 4979.715 ;
        RECT 698.465 4979.435 700.385 4979.715 ;
        RECT 701.225 4979.435 703.605 4979.715 ;
        RECT 704.445 4979.435 706.825 4979.715 ;
        RECT 707.665 4979.435 709.585 4979.715 ;
        RECT 710.425 4979.435 712.805 4979.715 ;
        RECT 713.645 4979.435 716.025 4979.715 ;
        RECT 716.865 4979.435 717.915 4979.715 ;
        RECT 895.210 4979.715 974.915 5188.000 ;
        RECT 895.210 4979.435 896.205 4979.715 ;
        RECT 897.045 4979.435 898.965 4979.715 ;
        RECT 899.805 4979.435 902.185 4979.715 ;
        RECT 903.025 4979.435 905.405 4979.715 ;
        RECT 906.245 4979.435 908.165 4979.715 ;
        RECT 909.005 4979.435 911.385 4979.715 ;
        RECT 912.225 4979.435 914.605 4979.715 ;
        RECT 915.445 4979.435 917.365 4979.715 ;
        RECT 918.205 4979.435 920.585 4979.715 ;
        RECT 921.425 4979.435 923.805 4979.715 ;
        RECT 924.645 4979.435 926.565 4979.715 ;
        RECT 927.405 4979.435 929.785 4979.715 ;
        RECT 930.625 4979.435 933.005 4979.715 ;
        RECT 933.845 4979.435 936.225 4979.715 ;
        RECT 937.065 4979.435 938.985 4979.715 ;
        RECT 939.825 4979.435 942.205 4979.715 ;
        RECT 943.045 4979.435 945.425 4979.715 ;
        RECT 946.265 4979.435 948.185 4979.715 ;
        RECT 949.025 4979.435 951.405 4979.715 ;
        RECT 952.245 4979.435 954.625 4979.715 ;
        RECT 955.465 4979.435 957.385 4979.715 ;
        RECT 958.225 4979.435 960.605 4979.715 ;
        RECT 961.445 4979.435 963.825 4979.715 ;
        RECT 964.665 4979.435 966.585 4979.715 ;
        RECT 967.425 4979.435 969.805 4979.715 ;
        RECT 970.645 4979.435 973.025 4979.715 ;
        RECT 973.865 4979.435 974.915 4979.715 ;
        RECT 1152.210 4979.715 1231.915 5188.000 ;
        RECT 1152.210 4979.435 1153.205 4979.715 ;
        RECT 1154.045 4979.435 1155.965 4979.715 ;
        RECT 1156.805 4979.435 1159.185 4979.715 ;
        RECT 1160.025 4979.435 1162.405 4979.715 ;
        RECT 1163.245 4979.435 1165.165 4979.715 ;
        RECT 1166.005 4979.435 1168.385 4979.715 ;
        RECT 1169.225 4979.435 1171.605 4979.715 ;
        RECT 1172.445 4979.435 1174.365 4979.715 ;
        RECT 1175.205 4979.435 1177.585 4979.715 ;
        RECT 1178.425 4979.435 1180.805 4979.715 ;
        RECT 1181.645 4979.435 1183.565 4979.715 ;
        RECT 1184.405 4979.435 1186.785 4979.715 ;
        RECT 1187.625 4979.435 1190.005 4979.715 ;
        RECT 1190.845 4979.435 1193.225 4979.715 ;
        RECT 1194.065 4979.435 1195.985 4979.715 ;
        RECT 1196.825 4979.435 1199.205 4979.715 ;
        RECT 1200.045 4979.435 1202.425 4979.715 ;
        RECT 1203.265 4979.435 1205.185 4979.715 ;
        RECT 1206.025 4979.435 1208.405 4979.715 ;
        RECT 1209.245 4979.435 1211.625 4979.715 ;
        RECT 1212.465 4979.435 1214.385 4979.715 ;
        RECT 1215.225 4979.435 1217.605 4979.715 ;
        RECT 1218.445 4979.435 1220.825 4979.715 ;
        RECT 1221.665 4979.435 1223.585 4979.715 ;
        RECT 1224.425 4979.435 1226.805 4979.715 ;
        RECT 1227.645 4979.435 1230.025 4979.715 ;
        RECT 1230.865 4979.435 1231.915 4979.715 ;
        RECT 1410.210 4979.715 1489.915 5188.000 ;
        RECT 1667.265 4990.035 1741.290 5183.075 ;
        RECT 1667.495 4988.000 1691.395 4990.035 ;
        RECT 1692.895 4988.000 1694.895 4989.920 ;
        RECT 1717.390 4988.000 1741.290 4990.035 ;
        RECT 1410.210 4979.435 1411.205 4979.715 ;
        RECT 1412.045 4979.435 1413.965 4979.715 ;
        RECT 1414.805 4979.435 1417.185 4979.715 ;
        RECT 1418.025 4979.435 1420.405 4979.715 ;
        RECT 1421.245 4979.435 1423.165 4979.715 ;
        RECT 1424.005 4979.435 1426.385 4979.715 ;
        RECT 1427.225 4979.435 1429.605 4979.715 ;
        RECT 1430.445 4979.435 1432.365 4979.715 ;
        RECT 1433.205 4979.435 1435.585 4979.715 ;
        RECT 1436.425 4979.435 1438.805 4979.715 ;
        RECT 1439.645 4979.435 1441.565 4979.715 ;
        RECT 1442.405 4979.435 1444.785 4979.715 ;
        RECT 1445.625 4979.435 1448.005 4979.715 ;
        RECT 1448.845 4979.435 1451.225 4979.715 ;
        RECT 1452.065 4979.435 1453.985 4979.715 ;
        RECT 1454.825 4979.435 1457.205 4979.715 ;
        RECT 1458.045 4979.435 1460.425 4979.715 ;
        RECT 1461.265 4979.435 1463.185 4979.715 ;
        RECT 1464.025 4979.435 1466.405 4979.715 ;
        RECT 1467.245 4979.435 1469.625 4979.715 ;
        RECT 1470.465 4979.435 1472.385 4979.715 ;
        RECT 1473.225 4979.435 1475.605 4979.715 ;
        RECT 1476.445 4979.435 1478.825 4979.715 ;
        RECT 1479.665 4979.435 1481.585 4979.715 ;
        RECT 1482.425 4979.435 1484.805 4979.715 ;
        RECT 1485.645 4979.435 1488.025 4979.715 ;
        RECT 1488.865 4979.435 1489.915 4979.715 ;
        RECT 1919.210 4979.715 1998.915 5188.000 ;
        RECT 1919.210 4979.435 1920.205 4979.715 ;
        RECT 1921.045 4979.435 1922.965 4979.715 ;
        RECT 1923.805 4979.435 1926.185 4979.715 ;
        RECT 1927.025 4979.435 1929.405 4979.715 ;
        RECT 1930.245 4979.435 1932.165 4979.715 ;
        RECT 1933.005 4979.435 1935.385 4979.715 ;
        RECT 1936.225 4979.435 1938.605 4979.715 ;
        RECT 1939.445 4979.435 1941.365 4979.715 ;
        RECT 1942.205 4979.435 1944.585 4979.715 ;
        RECT 1945.425 4979.435 1947.805 4979.715 ;
        RECT 1948.645 4979.435 1950.565 4979.715 ;
        RECT 1951.405 4979.435 1953.785 4979.715 ;
        RECT 1954.625 4979.435 1957.005 4979.715 ;
        RECT 1957.845 4979.435 1960.225 4979.715 ;
        RECT 1961.065 4979.435 1962.985 4979.715 ;
        RECT 1963.825 4979.435 1966.205 4979.715 ;
        RECT 1967.045 4979.435 1969.425 4979.715 ;
        RECT 1970.265 4979.435 1972.185 4979.715 ;
        RECT 1973.025 4979.435 1975.405 4979.715 ;
        RECT 1976.245 4979.435 1978.625 4979.715 ;
        RECT 1979.465 4979.435 1981.385 4979.715 ;
        RECT 1982.225 4979.435 1984.605 4979.715 ;
        RECT 1985.445 4979.435 1987.825 4979.715 ;
        RECT 1988.665 4979.435 1990.585 4979.715 ;
        RECT 1991.425 4979.435 1993.805 4979.715 ;
        RECT 1994.645 4979.435 1997.025 4979.715 ;
        RECT 1997.865 4979.435 1998.915 4979.715 ;
        RECT 2364.210 4979.715 2443.915 5188.000 ;
        RECT 2364.210 4979.435 2365.205 4979.715 ;
        RECT 2366.045 4979.435 2367.965 4979.715 ;
        RECT 2368.805 4979.435 2371.185 4979.715 ;
        RECT 2372.025 4979.435 2374.405 4979.715 ;
        RECT 2375.245 4979.435 2377.165 4979.715 ;
        RECT 2378.005 4979.435 2380.385 4979.715 ;
        RECT 2381.225 4979.435 2383.605 4979.715 ;
        RECT 2384.445 4979.435 2386.365 4979.715 ;
        RECT 2387.205 4979.435 2389.585 4979.715 ;
        RECT 2390.425 4979.435 2392.805 4979.715 ;
        RECT 2393.645 4979.435 2395.565 4979.715 ;
        RECT 2396.405 4979.435 2398.785 4979.715 ;
        RECT 2399.625 4979.435 2402.005 4979.715 ;
        RECT 2402.845 4979.435 2405.225 4979.715 ;
        RECT 2406.065 4979.435 2407.985 4979.715 ;
        RECT 2408.825 4979.435 2411.205 4979.715 ;
        RECT 2412.045 4979.435 2414.425 4979.715 ;
        RECT 2415.265 4979.435 2417.185 4979.715 ;
        RECT 2418.025 4979.435 2420.405 4979.715 ;
        RECT 2421.245 4979.435 2423.625 4979.715 ;
        RECT 2424.465 4979.435 2426.385 4979.715 ;
        RECT 2427.225 4979.435 2429.605 4979.715 ;
        RECT 2430.445 4979.435 2432.825 4979.715 ;
        RECT 2433.665 4979.435 2435.585 4979.715 ;
        RECT 2436.425 4979.435 2438.805 4979.715 ;
        RECT 2439.645 4979.435 2442.025 4979.715 ;
        RECT 2442.865 4979.435 2443.915 4979.715 ;
        RECT 2621.210 4979.715 2700.915 5188.000 ;
        RECT 2878.265 4990.035 2952.290 5183.075 ;
        RECT 2878.495 4988.000 2902.395 4990.035 ;
        RECT 2903.895 4988.000 2905.895 4989.920 ;
        RECT 2928.390 4988.000 2952.290 4990.035 ;
        RECT 2621.210 4979.435 2622.205 4979.715 ;
        RECT 2623.045 4979.435 2624.965 4979.715 ;
        RECT 2625.805 4979.435 2628.185 4979.715 ;
        RECT 2629.025 4979.435 2631.405 4979.715 ;
        RECT 2632.245 4979.435 2634.165 4979.715 ;
        RECT 2635.005 4979.435 2637.385 4979.715 ;
        RECT 2638.225 4979.435 2640.605 4979.715 ;
        RECT 2641.445 4979.435 2643.365 4979.715 ;
        RECT 2644.205 4979.435 2646.585 4979.715 ;
        RECT 2647.425 4979.435 2649.805 4979.715 ;
        RECT 2650.645 4979.435 2652.565 4979.715 ;
        RECT 2653.405 4979.435 2655.785 4979.715 ;
        RECT 2656.625 4979.435 2659.005 4979.715 ;
        RECT 2659.845 4979.435 2662.225 4979.715 ;
        RECT 2663.065 4979.435 2664.985 4979.715 ;
        RECT 2665.825 4979.435 2668.205 4979.715 ;
        RECT 2669.045 4979.435 2671.425 4979.715 ;
        RECT 2672.265 4979.435 2674.185 4979.715 ;
        RECT 2675.025 4979.435 2677.405 4979.715 ;
        RECT 2678.245 4979.435 2680.625 4979.715 ;
        RECT 2681.465 4979.435 2683.385 4979.715 ;
        RECT 2684.225 4979.435 2686.605 4979.715 ;
        RECT 2687.445 4979.435 2689.825 4979.715 ;
        RECT 2690.665 4979.435 2692.585 4979.715 ;
        RECT 2693.425 4979.435 2695.805 4979.715 ;
        RECT 2696.645 4979.435 2699.025 4979.715 ;
        RECT 2699.865 4979.435 2700.915 4979.715 ;
        RECT 3130.210 4979.715 3209.915 5188.000 ;
        RECT 3130.210 4979.435 3131.205 4979.715 ;
        RECT 3132.045 4979.435 3133.965 4979.715 ;
        RECT 3134.805 4979.435 3137.185 4979.715 ;
        RECT 3138.025 4979.435 3140.405 4979.715 ;
        RECT 3141.245 4979.435 3143.165 4979.715 ;
        RECT 3144.005 4979.435 3146.385 4979.715 ;
        RECT 3147.225 4979.435 3149.605 4979.715 ;
        RECT 3150.445 4979.435 3152.365 4979.715 ;
        RECT 3153.205 4979.435 3155.585 4979.715 ;
        RECT 3156.425 4979.435 3158.805 4979.715 ;
        RECT 3159.645 4979.435 3161.565 4979.715 ;
        RECT 3162.405 4979.435 3164.785 4979.715 ;
        RECT 3165.625 4979.435 3168.005 4979.715 ;
        RECT 3168.845 4979.435 3171.225 4979.715 ;
        RECT 3172.065 4979.435 3173.985 4979.715 ;
        RECT 3174.825 4979.435 3177.205 4979.715 ;
        RECT 3178.045 4979.435 3180.425 4979.715 ;
        RECT 3181.265 4979.435 3183.185 4979.715 ;
        RECT 3184.025 4979.435 3186.405 4979.715 ;
        RECT 3187.245 4979.435 3189.625 4979.715 ;
        RECT 3190.465 4979.435 3192.385 4979.715 ;
        RECT 3193.225 4979.435 3195.605 4979.715 ;
        RECT 3196.445 4979.435 3198.825 4979.715 ;
        RECT 3199.665 4979.435 3201.585 4979.715 ;
        RECT 3202.425 4979.435 3204.805 4979.715 ;
        RECT 3205.645 4979.435 3208.025 4979.715 ;
        RECT 3208.865 4979.435 3209.915 4979.715 ;
      LAYER met2 ;
        RECT 382.485 4977.035 382.765 4979.435 ;
        RECT 419.285 4977.330 419.565 4979.435 ;
        RECT 420.080 4977.950 420.340 4978.270 ;
        RECT 420.140 4977.330 420.280 4977.950 ;
        RECT 419.285 4977.190 420.280 4977.330 ;
        RECT 419.285 4977.035 419.565 4977.190 ;
        RECT 434.465 4977.035 434.745 4979.435 ;
        RECT 440.905 4977.035 441.185 4979.435 ;
        RECT 452.865 4977.035 453.145 4979.435 ;
        RECT 458.720 4977.950 458.980 4978.270 ;
        RECT 458.780 4977.330 458.920 4977.950 ;
        RECT 459.305 4977.330 459.585 4979.435 ;
        RECT 458.780 4977.190 459.585 4977.330 ;
        RECT 459.305 4977.035 459.585 4977.190 ;
        RECT 639.485 4977.035 639.765 4979.435 ;
        RECT 676.285 4977.330 676.565 4979.435 ;
        RECT 676.760 4977.330 677.020 4977.590 ;
        RECT 676.285 4977.270 677.020 4977.330 ;
        RECT 676.285 4977.190 676.960 4977.270 ;
        RECT 676.285 4977.035 676.565 4977.190 ;
        RECT 691.465 4977.035 691.745 4979.435 ;
        RECT 697.905 4977.035 698.185 4979.435 ;
        RECT 709.865 4977.035 710.145 4979.435 ;
        RECT 715.860 4977.330 716.120 4977.590 ;
        RECT 716.305 4977.330 716.585 4979.435 ;
        RECT 715.860 4977.270 716.585 4977.330 ;
        RECT 715.920 4977.190 716.585 4977.270 ;
        RECT 716.305 4977.035 716.585 4977.190 ;
        RECT 896.485 4977.035 896.765 4979.435 ;
        RECT 933.285 4977.330 933.565 4979.435 ;
        RECT 933.285 4977.035 933.640 4977.330 ;
        RECT 948.465 4977.035 948.745 4979.435 ;
        RECT 954.905 4977.035 955.185 4979.435 ;
        RECT 966.865 4977.035 967.145 4979.435 ;
        RECT 973.305 4977.330 973.585 4979.435 ;
        RECT 973.305 4977.035 973.660 4977.330 ;
        RECT 1153.485 4977.035 1153.765 4979.435 ;
        RECT 1190.285 4977.330 1190.565 4979.435 ;
        RECT 1191.040 4977.950 1191.300 4978.270 ;
        RECT 1191.100 4977.330 1191.240 4977.950 ;
        RECT 1190.285 4977.190 1191.240 4977.330 ;
        RECT 1190.285 4977.035 1190.565 4977.190 ;
        RECT 1205.465 4977.035 1205.745 4979.435 ;
        RECT 1211.905 4977.035 1212.185 4979.435 ;
        RECT 1223.865 4977.035 1224.145 4979.435 ;
        RECT 1229.680 4977.950 1229.940 4978.270 ;
        RECT 1229.740 4977.330 1229.880 4977.950 ;
        RECT 1230.305 4977.330 1230.585 4979.435 ;
        RECT 1229.740 4977.190 1230.585 4977.330 ;
        RECT 1230.305 4977.035 1230.585 4977.190 ;
        RECT 1411.485 4977.035 1411.765 4979.435 ;
        RECT 1448.285 4977.260 1448.565 4979.435 ;
        RECT 1448.240 4977.035 1448.565 4977.260 ;
        RECT 1463.465 4977.035 1463.745 4979.435 ;
        RECT 1469.905 4977.035 1470.185 4979.435 ;
        RECT 1481.865 4977.035 1482.145 4979.435 ;
        RECT 1488.305 4977.260 1488.585 4979.435 ;
        RECT 1488.260 4977.035 1488.585 4977.260 ;
        RECT 1920.485 4977.035 1920.765 4979.435 ;
        RECT 1957.285 4977.260 1957.565 4979.435 ;
        RECT 1957.285 4977.035 1957.600 4977.260 ;
        RECT 1972.465 4977.035 1972.745 4979.435 ;
        RECT 1978.905 4977.035 1979.185 4979.435 ;
        RECT 1990.865 4977.035 1991.145 4979.435 ;
        RECT 1997.305 4977.260 1997.585 4979.435 ;
        RECT 1997.305 4977.035 1997.620 4977.260 ;
        RECT 2365.485 4977.035 2365.765 4979.435 ;
        RECT 2402.285 4977.260 2402.565 4979.435 ;
        RECT 2402.280 4977.035 2402.565 4977.260 ;
        RECT 2417.465 4977.035 2417.745 4979.435 ;
        RECT 2423.905 4977.035 2424.185 4979.435 ;
        RECT 2435.865 4977.035 2436.145 4979.435 ;
        RECT 2442.305 4977.260 2442.585 4979.435 ;
        RECT 2442.300 4977.035 2442.585 4977.260 ;
        RECT 2622.485 4977.035 2622.765 4979.435 ;
        RECT 2659.285 4977.330 2659.565 4979.435 ;
        RECT 2659.820 4977.950 2660.080 4978.270 ;
        RECT 2659.880 4977.330 2660.020 4977.950 ;
        RECT 2659.285 4977.190 2660.020 4977.330 ;
        RECT 2659.285 4977.035 2659.565 4977.190 ;
        RECT 2674.465 4977.035 2674.745 4979.435 ;
        RECT 2680.905 4977.035 2681.185 4979.435 ;
        RECT 2692.865 4977.035 2693.145 4979.435 ;
        RECT 2698.460 4977.950 2698.720 4978.270 ;
        RECT 2698.520 4977.330 2698.660 4977.950 ;
        RECT 2699.305 4977.330 2699.585 4979.435 ;
        RECT 2698.520 4977.190 2699.585 4977.330 ;
        RECT 2699.305 4977.035 2699.585 4977.190 ;
        RECT 3131.485 4977.035 3131.765 4979.435 ;
        RECT 3168.285 4977.330 3168.565 4979.435 ;
        RECT 3169.040 4977.330 3169.300 4977.590 ;
        RECT 3168.285 4977.270 3169.300 4977.330 ;
        RECT 3168.285 4977.190 3169.240 4977.270 ;
        RECT 3168.285 4977.035 3168.565 4977.190 ;
        RECT 3183.465 4977.035 3183.745 4979.435 ;
        RECT 3189.905 4977.035 3190.185 4979.435 ;
        RECT 3201.865 4977.035 3202.145 4979.435 ;
        RECT 3207.680 4977.330 3207.940 4977.590 ;
        RECT 3208.305 4977.330 3208.585 4979.435 ;
        RECT 3207.680 4977.270 3208.585 4977.330 ;
        RECT 3207.740 4977.190 3208.585 4977.270 ;
        RECT 3208.305 4977.035 3208.585 4977.190 ;
        RECT 933.500 4953.110 933.640 4977.035 ;
        RECT 973.520 4953.110 973.660 4977.035 ;
        RECT 1448.240 4976.570 1448.380 4977.035 ;
        RECT 1488.260 4976.570 1488.400 4977.035 ;
        RECT 1957.460 4976.570 1957.600 4977.035 ;
        RECT 1997.480 4976.570 1997.620 4977.035 ;
        RECT 2402.280 4976.570 2402.420 4977.035 ;
        RECT 2442.300 4976.570 2442.440 4977.035 ;
        RECT 1448.180 4976.250 1448.440 4976.570 ;
        RECT 1488.200 4976.250 1488.460 4976.570 ;
        RECT 1957.400 4976.250 1957.660 4976.570 ;
        RECT 1997.420 4976.250 1997.680 4976.570 ;
        RECT 2402.220 4976.250 2402.480 4976.570 ;
        RECT 2442.240 4976.250 2442.500 4976.570 ;
        RECT 933.440 4952.790 933.700 4953.110 ;
        RECT 973.460 4952.790 973.720 4953.110 ;
      LAYER met2 ;
        RECT 0.000 4849.865 208.565 4850.915 ;
        RECT 0.000 4849.025 208.285 4849.865 ;
      LAYER met2 ;
        RECT 208.565 4849.305 210.965 4849.585 ;
      LAYER met2 ;
        RECT 0.000 4846.645 208.565 4849.025 ;
      LAYER met2 ;
        RECT 209.000 4847.030 209.140 4849.305 ;
        RECT 208.940 4846.710 209.200 4847.030 ;
        RECT 212.160 4846.710 212.420 4847.030 ;
      LAYER met2 ;
        RECT 0.000 4845.805 208.285 4846.645 ;
        RECT 0.000 4843.425 208.565 4845.805 ;
        RECT 0.000 4842.585 208.285 4843.425 ;
      LAYER met2 ;
        RECT 208.565 4842.865 210.965 4843.145 ;
      LAYER met2 ;
        RECT 0.000 4840.665 208.565 4842.585 ;
        RECT 0.000 4839.825 208.285 4840.665 ;
        RECT 0.000 4837.445 208.565 4839.825 ;
        RECT 0.000 4836.605 208.285 4837.445 ;
        RECT 0.000 4834.225 208.565 4836.605 ;
        RECT 0.000 4833.385 208.285 4834.225 ;
        RECT 0.000 4831.465 208.565 4833.385 ;
        RECT 0.000 4830.625 208.285 4831.465 ;
      LAYER met2 ;
        RECT 208.565 4830.905 210.965 4831.185 ;
      LAYER met2 ;
        RECT 0.000 4828.245 208.565 4830.625 ;
        RECT 0.000 4827.405 208.285 4828.245 ;
        RECT 0.000 4825.025 208.565 4827.405 ;
        RECT 0.000 4824.185 208.285 4825.025 ;
      LAYER met2 ;
        RECT 208.565 4824.465 210.965 4824.745 ;
      LAYER met2 ;
        RECT 0.000 4822.265 208.565 4824.185 ;
        RECT 0.000 4821.425 208.285 4822.265 ;
        RECT 0.000 4819.045 208.565 4821.425 ;
        RECT 0.000 4818.205 208.285 4819.045 ;
        RECT 0.000 4815.825 208.565 4818.205 ;
        RECT 0.000 4814.985 208.285 4815.825 ;
        RECT 0.000 4813.065 208.565 4814.985 ;
        RECT 0.000 4812.225 208.285 4813.065 ;
      LAYER met2 ;
        RECT 212.220 4812.350 212.360 4846.710 ;
      LAYER met2 ;
        RECT 3379.435 4836.795 3588.000 4837.790 ;
      LAYER met2 ;
        RECT 3377.035 4836.235 3379.435 4836.515 ;
      LAYER met2 ;
        RECT 3379.715 4835.955 3588.000 4836.795 ;
        RECT 3379.435 4834.035 3588.000 4835.955 ;
        RECT 3379.715 4833.195 3588.000 4834.035 ;
        RECT 3379.435 4830.815 3588.000 4833.195 ;
        RECT 3379.715 4829.975 3588.000 4830.815 ;
        RECT 3379.435 4827.595 3588.000 4829.975 ;
        RECT 3379.715 4826.755 3588.000 4827.595 ;
        RECT 3379.435 4824.835 3588.000 4826.755 ;
        RECT 3379.715 4823.995 3588.000 4824.835 ;
        RECT 3379.435 4821.615 3588.000 4823.995 ;
        RECT 3379.715 4820.775 3588.000 4821.615 ;
        RECT 3379.435 4818.395 3588.000 4820.775 ;
        RECT 3379.715 4817.555 3588.000 4818.395 ;
        RECT 3379.435 4815.635 3588.000 4817.555 ;
        RECT 3379.715 4814.795 3588.000 4815.635 ;
        RECT 3379.435 4812.415 3588.000 4814.795 ;
        RECT 0.000 4809.845 208.565 4812.225 ;
      LAYER met2 ;
        RECT 208.940 4812.030 209.200 4812.350 ;
        RECT 212.160 4812.030 212.420 4812.350 ;
      LAYER met2 ;
        RECT 0.000 4809.005 208.285 4809.845 ;
      LAYER met2 ;
        RECT 209.000 4809.565 209.140 4812.030 ;
      LAYER met2 ;
        RECT 3379.715 4811.575 3588.000 4812.415 ;
      LAYER met2 ;
        RECT 208.565 4809.285 210.965 4809.565 ;
      LAYER met2 ;
        RECT 3379.435 4809.195 3588.000 4811.575 ;
        RECT 0.000 4806.625 208.565 4809.005 ;
        RECT 3379.715 4808.355 3588.000 4809.195 ;
        RECT 0.000 4805.785 208.285 4806.625 ;
        RECT 3379.435 4806.435 3588.000 4808.355 ;
        RECT 0.000 4803.405 208.565 4805.785 ;
        RECT 3379.715 4805.595 3588.000 4806.435 ;
        RECT 0.000 4802.565 208.285 4803.405 ;
        RECT 3379.435 4803.215 3588.000 4805.595 ;
        RECT 0.000 4800.645 208.565 4802.565 ;
        RECT 3379.715 4802.375 3588.000 4803.215 ;
        RECT 0.000 4799.805 208.285 4800.645 ;
        RECT 3379.435 4799.995 3588.000 4802.375 ;
        RECT 0.000 4797.425 208.565 4799.805 ;
      LAYER met2 ;
        RECT 3377.035 4799.645 3379.435 4799.715 ;
        RECT 3376.560 4799.505 3379.435 4799.645 ;
      LAYER met2 ;
        RECT 0.000 4796.585 208.285 4797.425 ;
        RECT 0.000 4794.205 208.565 4796.585 ;
        RECT 0.000 4793.365 208.285 4794.205 ;
        RECT 0.000 4791.445 208.565 4793.365 ;
        RECT 0.000 4790.605 208.285 4791.445 ;
        RECT 0.000 4788.225 208.565 4790.605 ;
        RECT 0.000 4787.385 208.285 4788.225 ;
        RECT 0.000 4785.005 208.565 4787.385 ;
        RECT 0.000 4784.165 208.285 4785.005 ;
        RECT 0.000 4782.245 208.565 4784.165 ;
        RECT 0.000 4781.405 208.285 4782.245 ;
        RECT 0.000 4779.025 208.565 4781.405 ;
        RECT 0.000 4778.185 208.285 4779.025 ;
        RECT 0.000 4775.805 208.565 4778.185 ;
        RECT 0.000 4774.965 208.285 4775.805 ;
        RECT 0.000 4773.045 208.565 4774.965 ;
        RECT 0.000 4772.205 208.285 4773.045 ;
      LAYER met2 ;
        RECT 208.565 4772.485 210.965 4772.765 ;
      LAYER met2 ;
        RECT 0.000 4771.210 208.565 4772.205 ;
      LAYER met2 ;
        RECT 3376.560 4759.050 3376.700 4799.505 ;
        RECT 3377.035 4799.435 3379.435 4799.505 ;
      LAYER met2 ;
        RECT 3379.715 4799.155 3588.000 4799.995 ;
        RECT 3379.435 4796.775 3588.000 4799.155 ;
        RECT 3379.715 4795.935 3588.000 4796.775 ;
        RECT 3379.435 4794.015 3588.000 4795.935 ;
        RECT 3379.715 4793.175 3588.000 4794.015 ;
        RECT 3379.435 4790.795 3588.000 4793.175 ;
        RECT 3379.715 4789.955 3588.000 4790.795 ;
        RECT 3379.435 4787.575 3588.000 4789.955 ;
        RECT 3379.715 4786.735 3588.000 4787.575 ;
        RECT 3379.435 4784.815 3588.000 4786.735 ;
      LAYER met2 ;
        RECT 3377.035 4784.255 3379.435 4784.535 ;
      LAYER met2 ;
        RECT 3379.715 4783.975 3588.000 4784.815 ;
        RECT 3379.435 4781.595 3588.000 4783.975 ;
        RECT 3379.715 4780.755 3588.000 4781.595 ;
        RECT 3379.435 4778.375 3588.000 4780.755 ;
      LAYER met2 ;
        RECT 3377.035 4777.815 3379.435 4778.095 ;
      LAYER met2 ;
        RECT 3379.715 4777.535 3588.000 4778.375 ;
        RECT 3379.435 4775.615 3588.000 4777.535 ;
        RECT 3379.715 4774.775 3588.000 4775.615 ;
        RECT 3379.435 4772.395 3588.000 4774.775 ;
        RECT 3379.715 4771.555 3588.000 4772.395 ;
        RECT 3379.435 4769.175 3588.000 4771.555 ;
        RECT 3379.715 4768.335 3588.000 4769.175 ;
        RECT 3379.435 4766.415 3588.000 4768.335 ;
      LAYER met2 ;
        RECT 3377.035 4765.855 3379.435 4766.135 ;
      LAYER met2 ;
        RECT 3379.715 4765.575 3588.000 4766.415 ;
        RECT 3379.435 4763.195 3588.000 4765.575 ;
        RECT 3379.715 4762.355 3588.000 4763.195 ;
        RECT 3379.435 4759.975 3588.000 4762.355 ;
      LAYER met2 ;
        RECT 3377.035 4759.660 3379.435 4759.695 ;
        RECT 3377.020 4759.415 3379.435 4759.660 ;
        RECT 3377.020 4759.050 3377.160 4759.415 ;
      LAYER met2 ;
        RECT 3379.715 4759.135 3588.000 4759.975 ;
      LAYER met2 ;
        RECT 3376.560 4758.910 3377.160 4759.050 ;
      LAYER met2 ;
        RECT 3379.435 4758.085 3588.000 4759.135 ;
        RECT 153.765 4635.000 158.415 4646.140 ;
        RECT 159.640 4635.245 163.510 4646.195 ;
        RECT 3.570 4634.700 197.965 4635.000 ;
        RECT 3.570 4614.095 198.000 4634.700 ;
        RECT 3.570 4613.535 197.965 4614.095 ;
        RECT 3.570 4580.925 198.000 4613.535 ;
        RECT 3390.035 4612.500 3584.430 4612.510 ;
        RECT 3390.000 4592.505 3584.430 4612.500 ;
        RECT 3390.035 4592.075 3584.430 4592.505 ;
        RECT 3.570 4580.495 197.965 4580.925 ;
        RECT 3.570 4560.500 198.000 4580.495 ;
        RECT 3.570 4560.490 197.965 4560.500 ;
        RECT 3390.000 4559.465 3584.430 4592.075 ;
        RECT 3390.035 4558.905 3584.430 4559.465 ;
        RECT 3390.000 4538.300 3584.430 4558.905 ;
        RECT 3390.035 4538.000 3584.430 4538.300 ;
        RECT 3424.490 4526.805 3428.360 4537.755 ;
        RECT 3429.585 4526.860 3434.235 4538.000 ;
        RECT 4.925 4399.390 200.000 4423.290 ;
        RECT 4.925 4373.395 197.965 4399.390 ;
        RECT 3379.435 4390.795 3588.000 4391.790 ;
      LAYER met2 ;
        RECT 3377.035 4390.235 3379.435 4390.515 ;
      LAYER met2 ;
        RECT 3379.715 4389.955 3588.000 4390.795 ;
        RECT 3379.435 4388.035 3588.000 4389.955 ;
        RECT 3379.715 4387.195 3588.000 4388.035 ;
        RECT 3379.435 4384.815 3588.000 4387.195 ;
        RECT 3379.715 4383.975 3588.000 4384.815 ;
        RECT 3379.435 4381.595 3588.000 4383.975 ;
        RECT 3379.715 4380.755 3588.000 4381.595 ;
        RECT 3379.435 4378.835 3588.000 4380.755 ;
        RECT 3379.715 4377.995 3588.000 4378.835 ;
        RECT 198.080 4374.895 200.000 4376.895 ;
        RECT 3379.435 4375.615 3588.000 4377.995 ;
        RECT 3379.715 4374.775 3588.000 4375.615 ;
        RECT 4.925 4349.495 200.000 4373.395 ;
        RECT 3379.435 4372.395 3588.000 4374.775 ;
        RECT 3379.715 4371.555 3588.000 4372.395 ;
        RECT 3379.435 4369.635 3588.000 4371.555 ;
        RECT 3379.715 4368.795 3588.000 4369.635 ;
        RECT 3379.435 4366.415 3588.000 4368.795 ;
        RECT 3379.715 4365.575 3588.000 4366.415 ;
        RECT 3379.435 4363.195 3588.000 4365.575 ;
        RECT 3379.715 4362.355 3588.000 4363.195 ;
        RECT 3379.435 4360.435 3588.000 4362.355 ;
        RECT 3379.715 4359.595 3588.000 4360.435 ;
        RECT 3379.435 4357.215 3588.000 4359.595 ;
        RECT 3379.715 4356.375 3588.000 4357.215 ;
        RECT 3379.435 4353.995 3588.000 4356.375 ;
      LAYER met2 ;
        RECT 3377.035 4353.700 3379.435 4353.715 ;
        RECT 3377.020 4353.435 3379.435 4353.700 ;
        RECT 3377.020 4350.970 3377.160 4353.435 ;
      LAYER met2 ;
        RECT 3379.715 4353.155 3588.000 4353.995 ;
      LAYER met2 ;
        RECT 3368.680 4350.650 3368.940 4350.970 ;
        RECT 3376.960 4350.650 3377.220 4350.970 ;
      LAYER met2 ;
        RECT 3379.435 4350.775 3588.000 4353.155 ;
        RECT 4.925 4349.265 197.965 4349.495 ;
      LAYER met2 ;
        RECT 3368.740 4316.290 3368.880 4350.650 ;
      LAYER met2 ;
        RECT 3379.715 4349.935 3588.000 4350.775 ;
        RECT 3379.435 4348.015 3588.000 4349.935 ;
        RECT 3379.715 4347.175 3588.000 4348.015 ;
        RECT 3379.435 4344.795 3588.000 4347.175 ;
        RECT 3379.715 4343.955 3588.000 4344.795 ;
        RECT 3379.435 4341.575 3588.000 4343.955 ;
        RECT 3379.715 4340.735 3588.000 4341.575 ;
        RECT 3379.435 4338.815 3588.000 4340.735 ;
      LAYER met2 ;
        RECT 3377.035 4338.255 3379.435 4338.535 ;
      LAYER met2 ;
        RECT 3379.715 4337.975 3588.000 4338.815 ;
        RECT 3379.435 4335.595 3588.000 4337.975 ;
        RECT 3379.715 4334.755 3588.000 4335.595 ;
        RECT 3379.435 4332.375 3588.000 4334.755 ;
      LAYER met2 ;
        RECT 3377.035 4331.815 3379.435 4332.095 ;
      LAYER met2 ;
        RECT 3379.715 4331.535 3588.000 4332.375 ;
        RECT 3379.435 4329.615 3588.000 4331.535 ;
        RECT 3379.715 4328.775 3588.000 4329.615 ;
        RECT 3379.435 4326.395 3588.000 4328.775 ;
        RECT 3379.715 4325.555 3588.000 4326.395 ;
        RECT 3379.435 4323.175 3588.000 4325.555 ;
        RECT 3379.715 4322.335 3588.000 4323.175 ;
        RECT 3379.435 4320.415 3588.000 4322.335 ;
      LAYER met2 ;
        RECT 3377.035 4319.855 3379.435 4320.135 ;
      LAYER met2 ;
        RECT 3379.715 4319.575 3588.000 4320.415 ;
        RECT 3379.435 4317.195 3588.000 4319.575 ;
        RECT 3379.715 4316.355 3588.000 4317.195 ;
      LAYER met2 ;
        RECT 3368.680 4315.970 3368.940 4316.290 ;
        RECT 3376.960 4315.970 3377.220 4316.290 ;
        RECT 3377.020 4313.695 3377.160 4315.970 ;
      LAYER met2 ;
        RECT 3379.435 4313.975 3588.000 4316.355 ;
      LAYER met2 ;
        RECT 3377.020 4313.580 3379.435 4313.695 ;
        RECT 3377.035 4313.415 3379.435 4313.580 ;
      LAYER met2 ;
        RECT 3379.715 4313.135 3588.000 4313.975 ;
        RECT 3379.435 4312.085 3588.000 4313.135 ;
        RECT 4.925 4188.390 200.000 4212.290 ;
        RECT 4.925 4162.395 197.965 4188.390 ;
        RECT 3390.035 4166.505 3583.075 4166.735 ;
        RECT 198.080 4163.895 200.000 4165.895 ;
        RECT 4.925 4138.495 200.000 4162.395 ;
        RECT 3388.000 4142.605 3583.075 4166.505 ;
        RECT 3388.000 4139.105 3389.920 4141.105 ;
        RECT 4.925 4138.265 197.965 4138.495 ;
        RECT 3390.035 4116.610 3583.075 4142.605 ;
        RECT 3388.000 4092.710 3583.075 4116.610 ;
        RECT 0.000 4000.865 208.565 4001.915 ;
        RECT 0.000 4000.025 208.285 4000.865 ;
      LAYER met2 ;
        RECT 208.565 4000.305 210.965 4000.585 ;
      LAYER met2 ;
        RECT 0.000 3997.645 208.565 4000.025 ;
      LAYER met2 ;
        RECT 209.000 3998.050 209.140 4000.305 ;
        RECT 208.940 3997.730 209.200 3998.050 ;
        RECT 211.700 3997.730 211.960 3998.050 ;
      LAYER met2 ;
        RECT 0.000 3996.805 208.285 3997.645 ;
        RECT 0.000 3994.425 208.565 3996.805 ;
        RECT 0.000 3993.585 208.285 3994.425 ;
      LAYER met2 ;
        RECT 208.565 3993.865 210.965 3994.145 ;
      LAYER met2 ;
        RECT 0.000 3991.665 208.565 3993.585 ;
        RECT 0.000 3990.825 208.285 3991.665 ;
        RECT 0.000 3988.445 208.565 3990.825 ;
        RECT 0.000 3987.605 208.285 3988.445 ;
        RECT 0.000 3985.225 208.565 3987.605 ;
        RECT 0.000 3984.385 208.285 3985.225 ;
        RECT 0.000 3982.465 208.565 3984.385 ;
        RECT 0.000 3981.625 208.285 3982.465 ;
      LAYER met2 ;
        RECT 208.565 3981.905 210.965 3982.185 ;
      LAYER met2 ;
        RECT 0.000 3979.245 208.565 3981.625 ;
        RECT 0.000 3978.405 208.285 3979.245 ;
        RECT 0.000 3976.025 208.565 3978.405 ;
        RECT 0.000 3975.185 208.285 3976.025 ;
      LAYER met2 ;
        RECT 208.565 3975.465 210.965 3975.745 ;
      LAYER met2 ;
        RECT 0.000 3973.265 208.565 3975.185 ;
        RECT 0.000 3972.425 208.285 3973.265 ;
        RECT 0.000 3970.045 208.565 3972.425 ;
        RECT 0.000 3969.205 208.285 3970.045 ;
        RECT 0.000 3966.825 208.565 3969.205 ;
        RECT 0.000 3965.985 208.285 3966.825 ;
        RECT 0.000 3964.065 208.565 3965.985 ;
        RECT 0.000 3963.225 208.285 3964.065 ;
        RECT 0.000 3960.845 208.565 3963.225 ;
      LAYER met2 ;
        RECT 211.760 3963.030 211.900 3997.730 ;
        RECT 208.940 3962.710 209.200 3963.030 ;
        RECT 211.700 3962.710 211.960 3963.030 ;
      LAYER met2 ;
        RECT 0.000 3960.005 208.285 3960.845 ;
      LAYER met2 ;
        RECT 209.000 3960.565 209.140 3962.710 ;
        RECT 208.565 3960.285 210.965 3960.565 ;
      LAYER met2 ;
        RECT 0.000 3957.625 208.565 3960.005 ;
        RECT 0.000 3956.785 208.285 3957.625 ;
        RECT 0.000 3954.405 208.565 3956.785 ;
        RECT 0.000 3953.565 208.285 3954.405 ;
        RECT 0.000 3951.645 208.565 3953.565 ;
        RECT 0.000 3950.805 208.285 3951.645 ;
        RECT 0.000 3948.425 208.565 3950.805 ;
        RECT 0.000 3947.585 208.285 3948.425 ;
        RECT 0.000 3945.205 208.565 3947.585 ;
        RECT 0.000 3944.365 208.285 3945.205 ;
        RECT 3379.435 3944.795 3588.000 3945.790 ;
        RECT 0.000 3942.445 208.565 3944.365 ;
      LAYER met2 ;
        RECT 3377.035 3944.235 3379.435 3944.515 ;
      LAYER met2 ;
        RECT 3379.715 3943.955 3588.000 3944.795 ;
        RECT 0.000 3941.605 208.285 3942.445 ;
        RECT 3379.435 3942.035 3588.000 3943.955 ;
        RECT 0.000 3939.225 208.565 3941.605 ;
        RECT 3379.715 3941.195 3588.000 3942.035 ;
        RECT 0.000 3938.385 208.285 3939.225 ;
        RECT 3379.435 3938.815 3588.000 3941.195 ;
        RECT 0.000 3936.005 208.565 3938.385 ;
        RECT 3379.715 3937.975 3588.000 3938.815 ;
        RECT 0.000 3935.165 208.285 3936.005 ;
        RECT 3379.435 3935.595 3588.000 3937.975 ;
        RECT 0.000 3933.245 208.565 3935.165 ;
        RECT 3379.715 3934.755 3588.000 3935.595 ;
        RECT 0.000 3932.405 208.285 3933.245 ;
        RECT 3379.435 3932.835 3588.000 3934.755 ;
        RECT 0.000 3930.025 208.565 3932.405 ;
        RECT 3379.715 3931.995 3588.000 3932.835 ;
        RECT 0.000 3929.185 208.285 3930.025 ;
        RECT 3379.435 3929.615 3588.000 3931.995 ;
        RECT 0.000 3926.805 208.565 3929.185 ;
        RECT 3379.715 3928.775 3588.000 3929.615 ;
        RECT 0.000 3925.965 208.285 3926.805 ;
        RECT 3379.435 3926.395 3588.000 3928.775 ;
        RECT 0.000 3924.045 208.565 3925.965 ;
        RECT 3379.715 3925.555 3588.000 3926.395 ;
        RECT 0.000 3923.205 208.285 3924.045 ;
      LAYER met2 ;
        RECT 208.565 3923.485 210.965 3923.765 ;
      LAYER met2 ;
        RECT 3379.435 3923.635 3588.000 3925.555 ;
        RECT 0.000 3922.210 208.565 3923.205 ;
        RECT 3379.715 3922.795 3588.000 3923.635 ;
        RECT 3379.435 3920.415 3588.000 3922.795 ;
        RECT 3379.715 3919.575 3588.000 3920.415 ;
        RECT 3379.435 3917.195 3588.000 3919.575 ;
        RECT 3379.715 3916.355 3588.000 3917.195 ;
        RECT 3379.435 3914.435 3588.000 3916.355 ;
        RECT 3379.715 3913.595 3588.000 3914.435 ;
        RECT 3379.435 3911.215 3588.000 3913.595 ;
        RECT 3379.715 3910.375 3588.000 3911.215 ;
        RECT 3379.435 3907.995 3588.000 3910.375 ;
      LAYER met2 ;
        RECT 3377.035 3907.690 3379.435 3907.715 ;
        RECT 3376.100 3907.550 3379.435 3907.690 ;
        RECT 3376.100 3870.210 3376.240 3907.550 ;
        RECT 3377.035 3907.435 3379.435 3907.550 ;
      LAYER met2 ;
        RECT 3379.715 3907.155 3588.000 3907.995 ;
        RECT 3379.435 3904.775 3588.000 3907.155 ;
        RECT 3379.715 3903.935 3588.000 3904.775 ;
        RECT 3379.435 3902.015 3588.000 3903.935 ;
        RECT 3379.715 3901.175 3588.000 3902.015 ;
        RECT 3379.435 3898.795 3588.000 3901.175 ;
        RECT 3379.715 3897.955 3588.000 3898.795 ;
        RECT 3379.435 3895.575 3588.000 3897.955 ;
        RECT 3379.715 3894.735 3588.000 3895.575 ;
        RECT 3379.435 3892.815 3588.000 3894.735 ;
      LAYER met2 ;
        RECT 3377.035 3892.255 3379.435 3892.535 ;
      LAYER met2 ;
        RECT 3379.715 3891.975 3588.000 3892.815 ;
        RECT 3379.435 3889.595 3588.000 3891.975 ;
        RECT 3379.715 3888.755 3588.000 3889.595 ;
        RECT 3379.435 3886.375 3588.000 3888.755 ;
      LAYER met2 ;
        RECT 3377.035 3885.815 3379.435 3886.095 ;
      LAYER met2 ;
        RECT 3379.715 3885.535 3588.000 3886.375 ;
        RECT 3379.435 3883.615 3588.000 3885.535 ;
        RECT 3379.715 3882.775 3588.000 3883.615 ;
        RECT 3379.435 3880.395 3588.000 3882.775 ;
        RECT 3379.715 3879.555 3588.000 3880.395 ;
        RECT 3379.435 3877.175 3588.000 3879.555 ;
        RECT 3379.715 3876.335 3588.000 3877.175 ;
        RECT 3379.435 3874.415 3588.000 3876.335 ;
      LAYER met2 ;
        RECT 3377.035 3873.855 3379.435 3874.135 ;
      LAYER met2 ;
        RECT 3379.715 3873.575 3588.000 3874.415 ;
        RECT 3379.435 3871.195 3588.000 3873.575 ;
        RECT 3379.715 3870.355 3588.000 3871.195 ;
      LAYER met2 ;
        RECT 3376.040 3869.890 3376.300 3870.210 ;
        RECT 3376.960 3869.890 3377.220 3870.210 ;
        RECT 3377.020 3867.695 3377.160 3869.890 ;
      LAYER met2 ;
        RECT 3379.435 3867.975 3588.000 3870.355 ;
      LAYER met2 ;
        RECT 3377.020 3867.500 3379.435 3867.695 ;
        RECT 3377.035 3867.415 3379.435 3867.500 ;
      LAYER met2 ;
        RECT 3379.715 3867.135 3588.000 3867.975 ;
        RECT 3379.435 3866.085 3588.000 3867.135 ;
        RECT 0.000 3784.865 208.565 3785.915 ;
        RECT 0.000 3784.025 208.285 3784.865 ;
      LAYER met2 ;
        RECT 208.610 3784.585 209.140 3784.610 ;
        RECT 208.565 3784.305 210.965 3784.585 ;
      LAYER met2 ;
        RECT 0.000 3781.645 208.565 3784.025 ;
      LAYER met2 ;
        RECT 209.000 3782.150 209.140 3784.305 ;
        RECT 208.940 3781.830 209.200 3782.150 ;
        RECT 211.700 3781.830 211.960 3782.150 ;
      LAYER met2 ;
        RECT 0.000 3780.805 208.285 3781.645 ;
        RECT 0.000 3778.425 208.565 3780.805 ;
        RECT 0.000 3777.585 208.285 3778.425 ;
      LAYER met2 ;
        RECT 208.565 3777.865 210.965 3778.145 ;
      LAYER met2 ;
        RECT 0.000 3775.665 208.565 3777.585 ;
        RECT 0.000 3774.825 208.285 3775.665 ;
        RECT 0.000 3772.445 208.565 3774.825 ;
        RECT 0.000 3771.605 208.285 3772.445 ;
        RECT 0.000 3769.225 208.565 3771.605 ;
        RECT 0.000 3768.385 208.285 3769.225 ;
        RECT 0.000 3766.465 208.565 3768.385 ;
        RECT 0.000 3765.625 208.285 3766.465 ;
      LAYER met2 ;
        RECT 208.565 3765.905 210.965 3766.185 ;
      LAYER met2 ;
        RECT 0.000 3763.245 208.565 3765.625 ;
        RECT 0.000 3762.405 208.285 3763.245 ;
        RECT 0.000 3760.025 208.565 3762.405 ;
        RECT 0.000 3759.185 208.285 3760.025 ;
      LAYER met2 ;
        RECT 208.565 3759.465 210.965 3759.745 ;
      LAYER met2 ;
        RECT 0.000 3757.265 208.565 3759.185 ;
        RECT 0.000 3756.425 208.285 3757.265 ;
        RECT 0.000 3754.045 208.565 3756.425 ;
        RECT 0.000 3753.205 208.285 3754.045 ;
        RECT 0.000 3750.825 208.565 3753.205 ;
        RECT 0.000 3749.985 208.285 3750.825 ;
        RECT 0.000 3748.065 208.565 3749.985 ;
        RECT 0.000 3747.225 208.285 3748.065 ;
        RECT 0.000 3744.845 208.565 3747.225 ;
      LAYER met2 ;
        RECT 211.760 3747.130 211.900 3781.830 ;
        RECT 208.940 3746.810 209.200 3747.130 ;
        RECT 211.700 3746.810 211.960 3747.130 ;
      LAYER met2 ;
        RECT 0.000 3744.005 208.285 3744.845 ;
      LAYER met2 ;
        RECT 209.000 3744.565 209.140 3746.810 ;
        RECT 208.565 3744.285 210.965 3744.565 ;
      LAYER met2 ;
        RECT 0.000 3741.625 208.565 3744.005 ;
        RECT 0.000 3740.785 208.285 3741.625 ;
        RECT 0.000 3738.405 208.565 3740.785 ;
        RECT 0.000 3737.565 208.285 3738.405 ;
        RECT 0.000 3735.645 208.565 3737.565 ;
        RECT 0.000 3734.805 208.285 3735.645 ;
        RECT 0.000 3732.425 208.565 3734.805 ;
        RECT 0.000 3731.585 208.285 3732.425 ;
        RECT 0.000 3729.205 208.565 3731.585 ;
        RECT 0.000 3728.365 208.285 3729.205 ;
        RECT 0.000 3726.445 208.565 3728.365 ;
        RECT 0.000 3725.605 208.285 3726.445 ;
        RECT 0.000 3723.225 208.565 3725.605 ;
        RECT 0.000 3722.385 208.285 3723.225 ;
        RECT 0.000 3720.005 208.565 3722.385 ;
        RECT 0.000 3719.165 208.285 3720.005 ;
        RECT 3379.435 3719.795 3588.000 3720.790 ;
      LAYER met2 ;
        RECT 3377.035 3719.235 3379.435 3719.515 ;
      LAYER met2 ;
        RECT 0.000 3717.245 208.565 3719.165 ;
        RECT 3379.715 3718.955 3588.000 3719.795 ;
        RECT 0.000 3716.405 208.285 3717.245 ;
        RECT 3379.435 3717.035 3588.000 3718.955 ;
        RECT 0.000 3714.025 208.565 3716.405 ;
        RECT 3379.715 3716.195 3588.000 3717.035 ;
        RECT 0.000 3713.185 208.285 3714.025 ;
        RECT 3379.435 3713.815 3588.000 3716.195 ;
        RECT 0.000 3710.805 208.565 3713.185 ;
        RECT 3379.715 3712.975 3588.000 3713.815 ;
        RECT 0.000 3709.965 208.285 3710.805 ;
        RECT 3379.435 3710.595 3588.000 3712.975 ;
        RECT 0.000 3708.045 208.565 3709.965 ;
        RECT 3379.715 3709.755 3588.000 3710.595 ;
        RECT 0.000 3707.205 208.285 3708.045 ;
        RECT 3379.435 3707.835 3588.000 3709.755 ;
      LAYER met2 ;
        RECT 208.565 3707.485 210.965 3707.765 ;
      LAYER met2 ;
        RECT 0.000 3706.210 208.565 3707.205 ;
        RECT 3379.715 3706.995 3588.000 3707.835 ;
        RECT 3379.435 3704.615 3588.000 3706.995 ;
        RECT 3379.715 3703.775 3588.000 3704.615 ;
        RECT 3379.435 3701.395 3588.000 3703.775 ;
        RECT 3379.715 3700.555 3588.000 3701.395 ;
        RECT 3379.435 3698.635 3588.000 3700.555 ;
        RECT 3379.715 3697.795 3588.000 3698.635 ;
        RECT 3379.435 3695.415 3588.000 3697.795 ;
        RECT 3379.715 3694.575 3588.000 3695.415 ;
        RECT 3379.435 3692.195 3588.000 3694.575 ;
        RECT 3379.715 3691.355 3588.000 3692.195 ;
        RECT 3379.435 3689.435 3588.000 3691.355 ;
        RECT 3379.715 3688.595 3588.000 3689.435 ;
        RECT 3379.435 3686.215 3588.000 3688.595 ;
        RECT 3379.715 3685.375 3588.000 3686.215 ;
        RECT 3379.435 3682.995 3588.000 3685.375 ;
      LAYER met2 ;
        RECT 3377.035 3682.610 3379.435 3682.715 ;
        RECT 3376.560 3682.470 3379.435 3682.610 ;
        RECT 3376.560 3645.210 3376.700 3682.470 ;
        RECT 3377.035 3682.435 3379.435 3682.470 ;
      LAYER met2 ;
        RECT 3379.715 3682.155 3588.000 3682.995 ;
        RECT 3379.435 3679.775 3588.000 3682.155 ;
        RECT 3379.715 3678.935 3588.000 3679.775 ;
        RECT 3379.435 3677.015 3588.000 3678.935 ;
        RECT 3379.715 3676.175 3588.000 3677.015 ;
        RECT 3379.435 3673.795 3588.000 3676.175 ;
        RECT 3379.715 3672.955 3588.000 3673.795 ;
        RECT 3379.435 3670.575 3588.000 3672.955 ;
        RECT 3379.715 3669.735 3588.000 3670.575 ;
        RECT 3379.435 3667.815 3588.000 3669.735 ;
      LAYER met2 ;
        RECT 3377.035 3667.255 3379.435 3667.535 ;
      LAYER met2 ;
        RECT 3379.715 3666.975 3588.000 3667.815 ;
        RECT 3379.435 3664.595 3588.000 3666.975 ;
        RECT 3379.715 3663.755 3588.000 3664.595 ;
        RECT 3379.435 3661.375 3588.000 3663.755 ;
      LAYER met2 ;
        RECT 3377.035 3660.815 3379.435 3661.095 ;
      LAYER met2 ;
        RECT 3379.715 3660.535 3588.000 3661.375 ;
        RECT 3379.435 3658.615 3588.000 3660.535 ;
        RECT 3379.715 3657.775 3588.000 3658.615 ;
        RECT 3379.435 3655.395 3588.000 3657.775 ;
        RECT 3379.715 3654.555 3588.000 3655.395 ;
        RECT 3379.435 3652.175 3588.000 3654.555 ;
        RECT 3379.715 3651.335 3588.000 3652.175 ;
        RECT 3379.435 3649.415 3588.000 3651.335 ;
      LAYER met2 ;
        RECT 3377.035 3648.855 3379.435 3649.135 ;
      LAYER met2 ;
        RECT 3379.715 3648.575 3588.000 3649.415 ;
        RECT 3379.435 3646.195 3588.000 3648.575 ;
        RECT 3379.715 3645.355 3588.000 3646.195 ;
      LAYER met2 ;
        RECT 3376.560 3645.070 3377.160 3645.210 ;
        RECT 3377.020 3642.695 3377.160 3645.070 ;
      LAYER met2 ;
        RECT 3379.435 3642.975 3588.000 3645.355 ;
      LAYER met2 ;
        RECT 3377.020 3642.420 3379.435 3642.695 ;
        RECT 3377.035 3642.415 3379.435 3642.420 ;
      LAYER met2 ;
        RECT 3379.715 3642.135 3588.000 3642.975 ;
        RECT 3379.435 3641.085 3588.000 3642.135 ;
        RECT 0.000 3568.865 208.565 3569.915 ;
        RECT 0.000 3568.025 208.285 3568.865 ;
      LAYER met2 ;
        RECT 208.565 3568.305 210.965 3568.585 ;
      LAYER met2 ;
        RECT 0.000 3565.645 208.565 3568.025 ;
      LAYER met2 ;
        RECT 209.000 3565.910 209.140 3568.305 ;
      LAYER met2 ;
        RECT 0.000 3564.805 208.285 3565.645 ;
      LAYER met2 ;
        RECT 208.940 3565.590 209.200 3565.910 ;
        RECT 211.700 3565.590 211.960 3565.910 ;
      LAYER met2 ;
        RECT 0.000 3562.425 208.565 3564.805 ;
        RECT 0.000 3561.585 208.285 3562.425 ;
      LAYER met2 ;
        RECT 208.565 3561.865 210.965 3562.145 ;
      LAYER met2 ;
        RECT 0.000 3559.665 208.565 3561.585 ;
        RECT 0.000 3558.825 208.285 3559.665 ;
        RECT 0.000 3556.445 208.565 3558.825 ;
        RECT 0.000 3555.605 208.285 3556.445 ;
        RECT 0.000 3553.225 208.565 3555.605 ;
        RECT 0.000 3552.385 208.285 3553.225 ;
        RECT 0.000 3550.465 208.565 3552.385 ;
        RECT 0.000 3549.625 208.285 3550.465 ;
      LAYER met2 ;
        RECT 208.565 3549.905 210.965 3550.185 ;
      LAYER met2 ;
        RECT 0.000 3547.245 208.565 3549.625 ;
        RECT 0.000 3546.405 208.285 3547.245 ;
        RECT 0.000 3544.025 208.565 3546.405 ;
        RECT 0.000 3543.185 208.285 3544.025 ;
      LAYER met2 ;
        RECT 208.565 3543.465 210.965 3543.745 ;
      LAYER met2 ;
        RECT 0.000 3541.265 208.565 3543.185 ;
        RECT 0.000 3540.425 208.285 3541.265 ;
        RECT 0.000 3538.045 208.565 3540.425 ;
        RECT 0.000 3537.205 208.285 3538.045 ;
        RECT 0.000 3534.825 208.565 3537.205 ;
        RECT 0.000 3533.985 208.285 3534.825 ;
        RECT 0.000 3532.065 208.565 3533.985 ;
        RECT 0.000 3531.225 208.285 3532.065 ;
      LAYER met2 ;
        RECT 211.760 3531.230 211.900 3565.590 ;
      LAYER met2 ;
        RECT 0.000 3528.845 208.565 3531.225 ;
      LAYER met2 ;
        RECT 208.940 3530.910 209.200 3531.230 ;
        RECT 211.700 3530.910 211.960 3531.230 ;
      LAYER met2 ;
        RECT 0.000 3528.005 208.285 3528.845 ;
      LAYER met2 ;
        RECT 209.000 3528.565 209.140 3530.910 ;
        RECT 208.565 3528.285 210.965 3528.565 ;
      LAYER met2 ;
        RECT 0.000 3525.625 208.565 3528.005 ;
        RECT 0.000 3524.785 208.285 3525.625 ;
        RECT 0.000 3522.405 208.565 3524.785 ;
        RECT 0.000 3521.565 208.285 3522.405 ;
        RECT 0.000 3519.645 208.565 3521.565 ;
        RECT 0.000 3518.805 208.285 3519.645 ;
        RECT 0.000 3516.425 208.565 3518.805 ;
        RECT 0.000 3515.585 208.285 3516.425 ;
        RECT 0.000 3513.205 208.565 3515.585 ;
        RECT 0.000 3512.365 208.285 3513.205 ;
        RECT 0.000 3510.445 208.565 3512.365 ;
        RECT 0.000 3509.605 208.285 3510.445 ;
        RECT 0.000 3507.225 208.565 3509.605 ;
        RECT 0.000 3506.385 208.285 3507.225 ;
        RECT 0.000 3504.005 208.565 3506.385 ;
        RECT 0.000 3503.165 208.285 3504.005 ;
        RECT 0.000 3501.245 208.565 3503.165 ;
        RECT 0.000 3500.405 208.285 3501.245 ;
        RECT 0.000 3498.025 208.565 3500.405 ;
        RECT 0.000 3497.185 208.285 3498.025 ;
        RECT 0.000 3494.805 208.565 3497.185 ;
        RECT 0.000 3493.965 208.285 3494.805 ;
        RECT 3379.435 3494.795 3588.000 3495.790 ;
      LAYER met2 ;
        RECT 3377.035 3494.235 3379.435 3494.515 ;
      LAYER met2 ;
        RECT 0.000 3492.045 208.565 3493.965 ;
        RECT 3379.715 3493.955 3588.000 3494.795 ;
        RECT 0.000 3491.205 208.285 3492.045 ;
        RECT 3379.435 3492.035 3588.000 3493.955 ;
      LAYER met2 ;
        RECT 208.565 3491.485 210.965 3491.765 ;
      LAYER met2 ;
        RECT 0.000 3490.210 208.565 3491.205 ;
        RECT 3379.715 3491.195 3588.000 3492.035 ;
        RECT 3379.435 3488.815 3588.000 3491.195 ;
        RECT 3379.715 3487.975 3588.000 3488.815 ;
        RECT 3379.435 3485.595 3588.000 3487.975 ;
        RECT 3379.715 3484.755 3588.000 3485.595 ;
        RECT 3379.435 3482.835 3588.000 3484.755 ;
        RECT 3379.715 3481.995 3588.000 3482.835 ;
        RECT 3379.435 3479.615 3588.000 3481.995 ;
        RECT 3379.715 3478.775 3588.000 3479.615 ;
        RECT 3379.435 3476.395 3588.000 3478.775 ;
        RECT 3379.715 3475.555 3588.000 3476.395 ;
        RECT 3379.435 3473.635 3588.000 3475.555 ;
        RECT 3379.715 3472.795 3588.000 3473.635 ;
        RECT 3379.435 3470.415 3588.000 3472.795 ;
        RECT 3379.715 3469.575 3588.000 3470.415 ;
        RECT 3379.435 3467.195 3588.000 3469.575 ;
        RECT 3379.715 3466.355 3588.000 3467.195 ;
        RECT 3379.435 3464.435 3588.000 3466.355 ;
        RECT 3379.715 3463.595 3588.000 3464.435 ;
        RECT 3379.435 3461.215 3588.000 3463.595 ;
        RECT 3379.715 3460.375 3588.000 3461.215 ;
        RECT 3379.435 3457.995 3588.000 3460.375 ;
      LAYER met2 ;
        RECT 3377.035 3457.435 3379.435 3457.715 ;
        RECT 3377.090 3457.390 3377.620 3457.435 ;
        RECT 3377.480 3454.810 3377.620 3457.390 ;
      LAYER met2 ;
        RECT 3379.715 3457.155 3588.000 3457.995 ;
      LAYER met2 ;
        RECT 3376.560 3454.670 3377.620 3454.810 ;
      LAYER met2 ;
        RECT 3379.435 3454.775 3588.000 3457.155 ;
      LAYER met2 ;
        RECT 3376.560 3417.625 3376.700 3454.670 ;
      LAYER met2 ;
        RECT 3379.715 3453.935 3588.000 3454.775 ;
        RECT 3379.435 3452.015 3588.000 3453.935 ;
        RECT 3379.715 3451.175 3588.000 3452.015 ;
        RECT 3379.435 3448.795 3588.000 3451.175 ;
        RECT 3379.715 3447.955 3588.000 3448.795 ;
        RECT 3379.435 3445.575 3588.000 3447.955 ;
        RECT 3379.715 3444.735 3588.000 3445.575 ;
        RECT 3379.435 3442.815 3588.000 3444.735 ;
      LAYER met2 ;
        RECT 3377.035 3442.255 3379.435 3442.535 ;
      LAYER met2 ;
        RECT 3379.715 3441.975 3588.000 3442.815 ;
        RECT 3379.435 3439.595 3588.000 3441.975 ;
        RECT 3379.715 3438.755 3588.000 3439.595 ;
        RECT 3379.435 3436.375 3588.000 3438.755 ;
      LAYER met2 ;
        RECT 3377.035 3435.815 3379.435 3436.095 ;
      LAYER met2 ;
        RECT 3379.715 3435.535 3588.000 3436.375 ;
        RECT 3379.435 3433.615 3588.000 3435.535 ;
        RECT 3379.715 3432.775 3588.000 3433.615 ;
        RECT 3379.435 3430.395 3588.000 3432.775 ;
        RECT 3379.715 3429.555 3588.000 3430.395 ;
        RECT 3379.435 3427.175 3588.000 3429.555 ;
        RECT 3379.715 3426.335 3588.000 3427.175 ;
        RECT 3379.435 3424.415 3588.000 3426.335 ;
      LAYER met2 ;
        RECT 3377.035 3423.855 3379.435 3424.135 ;
      LAYER met2 ;
        RECT 3379.715 3423.575 3588.000 3424.415 ;
        RECT 3379.435 3421.195 3588.000 3423.575 ;
        RECT 3379.715 3420.355 3588.000 3421.195 ;
        RECT 3379.435 3417.975 3588.000 3420.355 ;
      LAYER met2 ;
        RECT 3377.035 3417.625 3379.435 3417.695 ;
        RECT 3376.560 3417.485 3379.435 3417.625 ;
        RECT 3377.035 3417.415 3379.435 3417.485 ;
      LAYER met2 ;
        RECT 3379.715 3417.135 3588.000 3417.975 ;
        RECT 3379.435 3416.085 3588.000 3417.135 ;
        RECT 0.000 3352.865 208.565 3353.915 ;
        RECT 0.000 3352.025 208.285 3352.865 ;
      LAYER met2 ;
        RECT 208.565 3352.305 210.965 3352.585 ;
      LAYER met2 ;
        RECT 0.000 3349.645 208.565 3352.025 ;
      LAYER met2 ;
        RECT 209.000 3350.010 209.140 3352.305 ;
        RECT 208.940 3349.690 209.200 3350.010 ;
        RECT 211.700 3349.690 211.960 3350.010 ;
      LAYER met2 ;
        RECT 0.000 3348.805 208.285 3349.645 ;
        RECT 0.000 3346.425 208.565 3348.805 ;
        RECT 0.000 3345.585 208.285 3346.425 ;
      LAYER met2 ;
        RECT 208.565 3345.865 210.965 3346.145 ;
      LAYER met2 ;
        RECT 0.000 3343.665 208.565 3345.585 ;
        RECT 0.000 3342.825 208.285 3343.665 ;
        RECT 0.000 3340.445 208.565 3342.825 ;
        RECT 0.000 3339.605 208.285 3340.445 ;
        RECT 0.000 3337.225 208.565 3339.605 ;
        RECT 0.000 3336.385 208.285 3337.225 ;
        RECT 0.000 3334.465 208.565 3336.385 ;
        RECT 0.000 3333.625 208.285 3334.465 ;
      LAYER met2 ;
        RECT 208.565 3333.905 210.965 3334.185 ;
      LAYER met2 ;
        RECT 0.000 3331.245 208.565 3333.625 ;
        RECT 0.000 3330.405 208.285 3331.245 ;
        RECT 0.000 3328.025 208.565 3330.405 ;
        RECT 0.000 3327.185 208.285 3328.025 ;
      LAYER met2 ;
        RECT 208.565 3327.465 210.965 3327.745 ;
      LAYER met2 ;
        RECT 0.000 3325.265 208.565 3327.185 ;
        RECT 0.000 3324.425 208.285 3325.265 ;
        RECT 0.000 3322.045 208.565 3324.425 ;
        RECT 0.000 3321.205 208.285 3322.045 ;
        RECT 0.000 3318.825 208.565 3321.205 ;
        RECT 0.000 3317.985 208.285 3318.825 ;
        RECT 0.000 3316.065 208.565 3317.985 ;
        RECT 0.000 3315.225 208.285 3316.065 ;
      LAYER met2 ;
        RECT 211.760 3315.330 211.900 3349.690 ;
      LAYER met2 ;
        RECT 0.000 3312.845 208.565 3315.225 ;
      LAYER met2 ;
        RECT 208.940 3315.010 209.200 3315.330 ;
        RECT 211.700 3315.010 211.960 3315.330 ;
      LAYER met2 ;
        RECT 0.000 3312.005 208.285 3312.845 ;
      LAYER met2 ;
        RECT 209.000 3312.565 209.140 3315.010 ;
        RECT 208.565 3312.285 210.965 3312.565 ;
      LAYER met2 ;
        RECT 0.000 3309.625 208.565 3312.005 ;
        RECT 0.000 3308.785 208.285 3309.625 ;
        RECT 0.000 3306.405 208.565 3308.785 ;
        RECT 0.000 3305.565 208.285 3306.405 ;
        RECT 0.000 3303.645 208.565 3305.565 ;
        RECT 0.000 3302.805 208.285 3303.645 ;
        RECT 0.000 3300.425 208.565 3302.805 ;
        RECT 0.000 3299.585 208.285 3300.425 ;
        RECT 0.000 3297.205 208.565 3299.585 ;
        RECT 0.000 3296.365 208.285 3297.205 ;
        RECT 0.000 3294.445 208.565 3296.365 ;
        RECT 0.000 3293.605 208.285 3294.445 ;
        RECT 0.000 3291.225 208.565 3293.605 ;
        RECT 0.000 3290.385 208.285 3291.225 ;
        RECT 0.000 3288.005 208.565 3290.385 ;
        RECT 0.000 3287.165 208.285 3288.005 ;
        RECT 0.000 3285.245 208.565 3287.165 ;
        RECT 0.000 3284.405 208.285 3285.245 ;
        RECT 0.000 3282.025 208.565 3284.405 ;
        RECT 0.000 3281.185 208.285 3282.025 ;
        RECT 0.000 3278.805 208.565 3281.185 ;
        RECT 0.000 3277.965 208.285 3278.805 ;
        RECT 0.000 3276.045 208.565 3277.965 ;
        RECT 0.000 3275.205 208.285 3276.045 ;
      LAYER met2 ;
        RECT 208.565 3275.485 210.965 3275.765 ;
      LAYER met2 ;
        RECT 0.000 3274.210 208.565 3275.205 ;
        RECT 3379.435 3268.795 3588.000 3269.790 ;
      LAYER met2 ;
        RECT 3377.035 3268.235 3379.435 3268.515 ;
      LAYER met2 ;
        RECT 3379.715 3267.955 3588.000 3268.795 ;
        RECT 3379.435 3266.035 3588.000 3267.955 ;
        RECT 3379.715 3265.195 3588.000 3266.035 ;
        RECT 3379.435 3262.815 3588.000 3265.195 ;
        RECT 3379.715 3261.975 3588.000 3262.815 ;
        RECT 3379.435 3259.595 3588.000 3261.975 ;
        RECT 3379.715 3258.755 3588.000 3259.595 ;
        RECT 3379.435 3256.835 3588.000 3258.755 ;
        RECT 3379.715 3255.995 3588.000 3256.835 ;
        RECT 3379.435 3253.615 3588.000 3255.995 ;
        RECT 3379.715 3252.775 3588.000 3253.615 ;
        RECT 3379.435 3250.395 3588.000 3252.775 ;
        RECT 3379.715 3249.555 3588.000 3250.395 ;
        RECT 3379.435 3247.635 3588.000 3249.555 ;
        RECT 3379.715 3246.795 3588.000 3247.635 ;
        RECT 3379.435 3244.415 3588.000 3246.795 ;
        RECT 3379.715 3243.575 3588.000 3244.415 ;
        RECT 3379.435 3241.195 3588.000 3243.575 ;
        RECT 3379.715 3240.355 3588.000 3241.195 ;
        RECT 3379.435 3238.435 3588.000 3240.355 ;
        RECT 3379.715 3237.595 3588.000 3238.435 ;
        RECT 3379.435 3235.215 3588.000 3237.595 ;
        RECT 3379.715 3234.375 3588.000 3235.215 ;
        RECT 3379.435 3231.995 3588.000 3234.375 ;
      LAYER met2 ;
        RECT 3377.035 3231.700 3379.435 3231.715 ;
        RECT 3377.020 3231.435 3379.435 3231.700 ;
        RECT 3377.020 3229.730 3377.160 3231.435 ;
      LAYER met2 ;
        RECT 3379.715 3231.155 3588.000 3231.995 ;
      LAYER met2 ;
        RECT 3376.100 3229.590 3377.160 3229.730 ;
        RECT 3376.100 3194.290 3376.240 3229.590 ;
      LAYER met2 ;
        RECT 3379.435 3228.775 3588.000 3231.155 ;
        RECT 3379.715 3227.935 3588.000 3228.775 ;
        RECT 3379.435 3226.015 3588.000 3227.935 ;
        RECT 3379.715 3225.175 3588.000 3226.015 ;
        RECT 3379.435 3222.795 3588.000 3225.175 ;
        RECT 3379.715 3221.955 3588.000 3222.795 ;
        RECT 3379.435 3219.575 3588.000 3221.955 ;
        RECT 3379.715 3218.735 3588.000 3219.575 ;
        RECT 3379.435 3216.815 3588.000 3218.735 ;
      LAYER met2 ;
        RECT 3377.035 3216.255 3379.435 3216.535 ;
      LAYER met2 ;
        RECT 3379.715 3215.975 3588.000 3216.815 ;
        RECT 3379.435 3213.595 3588.000 3215.975 ;
        RECT 3379.715 3212.755 3588.000 3213.595 ;
        RECT 3379.435 3210.375 3588.000 3212.755 ;
      LAYER met2 ;
        RECT 3377.035 3209.815 3379.435 3210.095 ;
      LAYER met2 ;
        RECT 3379.715 3209.535 3588.000 3210.375 ;
        RECT 3379.435 3207.615 3588.000 3209.535 ;
        RECT 3379.715 3206.775 3588.000 3207.615 ;
        RECT 3379.435 3204.395 3588.000 3206.775 ;
        RECT 3379.715 3203.555 3588.000 3204.395 ;
        RECT 3379.435 3201.175 3588.000 3203.555 ;
        RECT 3379.715 3200.335 3588.000 3201.175 ;
        RECT 3379.435 3198.415 3588.000 3200.335 ;
      LAYER met2 ;
        RECT 3377.035 3197.855 3379.435 3198.135 ;
      LAYER met2 ;
        RECT 3379.715 3197.575 3588.000 3198.415 ;
        RECT 3379.435 3195.195 3588.000 3197.575 ;
        RECT 3379.715 3194.355 3588.000 3195.195 ;
      LAYER met2 ;
        RECT 3376.040 3193.970 3376.300 3194.290 ;
        RECT 3376.960 3193.970 3377.220 3194.290 ;
        RECT 3377.020 3191.695 3377.160 3193.970 ;
      LAYER met2 ;
        RECT 3379.435 3191.975 3588.000 3194.355 ;
      LAYER met2 ;
        RECT 3377.020 3191.580 3379.435 3191.695 ;
        RECT 3377.035 3191.415 3379.435 3191.580 ;
      LAYER met2 ;
        RECT 3379.715 3191.135 3588.000 3191.975 ;
        RECT 3379.435 3190.085 3588.000 3191.135 ;
        RECT 0.000 3136.865 208.565 3137.915 ;
        RECT 0.000 3136.025 208.285 3136.865 ;
      LAYER met2 ;
        RECT 208.565 3136.305 210.965 3136.585 ;
      LAYER met2 ;
        RECT 0.000 3133.645 208.565 3136.025 ;
      LAYER met2 ;
        RECT 209.000 3134.110 209.140 3136.305 ;
        RECT 208.940 3133.790 209.200 3134.110 ;
        RECT 211.700 3133.790 211.960 3134.110 ;
      LAYER met2 ;
        RECT 0.000 3132.805 208.285 3133.645 ;
        RECT 0.000 3130.425 208.565 3132.805 ;
        RECT 0.000 3129.585 208.285 3130.425 ;
      LAYER met2 ;
        RECT 208.565 3129.865 210.965 3130.145 ;
      LAYER met2 ;
        RECT 0.000 3127.665 208.565 3129.585 ;
        RECT 0.000 3126.825 208.285 3127.665 ;
        RECT 0.000 3124.445 208.565 3126.825 ;
        RECT 0.000 3123.605 208.285 3124.445 ;
        RECT 0.000 3121.225 208.565 3123.605 ;
        RECT 0.000 3120.385 208.285 3121.225 ;
        RECT 0.000 3118.465 208.565 3120.385 ;
        RECT 0.000 3117.625 208.285 3118.465 ;
      LAYER met2 ;
        RECT 208.565 3117.905 210.965 3118.185 ;
      LAYER met2 ;
        RECT 0.000 3115.245 208.565 3117.625 ;
        RECT 0.000 3114.405 208.285 3115.245 ;
        RECT 0.000 3112.025 208.565 3114.405 ;
        RECT 0.000 3111.185 208.285 3112.025 ;
      LAYER met2 ;
        RECT 208.565 3111.465 210.965 3111.745 ;
      LAYER met2 ;
        RECT 0.000 3109.265 208.565 3111.185 ;
        RECT 0.000 3108.425 208.285 3109.265 ;
        RECT 0.000 3106.045 208.565 3108.425 ;
        RECT 0.000 3105.205 208.285 3106.045 ;
        RECT 0.000 3102.825 208.565 3105.205 ;
        RECT 0.000 3101.985 208.285 3102.825 ;
        RECT 0.000 3100.065 208.565 3101.985 ;
        RECT 0.000 3099.225 208.285 3100.065 ;
        RECT 0.000 3096.845 208.565 3099.225 ;
      LAYER met2 ;
        RECT 211.760 3099.090 211.900 3133.790 ;
        RECT 208.940 3098.770 209.200 3099.090 ;
        RECT 211.700 3098.770 211.960 3099.090 ;
      LAYER met2 ;
        RECT 0.000 3096.005 208.285 3096.845 ;
      LAYER met2 ;
        RECT 209.000 3096.565 209.140 3098.770 ;
        RECT 208.565 3096.285 210.965 3096.565 ;
      LAYER met2 ;
        RECT 0.000 3093.625 208.565 3096.005 ;
        RECT 0.000 3092.785 208.285 3093.625 ;
        RECT 0.000 3090.405 208.565 3092.785 ;
        RECT 0.000 3089.565 208.285 3090.405 ;
        RECT 0.000 3087.645 208.565 3089.565 ;
        RECT 0.000 3086.805 208.285 3087.645 ;
        RECT 0.000 3084.425 208.565 3086.805 ;
        RECT 0.000 3083.585 208.285 3084.425 ;
        RECT 0.000 3081.205 208.565 3083.585 ;
        RECT 0.000 3080.365 208.285 3081.205 ;
        RECT 0.000 3078.445 208.565 3080.365 ;
        RECT 0.000 3077.605 208.285 3078.445 ;
        RECT 0.000 3075.225 208.565 3077.605 ;
        RECT 0.000 3074.385 208.285 3075.225 ;
        RECT 0.000 3072.005 208.565 3074.385 ;
        RECT 0.000 3071.165 208.285 3072.005 ;
        RECT 0.000 3069.245 208.565 3071.165 ;
        RECT 0.000 3068.405 208.285 3069.245 ;
        RECT 0.000 3066.025 208.565 3068.405 ;
        RECT 0.000 3065.185 208.285 3066.025 ;
        RECT 0.000 3062.805 208.565 3065.185 ;
        RECT 0.000 3061.965 208.285 3062.805 ;
        RECT 0.000 3060.045 208.565 3061.965 ;
        RECT 0.000 3059.205 208.285 3060.045 ;
      LAYER met2 ;
        RECT 208.565 3059.485 210.965 3059.765 ;
      LAYER met2 ;
        RECT 0.000 3058.210 208.565 3059.205 ;
        RECT 3379.435 3043.795 3588.000 3044.790 ;
      LAYER met2 ;
        RECT 3377.035 3043.235 3379.435 3043.515 ;
      LAYER met2 ;
        RECT 3379.715 3042.955 3588.000 3043.795 ;
        RECT 3379.435 3041.035 3588.000 3042.955 ;
        RECT 3379.715 3040.195 3588.000 3041.035 ;
        RECT 3379.435 3037.815 3588.000 3040.195 ;
        RECT 3379.715 3036.975 3588.000 3037.815 ;
        RECT 3379.435 3034.595 3588.000 3036.975 ;
        RECT 3379.715 3033.755 3588.000 3034.595 ;
        RECT 3379.435 3031.835 3588.000 3033.755 ;
        RECT 3379.715 3030.995 3588.000 3031.835 ;
        RECT 3379.435 3028.615 3588.000 3030.995 ;
        RECT 3379.715 3027.775 3588.000 3028.615 ;
        RECT 3379.435 3025.395 3588.000 3027.775 ;
        RECT 3379.715 3024.555 3588.000 3025.395 ;
        RECT 3379.435 3022.635 3588.000 3024.555 ;
        RECT 3379.715 3021.795 3588.000 3022.635 ;
        RECT 3379.435 3019.415 3588.000 3021.795 ;
        RECT 3379.715 3018.575 3588.000 3019.415 ;
        RECT 3379.435 3016.195 3588.000 3018.575 ;
        RECT 3379.715 3015.355 3588.000 3016.195 ;
        RECT 3379.435 3013.435 3588.000 3015.355 ;
        RECT 3379.715 3012.595 3588.000 3013.435 ;
        RECT 3379.435 3010.215 3588.000 3012.595 ;
        RECT 3379.715 3009.375 3588.000 3010.215 ;
        RECT 3379.435 3006.995 3588.000 3009.375 ;
      LAYER met2 ;
        RECT 3377.035 3006.620 3379.435 3006.715 ;
        RECT 3377.020 3006.435 3379.435 3006.620 ;
        RECT 3377.020 3004.230 3377.160 3006.435 ;
      LAYER met2 ;
        RECT 3379.715 3006.155 3588.000 3006.995 ;
      LAYER met2 ;
        RECT 3376.040 3003.910 3376.300 3004.230 ;
        RECT 3376.960 3003.910 3377.220 3004.230 ;
        RECT 3376.100 2966.570 3376.240 3003.910 ;
      LAYER met2 ;
        RECT 3379.435 3003.775 3588.000 3006.155 ;
        RECT 3379.715 3002.935 3588.000 3003.775 ;
        RECT 3379.435 3001.015 3588.000 3002.935 ;
        RECT 3379.715 3000.175 3588.000 3001.015 ;
        RECT 3379.435 2997.795 3588.000 3000.175 ;
        RECT 3379.715 2996.955 3588.000 2997.795 ;
        RECT 3379.435 2994.575 3588.000 2996.955 ;
        RECT 3379.715 2993.735 3588.000 2994.575 ;
        RECT 3379.435 2991.815 3588.000 2993.735 ;
      LAYER met2 ;
        RECT 3377.035 2991.255 3379.435 2991.535 ;
      LAYER met2 ;
        RECT 3379.715 2990.975 3588.000 2991.815 ;
        RECT 3379.435 2988.595 3588.000 2990.975 ;
        RECT 3379.715 2987.755 3588.000 2988.595 ;
        RECT 3379.435 2985.375 3588.000 2987.755 ;
      LAYER met2 ;
        RECT 3377.035 2984.815 3379.435 2985.095 ;
      LAYER met2 ;
        RECT 3379.715 2984.535 3588.000 2985.375 ;
        RECT 3379.435 2982.615 3588.000 2984.535 ;
        RECT 3379.715 2981.775 3588.000 2982.615 ;
        RECT 3379.435 2979.395 3588.000 2981.775 ;
        RECT 3379.715 2978.555 3588.000 2979.395 ;
        RECT 3379.435 2976.175 3588.000 2978.555 ;
        RECT 3379.715 2975.335 3588.000 2976.175 ;
        RECT 3379.435 2973.415 3588.000 2975.335 ;
      LAYER met2 ;
        RECT 3377.035 2972.855 3379.435 2973.135 ;
      LAYER met2 ;
        RECT 3379.715 2972.575 3588.000 2973.415 ;
        RECT 3379.435 2970.195 3588.000 2972.575 ;
        RECT 3379.715 2969.355 3588.000 2970.195 ;
        RECT 3379.435 2966.975 3588.000 2969.355 ;
      LAYER met2 ;
        RECT 3377.035 2966.570 3379.435 2966.695 ;
        RECT 3376.100 2966.430 3379.435 2966.570 ;
        RECT 3377.035 2966.415 3379.435 2966.430 ;
      LAYER met2 ;
        RECT 3379.715 2966.135 3588.000 2966.975 ;
        RECT 3379.435 2965.085 3588.000 2966.135 ;
        RECT 0.000 2920.865 208.565 2921.915 ;
        RECT 0.000 2920.025 208.285 2920.865 ;
      LAYER met2 ;
        RECT 208.565 2920.305 210.965 2920.585 ;
      LAYER met2 ;
        RECT 0.000 2917.645 208.565 2920.025 ;
      LAYER met2 ;
        RECT 209.000 2917.870 209.140 2920.305 ;
      LAYER met2 ;
        RECT 0.000 2916.805 208.285 2917.645 ;
      LAYER met2 ;
        RECT 208.940 2917.550 209.200 2917.870 ;
        RECT 211.700 2917.550 211.960 2917.870 ;
      LAYER met2 ;
        RECT 0.000 2914.425 208.565 2916.805 ;
        RECT 0.000 2913.585 208.285 2914.425 ;
      LAYER met2 ;
        RECT 208.565 2913.865 210.965 2914.145 ;
      LAYER met2 ;
        RECT 0.000 2911.665 208.565 2913.585 ;
        RECT 0.000 2910.825 208.285 2911.665 ;
        RECT 0.000 2908.445 208.565 2910.825 ;
        RECT 0.000 2907.605 208.285 2908.445 ;
        RECT 0.000 2905.225 208.565 2907.605 ;
        RECT 0.000 2904.385 208.285 2905.225 ;
        RECT 0.000 2902.465 208.565 2904.385 ;
        RECT 0.000 2901.625 208.285 2902.465 ;
      LAYER met2 ;
        RECT 208.565 2901.905 210.965 2902.185 ;
      LAYER met2 ;
        RECT 0.000 2899.245 208.565 2901.625 ;
        RECT 0.000 2898.405 208.285 2899.245 ;
        RECT 0.000 2896.025 208.565 2898.405 ;
        RECT 0.000 2895.185 208.285 2896.025 ;
      LAYER met2 ;
        RECT 208.565 2895.465 210.965 2895.745 ;
      LAYER met2 ;
        RECT 0.000 2893.265 208.565 2895.185 ;
        RECT 0.000 2892.425 208.285 2893.265 ;
        RECT 0.000 2890.045 208.565 2892.425 ;
        RECT 0.000 2889.205 208.285 2890.045 ;
        RECT 0.000 2886.825 208.565 2889.205 ;
        RECT 0.000 2885.985 208.285 2886.825 ;
        RECT 0.000 2884.065 208.565 2885.985 ;
        RECT 0.000 2883.225 208.285 2884.065 ;
        RECT 0.000 2880.845 208.565 2883.225 ;
      LAYER met2 ;
        RECT 211.760 2883.190 211.900 2917.550 ;
        RECT 208.940 2882.870 209.200 2883.190 ;
        RECT 211.700 2882.870 211.960 2883.190 ;
      LAYER met2 ;
        RECT 0.000 2880.005 208.285 2880.845 ;
      LAYER met2 ;
        RECT 209.000 2880.565 209.140 2882.870 ;
        RECT 208.565 2880.285 210.965 2880.565 ;
      LAYER met2 ;
        RECT 0.000 2877.625 208.565 2880.005 ;
        RECT 0.000 2876.785 208.285 2877.625 ;
        RECT 0.000 2874.405 208.565 2876.785 ;
        RECT 0.000 2873.565 208.285 2874.405 ;
        RECT 0.000 2871.645 208.565 2873.565 ;
        RECT 0.000 2870.805 208.285 2871.645 ;
        RECT 0.000 2868.425 208.565 2870.805 ;
        RECT 0.000 2867.585 208.285 2868.425 ;
        RECT 0.000 2865.205 208.565 2867.585 ;
        RECT 0.000 2864.365 208.285 2865.205 ;
        RECT 0.000 2862.445 208.565 2864.365 ;
        RECT 0.000 2861.605 208.285 2862.445 ;
        RECT 0.000 2859.225 208.565 2861.605 ;
        RECT 0.000 2858.385 208.285 2859.225 ;
        RECT 0.000 2856.005 208.565 2858.385 ;
        RECT 0.000 2855.165 208.285 2856.005 ;
        RECT 0.000 2853.245 208.565 2855.165 ;
        RECT 0.000 2852.405 208.285 2853.245 ;
        RECT 0.000 2850.025 208.565 2852.405 ;
        RECT 0.000 2849.185 208.285 2850.025 ;
        RECT 0.000 2846.805 208.565 2849.185 ;
        RECT 0.000 2845.965 208.285 2846.805 ;
        RECT 0.000 2844.045 208.565 2845.965 ;
        RECT 0.000 2843.205 208.285 2844.045 ;
      LAYER met2 ;
        RECT 208.565 2843.485 210.965 2843.765 ;
      LAYER met2 ;
        RECT 0.000 2842.210 208.565 2843.205 ;
        RECT 3379.435 2817.795 3588.000 2818.790 ;
      LAYER met2 ;
        RECT 3377.035 2817.235 3379.435 2817.515 ;
      LAYER met2 ;
        RECT 3379.715 2816.955 3588.000 2817.795 ;
        RECT 3379.435 2815.035 3588.000 2816.955 ;
        RECT 3379.715 2814.195 3588.000 2815.035 ;
        RECT 3379.435 2811.815 3588.000 2814.195 ;
        RECT 3379.715 2810.975 3588.000 2811.815 ;
        RECT 3379.435 2808.595 3588.000 2810.975 ;
        RECT 3379.715 2807.755 3588.000 2808.595 ;
        RECT 3379.435 2805.835 3588.000 2807.755 ;
        RECT 3379.715 2804.995 3588.000 2805.835 ;
        RECT 3379.435 2802.615 3588.000 2804.995 ;
        RECT 3379.715 2801.775 3588.000 2802.615 ;
        RECT 3379.435 2799.395 3588.000 2801.775 ;
        RECT 3379.715 2798.555 3588.000 2799.395 ;
        RECT 3379.435 2796.635 3588.000 2798.555 ;
        RECT 3379.715 2795.795 3588.000 2796.635 ;
        RECT 3379.435 2793.415 3588.000 2795.795 ;
        RECT 3379.715 2792.575 3588.000 2793.415 ;
        RECT 3379.435 2790.195 3588.000 2792.575 ;
        RECT 3379.715 2789.355 3588.000 2790.195 ;
        RECT 3379.435 2787.435 3588.000 2789.355 ;
        RECT 3379.715 2786.595 3588.000 2787.435 ;
        RECT 3379.435 2784.215 3588.000 2786.595 ;
        RECT 3379.715 2783.375 3588.000 2784.215 ;
        RECT 3379.435 2780.995 3588.000 2783.375 ;
      LAYER met2 ;
        RECT 3377.035 2780.645 3379.435 2780.715 ;
        RECT 3376.560 2780.505 3379.435 2780.645 ;
        RECT 3376.560 2742.850 3376.700 2780.505 ;
        RECT 3377.035 2780.435 3379.435 2780.505 ;
      LAYER met2 ;
        RECT 3379.715 2780.155 3588.000 2780.995 ;
        RECT 3379.435 2777.775 3588.000 2780.155 ;
        RECT 3379.715 2776.935 3588.000 2777.775 ;
        RECT 3379.435 2775.015 3588.000 2776.935 ;
        RECT 3379.715 2774.175 3588.000 2775.015 ;
        RECT 3379.435 2771.795 3588.000 2774.175 ;
        RECT 3379.715 2770.955 3588.000 2771.795 ;
        RECT 3379.435 2768.575 3588.000 2770.955 ;
        RECT 3379.715 2767.735 3588.000 2768.575 ;
        RECT 3379.435 2765.815 3588.000 2767.735 ;
      LAYER met2 ;
        RECT 3377.035 2765.255 3379.435 2765.535 ;
      LAYER met2 ;
        RECT 3379.715 2764.975 3588.000 2765.815 ;
        RECT 3379.435 2762.595 3588.000 2764.975 ;
        RECT 3379.715 2761.755 3588.000 2762.595 ;
        RECT 3379.435 2759.375 3588.000 2761.755 ;
      LAYER met2 ;
        RECT 3377.035 2758.815 3379.435 2759.095 ;
      LAYER met2 ;
        RECT 3379.715 2758.535 3588.000 2759.375 ;
        RECT 3379.435 2756.615 3588.000 2758.535 ;
        RECT 3379.715 2755.775 3588.000 2756.615 ;
        RECT 3379.435 2753.395 3588.000 2755.775 ;
        RECT 3379.715 2752.555 3588.000 2753.395 ;
        RECT 3379.435 2750.175 3588.000 2752.555 ;
        RECT 3379.715 2749.335 3588.000 2750.175 ;
        RECT 3379.435 2747.415 3588.000 2749.335 ;
      LAYER met2 ;
        RECT 3377.035 2746.855 3379.435 2747.135 ;
      LAYER met2 ;
        RECT 3379.715 2746.575 3588.000 2747.415 ;
        RECT 3379.435 2744.195 3588.000 2746.575 ;
        RECT 3379.715 2743.355 3588.000 2744.195 ;
      LAYER met2 ;
        RECT 3376.560 2742.710 3377.160 2742.850 ;
        RECT 3377.020 2740.695 3377.160 2742.710 ;
      LAYER met2 ;
        RECT 3379.435 2740.975 3588.000 2743.355 ;
      LAYER met2 ;
        RECT 3377.020 2740.555 3379.435 2740.695 ;
        RECT 3377.035 2740.415 3379.435 2740.555 ;
      LAYER met2 ;
        RECT 3379.715 2740.135 3588.000 2740.975 ;
        RECT 3379.435 2739.085 3588.000 2740.135 ;
        RECT 0.000 2704.865 208.565 2705.915 ;
        RECT 0.000 2704.025 208.285 2704.865 ;
      LAYER met2 ;
        RECT 208.565 2704.305 210.965 2704.585 ;
      LAYER met2 ;
        RECT 0.000 2701.645 208.565 2704.025 ;
      LAYER met2 ;
        RECT 209.000 2701.970 209.140 2704.305 ;
        RECT 208.940 2701.650 209.200 2701.970 ;
        RECT 211.700 2701.650 211.960 2701.970 ;
      LAYER met2 ;
        RECT 0.000 2700.805 208.285 2701.645 ;
        RECT 0.000 2698.425 208.565 2700.805 ;
        RECT 0.000 2697.585 208.285 2698.425 ;
      LAYER met2 ;
        RECT 208.565 2697.865 210.965 2698.145 ;
      LAYER met2 ;
        RECT 0.000 2695.665 208.565 2697.585 ;
        RECT 0.000 2694.825 208.285 2695.665 ;
        RECT 0.000 2692.445 208.565 2694.825 ;
        RECT 0.000 2691.605 208.285 2692.445 ;
        RECT 0.000 2689.225 208.565 2691.605 ;
        RECT 0.000 2688.385 208.285 2689.225 ;
        RECT 0.000 2686.465 208.565 2688.385 ;
        RECT 0.000 2685.625 208.285 2686.465 ;
      LAYER met2 ;
        RECT 208.565 2685.905 210.965 2686.185 ;
      LAYER met2 ;
        RECT 0.000 2683.245 208.565 2685.625 ;
        RECT 0.000 2682.405 208.285 2683.245 ;
        RECT 0.000 2680.025 208.565 2682.405 ;
        RECT 0.000 2679.185 208.285 2680.025 ;
      LAYER met2 ;
        RECT 208.565 2679.465 210.965 2679.745 ;
      LAYER met2 ;
        RECT 0.000 2677.265 208.565 2679.185 ;
        RECT 0.000 2676.425 208.285 2677.265 ;
        RECT 0.000 2674.045 208.565 2676.425 ;
        RECT 0.000 2673.205 208.285 2674.045 ;
        RECT 0.000 2670.825 208.565 2673.205 ;
        RECT 0.000 2669.985 208.285 2670.825 ;
        RECT 0.000 2668.065 208.565 2669.985 ;
        RECT 0.000 2667.225 208.285 2668.065 ;
      LAYER met2 ;
        RECT 211.760 2667.290 211.900 2701.650 ;
      LAYER met2 ;
        RECT 0.000 2664.845 208.565 2667.225 ;
      LAYER met2 ;
        RECT 208.940 2666.970 209.200 2667.290 ;
        RECT 211.700 2666.970 211.960 2667.290 ;
      LAYER met2 ;
        RECT 0.000 2664.005 208.285 2664.845 ;
      LAYER met2 ;
        RECT 209.000 2664.565 209.140 2666.970 ;
        RECT 208.565 2664.285 210.965 2664.565 ;
      LAYER met2 ;
        RECT 0.000 2661.625 208.565 2664.005 ;
        RECT 0.000 2660.785 208.285 2661.625 ;
        RECT 0.000 2658.405 208.565 2660.785 ;
        RECT 0.000 2657.565 208.285 2658.405 ;
        RECT 0.000 2655.645 208.565 2657.565 ;
        RECT 0.000 2654.805 208.285 2655.645 ;
        RECT 0.000 2652.425 208.565 2654.805 ;
        RECT 0.000 2651.585 208.285 2652.425 ;
        RECT 0.000 2649.205 208.565 2651.585 ;
        RECT 0.000 2648.365 208.285 2649.205 ;
        RECT 0.000 2646.445 208.565 2648.365 ;
        RECT 0.000 2645.605 208.285 2646.445 ;
        RECT 0.000 2643.225 208.565 2645.605 ;
        RECT 0.000 2642.385 208.285 2643.225 ;
        RECT 0.000 2640.005 208.565 2642.385 ;
        RECT 0.000 2639.165 208.285 2640.005 ;
        RECT 0.000 2637.245 208.565 2639.165 ;
        RECT 0.000 2636.405 208.285 2637.245 ;
        RECT 0.000 2634.025 208.565 2636.405 ;
        RECT 0.000 2633.185 208.285 2634.025 ;
        RECT 0.000 2630.805 208.565 2633.185 ;
        RECT 0.000 2629.965 208.285 2630.805 ;
        RECT 0.000 2628.045 208.565 2629.965 ;
        RECT 0.000 2627.205 208.285 2628.045 ;
      LAYER met2 ;
        RECT 208.565 2627.485 210.965 2627.765 ;
      LAYER met2 ;
        RECT 0.000 2626.210 208.565 2627.205 ;
        RECT 3390.035 2593.505 3583.075 2593.735 ;
        RECT 3388.000 2569.605 3583.075 2593.505 ;
        RECT 3388.000 2566.105 3389.920 2568.105 ;
        RECT 3390.035 2543.610 3583.075 2569.605 ;
        RECT 3388.000 2519.710 3583.075 2543.610 ;
        RECT 4.925 2465.390 200.000 2489.290 ;
        RECT 4.925 2439.395 197.965 2465.390 ;
        RECT 198.080 2440.895 200.000 2442.895 ;
        RECT 4.925 2415.495 200.000 2439.395 ;
        RECT 4.925 2415.265 197.965 2415.495 ;
        RECT 3390.000 2353.505 3584.430 2373.500 ;
        RECT 3390.035 2353.075 3584.430 2353.505 ;
        RECT 3390.000 2320.465 3584.430 2353.075 ;
        RECT 3390.035 2319.905 3584.430 2320.465 ;
        RECT 3390.000 2299.300 3584.430 2319.905 ;
        RECT 3390.035 2299.000 3584.430 2299.300 ;
        RECT 153.765 2279.000 158.415 2290.140 ;
        RECT 159.640 2279.245 163.510 2290.195 ;
        RECT 3424.490 2287.805 3428.360 2298.755 ;
        RECT 3429.585 2287.860 3434.235 2299.000 ;
        RECT 3.570 2278.700 197.965 2279.000 ;
        RECT 3.570 2258.095 198.000 2278.700 ;
        RECT 3.570 2257.535 197.965 2258.095 ;
        RECT 3.570 2224.925 198.000 2257.535 ;
        RECT 3.570 2224.495 197.965 2224.925 ;
        RECT 3.570 2204.500 198.000 2224.495 ;
        RECT 3390.035 2152.505 3583.075 2152.735 ;
        RECT 3388.000 2128.605 3583.075 2152.505 ;
        RECT 3388.000 2125.105 3389.920 2127.105 ;
        RECT 3390.035 2102.610 3583.075 2128.605 ;
        RECT 3388.000 2078.710 3583.075 2102.610 ;
        RECT 0.000 2066.865 208.565 2067.915 ;
        RECT 0.000 2066.025 208.285 2066.865 ;
      LAYER met2 ;
        RECT 208.565 2066.305 210.965 2066.585 ;
      LAYER met2 ;
        RECT 0.000 2063.645 208.565 2066.025 ;
      LAYER met2 ;
        RECT 209.000 2064.130 209.140 2066.305 ;
        RECT 208.940 2063.810 209.200 2064.130 ;
        RECT 211.700 2063.810 211.960 2064.130 ;
      LAYER met2 ;
        RECT 0.000 2062.805 208.285 2063.645 ;
        RECT 0.000 2060.425 208.565 2062.805 ;
        RECT 0.000 2059.585 208.285 2060.425 ;
      LAYER met2 ;
        RECT 208.565 2059.865 210.965 2060.145 ;
      LAYER met2 ;
        RECT 0.000 2057.665 208.565 2059.585 ;
        RECT 0.000 2056.825 208.285 2057.665 ;
        RECT 0.000 2054.445 208.565 2056.825 ;
        RECT 0.000 2053.605 208.285 2054.445 ;
        RECT 0.000 2051.225 208.565 2053.605 ;
        RECT 0.000 2050.385 208.285 2051.225 ;
        RECT 0.000 2048.465 208.565 2050.385 ;
        RECT 0.000 2047.625 208.285 2048.465 ;
      LAYER met2 ;
        RECT 208.565 2047.905 210.965 2048.185 ;
      LAYER met2 ;
        RECT 0.000 2045.245 208.565 2047.625 ;
        RECT 0.000 2044.405 208.285 2045.245 ;
        RECT 0.000 2042.025 208.565 2044.405 ;
        RECT 0.000 2041.185 208.285 2042.025 ;
      LAYER met2 ;
        RECT 208.565 2041.465 210.965 2041.745 ;
      LAYER met2 ;
        RECT 0.000 2039.265 208.565 2041.185 ;
        RECT 0.000 2038.425 208.285 2039.265 ;
        RECT 0.000 2036.045 208.565 2038.425 ;
        RECT 0.000 2035.205 208.285 2036.045 ;
        RECT 0.000 2032.825 208.565 2035.205 ;
        RECT 0.000 2031.985 208.285 2032.825 ;
        RECT 0.000 2030.065 208.565 2031.985 ;
        RECT 0.000 2029.225 208.285 2030.065 ;
        RECT 0.000 2026.845 208.565 2029.225 ;
      LAYER met2 ;
        RECT 211.760 2029.110 211.900 2063.810 ;
        RECT 208.940 2028.790 209.200 2029.110 ;
        RECT 211.700 2028.790 211.960 2029.110 ;
      LAYER met2 ;
        RECT 0.000 2026.005 208.285 2026.845 ;
      LAYER met2 ;
        RECT 209.000 2026.565 209.140 2028.790 ;
        RECT 208.565 2026.285 210.965 2026.565 ;
      LAYER met2 ;
        RECT 0.000 2023.625 208.565 2026.005 ;
        RECT 0.000 2022.785 208.285 2023.625 ;
        RECT 0.000 2020.405 208.565 2022.785 ;
        RECT 0.000 2019.565 208.285 2020.405 ;
        RECT 0.000 2017.645 208.565 2019.565 ;
        RECT 0.000 2016.805 208.285 2017.645 ;
        RECT 0.000 2014.425 208.565 2016.805 ;
        RECT 0.000 2013.585 208.285 2014.425 ;
        RECT 0.000 2011.205 208.565 2013.585 ;
        RECT 0.000 2010.365 208.285 2011.205 ;
        RECT 0.000 2008.445 208.565 2010.365 ;
        RECT 0.000 2007.605 208.285 2008.445 ;
        RECT 0.000 2005.225 208.565 2007.605 ;
        RECT 0.000 2004.385 208.285 2005.225 ;
        RECT 0.000 2002.005 208.565 2004.385 ;
        RECT 0.000 2001.165 208.285 2002.005 ;
        RECT 0.000 1999.245 208.565 2001.165 ;
        RECT 0.000 1998.405 208.285 1999.245 ;
        RECT 0.000 1996.025 208.565 1998.405 ;
        RECT 0.000 1995.185 208.285 1996.025 ;
        RECT 0.000 1992.805 208.565 1995.185 ;
        RECT 0.000 1991.965 208.285 1992.805 ;
        RECT 0.000 1990.045 208.565 1991.965 ;
        RECT 0.000 1989.205 208.285 1990.045 ;
      LAYER met2 ;
        RECT 208.565 1989.485 210.965 1989.765 ;
      LAYER met2 ;
        RECT 0.000 1988.210 208.565 1989.205 ;
        RECT 3379.435 1931.795 3588.000 1932.790 ;
      LAYER met2 ;
        RECT 3377.035 1931.235 3379.435 1931.515 ;
      LAYER met2 ;
        RECT 3379.715 1930.955 3588.000 1931.795 ;
        RECT 3379.435 1929.035 3588.000 1930.955 ;
        RECT 3379.715 1928.195 3588.000 1929.035 ;
        RECT 3379.435 1925.815 3588.000 1928.195 ;
        RECT 3379.715 1924.975 3588.000 1925.815 ;
        RECT 3379.435 1922.595 3588.000 1924.975 ;
        RECT 3379.715 1921.755 3588.000 1922.595 ;
        RECT 3379.435 1919.835 3588.000 1921.755 ;
        RECT 3379.715 1918.995 3588.000 1919.835 ;
        RECT 3379.435 1916.615 3588.000 1918.995 ;
        RECT 3379.715 1915.775 3588.000 1916.615 ;
        RECT 3379.435 1913.395 3588.000 1915.775 ;
        RECT 3379.715 1912.555 3588.000 1913.395 ;
        RECT 3379.435 1910.635 3588.000 1912.555 ;
        RECT 3379.715 1909.795 3588.000 1910.635 ;
        RECT 3379.435 1907.415 3588.000 1909.795 ;
        RECT 3379.715 1906.575 3588.000 1907.415 ;
        RECT 3379.435 1904.195 3588.000 1906.575 ;
        RECT 3379.715 1903.355 3588.000 1904.195 ;
        RECT 3379.435 1901.435 3588.000 1903.355 ;
        RECT 3379.715 1900.595 3588.000 1901.435 ;
        RECT 3379.435 1898.215 3588.000 1900.595 ;
        RECT 3379.715 1897.375 3588.000 1898.215 ;
        RECT 3379.435 1894.995 3588.000 1897.375 ;
      LAYER met2 ;
        RECT 3377.035 1894.645 3379.435 1894.715 ;
        RECT 3376.560 1894.505 3379.435 1894.645 ;
        RECT 3376.560 1854.625 3376.700 1894.505 ;
        RECT 3377.035 1894.435 3379.435 1894.505 ;
      LAYER met2 ;
        RECT 3379.715 1894.155 3588.000 1894.995 ;
        RECT 3379.435 1891.775 3588.000 1894.155 ;
        RECT 3379.715 1890.935 3588.000 1891.775 ;
        RECT 3379.435 1889.015 3588.000 1890.935 ;
        RECT 3379.715 1888.175 3588.000 1889.015 ;
        RECT 3379.435 1885.795 3588.000 1888.175 ;
        RECT 3379.715 1884.955 3588.000 1885.795 ;
        RECT 3379.435 1882.575 3588.000 1884.955 ;
        RECT 3379.715 1881.735 3588.000 1882.575 ;
        RECT 3379.435 1879.815 3588.000 1881.735 ;
      LAYER met2 ;
        RECT 3377.035 1879.255 3379.435 1879.535 ;
      LAYER met2 ;
        RECT 3379.715 1878.975 3588.000 1879.815 ;
        RECT 3379.435 1876.595 3588.000 1878.975 ;
        RECT 3379.715 1875.755 3588.000 1876.595 ;
        RECT 3379.435 1873.375 3588.000 1875.755 ;
      LAYER met2 ;
        RECT 3377.035 1872.815 3379.435 1873.095 ;
      LAYER met2 ;
        RECT 3379.715 1872.535 3588.000 1873.375 ;
        RECT 3379.435 1870.615 3588.000 1872.535 ;
      LAYER met2 ;
        RECT 3377.035 1870.055 3379.435 1870.335 ;
      LAYER met2 ;
        RECT 3379.715 1869.775 3588.000 1870.615 ;
        RECT 3379.435 1867.395 3588.000 1869.775 ;
        RECT 3379.715 1866.555 3588.000 1867.395 ;
        RECT 3379.435 1864.175 3588.000 1866.555 ;
        RECT 3379.715 1863.335 3588.000 1864.175 ;
        RECT 3379.435 1861.415 3588.000 1863.335 ;
      LAYER met2 ;
        RECT 3377.035 1860.855 3379.435 1861.135 ;
      LAYER met2 ;
        RECT 3379.715 1860.575 3588.000 1861.415 ;
        RECT 3379.435 1858.195 3588.000 1860.575 ;
        RECT 3379.715 1857.355 3588.000 1858.195 ;
        RECT 3379.435 1854.975 3588.000 1857.355 ;
      LAYER met2 ;
        RECT 3377.035 1854.625 3379.435 1854.695 ;
        RECT 3376.560 1854.485 3379.435 1854.625 ;
        RECT 3377.035 1854.415 3379.435 1854.485 ;
      LAYER met2 ;
        RECT 3379.715 1854.135 3588.000 1854.975 ;
        RECT 3379.435 1853.085 3588.000 1854.135 ;
        RECT 0.000 1850.865 208.565 1851.915 ;
        RECT 0.000 1850.025 208.285 1850.865 ;
      LAYER met2 ;
        RECT 208.565 1850.305 210.965 1850.585 ;
      LAYER met2 ;
        RECT 0.000 1847.645 208.565 1850.025 ;
      LAYER met2 ;
        RECT 209.000 1847.890 209.140 1850.305 ;
      LAYER met2 ;
        RECT 0.000 1846.805 208.285 1847.645 ;
      LAYER met2 ;
        RECT 208.940 1847.570 209.200 1847.890 ;
        RECT 211.700 1847.570 211.960 1847.890 ;
      LAYER met2 ;
        RECT 0.000 1844.425 208.565 1846.805 ;
        RECT 0.000 1843.585 208.285 1844.425 ;
      LAYER met2 ;
        RECT 208.565 1843.865 210.965 1844.145 ;
      LAYER met2 ;
        RECT 0.000 1841.665 208.565 1843.585 ;
        RECT 0.000 1840.825 208.285 1841.665 ;
        RECT 0.000 1838.445 208.565 1840.825 ;
        RECT 0.000 1837.605 208.285 1838.445 ;
        RECT 0.000 1835.225 208.565 1837.605 ;
        RECT 0.000 1834.385 208.285 1835.225 ;
        RECT 0.000 1832.465 208.565 1834.385 ;
        RECT 0.000 1831.625 208.285 1832.465 ;
      LAYER met2 ;
        RECT 208.565 1831.905 210.965 1832.185 ;
      LAYER met2 ;
        RECT 0.000 1829.245 208.565 1831.625 ;
        RECT 0.000 1828.405 208.285 1829.245 ;
        RECT 0.000 1826.025 208.565 1828.405 ;
        RECT 0.000 1825.185 208.285 1826.025 ;
      LAYER met2 ;
        RECT 208.565 1825.465 210.965 1825.745 ;
      LAYER met2 ;
        RECT 0.000 1823.265 208.565 1825.185 ;
        RECT 0.000 1822.425 208.285 1823.265 ;
        RECT 0.000 1820.045 208.565 1822.425 ;
        RECT 0.000 1819.205 208.285 1820.045 ;
        RECT 0.000 1816.825 208.565 1819.205 ;
        RECT 0.000 1815.985 208.285 1816.825 ;
        RECT 0.000 1814.065 208.565 1815.985 ;
        RECT 0.000 1813.225 208.285 1814.065 ;
        RECT 0.000 1810.845 208.565 1813.225 ;
      LAYER met2 ;
        RECT 211.760 1813.210 211.900 1847.570 ;
        RECT 208.940 1812.890 209.200 1813.210 ;
        RECT 211.700 1812.890 211.960 1813.210 ;
      LAYER met2 ;
        RECT 0.000 1810.005 208.285 1810.845 ;
      LAYER met2 ;
        RECT 209.000 1810.565 209.140 1812.890 ;
        RECT 208.565 1810.285 210.965 1810.565 ;
      LAYER met2 ;
        RECT 0.000 1807.625 208.565 1810.005 ;
        RECT 0.000 1806.785 208.285 1807.625 ;
        RECT 0.000 1804.405 208.565 1806.785 ;
        RECT 0.000 1803.565 208.285 1804.405 ;
        RECT 0.000 1801.645 208.565 1803.565 ;
        RECT 0.000 1800.805 208.285 1801.645 ;
        RECT 0.000 1798.425 208.565 1800.805 ;
        RECT 0.000 1797.585 208.285 1798.425 ;
        RECT 0.000 1795.205 208.565 1797.585 ;
        RECT 0.000 1794.365 208.285 1795.205 ;
        RECT 0.000 1792.445 208.565 1794.365 ;
        RECT 0.000 1791.605 208.285 1792.445 ;
        RECT 0.000 1789.225 208.565 1791.605 ;
        RECT 0.000 1788.385 208.285 1789.225 ;
        RECT 0.000 1786.005 208.565 1788.385 ;
        RECT 0.000 1785.165 208.285 1786.005 ;
        RECT 0.000 1783.245 208.565 1785.165 ;
        RECT 0.000 1782.405 208.285 1783.245 ;
        RECT 0.000 1780.025 208.565 1782.405 ;
        RECT 0.000 1779.185 208.285 1780.025 ;
        RECT 0.000 1776.805 208.565 1779.185 ;
        RECT 0.000 1775.965 208.285 1776.805 ;
        RECT 0.000 1774.045 208.565 1775.965 ;
        RECT 0.000 1773.205 208.285 1774.045 ;
      LAYER met2 ;
        RECT 208.565 1773.485 210.965 1773.765 ;
      LAYER met2 ;
        RECT 0.000 1772.210 208.565 1773.205 ;
        RECT 3379.435 1705.795 3588.000 1706.790 ;
      LAYER met2 ;
        RECT 3377.035 1705.235 3379.435 1705.515 ;
      LAYER met2 ;
        RECT 3379.715 1704.955 3588.000 1705.795 ;
        RECT 3379.435 1703.035 3588.000 1704.955 ;
        RECT 3379.715 1702.195 3588.000 1703.035 ;
        RECT 3379.435 1699.815 3588.000 1702.195 ;
        RECT 3379.715 1698.975 3588.000 1699.815 ;
        RECT 3379.435 1696.595 3588.000 1698.975 ;
        RECT 3379.715 1695.755 3588.000 1696.595 ;
        RECT 3379.435 1693.835 3588.000 1695.755 ;
        RECT 3379.715 1692.995 3588.000 1693.835 ;
        RECT 3379.435 1690.615 3588.000 1692.995 ;
        RECT 3379.715 1689.775 3588.000 1690.615 ;
        RECT 3379.435 1687.395 3588.000 1689.775 ;
        RECT 3379.715 1686.555 3588.000 1687.395 ;
        RECT 3379.435 1684.635 3588.000 1686.555 ;
        RECT 3379.715 1683.795 3588.000 1684.635 ;
        RECT 3379.435 1681.415 3588.000 1683.795 ;
        RECT 3379.715 1680.575 3588.000 1681.415 ;
        RECT 3379.435 1678.195 3588.000 1680.575 ;
        RECT 3379.715 1677.355 3588.000 1678.195 ;
        RECT 3379.435 1675.435 3588.000 1677.355 ;
        RECT 3379.715 1674.595 3588.000 1675.435 ;
        RECT 3379.435 1672.215 3588.000 1674.595 ;
        RECT 3379.715 1671.375 3588.000 1672.215 ;
        RECT 3379.435 1668.995 3588.000 1671.375 ;
      LAYER met2 ;
        RECT 3377.035 1668.645 3379.435 1668.715 ;
        RECT 3376.560 1668.505 3379.435 1668.645 ;
      LAYER met2 ;
        RECT 0.000 1634.865 208.565 1635.915 ;
        RECT 0.000 1634.025 208.285 1634.865 ;
      LAYER met2 ;
        RECT 208.565 1634.305 210.965 1634.585 ;
      LAYER met2 ;
        RECT 0.000 1631.645 208.565 1634.025 ;
      LAYER met2 ;
        RECT 209.000 1631.990 209.140 1634.305 ;
        RECT 208.940 1631.670 209.200 1631.990 ;
        RECT 211.700 1631.670 211.960 1631.990 ;
      LAYER met2 ;
        RECT 0.000 1630.805 208.285 1631.645 ;
        RECT 0.000 1628.425 208.565 1630.805 ;
        RECT 0.000 1627.585 208.285 1628.425 ;
      LAYER met2 ;
        RECT 208.565 1627.865 210.965 1628.145 ;
      LAYER met2 ;
        RECT 0.000 1625.665 208.565 1627.585 ;
        RECT 0.000 1624.825 208.285 1625.665 ;
        RECT 0.000 1622.445 208.565 1624.825 ;
        RECT 0.000 1621.605 208.285 1622.445 ;
        RECT 0.000 1619.225 208.565 1621.605 ;
        RECT 0.000 1618.385 208.285 1619.225 ;
        RECT 0.000 1616.465 208.565 1618.385 ;
        RECT 0.000 1615.625 208.285 1616.465 ;
      LAYER met2 ;
        RECT 208.565 1615.905 210.965 1616.185 ;
      LAYER met2 ;
        RECT 0.000 1613.245 208.565 1615.625 ;
        RECT 0.000 1612.405 208.285 1613.245 ;
        RECT 0.000 1610.025 208.565 1612.405 ;
        RECT 0.000 1609.185 208.285 1610.025 ;
      LAYER met2 ;
        RECT 208.565 1609.465 210.965 1609.745 ;
      LAYER met2 ;
        RECT 0.000 1607.265 208.565 1609.185 ;
        RECT 0.000 1606.425 208.285 1607.265 ;
        RECT 0.000 1604.045 208.565 1606.425 ;
        RECT 0.000 1603.205 208.285 1604.045 ;
        RECT 0.000 1600.825 208.565 1603.205 ;
        RECT 0.000 1599.985 208.285 1600.825 ;
        RECT 0.000 1598.065 208.565 1599.985 ;
        RECT 0.000 1597.225 208.285 1598.065 ;
      LAYER met2 ;
        RECT 211.760 1597.310 211.900 1631.670 ;
        RECT 3376.560 1628.625 3376.700 1668.505 ;
        RECT 3377.035 1668.435 3379.435 1668.505 ;
      LAYER met2 ;
        RECT 3379.715 1668.155 3588.000 1668.995 ;
        RECT 3379.435 1665.775 3588.000 1668.155 ;
        RECT 3379.715 1664.935 3588.000 1665.775 ;
        RECT 3379.435 1663.015 3588.000 1664.935 ;
        RECT 3379.715 1662.175 3588.000 1663.015 ;
        RECT 3379.435 1659.795 3588.000 1662.175 ;
        RECT 3379.715 1658.955 3588.000 1659.795 ;
        RECT 3379.435 1656.575 3588.000 1658.955 ;
        RECT 3379.715 1655.735 3588.000 1656.575 ;
        RECT 3379.435 1653.815 3588.000 1655.735 ;
      LAYER met2 ;
        RECT 3377.035 1653.255 3379.435 1653.535 ;
      LAYER met2 ;
        RECT 3379.715 1652.975 3588.000 1653.815 ;
        RECT 3379.435 1650.595 3588.000 1652.975 ;
        RECT 3379.715 1649.755 3588.000 1650.595 ;
        RECT 3379.435 1647.375 3588.000 1649.755 ;
      LAYER met2 ;
        RECT 3377.035 1646.815 3379.435 1647.095 ;
      LAYER met2 ;
        RECT 3379.715 1646.535 3588.000 1647.375 ;
        RECT 3379.435 1644.615 3588.000 1646.535 ;
      LAYER met2 ;
        RECT 3377.035 1644.055 3379.435 1644.335 ;
      LAYER met2 ;
        RECT 3379.715 1643.775 3588.000 1644.615 ;
        RECT 3379.435 1641.395 3588.000 1643.775 ;
        RECT 3379.715 1640.555 3588.000 1641.395 ;
        RECT 3379.435 1638.175 3588.000 1640.555 ;
        RECT 3379.715 1637.335 3588.000 1638.175 ;
        RECT 3379.435 1635.415 3588.000 1637.335 ;
      LAYER met2 ;
        RECT 3377.035 1634.855 3379.435 1635.135 ;
      LAYER met2 ;
        RECT 3379.715 1634.575 3588.000 1635.415 ;
        RECT 3379.435 1632.195 3588.000 1634.575 ;
        RECT 3379.715 1631.355 3588.000 1632.195 ;
        RECT 3379.435 1628.975 3588.000 1631.355 ;
      LAYER met2 ;
        RECT 3377.035 1628.625 3379.435 1628.695 ;
        RECT 3376.560 1628.485 3379.435 1628.625 ;
        RECT 3377.035 1628.415 3379.435 1628.485 ;
      LAYER met2 ;
        RECT 3379.715 1628.135 3588.000 1628.975 ;
        RECT 3379.435 1627.085 3588.000 1628.135 ;
        RECT 0.000 1594.845 208.565 1597.225 ;
      LAYER met2 ;
        RECT 208.940 1596.990 209.200 1597.310 ;
        RECT 211.700 1596.990 211.960 1597.310 ;
      LAYER met2 ;
        RECT 0.000 1594.005 208.285 1594.845 ;
      LAYER met2 ;
        RECT 209.000 1594.565 209.140 1596.990 ;
        RECT 208.565 1594.285 210.965 1594.565 ;
      LAYER met2 ;
        RECT 0.000 1591.625 208.565 1594.005 ;
        RECT 0.000 1590.785 208.285 1591.625 ;
        RECT 0.000 1588.405 208.565 1590.785 ;
        RECT 0.000 1587.565 208.285 1588.405 ;
        RECT 0.000 1585.645 208.565 1587.565 ;
        RECT 0.000 1584.805 208.285 1585.645 ;
        RECT 0.000 1582.425 208.565 1584.805 ;
        RECT 0.000 1581.585 208.285 1582.425 ;
        RECT 0.000 1579.205 208.565 1581.585 ;
        RECT 0.000 1578.365 208.285 1579.205 ;
        RECT 0.000 1576.445 208.565 1578.365 ;
        RECT 0.000 1575.605 208.285 1576.445 ;
        RECT 0.000 1573.225 208.565 1575.605 ;
        RECT 0.000 1572.385 208.285 1573.225 ;
        RECT 0.000 1570.005 208.565 1572.385 ;
        RECT 0.000 1569.165 208.285 1570.005 ;
        RECT 0.000 1567.245 208.565 1569.165 ;
        RECT 0.000 1566.405 208.285 1567.245 ;
        RECT 0.000 1564.025 208.565 1566.405 ;
        RECT 0.000 1563.185 208.285 1564.025 ;
        RECT 0.000 1560.805 208.565 1563.185 ;
        RECT 0.000 1559.965 208.285 1560.805 ;
        RECT 0.000 1558.045 208.565 1559.965 ;
        RECT 0.000 1557.205 208.285 1558.045 ;
      LAYER met2 ;
        RECT 208.565 1557.485 210.965 1557.765 ;
      LAYER met2 ;
        RECT 0.000 1556.210 208.565 1557.205 ;
        RECT 3379.435 1480.795 3588.000 1481.790 ;
      LAYER met2 ;
        RECT 3377.035 1480.235 3379.435 1480.515 ;
      LAYER met2 ;
        RECT 3379.715 1479.955 3588.000 1480.795 ;
        RECT 3379.435 1478.035 3588.000 1479.955 ;
        RECT 3379.715 1477.195 3588.000 1478.035 ;
        RECT 3379.435 1474.815 3588.000 1477.195 ;
        RECT 3379.715 1473.975 3588.000 1474.815 ;
        RECT 3379.435 1471.595 3588.000 1473.975 ;
        RECT 3379.715 1470.755 3588.000 1471.595 ;
        RECT 3379.435 1468.835 3588.000 1470.755 ;
        RECT 3379.715 1467.995 3588.000 1468.835 ;
        RECT 3379.435 1465.615 3588.000 1467.995 ;
        RECT 3379.715 1464.775 3588.000 1465.615 ;
        RECT 3379.435 1462.395 3588.000 1464.775 ;
        RECT 3379.715 1461.555 3588.000 1462.395 ;
        RECT 3379.435 1459.635 3588.000 1461.555 ;
        RECT 3379.715 1458.795 3588.000 1459.635 ;
        RECT 3379.435 1456.415 3588.000 1458.795 ;
        RECT 3379.715 1455.575 3588.000 1456.415 ;
        RECT 3379.435 1453.195 3588.000 1455.575 ;
        RECT 3379.715 1452.355 3588.000 1453.195 ;
        RECT 3379.435 1450.435 3588.000 1452.355 ;
        RECT 3379.715 1449.595 3588.000 1450.435 ;
        RECT 3379.435 1447.215 3588.000 1449.595 ;
        RECT 3379.715 1446.375 3588.000 1447.215 ;
        RECT 3379.435 1443.995 3588.000 1446.375 ;
      LAYER met2 ;
        RECT 3377.035 1443.645 3379.435 1443.715 ;
        RECT 3376.560 1443.505 3379.435 1443.645 ;
      LAYER met2 ;
        RECT 0.000 1418.865 208.565 1419.915 ;
        RECT 0.000 1418.025 208.285 1418.865 ;
      LAYER met2 ;
        RECT 208.565 1418.305 210.965 1418.585 ;
      LAYER met2 ;
        RECT 0.000 1415.645 208.565 1418.025 ;
      LAYER met2 ;
        RECT 209.000 1416.090 209.140 1418.305 ;
        RECT 208.940 1415.770 209.200 1416.090 ;
        RECT 211.700 1415.770 211.960 1416.090 ;
      LAYER met2 ;
        RECT 0.000 1414.805 208.285 1415.645 ;
        RECT 0.000 1412.425 208.565 1414.805 ;
        RECT 0.000 1411.585 208.285 1412.425 ;
      LAYER met2 ;
        RECT 208.565 1411.865 210.965 1412.145 ;
      LAYER met2 ;
        RECT 0.000 1409.665 208.565 1411.585 ;
        RECT 0.000 1408.825 208.285 1409.665 ;
        RECT 0.000 1406.445 208.565 1408.825 ;
        RECT 0.000 1405.605 208.285 1406.445 ;
        RECT 0.000 1403.225 208.565 1405.605 ;
        RECT 0.000 1402.385 208.285 1403.225 ;
        RECT 0.000 1400.465 208.565 1402.385 ;
        RECT 0.000 1399.625 208.285 1400.465 ;
      LAYER met2 ;
        RECT 208.565 1399.905 210.965 1400.185 ;
      LAYER met2 ;
        RECT 0.000 1397.245 208.565 1399.625 ;
        RECT 0.000 1396.405 208.285 1397.245 ;
        RECT 0.000 1394.025 208.565 1396.405 ;
        RECT 0.000 1393.185 208.285 1394.025 ;
      LAYER met2 ;
        RECT 208.565 1393.465 210.965 1393.745 ;
      LAYER met2 ;
        RECT 0.000 1391.265 208.565 1393.185 ;
        RECT 0.000 1390.425 208.285 1391.265 ;
        RECT 0.000 1388.045 208.565 1390.425 ;
        RECT 0.000 1387.205 208.285 1388.045 ;
        RECT 0.000 1384.825 208.565 1387.205 ;
        RECT 0.000 1383.985 208.285 1384.825 ;
        RECT 0.000 1382.065 208.565 1383.985 ;
        RECT 0.000 1381.225 208.285 1382.065 ;
        RECT 0.000 1378.845 208.565 1381.225 ;
      LAYER met2 ;
        RECT 211.760 1381.070 211.900 1415.770 ;
        RECT 3376.560 1403.625 3376.700 1443.505 ;
        RECT 3377.035 1443.435 3379.435 1443.505 ;
      LAYER met2 ;
        RECT 3379.715 1443.155 3588.000 1443.995 ;
        RECT 3379.435 1440.775 3588.000 1443.155 ;
        RECT 3379.715 1439.935 3588.000 1440.775 ;
        RECT 3379.435 1438.015 3588.000 1439.935 ;
        RECT 3379.715 1437.175 3588.000 1438.015 ;
        RECT 3379.435 1434.795 3588.000 1437.175 ;
        RECT 3379.715 1433.955 3588.000 1434.795 ;
        RECT 3379.435 1431.575 3588.000 1433.955 ;
        RECT 3379.715 1430.735 3588.000 1431.575 ;
        RECT 3379.435 1428.815 3588.000 1430.735 ;
      LAYER met2 ;
        RECT 3377.035 1428.255 3379.435 1428.535 ;
      LAYER met2 ;
        RECT 3379.715 1427.975 3588.000 1428.815 ;
        RECT 3379.435 1425.595 3588.000 1427.975 ;
        RECT 3379.715 1424.755 3588.000 1425.595 ;
        RECT 3379.435 1422.375 3588.000 1424.755 ;
      LAYER met2 ;
        RECT 3377.035 1421.815 3379.435 1422.095 ;
      LAYER met2 ;
        RECT 3379.715 1421.535 3588.000 1422.375 ;
        RECT 3379.435 1419.615 3588.000 1421.535 ;
      LAYER met2 ;
        RECT 3377.035 1419.055 3379.435 1419.335 ;
      LAYER met2 ;
        RECT 3379.715 1418.775 3588.000 1419.615 ;
        RECT 3379.435 1416.395 3588.000 1418.775 ;
        RECT 3379.715 1415.555 3588.000 1416.395 ;
        RECT 3379.435 1413.175 3588.000 1415.555 ;
        RECT 3379.715 1412.335 3588.000 1413.175 ;
        RECT 3379.435 1410.415 3588.000 1412.335 ;
      LAYER met2 ;
        RECT 3377.035 1409.855 3379.435 1410.135 ;
      LAYER met2 ;
        RECT 3379.715 1409.575 3588.000 1410.415 ;
        RECT 3379.435 1407.195 3588.000 1409.575 ;
        RECT 3379.715 1406.355 3588.000 1407.195 ;
        RECT 3379.435 1403.975 3588.000 1406.355 ;
      LAYER met2 ;
        RECT 3377.035 1403.625 3379.435 1403.695 ;
        RECT 3376.560 1403.485 3379.435 1403.625 ;
        RECT 3377.035 1403.415 3379.435 1403.485 ;
      LAYER met2 ;
        RECT 3379.715 1403.135 3588.000 1403.975 ;
        RECT 3379.435 1402.085 3588.000 1403.135 ;
      LAYER met2 ;
        RECT 208.940 1380.750 209.200 1381.070 ;
        RECT 211.700 1380.750 211.960 1381.070 ;
      LAYER met2 ;
        RECT 0.000 1378.005 208.285 1378.845 ;
      LAYER met2 ;
        RECT 209.000 1378.565 209.140 1380.750 ;
        RECT 208.565 1378.285 210.965 1378.565 ;
      LAYER met2 ;
        RECT 0.000 1375.625 208.565 1378.005 ;
        RECT 0.000 1374.785 208.285 1375.625 ;
        RECT 0.000 1372.405 208.565 1374.785 ;
        RECT 0.000 1371.565 208.285 1372.405 ;
        RECT 0.000 1369.645 208.565 1371.565 ;
        RECT 0.000 1368.805 208.285 1369.645 ;
        RECT 0.000 1366.425 208.565 1368.805 ;
        RECT 0.000 1365.585 208.285 1366.425 ;
        RECT 0.000 1363.205 208.565 1365.585 ;
        RECT 0.000 1362.365 208.285 1363.205 ;
        RECT 0.000 1360.445 208.565 1362.365 ;
        RECT 0.000 1359.605 208.285 1360.445 ;
        RECT 0.000 1357.225 208.565 1359.605 ;
        RECT 0.000 1356.385 208.285 1357.225 ;
        RECT 0.000 1354.005 208.565 1356.385 ;
        RECT 0.000 1353.165 208.285 1354.005 ;
        RECT 0.000 1351.245 208.565 1353.165 ;
        RECT 0.000 1350.405 208.285 1351.245 ;
        RECT 0.000 1348.025 208.565 1350.405 ;
        RECT 0.000 1347.185 208.285 1348.025 ;
        RECT 0.000 1344.805 208.565 1347.185 ;
        RECT 0.000 1343.965 208.285 1344.805 ;
        RECT 0.000 1342.045 208.565 1343.965 ;
        RECT 0.000 1341.205 208.285 1342.045 ;
      LAYER met2 ;
        RECT 208.565 1341.485 210.965 1341.765 ;
      LAYER met2 ;
        RECT 0.000 1340.210 208.565 1341.205 ;
        RECT 3379.435 1255.795 3588.000 1256.790 ;
      LAYER met2 ;
        RECT 3377.035 1255.235 3379.435 1255.515 ;
      LAYER met2 ;
        RECT 3379.715 1254.955 3588.000 1255.795 ;
        RECT 3379.435 1253.035 3588.000 1254.955 ;
        RECT 3379.715 1252.195 3588.000 1253.035 ;
        RECT 3379.435 1249.815 3588.000 1252.195 ;
        RECT 3379.715 1248.975 3588.000 1249.815 ;
        RECT 3379.435 1246.595 3588.000 1248.975 ;
        RECT 3379.715 1245.755 3588.000 1246.595 ;
        RECT 3379.435 1243.835 3588.000 1245.755 ;
        RECT 3379.715 1242.995 3588.000 1243.835 ;
        RECT 3379.435 1240.615 3588.000 1242.995 ;
        RECT 3379.715 1239.775 3588.000 1240.615 ;
        RECT 3379.435 1237.395 3588.000 1239.775 ;
        RECT 3379.715 1236.555 3588.000 1237.395 ;
        RECT 3379.435 1234.635 3588.000 1236.555 ;
        RECT 3379.715 1233.795 3588.000 1234.635 ;
        RECT 3379.435 1231.415 3588.000 1233.795 ;
        RECT 3379.715 1230.575 3588.000 1231.415 ;
        RECT 3379.435 1228.195 3588.000 1230.575 ;
        RECT 3379.715 1227.355 3588.000 1228.195 ;
        RECT 3379.435 1225.435 3588.000 1227.355 ;
        RECT 3379.715 1224.595 3588.000 1225.435 ;
        RECT 3379.435 1222.215 3588.000 1224.595 ;
        RECT 3379.715 1221.375 3588.000 1222.215 ;
        RECT 3379.435 1218.995 3588.000 1221.375 ;
      LAYER met2 ;
        RECT 3377.035 1218.645 3379.435 1218.715 ;
        RECT 3376.560 1218.505 3379.435 1218.645 ;
      LAYER met2 ;
        RECT 0.000 1202.865 208.565 1203.915 ;
        RECT 0.000 1202.025 208.285 1202.865 ;
      LAYER met2 ;
        RECT 208.610 1202.585 209.140 1202.650 ;
        RECT 208.565 1202.305 210.965 1202.585 ;
      LAYER met2 ;
        RECT 0.000 1199.645 208.565 1202.025 ;
      LAYER met2 ;
        RECT 209.000 1199.850 209.140 1202.305 ;
      LAYER met2 ;
        RECT 0.000 1198.805 208.285 1199.645 ;
      LAYER met2 ;
        RECT 208.940 1199.530 209.200 1199.850 ;
        RECT 211.700 1199.530 211.960 1199.850 ;
      LAYER met2 ;
        RECT 0.000 1196.425 208.565 1198.805 ;
        RECT 0.000 1195.585 208.285 1196.425 ;
      LAYER met2 ;
        RECT 208.565 1195.865 210.965 1196.145 ;
      LAYER met2 ;
        RECT 0.000 1193.665 208.565 1195.585 ;
        RECT 0.000 1192.825 208.285 1193.665 ;
        RECT 0.000 1190.445 208.565 1192.825 ;
        RECT 0.000 1189.605 208.285 1190.445 ;
        RECT 0.000 1187.225 208.565 1189.605 ;
        RECT 0.000 1186.385 208.285 1187.225 ;
        RECT 0.000 1184.465 208.565 1186.385 ;
        RECT 0.000 1183.625 208.285 1184.465 ;
      LAYER met2 ;
        RECT 208.565 1183.905 210.965 1184.185 ;
      LAYER met2 ;
        RECT 0.000 1181.245 208.565 1183.625 ;
        RECT 0.000 1180.405 208.285 1181.245 ;
        RECT 0.000 1178.025 208.565 1180.405 ;
        RECT 0.000 1177.185 208.285 1178.025 ;
      LAYER met2 ;
        RECT 208.565 1177.465 210.965 1177.745 ;
      LAYER met2 ;
        RECT 0.000 1175.265 208.565 1177.185 ;
        RECT 0.000 1174.425 208.285 1175.265 ;
        RECT 0.000 1172.045 208.565 1174.425 ;
        RECT 0.000 1171.205 208.285 1172.045 ;
        RECT 0.000 1168.825 208.565 1171.205 ;
        RECT 0.000 1167.985 208.285 1168.825 ;
        RECT 0.000 1166.065 208.565 1167.985 ;
        RECT 0.000 1165.225 208.285 1166.065 ;
        RECT 0.000 1162.845 208.565 1165.225 ;
      LAYER met2 ;
        RECT 211.760 1165.170 211.900 1199.530 ;
        RECT 3376.560 1178.625 3376.700 1218.505 ;
        RECT 3377.035 1218.435 3379.435 1218.505 ;
      LAYER met2 ;
        RECT 3379.715 1218.155 3588.000 1218.995 ;
        RECT 3379.435 1215.775 3588.000 1218.155 ;
        RECT 3379.715 1214.935 3588.000 1215.775 ;
        RECT 3379.435 1213.015 3588.000 1214.935 ;
        RECT 3379.715 1212.175 3588.000 1213.015 ;
        RECT 3379.435 1209.795 3588.000 1212.175 ;
        RECT 3379.715 1208.955 3588.000 1209.795 ;
        RECT 3379.435 1206.575 3588.000 1208.955 ;
        RECT 3379.715 1205.735 3588.000 1206.575 ;
        RECT 3379.435 1203.815 3588.000 1205.735 ;
      LAYER met2 ;
        RECT 3377.035 1203.255 3379.435 1203.535 ;
      LAYER met2 ;
        RECT 3379.715 1202.975 3588.000 1203.815 ;
        RECT 3379.435 1200.595 3588.000 1202.975 ;
        RECT 3379.715 1199.755 3588.000 1200.595 ;
        RECT 3379.435 1197.375 3588.000 1199.755 ;
      LAYER met2 ;
        RECT 3377.035 1196.815 3379.435 1197.095 ;
      LAYER met2 ;
        RECT 3379.715 1196.535 3588.000 1197.375 ;
        RECT 3379.435 1194.615 3588.000 1196.535 ;
      LAYER met2 ;
        RECT 3377.035 1194.055 3379.435 1194.335 ;
      LAYER met2 ;
        RECT 3379.715 1193.775 3588.000 1194.615 ;
        RECT 3379.435 1191.395 3588.000 1193.775 ;
        RECT 3379.715 1190.555 3588.000 1191.395 ;
        RECT 3379.435 1188.175 3588.000 1190.555 ;
        RECT 3379.715 1187.335 3588.000 1188.175 ;
        RECT 3379.435 1185.415 3588.000 1187.335 ;
      LAYER met2 ;
        RECT 3377.035 1184.855 3379.435 1185.135 ;
      LAYER met2 ;
        RECT 3379.715 1184.575 3588.000 1185.415 ;
        RECT 3379.435 1182.195 3588.000 1184.575 ;
        RECT 3379.715 1181.355 3588.000 1182.195 ;
        RECT 3379.435 1178.975 3588.000 1181.355 ;
      LAYER met2 ;
        RECT 3377.035 1178.625 3379.435 1178.695 ;
        RECT 3376.560 1178.485 3379.435 1178.625 ;
        RECT 3377.035 1178.415 3379.435 1178.485 ;
      LAYER met2 ;
        RECT 3379.715 1178.135 3588.000 1178.975 ;
        RECT 3379.435 1177.085 3588.000 1178.135 ;
      LAYER met2 ;
        RECT 208.940 1164.850 209.200 1165.170 ;
        RECT 211.700 1164.850 211.960 1165.170 ;
      LAYER met2 ;
        RECT 0.000 1162.005 208.285 1162.845 ;
      LAYER met2 ;
        RECT 209.000 1162.565 209.140 1164.850 ;
        RECT 208.565 1162.285 210.965 1162.565 ;
      LAYER met2 ;
        RECT 0.000 1159.625 208.565 1162.005 ;
        RECT 0.000 1158.785 208.285 1159.625 ;
        RECT 0.000 1156.405 208.565 1158.785 ;
        RECT 0.000 1155.565 208.285 1156.405 ;
        RECT 0.000 1153.645 208.565 1155.565 ;
        RECT 0.000 1152.805 208.285 1153.645 ;
        RECT 0.000 1150.425 208.565 1152.805 ;
        RECT 0.000 1149.585 208.285 1150.425 ;
        RECT 0.000 1147.205 208.565 1149.585 ;
        RECT 0.000 1146.365 208.285 1147.205 ;
        RECT 0.000 1144.445 208.565 1146.365 ;
        RECT 0.000 1143.605 208.285 1144.445 ;
        RECT 0.000 1141.225 208.565 1143.605 ;
        RECT 0.000 1140.385 208.285 1141.225 ;
        RECT 0.000 1138.005 208.565 1140.385 ;
        RECT 0.000 1137.165 208.285 1138.005 ;
        RECT 0.000 1135.245 208.565 1137.165 ;
        RECT 0.000 1134.405 208.285 1135.245 ;
        RECT 0.000 1132.025 208.565 1134.405 ;
        RECT 0.000 1131.185 208.285 1132.025 ;
        RECT 0.000 1128.805 208.565 1131.185 ;
        RECT 0.000 1127.965 208.285 1128.805 ;
        RECT 0.000 1126.045 208.565 1127.965 ;
        RECT 0.000 1125.205 208.285 1126.045 ;
      LAYER met2 ;
        RECT 208.565 1125.485 210.965 1125.765 ;
      LAYER met2 ;
        RECT 0.000 1124.210 208.565 1125.205 ;
        RECT 3379.435 1029.795 3588.000 1030.790 ;
      LAYER met2 ;
        RECT 3377.035 1029.235 3379.435 1029.515 ;
      LAYER met2 ;
        RECT 3379.715 1028.955 3588.000 1029.795 ;
        RECT 3379.435 1027.035 3588.000 1028.955 ;
        RECT 3379.715 1026.195 3588.000 1027.035 ;
        RECT 3379.435 1023.815 3588.000 1026.195 ;
        RECT 3379.715 1022.975 3588.000 1023.815 ;
        RECT 3379.435 1020.595 3588.000 1022.975 ;
        RECT 3379.715 1019.755 3588.000 1020.595 ;
        RECT 3379.435 1017.835 3588.000 1019.755 ;
        RECT 3379.715 1016.995 3588.000 1017.835 ;
        RECT 3379.435 1014.615 3588.000 1016.995 ;
        RECT 3379.715 1013.775 3588.000 1014.615 ;
        RECT 3379.435 1011.395 3588.000 1013.775 ;
        RECT 3379.715 1010.555 3588.000 1011.395 ;
        RECT 3379.435 1008.635 3588.000 1010.555 ;
        RECT 3379.715 1007.795 3588.000 1008.635 ;
        RECT 3379.435 1005.415 3588.000 1007.795 ;
        RECT 3379.715 1004.575 3588.000 1005.415 ;
        RECT 3379.435 1002.195 3588.000 1004.575 ;
        RECT 3379.715 1001.355 3588.000 1002.195 ;
        RECT 3379.435 999.435 3588.000 1001.355 ;
        RECT 3379.715 998.595 3588.000 999.435 ;
        RECT 3379.435 996.215 3588.000 998.595 ;
        RECT 3379.715 995.375 3588.000 996.215 ;
      LAYER met2 ;
        RECT 3376.560 993.070 3377.160 993.210 ;
      LAYER met2 ;
        RECT 0.000 986.865 208.565 987.915 ;
        RECT 0.000 986.025 208.285 986.865 ;
      LAYER met2 ;
        RECT 208.565 986.305 210.965 986.585 ;
      LAYER met2 ;
        RECT 0.000 983.645 208.565 986.025 ;
      LAYER met2 ;
        RECT 209.000 983.950 209.140 986.305 ;
      LAYER met2 ;
        RECT 0.000 982.805 208.285 983.645 ;
      LAYER met2 ;
        RECT 208.940 983.630 209.200 983.950 ;
        RECT 211.700 983.630 211.960 983.950 ;
      LAYER met2 ;
        RECT 0.000 980.425 208.565 982.805 ;
        RECT 0.000 979.585 208.285 980.425 ;
      LAYER met2 ;
        RECT 208.565 979.865 210.965 980.145 ;
      LAYER met2 ;
        RECT 0.000 977.665 208.565 979.585 ;
        RECT 0.000 976.825 208.285 977.665 ;
        RECT 0.000 974.445 208.565 976.825 ;
        RECT 0.000 973.605 208.285 974.445 ;
        RECT 0.000 971.225 208.565 973.605 ;
        RECT 0.000 970.385 208.285 971.225 ;
        RECT 0.000 968.465 208.565 970.385 ;
        RECT 0.000 967.625 208.285 968.465 ;
      LAYER met2 ;
        RECT 208.565 967.905 210.965 968.185 ;
      LAYER met2 ;
        RECT 0.000 965.245 208.565 967.625 ;
        RECT 0.000 964.405 208.285 965.245 ;
        RECT 0.000 962.025 208.565 964.405 ;
        RECT 0.000 961.185 208.285 962.025 ;
      LAYER met2 ;
        RECT 208.565 961.465 210.965 961.745 ;
      LAYER met2 ;
        RECT 0.000 959.265 208.565 961.185 ;
        RECT 0.000 958.425 208.285 959.265 ;
        RECT 0.000 956.045 208.565 958.425 ;
        RECT 0.000 955.205 208.285 956.045 ;
        RECT 0.000 952.825 208.565 955.205 ;
        RECT 0.000 951.985 208.285 952.825 ;
        RECT 0.000 950.065 208.565 951.985 ;
        RECT 0.000 949.225 208.285 950.065 ;
      LAYER met2 ;
        RECT 211.760 949.270 211.900 983.630 ;
        RECT 3376.560 952.625 3376.700 993.070 ;
        RECT 3377.020 992.715 3377.160 993.070 ;
      LAYER met2 ;
        RECT 3379.435 992.995 3588.000 995.375 ;
      LAYER met2 ;
        RECT 3377.020 992.460 3379.435 992.715 ;
        RECT 3377.035 992.435 3379.435 992.460 ;
      LAYER met2 ;
        RECT 3379.715 992.155 3588.000 992.995 ;
        RECT 3379.435 989.775 3588.000 992.155 ;
        RECT 3379.715 988.935 3588.000 989.775 ;
        RECT 3379.435 987.015 3588.000 988.935 ;
        RECT 3379.715 986.175 3588.000 987.015 ;
        RECT 3379.435 983.795 3588.000 986.175 ;
        RECT 3379.715 982.955 3588.000 983.795 ;
        RECT 3379.435 980.575 3588.000 982.955 ;
        RECT 3379.715 979.735 3588.000 980.575 ;
        RECT 3379.435 977.815 3588.000 979.735 ;
      LAYER met2 ;
        RECT 3377.035 977.255 3379.435 977.535 ;
      LAYER met2 ;
        RECT 3379.715 976.975 3588.000 977.815 ;
        RECT 3379.435 974.595 3588.000 976.975 ;
        RECT 3379.715 973.755 3588.000 974.595 ;
        RECT 3379.435 971.375 3588.000 973.755 ;
      LAYER met2 ;
        RECT 3377.035 970.815 3379.435 971.095 ;
      LAYER met2 ;
        RECT 3379.715 970.535 3588.000 971.375 ;
        RECT 3379.435 968.615 3588.000 970.535 ;
      LAYER met2 ;
        RECT 3377.035 968.055 3379.435 968.335 ;
      LAYER met2 ;
        RECT 3379.715 967.775 3588.000 968.615 ;
        RECT 3379.435 965.395 3588.000 967.775 ;
        RECT 3379.715 964.555 3588.000 965.395 ;
        RECT 3379.435 962.175 3588.000 964.555 ;
        RECT 3379.715 961.335 3588.000 962.175 ;
        RECT 3379.435 959.415 3588.000 961.335 ;
      LAYER met2 ;
        RECT 3377.035 958.855 3379.435 959.135 ;
      LAYER met2 ;
        RECT 3379.715 958.575 3588.000 959.415 ;
        RECT 3379.435 956.195 3588.000 958.575 ;
        RECT 3379.715 955.355 3588.000 956.195 ;
        RECT 3379.435 952.975 3588.000 955.355 ;
      LAYER met2 ;
        RECT 3377.035 952.625 3379.435 952.695 ;
        RECT 3376.560 952.485 3379.435 952.625 ;
        RECT 3377.035 952.415 3379.435 952.485 ;
      LAYER met2 ;
        RECT 3379.715 952.135 3588.000 952.975 ;
        RECT 3379.435 951.085 3588.000 952.135 ;
        RECT 0.000 946.845 208.565 949.225 ;
      LAYER met2 ;
        RECT 208.940 948.950 209.200 949.270 ;
        RECT 211.700 948.950 211.960 949.270 ;
      LAYER met2 ;
        RECT 0.000 946.005 208.285 946.845 ;
      LAYER met2 ;
        RECT 209.000 946.565 209.140 948.950 ;
        RECT 208.565 946.285 210.965 946.565 ;
      LAYER met2 ;
        RECT 0.000 943.625 208.565 946.005 ;
        RECT 0.000 942.785 208.285 943.625 ;
        RECT 0.000 940.405 208.565 942.785 ;
        RECT 0.000 939.565 208.285 940.405 ;
        RECT 0.000 937.645 208.565 939.565 ;
        RECT 0.000 936.805 208.285 937.645 ;
        RECT 0.000 934.425 208.565 936.805 ;
        RECT 0.000 933.585 208.285 934.425 ;
        RECT 0.000 931.205 208.565 933.585 ;
        RECT 0.000 930.365 208.285 931.205 ;
        RECT 0.000 928.445 208.565 930.365 ;
        RECT 0.000 927.605 208.285 928.445 ;
        RECT 0.000 925.225 208.565 927.605 ;
        RECT 0.000 924.385 208.285 925.225 ;
        RECT 0.000 922.005 208.565 924.385 ;
        RECT 0.000 921.165 208.285 922.005 ;
        RECT 0.000 919.245 208.565 921.165 ;
        RECT 0.000 918.405 208.285 919.245 ;
        RECT 0.000 916.025 208.565 918.405 ;
        RECT 0.000 915.185 208.285 916.025 ;
        RECT 0.000 912.805 208.565 915.185 ;
        RECT 0.000 911.965 208.285 912.805 ;
        RECT 0.000 910.045 208.565 911.965 ;
        RECT 0.000 909.205 208.285 910.045 ;
      LAYER met2 ;
        RECT 208.565 909.485 210.965 909.765 ;
      LAYER met2 ;
        RECT 0.000 908.210 208.565 909.205 ;
        RECT 3379.435 804.795 3588.000 805.790 ;
      LAYER met2 ;
        RECT 3377.035 804.235 3379.435 804.515 ;
      LAYER met2 ;
        RECT 3379.715 803.955 3588.000 804.795 ;
        RECT 3379.435 802.035 3588.000 803.955 ;
        RECT 3379.715 801.195 3588.000 802.035 ;
        RECT 3379.435 798.815 3588.000 801.195 ;
        RECT 3379.715 797.975 3588.000 798.815 ;
        RECT 3379.435 795.595 3588.000 797.975 ;
        RECT 3379.715 794.755 3588.000 795.595 ;
        RECT 3379.435 792.835 3588.000 794.755 ;
        RECT 3379.715 791.995 3588.000 792.835 ;
        RECT 3379.435 789.615 3588.000 791.995 ;
        RECT 3379.715 788.775 3588.000 789.615 ;
        RECT 3379.435 786.395 3588.000 788.775 ;
        RECT 3379.715 785.555 3588.000 786.395 ;
        RECT 3379.435 783.635 3588.000 785.555 ;
        RECT 3379.715 782.795 3588.000 783.635 ;
        RECT 3379.435 780.415 3588.000 782.795 ;
        RECT 3379.715 779.575 3588.000 780.415 ;
        RECT 3379.435 777.195 3588.000 779.575 ;
        RECT 3379.715 776.355 3588.000 777.195 ;
        RECT 3379.435 774.435 3588.000 776.355 ;
        RECT 3379.715 773.595 3588.000 774.435 ;
        RECT 3379.435 771.215 3588.000 773.595 ;
        RECT 3379.715 770.375 3588.000 771.215 ;
        RECT 3379.435 767.995 3588.000 770.375 ;
      LAYER met2 ;
        RECT 3377.035 767.645 3379.435 767.715 ;
        RECT 3376.560 767.505 3379.435 767.645 ;
        RECT 3376.560 727.625 3376.700 767.505 ;
        RECT 3377.035 767.435 3379.435 767.505 ;
      LAYER met2 ;
        RECT 3379.715 767.155 3588.000 767.995 ;
        RECT 3379.435 764.775 3588.000 767.155 ;
        RECT 3379.715 763.935 3588.000 764.775 ;
        RECT 3379.435 762.015 3588.000 763.935 ;
        RECT 3379.715 761.175 3588.000 762.015 ;
        RECT 3379.435 758.795 3588.000 761.175 ;
        RECT 3379.715 757.955 3588.000 758.795 ;
        RECT 3379.435 755.575 3588.000 757.955 ;
        RECT 3379.715 754.735 3588.000 755.575 ;
        RECT 3379.435 752.815 3588.000 754.735 ;
      LAYER met2 ;
        RECT 3377.035 752.255 3379.435 752.535 ;
      LAYER met2 ;
        RECT 3379.715 751.975 3588.000 752.815 ;
        RECT 3379.435 749.595 3588.000 751.975 ;
        RECT 3379.715 748.755 3588.000 749.595 ;
        RECT 3379.435 746.375 3588.000 748.755 ;
      LAYER met2 ;
        RECT 3377.035 745.815 3379.435 746.095 ;
      LAYER met2 ;
        RECT 3379.715 745.535 3588.000 746.375 ;
        RECT 3379.435 743.615 3588.000 745.535 ;
      LAYER met2 ;
        RECT 3377.035 743.055 3379.435 743.335 ;
      LAYER met2 ;
        RECT 3379.715 742.775 3588.000 743.615 ;
        RECT 3379.435 740.395 3588.000 742.775 ;
        RECT 3379.715 739.555 3588.000 740.395 ;
        RECT 3379.435 737.175 3588.000 739.555 ;
        RECT 3379.715 736.335 3588.000 737.175 ;
        RECT 3379.435 734.415 3588.000 736.335 ;
      LAYER met2 ;
        RECT 3377.035 733.855 3379.435 734.135 ;
      LAYER met2 ;
        RECT 3379.715 733.575 3588.000 734.415 ;
        RECT 3379.435 731.195 3588.000 733.575 ;
        RECT 3379.715 730.355 3588.000 731.195 ;
        RECT 3379.435 727.975 3588.000 730.355 ;
      LAYER met2 ;
        RECT 3377.035 727.625 3379.435 727.695 ;
        RECT 3376.560 727.485 3379.435 727.625 ;
        RECT 3377.035 727.415 3379.435 727.485 ;
      LAYER met2 ;
        RECT 3379.715 727.135 3588.000 727.975 ;
        RECT 3379.435 726.085 3588.000 727.135 ;
        RECT 4.925 601.390 200.000 625.290 ;
        RECT 4.925 575.395 197.965 601.390 ;
        RECT 198.080 576.895 200.000 578.895 ;
        RECT 3379.435 578.795 3588.000 579.790 ;
      LAYER met2 ;
        RECT 3377.035 578.235 3379.435 578.515 ;
      LAYER met2 ;
        RECT 3379.715 577.955 3588.000 578.795 ;
        RECT 3379.435 576.035 3588.000 577.955 ;
        RECT 4.925 551.495 200.000 575.395 ;
        RECT 3379.715 575.195 3588.000 576.035 ;
        RECT 3379.435 572.815 3588.000 575.195 ;
        RECT 3379.715 571.975 3588.000 572.815 ;
        RECT 3379.435 569.595 3588.000 571.975 ;
        RECT 3379.715 568.755 3588.000 569.595 ;
        RECT 3379.435 566.835 3588.000 568.755 ;
        RECT 3379.715 565.995 3588.000 566.835 ;
        RECT 3379.435 563.615 3588.000 565.995 ;
        RECT 3379.715 562.775 3588.000 563.615 ;
        RECT 3379.435 560.395 3588.000 562.775 ;
        RECT 3379.715 559.555 3588.000 560.395 ;
        RECT 3379.435 557.635 3588.000 559.555 ;
        RECT 3379.715 556.795 3588.000 557.635 ;
        RECT 3379.435 554.415 3588.000 556.795 ;
        RECT 3379.715 553.575 3588.000 554.415 ;
        RECT 4.925 551.265 197.965 551.495 ;
        RECT 3379.435 551.195 3588.000 553.575 ;
        RECT 3379.715 550.355 3588.000 551.195 ;
        RECT 3379.435 548.435 3588.000 550.355 ;
        RECT 3379.715 547.595 3588.000 548.435 ;
        RECT 3379.435 545.215 3588.000 547.595 ;
        RECT 3379.715 544.375 3588.000 545.215 ;
        RECT 3379.435 541.995 3588.000 544.375 ;
      LAYER met2 ;
        RECT 3377.035 541.690 3379.435 541.715 ;
        RECT 3376.560 541.550 3379.435 541.690 ;
        RECT 3376.560 501.570 3376.700 541.550 ;
        RECT 3377.035 541.435 3379.435 541.550 ;
      LAYER met2 ;
        RECT 3379.715 541.155 3588.000 541.995 ;
        RECT 3379.435 538.775 3588.000 541.155 ;
        RECT 3379.715 537.935 3588.000 538.775 ;
        RECT 3379.435 536.015 3588.000 537.935 ;
        RECT 3379.715 535.175 3588.000 536.015 ;
        RECT 3379.435 532.795 3588.000 535.175 ;
        RECT 3379.715 531.955 3588.000 532.795 ;
        RECT 3379.435 529.575 3588.000 531.955 ;
        RECT 3379.715 528.735 3588.000 529.575 ;
        RECT 3379.435 526.815 3588.000 528.735 ;
      LAYER met2 ;
        RECT 3377.035 526.255 3379.435 526.535 ;
      LAYER met2 ;
        RECT 3379.715 525.975 3588.000 526.815 ;
        RECT 3379.435 523.595 3588.000 525.975 ;
        RECT 3379.715 522.755 3588.000 523.595 ;
        RECT 3379.435 520.375 3588.000 522.755 ;
      LAYER met2 ;
        RECT 3377.035 519.815 3379.435 520.095 ;
      LAYER met2 ;
        RECT 3379.715 519.535 3588.000 520.375 ;
        RECT 3379.435 517.615 3588.000 519.535 ;
      LAYER met2 ;
        RECT 3377.035 517.055 3379.435 517.335 ;
      LAYER met2 ;
        RECT 3379.715 516.775 3588.000 517.615 ;
        RECT 3379.435 514.395 3588.000 516.775 ;
        RECT 3379.715 513.555 3588.000 514.395 ;
        RECT 3379.435 511.175 3588.000 513.555 ;
        RECT 3379.715 510.335 3588.000 511.175 ;
        RECT 3379.435 508.415 3588.000 510.335 ;
      LAYER met2 ;
        RECT 3377.035 507.855 3379.435 508.135 ;
      LAYER met2 ;
        RECT 3379.715 507.575 3588.000 508.415 ;
        RECT 3379.435 505.195 3588.000 507.575 ;
        RECT 3379.715 504.355 3588.000 505.195 ;
        RECT 3379.435 501.975 3588.000 504.355 ;
      LAYER met2 ;
        RECT 3377.035 501.570 3379.435 501.695 ;
        RECT 3376.560 501.430 3379.435 501.570 ;
        RECT 3377.035 501.415 3379.435 501.430 ;
      LAYER met2 ;
        RECT 3379.715 501.135 3588.000 501.975 ;
        RECT 3379.435 500.085 3588.000 501.135 ;
        RECT 0.035 416.200 151.405 425.935 ;
        RECT 153.765 415.000 158.415 426.140 ;
        RECT 160.165 416.200 174.575 425.935 ;
        RECT 0.035 414.700 197.965 415.000 ;
        RECT 0.035 394.095 198.000 414.700 ;
        RECT 0.035 393.535 197.965 394.095 ;
        RECT 0.035 360.925 198.000 393.535 ;
        RECT 0.035 360.495 197.965 360.925 ;
        RECT 0.035 340.500 198.000 360.495 ;
        RECT 0.035 340.000 197.965 340.500 ;
        RECT 153.800 329.025 158.450 340.000 ;
      LAYER met2 ;
        RECT 933.440 221.010 933.700 221.330 ;
        RECT 973.460 221.010 973.720 221.330 ;
        RECT 933.500 210.965 933.640 221.010 ;
        RECT 973.520 210.965 973.660 221.010 ;
        RECT 1476.240 220.670 1476.500 220.990 ;
        RECT 1516.260 220.670 1516.520 220.990 ;
        RECT 1750.400 220.670 1750.660 220.990 ;
        RECT 1790.420 220.670 1790.680 220.990 ;
        RECT 2024.560 220.670 2024.820 220.990 ;
        RECT 2064.580 220.670 2064.840 220.990 ;
        RECT 2298.260 220.670 2298.520 220.990 ;
        RECT 2338.280 220.670 2338.540 220.990 ;
        RECT 2572.420 220.670 2572.680 220.990 ;
        RECT 2612.440 220.670 2612.700 220.990 ;
        RECT 1476.300 210.965 1476.440 220.670 ;
        RECT 1516.320 210.965 1516.460 220.670 ;
        RECT 1750.460 210.965 1750.600 220.670 ;
        RECT 1790.480 210.965 1790.620 220.670 ;
        RECT 2024.620 210.965 2024.760 220.670 ;
        RECT 2064.640 210.965 2064.780 220.670 ;
        RECT 2298.320 210.965 2298.460 220.670 ;
        RECT 2338.340 210.965 2338.480 220.670 ;
        RECT 2572.480 210.965 2572.620 220.670 ;
        RECT 2612.500 210.965 2612.640 220.670 ;
        RECT 933.415 208.565 933.695 210.965 ;
        RECT 939.855 208.565 940.135 210.965 ;
        RECT 949.055 208.565 949.335 210.965 ;
        RECT 951.815 208.565 952.095 210.965 ;
        RECT 958.255 208.565 958.535 210.965 ;
        RECT 973.435 208.565 973.715 210.965 ;
        RECT 1010.235 208.565 1010.515 210.965 ;
        RECT 1476.300 209.030 1476.695 210.965 ;
        RECT 1476.415 208.565 1476.695 209.030 ;
        RECT 1479.635 208.565 1479.915 210.965 ;
        RECT 1482.855 208.565 1483.135 210.965 ;
        RECT 1492.055 208.565 1492.335 210.965 ;
        RECT 1494.815 208.565 1495.095 210.965 ;
        RECT 1501.255 208.565 1501.535 210.965 ;
        RECT 1516.320 209.030 1516.715 210.965 ;
        RECT 1516.435 208.565 1516.715 209.030 ;
        RECT 1553.235 208.565 1553.515 210.965 ;
        RECT 1750.415 208.565 1750.695 210.965 ;
        RECT 1753.635 208.565 1753.915 210.965 ;
        RECT 1756.855 208.565 1757.135 210.965 ;
        RECT 1766.055 208.565 1766.335 210.965 ;
        RECT 1768.815 208.565 1769.095 210.965 ;
        RECT 1775.255 208.565 1775.535 210.965 ;
        RECT 1790.435 208.565 1790.715 210.965 ;
        RECT 1827.235 208.565 1827.515 210.965 ;
        RECT 2024.415 209.100 2024.760 210.965 ;
        RECT 2024.415 208.565 2024.695 209.100 ;
        RECT 2030.855 208.565 2031.135 210.965 ;
        RECT 2040.055 208.565 2040.335 210.965 ;
        RECT 2042.815 208.565 2043.095 210.965 ;
        RECT 2049.255 208.565 2049.535 210.965 ;
        RECT 2064.435 209.100 2064.780 210.965 ;
        RECT 2064.435 208.565 2064.715 209.100 ;
        RECT 2101.235 208.565 2101.515 210.965 ;
        RECT 2298.320 209.030 2298.695 210.965 ;
        RECT 2298.415 208.565 2298.695 209.030 ;
        RECT 2304.855 208.565 2305.135 210.965 ;
        RECT 2314.055 208.565 2314.335 210.965 ;
        RECT 2316.815 208.565 2317.095 210.965 ;
        RECT 2323.255 208.565 2323.535 210.965 ;
        RECT 2338.340 209.030 2338.715 210.965 ;
        RECT 2338.435 208.565 2338.715 209.030 ;
        RECT 2375.235 208.565 2375.515 210.965 ;
        RECT 2572.415 208.565 2572.695 210.965 ;
        RECT 2578.855 208.565 2579.135 210.965 ;
        RECT 2588.055 208.565 2588.335 210.965 ;
        RECT 2590.815 208.565 2591.095 210.965 ;
        RECT 2597.255 208.565 2597.535 210.965 ;
        RECT 2612.435 208.565 2612.715 210.965 ;
        RECT 2649.235 208.565 2649.515 210.965 ;
      LAYER met2 ;
        RECT 932.085 208.285 933.135 208.565 ;
        RECT 933.975 208.285 936.355 208.565 ;
        RECT 937.195 208.285 939.575 208.565 ;
        RECT 940.415 208.285 942.335 208.565 ;
        RECT 943.175 208.285 945.555 208.565 ;
        RECT 946.395 208.285 948.775 208.565 ;
        RECT 949.615 208.285 951.535 208.565 ;
        RECT 952.375 208.285 954.755 208.565 ;
        RECT 955.595 208.285 957.975 208.565 ;
        RECT 958.815 208.285 960.735 208.565 ;
        RECT 961.575 208.285 963.955 208.565 ;
        RECT 964.795 208.285 967.175 208.565 ;
        RECT 968.015 208.285 969.935 208.565 ;
        RECT 970.775 208.285 973.155 208.565 ;
        RECT 973.995 208.285 976.375 208.565 ;
        RECT 977.215 208.285 979.595 208.565 ;
        RECT 980.435 208.285 982.355 208.565 ;
        RECT 983.195 208.285 985.575 208.565 ;
        RECT 986.415 208.285 988.795 208.565 ;
        RECT 989.635 208.285 991.555 208.565 ;
        RECT 992.395 208.285 994.775 208.565 ;
        RECT 995.615 208.285 997.995 208.565 ;
        RECT 998.835 208.285 1000.755 208.565 ;
        RECT 1001.595 208.285 1003.975 208.565 ;
        RECT 1004.815 208.285 1007.195 208.565 ;
        RECT 1008.035 208.285 1009.955 208.565 ;
        RECT 1010.795 208.285 1011.790 208.565 ;
      LAYER met2 ;
        RECT 675.840 201.125 676.100 201.270 ;
        RECT 717.700 201.125 717.960 201.270 ;
        RECT 675.830 200.755 676.110 201.125 ;
        RECT 717.690 200.755 717.970 201.125 ;
      LAYER met2 ;
        RECT 394.710 197.965 418.610 200.000 ;
        RECT 441.105 198.080 443.105 200.000 ;
        RECT 444.605 197.965 468.505 200.000 ;
        RECT 663.085 199.390 664.485 200.000 ;
      LAYER met2 ;
        RECT 664.765 199.670 665.785 200.000 ;
      LAYER met2 ;
        RECT 666.065 199.390 704.700 200.000 ;
        RECT 663.085 199.080 704.700 199.390 ;
        RECT 705.520 199.390 706.565 200.000 ;
      LAYER met2 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met2 ;
        RECT 707.775 199.390 708.055 200.000 ;
        RECT 709.345 199.390 709.490 200.000 ;
      LAYER met2 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met2 ;
        RECT 710.700 199.390 715.060 200.000 ;
        RECT 705.520 199.080 715.060 199.390 ;
        RECT 394.710 4.925 468.735 197.965 ;
        RECT 663.085 196.020 715.060 199.080 ;
        RECT 715.920 198.310 716.495 200.000 ;
      LAYER met2 ;
        RECT 716.775 198.590 717.925 200.000 ;
      LAYER met2 ;
        RECT 718.205 199.155 718.810 200.000 ;
      LAYER met2 ;
        RECT 719.090 199.435 720.755 200.000 ;
      LAYER met2 ;
        RECT 721.035 199.155 722.585 200.000 ;
        RECT 718.205 198.735 722.585 199.155 ;
        RECT 723.725 198.735 725.175 200.000 ;
        RECT 718.205 198.310 725.175 198.735 ;
        RECT 715.920 198.250 725.175 198.310 ;
        RECT 725.995 199.390 728.825 200.000 ;
      LAYER met2 ;
        RECT 729.105 199.670 729.575 200.000 ;
      LAYER met2 ;
        RECT 729.855 199.390 737.660 200.000 ;
        RECT 725.995 198.250 737.660 199.390 ;
        RECT 715.920 196.845 737.660 198.250 ;
        RECT 715.920 196.485 722.475 196.845 ;
        RECT 727.600 196.705 737.660 196.845 ;
        RECT 715.920 196.215 722.205 196.485 ;
        RECT 727.930 196.375 737.660 196.705 ;
        RECT 715.920 196.035 721.835 196.215 ;
        RECT 663.085 195.735 714.775 196.020 ;
        RECT 716.220 195.845 721.835 196.035 ;
        RECT 723.505 195.925 726.790 196.025 ;
        RECT 716.220 195.735 721.725 195.845 ;
        RECT 723.405 195.790 726.790 195.925 ;
      LAYER met2 ;
        RECT 727.305 195.955 727.625 196.070 ;
        RECT 727.650 195.955 727.995 196.095 ;
      LAYER met2 ;
        RECT 728.275 196.030 737.660 196.375 ;
      LAYER met2 ;
        RECT 727.305 195.815 727.995 195.955 ;
      LAYER met2 ;
        RECT 663.085 195.380 708.600 195.735 ;
        RECT 723.405 195.655 727.025 195.790 ;
      LAYER met2 ;
        RECT 727.305 195.750 727.625 195.815 ;
        RECT 727.650 195.750 727.995 195.815 ;
      LAYER met2 ;
        RECT 723.135 195.470 727.025 195.655 ;
      LAYER met2 ;
        RECT 727.625 195.675 727.955 195.750 ;
        RECT 727.995 195.675 728.265 195.750 ;
      LAYER met2 ;
        RECT 663.085 195.050 708.270 195.380 ;
        RECT 723.135 195.285 727.345 195.470 ;
      LAYER met2 ;
        RECT 727.625 195.425 728.265 195.675 ;
        RECT 727.625 195.420 727.955 195.425 ;
      LAYER met2 ;
        RECT 722.765 195.140 727.345 195.285 ;
        RECT 663.085 189.305 708.140 195.050 ;
        RECT 722.765 194.915 727.725 195.140 ;
        RECT 709.625 194.820 727.725 194.915 ;
        RECT 709.530 194.490 727.725 194.820 ;
        RECT 709.200 194.250 727.725 194.490 ;
        RECT 708.960 191.420 727.725 194.250 ;
        RECT 708.960 191.080 727.385 191.420 ;
      LAYER met2 ;
        RECT 728.005 191.140 728.265 195.425 ;
      LAYER met2 ;
        RECT 708.960 190.880 727.185 191.080 ;
      LAYER met2 ;
        RECT 727.665 190.890 728.265 191.140 ;
      LAYER met2 ;
        RECT 708.960 190.550 726.855 190.880 ;
      LAYER met2 ;
        RECT 727.665 190.800 728.005 190.890 ;
        RECT 728.035 190.800 728.265 190.890 ;
        RECT 727.465 190.750 727.665 190.800 ;
        RECT 727.835 190.750 728.035 190.800 ;
        RECT 727.465 190.680 728.035 190.750 ;
        RECT 727.465 190.600 727.665 190.680 ;
        RECT 727.835 190.600 728.035 190.680 ;
      LAYER met2 ;
        RECT 663.085 189.115 707.950 189.305 ;
        RECT 663.085 184.635 707.690 189.115 ;
        RECT 708.960 188.555 726.595 190.550 ;
      LAYER met2 ;
        RECT 727.135 190.540 727.465 190.600 ;
        RECT 727.505 190.540 727.835 190.600 ;
        RECT 727.135 190.400 727.835 190.540 ;
      LAYER met2 ;
        RECT 728.545 190.520 737.660 196.030 ;
      LAYER met2 ;
        RECT 727.135 190.270 727.465 190.400 ;
        RECT 727.505 190.270 727.835 190.400 ;
      LAYER met2 ;
        RECT 728.315 190.320 737.660 190.520 ;
        RECT 708.880 188.185 726.595 188.555 ;
        RECT 663.085 184.300 707.355 184.635 ;
        RECT 663.085 179.225 707.095 184.300 ;
        RECT 708.510 183.740 726.595 188.185 ;
        RECT 708.285 183.370 726.595 183.740 ;
        RECT 707.915 179.225 726.595 183.370 ;
        RECT 663.085 172.420 726.595 179.225 ;
      LAYER met2 ;
        RECT 726.875 189.900 727.505 190.270 ;
      LAYER met2 ;
        RECT 728.115 189.990 737.660 190.320 ;
      LAYER met2 ;
        RECT 726.875 173.390 727.135 189.900 ;
      LAYER met2 ;
        RECT 727.785 189.620 737.660 189.990 ;
        RECT 727.415 173.670 737.660 189.620 ;
      LAYER met2 ;
        RECT 726.875 172.700 727.350 173.390 ;
      LAYER met2 ;
        RECT 663.085 172.345 726.810 172.420 ;
        RECT 663.085 169.195 726.595 172.345 ;
      LAYER met2 ;
        RECT 727.090 172.065 727.350 172.700 ;
        RECT 726.875 171.855 727.350 172.065 ;
        RECT 726.875 171.850 727.090 171.855 ;
        RECT 726.875 171.375 727.350 171.850 ;
      LAYER met2 ;
        RECT 663.085 169.050 726.450 169.195 ;
        RECT 663.085 168.825 726.225 169.050 ;
      LAYER met2 ;
        RECT 726.875 168.915 727.135 171.375 ;
      LAYER met2 ;
        RECT 727.630 171.095 737.660 173.670 ;
        RECT 663.085 164.260 726.200 168.825 ;
      LAYER met2 ;
        RECT 726.730 168.770 727.135 168.915 ;
        RECT 726.505 168.735 726.730 168.770 ;
        RECT 726.875 168.735 727.135 168.770 ;
        RECT 726.505 168.665 727.135 168.735 ;
        RECT 726.505 168.545 726.730 168.665 ;
        RECT 726.875 168.545 727.135 168.665 ;
        RECT 726.480 168.520 726.505 168.545 ;
        RECT 726.740 168.520 726.875 168.545 ;
        RECT 726.480 168.410 726.875 168.520 ;
      LAYER met2 ;
        RECT 663.085 163.440 725.570 164.260 ;
      LAYER met2 ;
        RECT 726.480 163.980 726.740 168.410 ;
      LAYER met2 ;
        RECT 727.415 168.265 737.660 171.095 ;
        RECT 727.155 168.130 737.660 168.265 ;
      LAYER met2 ;
        RECT 725.850 163.720 726.740 163.980 ;
      LAYER met2 ;
        RECT 727.020 163.440 737.660 168.130 ;
        RECT 663.085 0.790 737.660 163.440 ;
        RECT 932.085 0.000 1011.790 208.285 ;
        RECT 1475.085 208.285 1476.135 208.565 ;
        RECT 1476.975 208.285 1479.355 208.565 ;
        RECT 1480.195 208.285 1482.575 208.565 ;
        RECT 1483.415 208.285 1485.335 208.565 ;
        RECT 1486.175 208.285 1488.555 208.565 ;
        RECT 1489.395 208.285 1491.775 208.565 ;
        RECT 1492.615 208.285 1494.535 208.565 ;
        RECT 1495.375 208.285 1497.755 208.565 ;
        RECT 1498.595 208.285 1500.975 208.565 ;
        RECT 1501.815 208.285 1503.735 208.565 ;
        RECT 1504.575 208.285 1506.955 208.565 ;
        RECT 1507.795 208.285 1510.175 208.565 ;
        RECT 1511.015 208.285 1512.935 208.565 ;
        RECT 1513.775 208.285 1516.155 208.565 ;
        RECT 1516.995 208.285 1519.375 208.565 ;
        RECT 1520.215 208.285 1522.595 208.565 ;
        RECT 1523.435 208.285 1525.355 208.565 ;
        RECT 1526.195 208.285 1528.575 208.565 ;
        RECT 1529.415 208.285 1531.795 208.565 ;
        RECT 1532.635 208.285 1534.555 208.565 ;
        RECT 1535.395 208.285 1537.775 208.565 ;
        RECT 1538.615 208.285 1540.995 208.565 ;
        RECT 1541.835 208.285 1543.755 208.565 ;
        RECT 1544.595 208.285 1546.975 208.565 ;
        RECT 1547.815 208.285 1550.195 208.565 ;
        RECT 1551.035 208.285 1552.955 208.565 ;
        RECT 1553.795 208.285 1554.790 208.565 ;
        RECT 1206.300 197.965 1226.905 198.000 ;
        RECT 1227.465 197.965 1260.075 198.000 ;
        RECT 1260.505 197.965 1280.500 198.000 ;
        RECT 1195.065 160.165 1204.800 174.575 ;
        RECT 1206.000 158.450 1281.000 197.965 ;
        RECT 1206.000 158.415 1291.975 158.450 ;
        RECT 1194.860 153.800 1291.975 158.415 ;
        RECT 1194.860 153.765 1281.000 153.800 ;
        RECT 1195.065 0.035 1204.800 151.405 ;
        RECT 1206.000 0.035 1281.000 153.765 ;
        RECT 1475.085 0.000 1554.790 208.285 ;
        RECT 1749.085 208.285 1750.135 208.565 ;
        RECT 1750.975 208.285 1753.355 208.565 ;
        RECT 1754.195 208.285 1756.575 208.565 ;
        RECT 1757.415 208.285 1759.335 208.565 ;
        RECT 1760.175 208.285 1762.555 208.565 ;
        RECT 1763.395 208.285 1765.775 208.565 ;
        RECT 1766.615 208.285 1768.535 208.565 ;
        RECT 1769.375 208.285 1771.755 208.565 ;
        RECT 1772.595 208.285 1774.975 208.565 ;
        RECT 1775.815 208.285 1777.735 208.565 ;
        RECT 1778.575 208.285 1780.955 208.565 ;
        RECT 1781.795 208.285 1784.175 208.565 ;
        RECT 1785.015 208.285 1786.935 208.565 ;
        RECT 1787.775 208.285 1790.155 208.565 ;
        RECT 1790.995 208.285 1793.375 208.565 ;
        RECT 1794.215 208.285 1796.595 208.565 ;
        RECT 1797.435 208.285 1799.355 208.565 ;
        RECT 1800.195 208.285 1802.575 208.565 ;
        RECT 1803.415 208.285 1805.795 208.565 ;
        RECT 1806.635 208.285 1808.555 208.565 ;
        RECT 1809.395 208.285 1811.775 208.565 ;
        RECT 1812.615 208.285 1814.995 208.565 ;
        RECT 1815.835 208.285 1817.755 208.565 ;
        RECT 1818.595 208.285 1820.975 208.565 ;
        RECT 1821.815 208.285 1824.195 208.565 ;
        RECT 1825.035 208.285 1826.955 208.565 ;
        RECT 1827.795 208.285 1828.790 208.565 ;
        RECT 1749.085 0.000 1828.790 208.285 ;
        RECT 2023.085 208.285 2024.135 208.565 ;
        RECT 2024.975 208.285 2027.355 208.565 ;
        RECT 2028.195 208.285 2030.575 208.565 ;
        RECT 2031.415 208.285 2033.335 208.565 ;
        RECT 2034.175 208.285 2036.555 208.565 ;
        RECT 2037.395 208.285 2039.775 208.565 ;
        RECT 2040.615 208.285 2042.535 208.565 ;
        RECT 2043.375 208.285 2045.755 208.565 ;
        RECT 2046.595 208.285 2048.975 208.565 ;
        RECT 2049.815 208.285 2051.735 208.565 ;
        RECT 2052.575 208.285 2054.955 208.565 ;
        RECT 2055.795 208.285 2058.175 208.565 ;
        RECT 2059.015 208.285 2060.935 208.565 ;
        RECT 2061.775 208.285 2064.155 208.565 ;
        RECT 2064.995 208.285 2067.375 208.565 ;
        RECT 2068.215 208.285 2070.595 208.565 ;
        RECT 2071.435 208.285 2073.355 208.565 ;
        RECT 2074.195 208.285 2076.575 208.565 ;
        RECT 2077.415 208.285 2079.795 208.565 ;
        RECT 2080.635 208.285 2082.555 208.565 ;
        RECT 2083.395 208.285 2085.775 208.565 ;
        RECT 2086.615 208.285 2088.995 208.565 ;
        RECT 2089.835 208.285 2091.755 208.565 ;
        RECT 2092.595 208.285 2094.975 208.565 ;
        RECT 2095.815 208.285 2098.195 208.565 ;
        RECT 2099.035 208.285 2100.955 208.565 ;
        RECT 2101.795 208.285 2102.790 208.565 ;
        RECT 2023.085 0.000 2102.790 208.285 ;
        RECT 2297.085 208.285 2298.135 208.565 ;
        RECT 2298.975 208.285 2301.355 208.565 ;
        RECT 2302.195 208.285 2304.575 208.565 ;
        RECT 2305.415 208.285 2307.335 208.565 ;
        RECT 2308.175 208.285 2310.555 208.565 ;
        RECT 2311.395 208.285 2313.775 208.565 ;
        RECT 2314.615 208.285 2316.535 208.565 ;
        RECT 2317.375 208.285 2319.755 208.565 ;
        RECT 2320.595 208.285 2322.975 208.565 ;
        RECT 2323.815 208.285 2325.735 208.565 ;
        RECT 2326.575 208.285 2328.955 208.565 ;
        RECT 2329.795 208.285 2332.175 208.565 ;
        RECT 2333.015 208.285 2334.935 208.565 ;
        RECT 2335.775 208.285 2338.155 208.565 ;
        RECT 2338.995 208.285 2341.375 208.565 ;
        RECT 2342.215 208.285 2344.595 208.565 ;
        RECT 2345.435 208.285 2347.355 208.565 ;
        RECT 2348.195 208.285 2350.575 208.565 ;
        RECT 2351.415 208.285 2353.795 208.565 ;
        RECT 2354.635 208.285 2356.555 208.565 ;
        RECT 2357.395 208.285 2359.775 208.565 ;
        RECT 2360.615 208.285 2362.995 208.565 ;
        RECT 2363.835 208.285 2365.755 208.565 ;
        RECT 2366.595 208.285 2368.975 208.565 ;
        RECT 2369.815 208.285 2372.195 208.565 ;
        RECT 2373.035 208.285 2374.955 208.565 ;
        RECT 2375.795 208.285 2376.790 208.565 ;
        RECT 2297.085 0.000 2376.790 208.285 ;
        RECT 2571.085 208.285 2572.135 208.565 ;
        RECT 2572.975 208.285 2575.355 208.565 ;
        RECT 2576.195 208.285 2578.575 208.565 ;
        RECT 2579.415 208.285 2581.335 208.565 ;
        RECT 2582.175 208.285 2584.555 208.565 ;
        RECT 2585.395 208.285 2587.775 208.565 ;
        RECT 2588.615 208.285 2590.535 208.565 ;
        RECT 2591.375 208.285 2593.755 208.565 ;
        RECT 2594.595 208.285 2596.975 208.565 ;
        RECT 2597.815 208.285 2599.735 208.565 ;
        RECT 2600.575 208.285 2602.955 208.565 ;
        RECT 2603.795 208.285 2606.175 208.565 ;
        RECT 2607.015 208.285 2608.935 208.565 ;
        RECT 2609.775 208.285 2612.155 208.565 ;
        RECT 2612.995 208.285 2615.375 208.565 ;
        RECT 2616.215 208.285 2618.595 208.565 ;
        RECT 2619.435 208.285 2621.355 208.565 ;
        RECT 2622.195 208.285 2624.575 208.565 ;
        RECT 2625.415 208.285 2627.795 208.565 ;
        RECT 2628.635 208.285 2630.555 208.565 ;
        RECT 2631.395 208.285 2633.775 208.565 ;
        RECT 2634.615 208.285 2636.995 208.565 ;
        RECT 2637.835 208.285 2639.755 208.565 ;
        RECT 2640.595 208.285 2642.975 208.565 ;
        RECT 2643.815 208.285 2646.195 208.565 ;
        RECT 2647.035 208.285 2648.955 208.565 ;
        RECT 2649.795 208.285 2650.790 208.565 ;
        RECT 2571.085 0.000 2650.790 208.285 ;
        RECT 2845.710 197.965 2869.610 200.000 ;
        RECT 2892.105 198.080 2894.105 200.000 ;
        RECT 2895.605 197.965 2919.505 200.000 ;
        RECT 3114.710 197.965 3138.610 200.000 ;
        RECT 3161.105 198.080 3163.105 200.000 ;
        RECT 3164.605 197.965 3188.505 200.000 ;
        RECT 2845.710 4.925 2919.735 197.965 ;
        RECT 3114.710 4.925 3188.735 197.965 ;
      LAYER via2 ;
        RECT 675.830 200.800 676.110 201.080 ;
        RECT 717.690 200.800 717.970 201.080 ;
      LAYER met3 ;
        RECT 381.310 4986.690 460.570 5188.000 ;
        RECT 638.310 4986.690 717.570 5188.000 ;
        RECT 895.310 4986.690 974.570 5188.000 ;
        RECT 1152.310 4986.690 1231.570 5188.000 ;
        RECT 1410.310 4986.690 1489.570 5188.000 ;
        RECT 1667.240 5014.250 1741.290 5188.000 ;
        RECT 1691.795 4990.035 1716.990 5014.250 ;
        RECT 1692.895 4988.000 1703.895 4990.035 ;
        RECT 1704.890 4988.000 1715.890 4990.035 ;
        RECT 1919.310 4986.690 1998.570 5188.000 ;
        RECT 2364.310 4986.690 2443.570 5188.000 ;
        RECT 2621.310 4986.690 2700.570 5188.000 ;
        RECT 2878.240 5025.160 2952.290 5183.100 ;
        RECT 2878.240 5020.915 2927.990 5025.160 ;
        RECT 2902.795 4990.035 2927.990 5020.915 ;
        RECT 2903.895 4988.000 2914.895 4990.035 ;
        RECT 2915.890 4988.000 2926.890 4990.035 ;
        RECT 3130.310 4986.690 3209.570 5188.000 ;
        RECT 0.000 4771.310 201.310 4850.570 ;
        RECT 3386.690 4758.430 3588.000 4837.690 ;
        RECT 153.765 4635.605 158.415 4646.140 ;
        RECT 159.805 4635.440 163.270 4646.140 ;
        RECT 4.395 4610.355 190.700 4635.000 ;
        RECT 4.395 4609.255 197.965 4610.355 ;
        RECT 4.395 4598.380 198.000 4609.255 ;
        RECT 4.395 4596.880 197.965 4598.380 ;
        RECT 4.395 4586.000 198.000 4596.880 ;
        RECT 3397.300 4588.100 3583.605 4612.510 ;
        RECT 3390.035 4587.000 3583.605 4588.100 ;
        RECT 4.395 4584.900 197.965 4586.000 ;
        RECT 4.395 4560.490 190.700 4584.900 ;
        RECT 3390.000 4576.120 3583.605 4587.000 ;
        RECT 3390.035 4574.620 3583.605 4576.120 ;
        RECT 3390.000 4563.745 3583.605 4574.620 ;
        RECT 3390.035 4562.645 3583.605 4563.745 ;
        RECT 3397.300 4538.000 3583.605 4562.645 ;
        RECT 3424.730 4526.860 3428.195 4537.560 ;
        RECT 3429.585 4526.860 3434.235 4537.395 ;
        RECT 0.000 4398.990 179.800 4423.290 ;
      LAYER met3 ;
        RECT 180.200 4399.390 200.000 4423.290 ;
      LAYER met3 ;
        RECT 0.000 4397.890 197.965 4398.990 ;
        RECT 0.000 4386.890 200.000 4397.890 ;
        RECT 0.000 4385.895 197.965 4386.890 ;
        RECT 0.000 4374.895 200.000 4385.895 ;
        RECT 0.000 4373.795 197.965 4374.895 ;
        RECT 0.000 4349.240 179.800 4373.795 ;
        RECT 3386.690 4312.430 3588.000 4391.690 ;
        RECT 4.900 4187.990 162.840 4212.290 ;
        RECT 4.900 4186.890 197.965 4187.990 ;
        RECT 4.900 4175.890 200.000 4186.890 ;
        RECT 4.900 4174.895 197.965 4175.890 ;
        RECT 4.900 4163.895 200.000 4174.895 ;
        RECT 4.900 4162.795 197.965 4163.895 ;
        RECT 4.900 4138.240 167.085 4162.795 ;
        RECT 3403.360 4142.205 3588.000 4166.760 ;
        RECT 3390.035 4141.105 3588.000 4142.205 ;
        RECT 3388.000 4130.105 3588.000 4141.105 ;
        RECT 3390.035 4129.110 3588.000 4130.105 ;
        RECT 3388.000 4118.110 3588.000 4129.110 ;
        RECT 3390.035 4117.010 3588.000 4118.110 ;
        RECT 3403.360 4092.710 3588.000 4117.010 ;
        RECT 0.000 3922.310 201.310 4001.570 ;
        RECT 3386.690 3866.430 3588.000 3945.690 ;
        RECT 0.000 3706.310 201.310 3785.570 ;
        RECT 3386.690 3641.430 3588.000 3720.690 ;
        RECT 0.000 3490.310 201.310 3569.570 ;
        RECT 3386.690 3416.430 3588.000 3495.690 ;
        RECT 0.000 3274.310 201.310 3353.570 ;
        RECT 3386.690 3190.430 3588.000 3269.690 ;
        RECT 0.000 3058.310 201.310 3137.570 ;
        RECT 3386.690 2965.430 3588.000 3044.690 ;
        RECT 0.000 2842.310 201.310 2921.570 ;
        RECT 3386.690 2739.430 3588.000 2818.690 ;
        RECT 0.000 2626.310 201.310 2705.570 ;
        RECT 3403.360 2569.205 3588.000 2593.760 ;
        RECT 3390.035 2568.105 3588.000 2569.205 ;
        RECT 3388.000 2557.105 3588.000 2568.105 ;
        RECT 3390.035 2556.110 3588.000 2557.105 ;
        RECT 3388.000 2545.110 3588.000 2556.110 ;
        RECT 3390.035 2544.010 3588.000 2545.110 ;
      LAYER met3 ;
        RECT 3403.360 2519.710 3588.000 2544.010 ;
        RECT 0.000 2464.990 184.640 2489.290 ;
        RECT 0.000 2463.890 197.965 2464.990 ;
        RECT 0.000 2452.890 200.000 2463.890 ;
        RECT 0.000 2451.895 197.965 2452.890 ;
        RECT 0.000 2440.895 200.000 2451.895 ;
        RECT 0.000 2439.795 197.965 2440.895 ;
        RECT 0.000 2415.240 184.640 2439.795 ;
        RECT 3430.000 2349.100 3583.605 2373.500 ;
        RECT 3390.035 2348.000 3583.605 2349.100 ;
        RECT 3390.000 2337.120 3583.605 2348.000 ;
        RECT 3390.035 2335.620 3583.605 2337.120 ;
        RECT 3390.000 2324.745 3583.605 2335.620 ;
        RECT 3390.035 2323.645 3583.605 2324.745 ;
        RECT 3430.000 2299.000 3583.605 2323.645 ;
        RECT 153.765 2279.605 158.415 2290.140 ;
        RECT 159.805 2279.440 163.270 2290.140 ;
        RECT 3424.730 2287.860 3428.195 2298.560 ;
        RECT 3429.585 2287.860 3434.235 2298.395 ;
        RECT 4.395 2254.355 158.000 2279.000 ;
        RECT 4.395 2253.255 197.965 2254.355 ;
        RECT 4.395 2242.380 198.000 2253.255 ;
        RECT 4.395 2240.880 197.965 2242.380 ;
        RECT 4.395 2230.000 198.000 2240.880 ;
        RECT 4.395 2228.900 197.965 2230.000 ;
        RECT 4.395 2204.500 158.000 2228.900 ;
        RECT 3420.915 2128.205 3583.100 2152.760 ;
        RECT 3390.035 2127.105 3583.100 2128.205 ;
        RECT 3388.000 2116.105 3583.100 2127.105 ;
        RECT 3390.035 2115.110 3583.100 2116.105 ;
        RECT 3388.000 2104.110 3583.100 2115.110 ;
        RECT 3390.035 2103.010 3583.100 2104.110 ;
      LAYER met3 ;
        RECT 3388.000 2078.710 3424.760 2102.610 ;
      LAYER met3 ;
        RECT 3425.160 2078.710 3583.100 2103.010 ;
        RECT 0.000 1988.310 201.310 2067.570 ;
        RECT 3386.690 1853.430 3588.000 1932.690 ;
        RECT 0.000 1772.310 201.310 1851.570 ;
        RECT 0.000 1556.310 201.310 1635.570 ;
        RECT 3386.690 1627.430 3588.000 1706.690 ;
        RECT 0.000 1340.310 201.310 1419.570 ;
        RECT 3386.690 1402.430 3588.000 1481.690 ;
        RECT 0.000 1124.310 201.310 1203.570 ;
        RECT 3386.690 1177.430 3588.000 1256.690 ;
        RECT 0.000 908.310 201.310 987.570 ;
        RECT 3386.690 951.430 3588.000 1030.690 ;
        RECT 3386.690 726.430 3588.000 805.690 ;
        RECT 0.000 600.990 179.800 625.290 ;
        RECT 0.000 599.890 197.965 600.990 ;
        RECT 0.000 588.890 200.000 599.890 ;
        RECT 0.000 587.895 197.965 588.890 ;
        RECT 0.000 576.895 200.000 587.895 ;
        RECT 0.000 575.795 197.965 576.895 ;
        RECT 0.000 551.240 179.800 575.795 ;
        RECT 3386.690 500.430 3588.000 579.690 ;
        RECT 0.035 416.200 24.250 425.935 ;
        RECT 153.765 415.605 158.415 426.140 ;
        RECT 169.550 416.200 174.200 425.935 ;
        RECT 0.035 390.355 190.700 415.000 ;
        RECT 0.035 389.255 197.965 390.355 ;
        RECT 0.035 378.380 198.000 389.255 ;
        RECT 0.035 376.880 197.965 378.380 ;
        RECT 0.035 366.000 198.000 376.880 ;
        RECT 0.035 364.900 197.965 366.000 ;
        RECT 0.035 340.100 190.700 364.900 ;
        RECT 0.035 340.000 197.965 340.100 ;
        RECT 153.800 329.025 158.450 339.105 ;
      LAYER met3 ;
        RECT 675.805 201.090 676.135 201.105 ;
        RECT 665.470 200.790 676.135 201.090 ;
        RECT 665.470 200.000 665.770 200.790 ;
        RECT 675.805 200.775 676.135 200.790 ;
        RECT 717.665 201.090 717.995 201.105 ;
        RECT 717.665 200.790 720.050 201.090 ;
        RECT 717.665 200.775 717.995 200.790 ;
        RECT 719.750 200.000 720.050 200.790 ;
      LAYER met3 ;
        RECT 420.110 197.965 431.110 200.000 ;
        RECT 432.105 197.965 443.105 200.000 ;
      LAYER met3 ;
        RECT 238.000 164.765 256.010 180.085 ;
        RECT 258.000 164.765 276.010 180.085 ;
        RECT 278.000 164.765 296.010 180.085 ;
        RECT 298.000 164.765 316.010 180.085 ;
        RECT 318.000 164.765 336.010 180.085 ;
        RECT 338.000 164.765 356.010 180.085 ;
      LAYER met3 ;
        RECT 419.010 167.085 444.205 197.965 ;
        RECT 419.010 162.840 468.760 167.085 ;
      LAYER met3 ;
        RECT 507.000 164.765 525.010 180.085 ;
        RECT 527.000 164.765 545.010 180.085 ;
        RECT 547.000 164.765 565.010 180.085 ;
        RECT 567.000 164.765 585.010 180.085 ;
        RECT 587.000 164.765 605.010 180.085 ;
        RECT 607.000 164.765 625.010 180.085 ;
      LAYER met3 ;
        RECT 394.710 4.900 468.760 162.840 ;
        RECT 663.300 151.080 664.340 199.375 ;
        RECT 663.300 133.400 663.675 151.080 ;
      LAYER met3 ;
        RECT 664.740 150.680 665.810 200.000 ;
        RECT 664.075 150.080 665.810 150.680 ;
      LAYER met3 ;
        RECT 666.210 188.690 707.935 199.375 ;
        RECT 709.465 193.730 716.375 199.375 ;
        RECT 718.325 196.465 718.690 199.375 ;
      LAYER met3 ;
        RECT 719.090 196.865 720.755 200.000 ;
      LAYER met3 ;
        RECT 721.155 196.465 728.680 199.375 ;
        RECT 709.465 192.265 714.910 193.730 ;
        RECT 709.465 191.985 714.630 192.265 ;
        RECT 709.465 190.555 713.550 191.985 ;
      LAYER met3 ;
        RECT 715.030 191.585 715.310 191.865 ;
      LAYER met3 ;
        RECT 709.765 190.255 713.550 190.555 ;
        RECT 666.210 184.830 708.700 188.690 ;
        RECT 710.230 187.335 713.550 190.255 ;
      LAYER met3 ;
        RECT 713.950 191.500 715.030 191.585 ;
        RECT 715.095 191.500 716.660 191.585 ;
        RECT 713.950 190.600 716.660 191.500 ;
      LAYER met3 ;
        RECT 718.325 191.465 728.680 196.465 ;
        RECT 717.340 191.185 728.680 191.465 ;
      LAYER met3 ;
        RECT 713.950 190.505 715.030 190.600 ;
        RECT 715.095 190.505 716.660 190.600 ;
        RECT 713.950 190.020 716.660 190.505 ;
        RECT 713.950 187.735 715.095 190.020 ;
      LAYER met3 ;
        RECT 717.060 189.620 728.680 191.185 ;
        RECT 715.495 187.335 728.680 189.620 ;
        RECT 710.230 184.830 728.680 187.335 ;
        RECT 666.210 183.015 728.680 184.830 ;
        RECT 730.000 184.615 737.035 199.375 ;
        RECT 730.210 184.405 737.035 184.615 ;
        RECT 730.660 183.955 737.035 184.405 ;
      LAYER met3 ;
        RECT 729.670 183.255 730.130 183.415 ;
        RECT 730.260 183.255 730.710 183.555 ;
      LAYER met3 ;
        RECT 731.110 183.505 737.035 183.955 ;
      LAYER met3 ;
        RECT 729.670 183.105 730.710 183.255 ;
      LAYER met3 ;
        RECT 666.210 182.555 729.270 183.015 ;
      LAYER met3 ;
        RECT 729.670 182.955 731.225 183.105 ;
        RECT 730.130 182.655 730.705 182.955 ;
        RECT 730.710 182.655 731.225 182.955 ;
      LAYER met3 ;
        RECT 666.210 181.980 729.730 182.555 ;
      LAYER met3 ;
        RECT 730.130 182.380 731.225 182.655 ;
      LAYER met3 ;
        RECT 666.210 169.105 730.305 181.980 ;
        RECT 666.210 168.520 729.720 169.105 ;
      LAYER met3 ;
        RECT 730.705 168.705 731.225 182.380 ;
      LAYER met3 ;
        RECT 666.210 167.805 729.005 168.520 ;
      LAYER met3 ;
        RECT 730.120 168.345 731.225 168.705 ;
        RECT 730.120 168.120 730.705 168.345 ;
        RECT 730.850 168.120 731.225 168.345 ;
        RECT 729.405 168.045 730.120 168.120 ;
        RECT 730.135 168.045 730.850 168.120 ;
      LAYER met3 ;
        RECT 666.210 167.220 728.420 167.805 ;
      LAYER met3 ;
        RECT 729.405 167.595 730.850 168.045 ;
      LAYER met3 ;
        RECT 731.625 167.720 737.035 183.505 ;
      LAYER met3 ;
        RECT 729.405 167.405 730.120 167.595 ;
        RECT 730.135 167.405 730.850 167.595 ;
        RECT 728.820 167.295 729.405 167.405 ;
        RECT 729.550 167.295 730.135 167.405 ;
      LAYER met3 ;
        RECT 666.210 167.005 728.205 167.220 ;
        RECT 666.210 165.475 715.325 167.005 ;
      LAYER met3 ;
        RECT 728.820 166.995 730.135 167.295 ;
      LAYER met3 ;
        RECT 731.250 167.005 737.035 167.720 ;
      LAYER met3 ;
        RECT 728.820 166.820 729.405 166.995 ;
        RECT 729.550 166.820 730.135 166.995 ;
        RECT 728.605 166.605 728.820 166.820 ;
        RECT 729.030 166.605 729.550 166.820 ;
        RECT 715.725 166.455 729.550 166.605 ;
        RECT 715.725 166.300 728.885 166.305 ;
        RECT 729.030 166.300 729.550 166.455 ;
      LAYER met3 ;
        RECT 730.535 166.420 737.035 167.005 ;
      LAYER met3 ;
        RECT 715.725 166.155 729.030 166.300 ;
        RECT 728.605 166.005 729.030 166.155 ;
        RECT 715.725 165.875 729.030 166.005 ;
      LAYER met3 ;
        RECT 729.950 165.900 737.035 166.420 ;
        RECT 729.430 165.475 737.035 165.900 ;
      LAYER met3 ;
        RECT 664.075 150.015 664.740 150.080 ;
        RECT 664.075 135.400 665.810 150.015 ;
      LAYER met3 ;
        RECT 666.210 135.800 737.035 165.475 ;
      LAYER met3 ;
        RECT 776.000 164.765 794.010 180.085 ;
        RECT 796.000 164.765 814.010 180.085 ;
        RECT 816.000 164.765 834.010 180.085 ;
        RECT 836.000 164.765 854.010 180.085 ;
        RECT 856.000 164.765 874.010 180.085 ;
        RECT 876.000 164.765 894.010 180.085 ;
        RECT 664.075 133.800 667.410 135.400 ;
      LAYER met3 ;
        RECT 667.810 134.200 737.035 135.800 ;
        RECT 663.300 131.800 665.410 133.400 ;
      LAYER met3 ;
        RECT 665.810 132.400 668.810 133.800 ;
      LAYER met3 ;
        RECT 669.210 132.800 737.035 134.200 ;
      LAYER met3 ;
        RECT 665.810 132.250 669.745 132.400 ;
        RECT 665.810 132.200 667.410 132.250 ;
        RECT 667.410 131.950 668.695 132.200 ;
        RECT 668.810 131.950 669.745 132.250 ;
      LAYER met3 ;
        RECT 663.300 130.515 667.010 131.800 ;
      LAYER met3 ;
        RECT 667.410 131.465 669.745 131.950 ;
      LAYER met3 ;
        RECT 670.145 131.865 737.035 132.800 ;
      LAYER met3 ;
        RECT 667.410 131.350 669.710 131.465 ;
        RECT 667.410 131.200 668.695 131.350 ;
        RECT 669.745 131.200 670.610 131.465 ;
        RECT 667.410 131.050 670.610 131.200 ;
        RECT 667.410 130.915 668.695 131.050 ;
        RECT 668.695 130.900 669.645 130.915 ;
        RECT 669.745 130.900 670.610 131.050 ;
      LAYER met3 ;
        RECT 671.010 131.000 737.035 131.865 ;
      LAYER met3 ;
        RECT 668.695 130.600 670.610 130.900 ;
      LAYER met3 ;
        RECT 663.300 129.565 668.295 130.515 ;
      LAYER met3 ;
        RECT 668.695 130.450 671.960 130.600 ;
        RECT 668.695 130.300 669.645 130.450 ;
        RECT 670.610 130.300 671.960 130.450 ;
        RECT 668.695 130.000 671.960 130.300 ;
        RECT 668.695 129.965 669.645 130.000 ;
        RECT 670.610 129.965 671.960 130.000 ;
      LAYER met3 ;
        RECT 663.300 128.600 669.245 129.565 ;
      LAYER met3 ;
        RECT 669.645 129.250 671.960 129.965 ;
      LAYER met3 ;
        RECT 672.360 129.650 737.035 131.000 ;
      LAYER met3 ;
        RECT 669.645 129.100 673.140 129.250 ;
        RECT 669.645 129.000 670.610 129.100 ;
        RECT 670.610 128.800 671.820 129.000 ;
        RECT 671.960 128.800 673.140 129.100 ;
      LAYER met3 ;
        RECT 663.300 127.390 670.210 128.600 ;
      LAYER met3 ;
        RECT 670.610 127.920 673.140 128.800 ;
        RECT 670.610 127.790 671.820 127.920 ;
        RECT 671.840 127.790 673.140 127.920 ;
        RECT 671.820 127.600 673.140 127.790 ;
      LAYER met3 ;
        RECT 663.300 127.200 671.420 127.390 ;
        RECT 663.300 104.955 671.610 127.200 ;
      LAYER met3 ;
        RECT 672.010 105.355 673.140 127.600 ;
      LAYER met3 ;
        RECT 673.540 104.955 737.035 129.650 ;
        RECT 663.300 0.000 737.035 104.955 ;
        RECT 932.430 0.000 1011.690 201.310 ;
        RECT 1231.745 197.965 1242.620 198.000 ;
        RECT 1244.120 197.965 1255.000 198.000 ;
      LAYER met3 ;
        RECT 1050.000 164.765 1068.010 180.085 ;
        RECT 1070.000 164.765 1088.010 180.085 ;
        RECT 1090.000 164.765 1108.010 180.085 ;
        RECT 1110.000 164.765 1128.010 180.085 ;
        RECT 1130.000 164.765 1148.010 180.085 ;
        RECT 1150.000 164.765 1168.010 180.085 ;
      LAYER met3 ;
        RECT 1195.065 169.550 1204.800 174.200 ;
        RECT 1194.860 153.765 1205.395 158.415 ;
        RECT 1230.645 158.000 1256.100 197.965 ;
        RECT 1280.900 158.000 1281.000 197.965 ;
      LAYER met3 ;
        RECT 1319.000 164.765 1337.010 180.085 ;
        RECT 1339.000 164.765 1357.010 180.085 ;
        RECT 1359.000 164.765 1377.010 180.085 ;
        RECT 1379.000 164.765 1397.010 180.085 ;
        RECT 1399.000 164.765 1417.010 180.085 ;
        RECT 1419.000 164.765 1437.010 180.085 ;
      LAYER met3 ;
        RECT 1195.065 0.035 1204.800 24.250 ;
        RECT 1206.000 0.035 1281.000 158.000 ;
        RECT 1281.895 153.800 1291.975 158.450 ;
        RECT 1475.430 0.000 1554.690 201.310 ;
      LAYER met3 ;
        RECT 1593.000 164.765 1611.010 180.085 ;
        RECT 1613.000 164.765 1631.010 180.085 ;
        RECT 1633.000 164.765 1651.010 180.085 ;
        RECT 1653.000 164.765 1671.010 180.085 ;
        RECT 1673.000 164.765 1691.010 180.085 ;
        RECT 1693.000 164.765 1711.010 180.085 ;
      LAYER met3 ;
        RECT 1749.430 0.000 1828.690 201.310 ;
      LAYER met3 ;
        RECT 1867.000 164.765 1885.010 180.085 ;
        RECT 1887.000 164.765 1905.010 180.085 ;
        RECT 1907.000 164.765 1925.010 180.085 ;
        RECT 1927.000 164.765 1945.010 180.085 ;
        RECT 1947.000 164.765 1965.010 180.085 ;
        RECT 1967.000 164.765 1985.010 180.085 ;
      LAYER met3 ;
        RECT 2023.430 0.000 2102.690 201.310 ;
      LAYER met3 ;
        RECT 2141.000 164.765 2159.010 180.085 ;
        RECT 2161.000 164.765 2179.010 180.085 ;
        RECT 2181.000 164.765 2199.010 180.085 ;
        RECT 2201.000 164.765 2219.010 180.085 ;
        RECT 2221.000 164.765 2239.010 180.085 ;
        RECT 2241.000 164.765 2259.010 180.085 ;
      LAYER met3 ;
        RECT 2297.430 0.000 2376.690 201.310 ;
      LAYER met3 ;
        RECT 2415.000 164.765 2433.010 180.085 ;
        RECT 2435.000 164.765 2453.010 180.085 ;
        RECT 2455.000 164.765 2473.010 180.085 ;
        RECT 2475.000 164.765 2493.010 180.085 ;
        RECT 2495.000 164.765 2513.010 180.085 ;
        RECT 2515.000 164.765 2533.010 180.085 ;
      LAYER met3 ;
        RECT 2571.430 0.000 2650.690 201.310 ;
        RECT 2871.110 197.965 2882.110 200.000 ;
        RECT 2883.105 197.965 2894.105 200.000 ;
        RECT 3140.110 197.965 3151.110 200.000 ;
        RECT 3152.105 197.965 3163.105 200.000 ;
      LAYER met3 ;
        RECT 2689.000 164.765 2707.010 180.085 ;
        RECT 2709.000 164.765 2727.010 180.085 ;
        RECT 2729.000 164.765 2747.010 180.085 ;
        RECT 2749.000 164.765 2767.010 180.085 ;
        RECT 2769.000 164.765 2787.010 180.085 ;
        RECT 2789.000 164.765 2807.010 180.085 ;
      LAYER met3 ;
        RECT 2870.010 173.750 2895.205 197.965 ;
        RECT 3139.010 184.640 3164.205 197.965 ;
        RECT 2845.710 0.000 2919.760 173.750 ;
      LAYER met3 ;
        RECT 2958.000 164.765 2976.010 180.085 ;
        RECT 2978.000 164.765 2996.010 180.085 ;
        RECT 2998.000 164.765 3016.010 180.085 ;
        RECT 3018.000 164.765 3036.010 180.085 ;
        RECT 3038.000 164.765 3056.010 180.085 ;
        RECT 3058.000 164.765 3076.010 180.085 ;
      LAYER met3 ;
        RECT 3114.710 0.000 3188.760 184.640 ;
      LAYER met3 ;
        RECT 3227.000 164.765 3245.010 180.085 ;
        RECT 3247.000 164.765 3265.010 180.085 ;
        RECT 3267.000 164.765 3285.010 180.085 ;
        RECT 3287.000 164.765 3305.010 180.085 ;
        RECT 3307.000 164.765 3325.010 180.085 ;
        RECT 3327.000 164.765 3345.010 180.085 ;
      LAYER via3 ;
        RECT 238.230 175.875 255.720 179.885 ;
        RECT 238.260 164.935 255.910 167.885 ;
        RECT 258.230 175.875 275.720 179.885 ;
        RECT 258.260 164.935 275.910 167.885 ;
        RECT 278.230 175.875 295.720 179.885 ;
        RECT 278.260 164.935 295.910 167.885 ;
        RECT 298.230 175.875 315.720 179.885 ;
        RECT 298.260 164.935 315.910 167.885 ;
        RECT 318.230 175.875 335.720 179.885 ;
        RECT 318.260 164.935 335.910 167.885 ;
        RECT 338.230 175.875 355.720 179.885 ;
        RECT 338.260 164.935 355.910 167.885 ;
        RECT 507.230 175.875 524.720 179.885 ;
        RECT 507.260 164.935 524.910 167.885 ;
        RECT 527.230 175.875 544.720 179.885 ;
        RECT 527.260 164.935 544.910 167.885 ;
        RECT 547.230 175.875 564.720 179.885 ;
        RECT 547.260 164.935 564.910 167.885 ;
        RECT 567.230 175.875 584.720 179.885 ;
        RECT 567.260 164.935 584.910 167.885 ;
        RECT 587.230 175.875 604.720 179.885 ;
        RECT 587.260 164.935 604.910 167.885 ;
        RECT 607.230 175.875 624.720 179.885 ;
        RECT 607.260 164.935 624.910 167.885 ;
        RECT 776.230 175.875 793.720 179.885 ;
        RECT 776.260 164.935 793.910 167.885 ;
        RECT 796.230 175.875 813.720 179.885 ;
        RECT 796.260 164.935 813.910 167.885 ;
        RECT 816.230 175.875 833.720 179.885 ;
        RECT 816.260 164.935 833.910 167.885 ;
        RECT 836.230 175.875 853.720 179.885 ;
        RECT 836.260 164.935 853.910 167.885 ;
        RECT 856.230 175.875 873.720 179.885 ;
        RECT 856.260 164.935 873.910 167.885 ;
        RECT 876.230 175.875 893.720 179.885 ;
        RECT 876.260 164.935 893.910 167.885 ;
        RECT 1050.230 175.875 1067.720 179.885 ;
        RECT 1050.260 164.935 1067.910 167.885 ;
        RECT 1070.230 175.875 1087.720 179.885 ;
        RECT 1070.260 164.935 1087.910 167.885 ;
        RECT 1090.230 175.875 1107.720 179.885 ;
        RECT 1090.260 164.935 1107.910 167.885 ;
        RECT 1110.230 175.875 1127.720 179.885 ;
        RECT 1110.260 164.935 1127.910 167.885 ;
        RECT 1130.230 175.875 1147.720 179.885 ;
        RECT 1130.260 164.935 1147.910 167.885 ;
        RECT 1150.230 175.875 1167.720 179.885 ;
        RECT 1150.260 164.935 1167.910 167.885 ;
        RECT 1319.230 175.875 1336.720 179.885 ;
        RECT 1319.260 164.935 1336.910 167.885 ;
        RECT 1339.230 175.875 1356.720 179.885 ;
        RECT 1339.260 164.935 1356.910 167.885 ;
        RECT 1359.230 175.875 1376.720 179.885 ;
        RECT 1359.260 164.935 1376.910 167.885 ;
        RECT 1379.230 175.875 1396.720 179.885 ;
        RECT 1379.260 164.935 1396.910 167.885 ;
        RECT 1399.230 175.875 1416.720 179.885 ;
        RECT 1399.260 164.935 1416.910 167.885 ;
        RECT 1419.230 175.875 1436.720 179.885 ;
        RECT 1419.260 164.935 1436.910 167.885 ;
        RECT 1593.230 175.875 1610.720 179.885 ;
        RECT 1593.260 164.935 1610.910 167.885 ;
        RECT 1613.230 175.875 1630.720 179.885 ;
        RECT 1613.260 164.935 1630.910 167.885 ;
        RECT 1633.230 175.875 1650.720 179.885 ;
        RECT 1633.260 164.935 1650.910 167.885 ;
        RECT 1653.230 175.875 1670.720 179.885 ;
        RECT 1653.260 164.935 1670.910 167.885 ;
        RECT 1673.230 175.875 1690.720 179.885 ;
        RECT 1673.260 164.935 1690.910 167.885 ;
        RECT 1693.230 175.875 1710.720 179.885 ;
        RECT 1693.260 164.935 1710.910 167.885 ;
        RECT 1867.230 175.875 1884.720 179.885 ;
        RECT 1867.260 164.935 1884.910 167.885 ;
        RECT 1887.230 175.875 1904.720 179.885 ;
        RECT 1887.260 164.935 1904.910 167.885 ;
        RECT 1907.230 175.875 1924.720 179.885 ;
        RECT 1907.260 164.935 1924.910 167.885 ;
        RECT 1927.230 175.875 1944.720 179.885 ;
        RECT 1927.260 164.935 1944.910 167.885 ;
        RECT 1947.230 175.875 1964.720 179.885 ;
        RECT 1947.260 164.935 1964.910 167.885 ;
        RECT 1967.230 175.875 1984.720 179.885 ;
        RECT 1967.260 164.935 1984.910 167.885 ;
        RECT 2141.230 175.875 2158.720 179.885 ;
        RECT 2141.260 164.935 2158.910 167.885 ;
        RECT 2161.230 175.875 2178.720 179.885 ;
        RECT 2161.260 164.935 2178.910 167.885 ;
        RECT 2181.230 175.875 2198.720 179.885 ;
        RECT 2181.260 164.935 2198.910 167.885 ;
        RECT 2201.230 175.875 2218.720 179.885 ;
        RECT 2201.260 164.935 2218.910 167.885 ;
        RECT 2221.230 175.875 2238.720 179.885 ;
        RECT 2221.260 164.935 2238.910 167.885 ;
        RECT 2241.230 175.875 2258.720 179.885 ;
        RECT 2241.260 164.935 2258.910 167.885 ;
        RECT 2415.230 175.875 2432.720 179.885 ;
        RECT 2415.260 164.935 2432.910 167.885 ;
        RECT 2435.230 175.875 2452.720 179.885 ;
        RECT 2435.260 164.935 2452.910 167.885 ;
        RECT 2455.230 175.875 2472.720 179.885 ;
        RECT 2455.260 164.935 2472.910 167.885 ;
        RECT 2475.230 175.875 2492.720 179.885 ;
        RECT 2475.260 164.935 2492.910 167.885 ;
        RECT 2495.230 175.875 2512.720 179.885 ;
        RECT 2495.260 164.935 2512.910 167.885 ;
        RECT 2515.230 175.875 2532.720 179.885 ;
        RECT 2515.260 164.935 2532.910 167.885 ;
        RECT 2689.230 175.875 2706.720 179.885 ;
        RECT 2689.260 164.935 2706.910 167.885 ;
        RECT 2709.230 175.875 2726.720 179.885 ;
        RECT 2709.260 164.935 2726.910 167.885 ;
        RECT 2729.230 175.875 2746.720 179.885 ;
        RECT 2729.260 164.935 2746.910 167.885 ;
        RECT 2749.230 175.875 2766.720 179.885 ;
        RECT 2749.260 164.935 2766.910 167.885 ;
        RECT 2769.230 175.875 2786.720 179.885 ;
        RECT 2769.260 164.935 2786.910 167.885 ;
        RECT 2789.230 175.875 2806.720 179.885 ;
        RECT 2958.230 175.875 2975.720 179.885 ;
        RECT 2789.260 164.935 2806.910 167.885 ;
        RECT 2958.260 164.935 2975.910 167.885 ;
        RECT 2978.230 175.875 2995.720 179.885 ;
        RECT 2978.260 164.935 2995.910 167.885 ;
        RECT 2998.230 175.875 3015.720 179.885 ;
        RECT 2998.260 164.935 3015.910 167.885 ;
        RECT 3018.230 175.875 3035.720 179.885 ;
        RECT 3018.260 164.935 3035.910 167.885 ;
        RECT 3038.230 175.875 3055.720 179.885 ;
        RECT 3038.260 164.935 3055.910 167.885 ;
        RECT 3058.230 175.875 3075.720 179.885 ;
        RECT 3058.260 164.935 3075.910 167.885 ;
        RECT 3227.230 175.875 3244.720 179.885 ;
        RECT 3227.260 164.935 3244.910 167.885 ;
        RECT 3247.230 175.875 3264.720 179.885 ;
        RECT 3247.260 164.935 3264.910 167.885 ;
        RECT 3267.230 175.875 3284.720 179.885 ;
        RECT 3267.260 164.935 3284.910 167.885 ;
        RECT 3287.230 175.875 3304.720 179.885 ;
        RECT 3287.260 164.935 3304.910 167.885 ;
        RECT 3307.230 175.875 3324.720 179.885 ;
        RECT 3307.260 164.935 3324.910 167.885 ;
        RECT 3327.230 175.875 3344.720 179.885 ;
        RECT 3327.260 164.935 3344.910 167.885 ;
      LAYER met4 ;
        RECT 0.000 5163.385 202.330 5188.000 ;
      LAYER met4 ;
        RECT 202.730 5163.785 204.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5083.400 202.745 5163.385 ;
        RECT 204.000 5162.035 381.000 5188.000 ;
      LAYER met4 ;
        RECT 381.000 5163.785 382.270 5188.000 ;
      LAYER met4 ;
        RECT 382.670 5163.385 459.330 5188.000 ;
      LAYER met4 ;
        RECT 459.730 5163.785 461.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5057.635 201.745 5083.400 ;
        RECT 204.000 5083.000 381.000 5085.035 ;
        RECT 381.965 5083.400 459.970 5163.385 ;
        RECT 461.000 5162.035 638.000 5188.000 ;
      LAYER met4 ;
        RECT 638.000 5163.785 639.270 5188.000 ;
      LAYER met4 ;
        RECT 639.670 5163.385 716.330 5188.000 ;
      LAYER met4 ;
        RECT 716.730 5163.785 718.000 5188.000 ;
        RECT 202.145 5058.035 205.000 5083.000 ;
      LAYER met4 ;
        RECT 205.000 5058.035 223.000 5083.000 ;
      LAYER met4 ;
        RECT 223.000 5058.035 225.000 5083.000 ;
      LAYER met4 ;
        RECT 225.000 5058.035 243.000 5083.000 ;
      LAYER met4 ;
        RECT 243.000 5058.035 245.000 5083.000 ;
      LAYER met4 ;
        RECT 245.000 5058.035 263.000 5083.000 ;
      LAYER met4 ;
        RECT 263.000 5058.035 265.000 5083.000 ;
      LAYER met4 ;
        RECT 265.000 5058.035 283.000 5083.000 ;
      LAYER met4 ;
        RECT 283.000 5058.035 285.000 5083.000 ;
      LAYER met4 ;
        RECT 285.000 5058.035 303.000 5083.000 ;
      LAYER met4 ;
        RECT 303.000 5058.035 305.000 5083.000 ;
      LAYER met4 ;
        RECT 305.000 5058.035 323.000 5083.000 ;
      LAYER met4 ;
        RECT 323.000 5058.035 325.000 5083.000 ;
      LAYER met4 ;
        RECT 325.000 5058.035 343.000 5083.000 ;
      LAYER met4 ;
        RECT 343.000 5058.035 345.000 5083.000 ;
      LAYER met4 ;
        RECT 345.000 5058.035 363.000 5083.000 ;
      LAYER met4 ;
        RECT 363.000 5058.035 365.000 5083.000 ;
      LAYER met4 ;
        RECT 365.000 5058.035 373.000 5083.000 ;
      LAYER met4 ;
        RECT 373.000 5058.035 375.000 5083.000 ;
      LAYER met4 ;
        RECT 375.000 5058.035 378.000 5083.000 ;
      LAYER met4 ;
        RECT 378.000 5058.035 382.270 5083.000 ;
      LAYER met4 ;
        RECT 0.000 5056.935 202.745 5057.635 ;
        RECT 204.000 5056.935 381.000 5058.035 ;
        RECT 382.670 5057.635 459.330 5083.400 ;
        RECT 461.000 5083.000 638.000 5085.035 ;
        RECT 638.965 5083.400 716.970 5163.385 ;
        RECT 718.000 5162.035 895.000 5188.000 ;
      LAYER met4 ;
        RECT 895.000 5163.785 896.270 5188.000 ;
      LAYER met4 ;
        RECT 896.670 5163.385 973.330 5188.000 ;
      LAYER met4 ;
        RECT 973.730 5163.785 975.000 5188.000 ;
        RECT 459.730 5058.035 462.000 5083.000 ;
      LAYER met4 ;
        RECT 462.000 5058.035 480.000 5083.000 ;
      LAYER met4 ;
        RECT 480.000 5058.035 482.000 5083.000 ;
      LAYER met4 ;
        RECT 482.000 5058.035 500.000 5083.000 ;
      LAYER met4 ;
        RECT 500.000 5058.035 502.000 5083.000 ;
      LAYER met4 ;
        RECT 502.000 5058.035 520.000 5083.000 ;
      LAYER met4 ;
        RECT 520.000 5058.035 522.000 5083.000 ;
      LAYER met4 ;
        RECT 522.000 5058.035 540.000 5083.000 ;
      LAYER met4 ;
        RECT 540.000 5058.035 542.000 5083.000 ;
      LAYER met4 ;
        RECT 542.000 5058.035 560.000 5083.000 ;
      LAYER met4 ;
        RECT 560.000 5058.035 562.000 5083.000 ;
      LAYER met4 ;
        RECT 562.000 5058.035 580.000 5083.000 ;
      LAYER met4 ;
        RECT 580.000 5058.035 582.000 5083.000 ;
      LAYER met4 ;
        RECT 582.000 5058.035 600.000 5083.000 ;
      LAYER met4 ;
        RECT 600.000 5058.035 602.000 5083.000 ;
      LAYER met4 ;
        RECT 602.000 5058.035 620.000 5083.000 ;
      LAYER met4 ;
        RECT 620.000 5058.035 622.000 5083.000 ;
      LAYER met4 ;
        RECT 622.000 5058.035 630.000 5083.000 ;
      LAYER met4 ;
        RECT 630.000 5058.035 632.000 5083.000 ;
      LAYER met4 ;
        RECT 632.000 5058.035 635.000 5083.000 ;
      LAYER met4 ;
        RECT 635.000 5058.035 639.270 5083.000 ;
      LAYER met4 ;
        RECT 381.965 5056.935 459.970 5057.635 ;
        RECT 461.000 5056.935 638.000 5058.035 ;
        RECT 639.670 5057.635 716.330 5083.400 ;
        RECT 718.000 5083.000 895.000 5085.035 ;
        RECT 895.965 5083.400 973.970 5163.385 ;
        RECT 975.000 5162.035 1152.000 5188.000 ;
      LAYER met4 ;
        RECT 1152.000 5163.785 1153.270 5188.000 ;
      LAYER met4 ;
        RECT 1153.670 5163.385 1230.330 5188.000 ;
      LAYER met4 ;
        RECT 1230.730 5163.785 1232.000 5188.000 ;
        RECT 716.730 5058.035 719.000 5083.000 ;
      LAYER met4 ;
        RECT 719.000 5058.035 737.000 5083.000 ;
      LAYER met4 ;
        RECT 737.000 5058.035 739.000 5083.000 ;
      LAYER met4 ;
        RECT 739.000 5058.035 757.000 5083.000 ;
      LAYER met4 ;
        RECT 757.000 5058.035 759.000 5083.000 ;
      LAYER met4 ;
        RECT 759.000 5058.035 777.000 5083.000 ;
      LAYER met4 ;
        RECT 777.000 5058.035 779.000 5083.000 ;
      LAYER met4 ;
        RECT 779.000 5058.035 797.000 5083.000 ;
      LAYER met4 ;
        RECT 797.000 5058.035 799.000 5083.000 ;
      LAYER met4 ;
        RECT 799.000 5058.035 817.000 5083.000 ;
      LAYER met4 ;
        RECT 817.000 5058.035 819.000 5083.000 ;
      LAYER met4 ;
        RECT 819.000 5058.035 837.000 5083.000 ;
      LAYER met4 ;
        RECT 837.000 5058.035 839.000 5083.000 ;
      LAYER met4 ;
        RECT 839.000 5058.035 857.000 5083.000 ;
      LAYER met4 ;
        RECT 857.000 5058.035 859.000 5083.000 ;
      LAYER met4 ;
        RECT 859.000 5058.035 877.000 5083.000 ;
      LAYER met4 ;
        RECT 877.000 5058.035 879.000 5083.000 ;
      LAYER met4 ;
        RECT 879.000 5058.035 887.000 5083.000 ;
      LAYER met4 ;
        RECT 887.000 5058.035 889.000 5083.000 ;
      LAYER met4 ;
        RECT 889.000 5058.035 892.000 5083.000 ;
      LAYER met4 ;
        RECT 892.000 5058.035 896.270 5083.000 ;
      LAYER met4 ;
        RECT 638.965 5056.935 716.970 5057.635 ;
        RECT 718.000 5056.935 895.000 5058.035 ;
        RECT 896.670 5057.635 973.330 5083.400 ;
        RECT 975.000 5083.000 1152.000 5085.035 ;
        RECT 1152.965 5083.400 1230.970 5163.385 ;
        RECT 1232.000 5162.035 1410.000 5188.000 ;
      LAYER met4 ;
        RECT 1410.000 5163.785 1411.270 5188.000 ;
      LAYER met4 ;
        RECT 1411.670 5163.385 1488.330 5188.000 ;
      LAYER met4 ;
        RECT 1488.730 5163.785 1490.000 5188.000 ;
        RECT 973.730 5058.035 976.000 5083.000 ;
      LAYER met4 ;
        RECT 976.000 5058.035 994.000 5083.000 ;
      LAYER met4 ;
        RECT 994.000 5058.035 996.000 5083.000 ;
      LAYER met4 ;
        RECT 996.000 5058.035 1014.000 5083.000 ;
      LAYER met4 ;
        RECT 1014.000 5058.035 1016.000 5083.000 ;
      LAYER met4 ;
        RECT 1016.000 5058.035 1034.000 5083.000 ;
      LAYER met4 ;
        RECT 1034.000 5058.035 1036.000 5083.000 ;
      LAYER met4 ;
        RECT 1036.000 5058.035 1054.000 5083.000 ;
      LAYER met4 ;
        RECT 1054.000 5058.035 1056.000 5083.000 ;
      LAYER met4 ;
        RECT 1056.000 5058.035 1074.000 5083.000 ;
      LAYER met4 ;
        RECT 1074.000 5058.035 1076.000 5083.000 ;
      LAYER met4 ;
        RECT 1076.000 5058.035 1094.000 5083.000 ;
      LAYER met4 ;
        RECT 1094.000 5058.035 1096.000 5083.000 ;
      LAYER met4 ;
        RECT 1096.000 5058.035 1114.000 5083.000 ;
      LAYER met4 ;
        RECT 1114.000 5058.035 1116.000 5083.000 ;
      LAYER met4 ;
        RECT 1116.000 5058.035 1134.000 5083.000 ;
      LAYER met4 ;
        RECT 1134.000 5058.035 1136.000 5083.000 ;
      LAYER met4 ;
        RECT 1136.000 5058.035 1144.000 5083.000 ;
      LAYER met4 ;
        RECT 1144.000 5058.035 1146.000 5083.000 ;
      LAYER met4 ;
        RECT 1146.000 5058.035 1149.000 5083.000 ;
      LAYER met4 ;
        RECT 1149.000 5058.035 1153.270 5083.000 ;
      LAYER met4 ;
        RECT 895.965 5056.935 973.970 5057.635 ;
        RECT 975.000 5056.935 1152.000 5058.035 ;
        RECT 1153.670 5057.635 1230.330 5083.400 ;
        RECT 1232.000 5083.000 1410.000 5085.035 ;
        RECT 1410.965 5083.400 1488.970 5163.385 ;
        RECT 1490.000 5162.035 1667.000 5188.000 ;
        RECT 1668.670 5163.385 1740.330 5188.000 ;
      LAYER met4 ;
        RECT 1230.730 5058.035 1233.000 5083.000 ;
      LAYER met4 ;
        RECT 1233.000 5058.035 1251.000 5083.000 ;
      LAYER met4 ;
        RECT 1251.000 5058.035 1253.000 5083.000 ;
      LAYER met4 ;
        RECT 1253.000 5058.035 1271.000 5083.000 ;
      LAYER met4 ;
        RECT 1271.000 5058.035 1273.000 5083.000 ;
      LAYER met4 ;
        RECT 1273.000 5058.035 1291.000 5083.000 ;
      LAYER met4 ;
        RECT 1291.000 5058.035 1293.000 5083.000 ;
      LAYER met4 ;
        RECT 1293.000 5058.035 1311.000 5083.000 ;
      LAYER met4 ;
        RECT 1311.000 5058.035 1313.000 5083.000 ;
      LAYER met4 ;
        RECT 1313.000 5058.035 1331.000 5083.000 ;
      LAYER met4 ;
        RECT 1331.000 5058.035 1333.000 5083.000 ;
      LAYER met4 ;
        RECT 1333.000 5058.035 1351.000 5083.000 ;
      LAYER met4 ;
        RECT 1351.000 5058.035 1353.000 5083.000 ;
      LAYER met4 ;
        RECT 1353.000 5058.035 1371.000 5083.000 ;
      LAYER met4 ;
        RECT 1371.000 5058.035 1373.000 5083.000 ;
      LAYER met4 ;
        RECT 1373.000 5058.035 1391.000 5083.000 ;
      LAYER met4 ;
        RECT 1391.000 5058.035 1393.000 5083.000 ;
      LAYER met4 ;
        RECT 1393.000 5058.035 1401.000 5083.000 ;
      LAYER met4 ;
        RECT 1401.000 5058.035 1403.000 5083.000 ;
      LAYER met4 ;
        RECT 1403.000 5058.035 1406.000 5083.000 ;
      LAYER met4 ;
        RECT 1406.000 5058.035 1411.270 5083.000 ;
      LAYER met4 ;
        RECT 1152.965 5056.935 1230.970 5057.635 ;
        RECT 1232.000 5056.935 1410.000 5058.035 ;
        RECT 1411.670 5057.635 1488.330 5083.400 ;
        RECT 1490.000 5083.000 1667.000 5085.035 ;
        RECT 1667.965 5083.400 1741.035 5163.385 ;
        RECT 1742.000 5162.035 1919.000 5188.000 ;
      LAYER met4 ;
        RECT 1919.000 5163.785 1920.270 5188.000 ;
      LAYER met4 ;
        RECT 1920.670 5163.385 1997.330 5188.000 ;
      LAYER met4 ;
        RECT 1997.730 5163.785 1999.000 5188.000 ;
      LAYER met4 ;
        RECT 1999.000 5163.785 2364.000 5188.000 ;
      LAYER met4 ;
        RECT 2364.000 5163.785 2365.270 5188.000 ;
        RECT 1488.730 5058.035 1491.000 5083.000 ;
      LAYER met4 ;
        RECT 1491.000 5058.035 1509.000 5083.000 ;
      LAYER met4 ;
        RECT 1509.000 5058.035 1511.000 5083.000 ;
      LAYER met4 ;
        RECT 1511.000 5058.035 1529.000 5083.000 ;
      LAYER met4 ;
        RECT 1529.000 5058.035 1531.000 5083.000 ;
      LAYER met4 ;
        RECT 1531.000 5058.035 1549.000 5083.000 ;
      LAYER met4 ;
        RECT 1549.000 5058.035 1551.000 5083.000 ;
      LAYER met4 ;
        RECT 1551.000 5058.035 1569.000 5083.000 ;
      LAYER met4 ;
        RECT 1569.000 5058.035 1571.000 5083.000 ;
      LAYER met4 ;
        RECT 1571.000 5058.035 1589.000 5083.000 ;
      LAYER met4 ;
        RECT 1589.000 5058.035 1591.000 5083.000 ;
      LAYER met4 ;
        RECT 1591.000 5058.035 1609.000 5083.000 ;
      LAYER met4 ;
        RECT 1609.000 5058.035 1611.000 5083.000 ;
      LAYER met4 ;
        RECT 1611.000 5058.035 1629.000 5083.000 ;
      LAYER met4 ;
        RECT 1629.000 5058.035 1631.000 5083.000 ;
      LAYER met4 ;
        RECT 1631.000 5058.035 1649.000 5083.000 ;
      LAYER met4 ;
        RECT 1649.000 5058.035 1651.000 5083.000 ;
      LAYER met4 ;
        RECT 1651.000 5058.035 1659.000 5083.000 ;
      LAYER met4 ;
        RECT 1659.000 5058.035 1661.000 5083.000 ;
      LAYER met4 ;
        RECT 1661.000 5058.035 1664.000 5083.000 ;
      LAYER met4 ;
        RECT 1664.000 5058.035 1668.270 5083.000 ;
      LAYER met4 ;
        RECT 1410.965 5056.935 1488.970 5057.635 ;
        RECT 1490.000 5056.935 1667.000 5058.035 ;
        RECT 1668.670 5057.635 1740.330 5083.400 ;
        RECT 1742.000 5083.000 1919.000 5085.035 ;
        RECT 1919.965 5083.400 1997.970 5163.385 ;
        RECT 1999.000 5162.035 2176.000 5163.785 ;
        RECT 2186.000 5162.035 2364.000 5163.785 ;
        RECT 2365.670 5163.385 2442.330 5188.000 ;
      LAYER met4 ;
        RECT 2442.730 5163.785 2444.000 5188.000 ;
        RECT 1740.730 5058.035 1743.000 5083.000 ;
      LAYER met4 ;
        RECT 1743.000 5058.035 1761.000 5083.000 ;
      LAYER met4 ;
        RECT 1761.000 5058.035 1763.000 5083.000 ;
      LAYER met4 ;
        RECT 1763.000 5058.035 1781.000 5083.000 ;
      LAYER met4 ;
        RECT 1781.000 5058.035 1783.000 5083.000 ;
      LAYER met4 ;
        RECT 1783.000 5058.035 1801.000 5083.000 ;
      LAYER met4 ;
        RECT 1801.000 5058.035 1803.000 5083.000 ;
      LAYER met4 ;
        RECT 1803.000 5058.035 1821.000 5083.000 ;
      LAYER met4 ;
        RECT 1821.000 5058.035 1823.000 5083.000 ;
      LAYER met4 ;
        RECT 1823.000 5058.035 1841.000 5083.000 ;
      LAYER met4 ;
        RECT 1841.000 5058.035 1843.000 5083.000 ;
      LAYER met4 ;
        RECT 1843.000 5058.035 1861.000 5083.000 ;
      LAYER met4 ;
        RECT 1861.000 5058.035 1863.000 5083.000 ;
      LAYER met4 ;
        RECT 1863.000 5058.035 1881.000 5083.000 ;
      LAYER met4 ;
        RECT 1881.000 5058.035 1883.000 5083.000 ;
      LAYER met4 ;
        RECT 1883.000 5058.035 1901.000 5083.000 ;
      LAYER met4 ;
        RECT 1901.000 5058.035 1903.000 5083.000 ;
      LAYER met4 ;
        RECT 1903.000 5058.035 1911.000 5083.000 ;
      LAYER met4 ;
        RECT 1911.000 5058.035 1913.000 5083.000 ;
      LAYER met4 ;
        RECT 1913.000 5058.035 1916.000 5083.000 ;
      LAYER met4 ;
        RECT 1916.000 5058.035 1920.270 5083.000 ;
      LAYER met4 ;
        RECT 1667.965 5056.935 1741.035 5057.635 ;
        RECT 1742.000 5056.935 1919.000 5058.035 ;
        RECT 1920.670 5057.635 1997.330 5083.400 ;
        RECT 1999.000 5083.000 2176.000 5085.035 ;
        RECT 2186.000 5083.000 2364.000 5085.035 ;
        RECT 2364.965 5083.400 2442.970 5163.385 ;
        RECT 2444.000 5162.035 2621.000 5188.000 ;
      LAYER met4 ;
        RECT 2621.000 5163.785 2622.270 5188.000 ;
      LAYER met4 ;
        RECT 2622.670 5163.385 2699.330 5188.000 ;
      LAYER met4 ;
        RECT 2699.730 5163.785 2701.000 5188.000 ;
        RECT 1997.730 5058.035 2000.000 5083.000 ;
      LAYER met4 ;
        RECT 2000.000 5058.035 2018.000 5083.000 ;
      LAYER met4 ;
        RECT 2018.000 5058.035 2020.000 5083.000 ;
      LAYER met4 ;
        RECT 2020.000 5058.035 2038.000 5083.000 ;
      LAYER met4 ;
        RECT 2038.000 5058.035 2040.000 5083.000 ;
      LAYER met4 ;
        RECT 2040.000 5058.035 2058.000 5083.000 ;
      LAYER met4 ;
        RECT 2058.000 5058.035 2060.000 5083.000 ;
      LAYER met4 ;
        RECT 2060.000 5058.035 2078.000 5083.000 ;
      LAYER met4 ;
        RECT 2078.000 5058.035 2080.000 5083.000 ;
      LAYER met4 ;
        RECT 2080.000 5058.035 2098.000 5083.000 ;
      LAYER met4 ;
        RECT 2098.000 5058.035 2100.000 5083.000 ;
      LAYER met4 ;
        RECT 2100.000 5058.035 2118.000 5083.000 ;
      LAYER met4 ;
        RECT 2118.000 5058.035 2120.000 5083.000 ;
      LAYER met4 ;
        RECT 2120.000 5058.035 2138.000 5083.000 ;
      LAYER met4 ;
        RECT 2138.000 5058.035 2140.000 5083.000 ;
      LAYER met4 ;
        RECT 2140.000 5058.035 2158.000 5083.000 ;
      LAYER met4 ;
        RECT 2158.000 5058.035 2160.000 5083.000 ;
      LAYER met4 ;
        RECT 2160.000 5058.035 2168.000 5083.000 ;
      LAYER met4 ;
        RECT 2168.000 5058.035 2170.000 5083.000 ;
      LAYER met4 ;
        RECT 2170.000 5058.035 2173.000 5083.000 ;
      LAYER met4 ;
        RECT 2173.000 5058.035 2187.000 5083.000 ;
      LAYER met4 ;
        RECT 2187.000 5058.035 2205.000 5083.000 ;
      LAYER met4 ;
        RECT 2205.000 5058.035 2207.000 5083.000 ;
      LAYER met4 ;
        RECT 2207.000 5058.035 2225.000 5083.000 ;
      LAYER met4 ;
        RECT 2225.000 5058.035 2227.000 5083.000 ;
      LAYER met4 ;
        RECT 2227.000 5058.035 2245.000 5083.000 ;
      LAYER met4 ;
        RECT 2245.000 5058.035 2247.000 5083.000 ;
      LAYER met4 ;
        RECT 2247.000 5058.035 2265.000 5083.000 ;
      LAYER met4 ;
        RECT 2265.000 5058.035 2267.000 5083.000 ;
      LAYER met4 ;
        RECT 2267.000 5058.035 2285.000 5083.000 ;
      LAYER met4 ;
        RECT 2285.000 5058.035 2287.000 5083.000 ;
      LAYER met4 ;
        RECT 2287.000 5058.035 2305.000 5083.000 ;
      LAYER met4 ;
        RECT 2305.000 5058.035 2307.000 5083.000 ;
      LAYER met4 ;
        RECT 2307.000 5058.035 2325.000 5083.000 ;
      LAYER met4 ;
        RECT 2325.000 5058.035 2327.000 5083.000 ;
      LAYER met4 ;
        RECT 2327.000 5058.035 2345.000 5083.000 ;
      LAYER met4 ;
        RECT 2345.000 5058.035 2347.000 5083.000 ;
      LAYER met4 ;
        RECT 2347.000 5058.035 2355.000 5083.000 ;
      LAYER met4 ;
        RECT 2355.000 5058.035 2357.000 5083.000 ;
      LAYER met4 ;
        RECT 2357.000 5058.035 2360.000 5083.000 ;
      LAYER met4 ;
        RECT 2360.000 5058.035 2365.270 5083.000 ;
      LAYER met4 ;
        RECT 1919.965 5056.935 1997.970 5057.635 ;
        RECT 1999.000 5056.935 2176.000 5058.035 ;
        RECT 2186.000 5056.935 2364.000 5058.035 ;
        RECT 2365.670 5057.635 2442.330 5083.400 ;
        RECT 2444.000 5083.000 2621.000 5085.035 ;
        RECT 2621.965 5083.400 2699.970 5163.385 ;
        RECT 2701.000 5162.035 2878.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.000 5163.785 2879.270 5188.000 ;
      LAYER met4 ;
        RECT 2879.670 5163.385 2951.330 5188.000 ;
      LAYER met4 ;
        RECT 2951.730 5163.785 2953.000 5188.000 ;
        RECT 2442.730 5058.035 2445.000 5083.000 ;
      LAYER met4 ;
        RECT 2445.000 5058.035 2463.000 5083.000 ;
      LAYER met4 ;
        RECT 2463.000 5058.035 2465.000 5083.000 ;
      LAYER met4 ;
        RECT 2465.000 5058.035 2483.000 5083.000 ;
      LAYER met4 ;
        RECT 2483.000 5058.035 2485.000 5083.000 ;
      LAYER met4 ;
        RECT 2485.000 5058.035 2503.000 5083.000 ;
      LAYER met4 ;
        RECT 2503.000 5058.035 2505.000 5083.000 ;
      LAYER met4 ;
        RECT 2505.000 5058.035 2523.000 5083.000 ;
      LAYER met4 ;
        RECT 2523.000 5058.035 2525.000 5083.000 ;
      LAYER met4 ;
        RECT 2525.000 5058.035 2543.000 5083.000 ;
      LAYER met4 ;
        RECT 2543.000 5058.035 2545.000 5083.000 ;
      LAYER met4 ;
        RECT 2545.000 5058.035 2563.000 5083.000 ;
      LAYER met4 ;
        RECT 2563.000 5058.035 2565.000 5083.000 ;
      LAYER met4 ;
        RECT 2565.000 5058.035 2583.000 5083.000 ;
      LAYER met4 ;
        RECT 2583.000 5058.035 2585.000 5083.000 ;
      LAYER met4 ;
        RECT 2585.000 5058.035 2603.000 5083.000 ;
      LAYER met4 ;
        RECT 2603.000 5058.035 2605.000 5083.000 ;
      LAYER met4 ;
        RECT 2605.000 5058.035 2613.000 5083.000 ;
      LAYER met4 ;
        RECT 2613.000 5058.035 2615.000 5083.000 ;
      LAYER met4 ;
        RECT 2615.000 5058.035 2618.000 5083.000 ;
      LAYER met4 ;
        RECT 2618.000 5058.035 2622.270 5083.000 ;
      LAYER met4 ;
        RECT 2364.965 5056.935 2442.970 5057.635 ;
        RECT 2444.000 5056.935 2621.000 5058.035 ;
        RECT 2622.670 5057.635 2699.330 5083.400 ;
        RECT 2701.000 5083.000 2878.000 5085.035 ;
        RECT 2878.965 5083.400 2952.035 5163.385 ;
        RECT 2953.000 5162.035 3130.000 5188.000 ;
      LAYER met4 ;
        RECT 3130.000 5163.785 3131.270 5188.000 ;
      LAYER met4 ;
        RECT 3131.670 5163.385 3208.330 5188.000 ;
      LAYER met4 ;
        RECT 3208.730 5163.785 3210.000 5188.000 ;
      LAYER met4 ;
        RECT 3210.000 5163.385 3388.000 5188.000 ;
      LAYER met4 ;
        RECT 3388.000 5163.785 3389.435 5188.000 ;
      LAYER met4 ;
        RECT 3389.835 5163.385 3588.000 5188.000 ;
      LAYER met4 ;
        RECT 2699.730 5058.035 2702.000 5083.000 ;
      LAYER met4 ;
        RECT 2702.000 5058.035 2720.000 5083.000 ;
      LAYER met4 ;
        RECT 2720.000 5058.035 2722.000 5083.000 ;
      LAYER met4 ;
        RECT 2722.000 5058.035 2740.000 5083.000 ;
      LAYER met4 ;
        RECT 2740.000 5058.035 2742.000 5083.000 ;
      LAYER met4 ;
        RECT 2742.000 5058.035 2760.000 5083.000 ;
      LAYER met4 ;
        RECT 2760.000 5058.035 2762.000 5083.000 ;
      LAYER met4 ;
        RECT 2762.000 5058.035 2780.000 5083.000 ;
      LAYER met4 ;
        RECT 2780.000 5058.035 2782.000 5083.000 ;
      LAYER met4 ;
        RECT 2782.000 5058.035 2800.000 5083.000 ;
      LAYER met4 ;
        RECT 2800.000 5058.035 2802.000 5083.000 ;
      LAYER met4 ;
        RECT 2802.000 5058.035 2820.000 5083.000 ;
      LAYER met4 ;
        RECT 2820.000 5058.035 2822.000 5083.000 ;
      LAYER met4 ;
        RECT 2822.000 5058.035 2840.000 5083.000 ;
      LAYER met4 ;
        RECT 2840.000 5058.035 2842.000 5083.000 ;
      LAYER met4 ;
        RECT 2842.000 5058.035 2860.000 5083.000 ;
      LAYER met4 ;
        RECT 2860.000 5058.035 2862.000 5083.000 ;
      LAYER met4 ;
        RECT 2862.000 5058.035 2870.000 5083.000 ;
      LAYER met4 ;
        RECT 2870.000 5058.035 2872.000 5083.000 ;
      LAYER met4 ;
        RECT 2872.000 5058.035 2875.000 5083.000 ;
      LAYER met4 ;
        RECT 2875.000 5058.035 2879.270 5083.000 ;
      LAYER met4 ;
        RECT 2621.965 5056.935 2699.970 5057.635 ;
        RECT 2701.000 5056.935 2878.000 5058.035 ;
        RECT 2879.670 5057.635 2951.330 5083.400 ;
        RECT 2953.000 5083.000 3130.000 5085.035 ;
        RECT 3130.965 5083.400 3208.970 5163.385 ;
        RECT 3210.000 5162.035 3588.000 5163.385 ;
        RECT 3388.000 5085.035 3588.000 5162.035 ;
        RECT 3210.000 5083.400 3588.000 5085.035 ;
      LAYER met4 ;
        RECT 2951.730 5058.035 2954.000 5083.000 ;
      LAYER met4 ;
        RECT 2954.000 5058.035 2972.000 5083.000 ;
      LAYER met4 ;
        RECT 2972.000 5058.035 2974.000 5083.000 ;
      LAYER met4 ;
        RECT 2974.000 5058.035 2992.000 5083.000 ;
      LAYER met4 ;
        RECT 2992.000 5058.035 2994.000 5083.000 ;
      LAYER met4 ;
        RECT 2994.000 5058.035 3012.000 5083.000 ;
      LAYER met4 ;
        RECT 3012.000 5058.035 3014.000 5083.000 ;
      LAYER met4 ;
        RECT 3014.000 5058.035 3032.000 5083.000 ;
      LAYER met4 ;
        RECT 3032.000 5058.035 3034.000 5083.000 ;
      LAYER met4 ;
        RECT 3034.000 5058.035 3052.000 5083.000 ;
      LAYER met4 ;
        RECT 3052.000 5058.035 3054.000 5083.000 ;
      LAYER met4 ;
        RECT 3054.000 5058.035 3072.000 5083.000 ;
      LAYER met4 ;
        RECT 3072.000 5058.035 3074.000 5083.000 ;
      LAYER met4 ;
        RECT 3074.000 5058.035 3092.000 5083.000 ;
      LAYER met4 ;
        RECT 3092.000 5058.035 3094.000 5083.000 ;
      LAYER met4 ;
        RECT 3094.000 5058.035 3112.000 5083.000 ;
      LAYER met4 ;
        RECT 3112.000 5058.035 3114.000 5083.000 ;
      LAYER met4 ;
        RECT 3114.000 5058.035 3122.000 5083.000 ;
      LAYER met4 ;
        RECT 3122.000 5058.035 3124.000 5083.000 ;
      LAYER met4 ;
        RECT 3124.000 5058.035 3127.000 5083.000 ;
      LAYER met4 ;
        RECT 3127.000 5058.035 3131.270 5083.000 ;
      LAYER met4 ;
        RECT 2878.965 5056.935 2952.035 5057.635 ;
        RECT 2953.000 5056.935 3130.000 5058.035 ;
        RECT 3131.670 5057.635 3208.330 5083.400 ;
        RECT 3210.000 5083.000 3388.000 5083.400 ;
      LAYER met4 ;
        RECT 3208.730 5058.035 3211.000 5083.000 ;
      LAYER met4 ;
        RECT 3211.000 5058.035 3229.000 5083.000 ;
      LAYER met4 ;
        RECT 3229.000 5058.035 3231.000 5083.000 ;
      LAYER met4 ;
        RECT 3231.000 5058.035 3249.000 5083.000 ;
      LAYER met4 ;
        RECT 3249.000 5058.035 3251.000 5083.000 ;
      LAYER met4 ;
        RECT 3251.000 5058.035 3269.000 5083.000 ;
      LAYER met4 ;
        RECT 3269.000 5058.035 3271.000 5083.000 ;
      LAYER met4 ;
        RECT 3271.000 5058.035 3289.000 5083.000 ;
      LAYER met4 ;
        RECT 3289.000 5058.035 3291.000 5083.000 ;
      LAYER met4 ;
        RECT 3291.000 5058.035 3309.000 5083.000 ;
      LAYER met4 ;
        RECT 3309.000 5058.035 3311.000 5083.000 ;
      LAYER met4 ;
        RECT 3311.000 5058.035 3329.000 5083.000 ;
      LAYER met4 ;
        RECT 3329.000 5058.035 3331.000 5083.000 ;
      LAYER met4 ;
        RECT 3331.000 5058.035 3349.000 5083.000 ;
      LAYER met4 ;
        RECT 3349.000 5058.035 3351.000 5083.000 ;
      LAYER met4 ;
        RECT 3351.000 5058.035 3369.000 5083.000 ;
      LAYER met4 ;
        RECT 3369.000 5058.035 3371.000 5083.000 ;
      LAYER met4 ;
        RECT 3371.000 5058.035 3379.000 5083.000 ;
      LAYER met4 ;
        RECT 3379.000 5058.035 3381.000 5083.000 ;
      LAYER met4 ;
        RECT 3381.000 5058.035 3384.000 5083.000 ;
      LAYER met4 ;
        RECT 3384.000 5058.035 3390.645 5083.000 ;
      LAYER met4 ;
        RECT 3210.000 5057.635 3388.000 5058.035 ;
        RECT 3391.045 5057.635 3588.000 5083.400 ;
        RECT 3130.965 5056.935 3208.970 5057.635 ;
        RECT 3210.000 5056.935 3588.000 5057.635 ;
        RECT 0.000 5051.685 202.330 5056.935 ;
      LAYER met4 ;
        RECT 202.730 5052.085 382.270 5056.535 ;
      LAYER met4 ;
        RECT 382.670 5051.685 459.330 5056.935 ;
      LAYER met4 ;
        RECT 459.730 5052.085 639.270 5056.535 ;
      LAYER met4 ;
        RECT 639.670 5051.685 716.330 5056.935 ;
      LAYER met4 ;
        RECT 716.730 5052.085 896.270 5056.535 ;
      LAYER met4 ;
        RECT 896.670 5051.685 973.330 5056.935 ;
      LAYER met4 ;
        RECT 973.730 5052.085 1153.270 5056.535 ;
      LAYER met4 ;
        RECT 1153.670 5051.685 1230.330 5056.935 ;
      LAYER met4 ;
        RECT 1230.730 5052.085 1411.270 5056.535 ;
      LAYER met4 ;
        RECT 1411.670 5051.685 1488.330 5056.935 ;
      LAYER met4 ;
        RECT 1488.730 5052.085 1668.270 5056.535 ;
      LAYER met4 ;
        RECT 1668.670 5051.685 1740.330 5056.935 ;
      LAYER met4 ;
        RECT 1740.730 5052.085 1920.270 5056.535 ;
      LAYER met4 ;
        RECT 1920.670 5051.685 1997.330 5056.935 ;
      LAYER met4 ;
        RECT 1997.730 5052.085 2365.270 5056.535 ;
      LAYER met4 ;
        RECT 2365.670 5051.685 2442.330 5056.935 ;
      LAYER met4 ;
        RECT 2442.730 5052.085 2622.270 5056.535 ;
      LAYER met4 ;
        RECT 2622.670 5051.685 2699.330 5056.935 ;
      LAYER met4 ;
        RECT 2699.730 5052.085 2879.270 5056.535 ;
      LAYER met4 ;
        RECT 2879.670 5051.685 2951.330 5056.935 ;
      LAYER met4 ;
        RECT 2951.730 5052.085 3131.270 5056.535 ;
      LAYER met4 ;
        RECT 3131.670 5051.685 3208.330 5056.935 ;
      LAYER met4 ;
        RECT 3208.730 5052.085 3389.480 5056.535 ;
      LAYER met4 ;
        RECT 3389.880 5051.685 3588.000 5056.935 ;
        RECT 0.000 5051.085 202.745 5051.685 ;
        RECT 204.000 5051.085 379.000 5051.685 ;
        RECT 381.965 5051.085 459.970 5051.685 ;
        RECT 461.000 5051.085 636.000 5051.685 ;
        RECT 638.965 5051.085 716.970 5051.685 ;
        RECT 718.000 5051.085 893.000 5051.685 ;
        RECT 895.965 5051.085 973.970 5051.685 ;
        RECT 975.000 5051.085 1150.000 5051.685 ;
        RECT 1152.965 5051.085 1230.970 5051.685 ;
        RECT 1232.000 5051.085 1407.000 5051.685 ;
        RECT 1410.965 5051.085 1488.970 5051.685 ;
        RECT 1490.000 5051.085 1665.000 5051.685 ;
        RECT 1667.965 5051.085 1741.035 5051.685 ;
        RECT 1742.000 5051.085 1917.000 5051.685 ;
        RECT 1919.965 5051.085 1997.970 5051.685 ;
        RECT 1999.000 5051.085 2174.000 5051.685 ;
        RECT 2186.000 5051.085 2361.000 5051.685 ;
        RECT 2364.965 5051.085 2442.970 5051.685 ;
        RECT 2444.000 5051.085 2619.000 5051.685 ;
        RECT 2621.965 5051.085 2699.970 5051.685 ;
        RECT 2701.000 5051.085 2876.000 5051.685 ;
        RECT 2878.965 5051.085 2952.035 5051.685 ;
        RECT 2953.000 5051.085 3128.000 5051.685 ;
        RECT 3130.965 5051.085 3208.970 5051.685 ;
        RECT 3210.000 5051.085 3385.000 5051.685 ;
        RECT 3388.000 5051.085 3588.000 5051.685 ;
        RECT 0.000 5045.835 202.330 5051.085 ;
      LAYER met4 ;
        RECT 202.730 5046.235 382.270 5050.685 ;
      LAYER met4 ;
        RECT 382.670 5045.835 459.330 5051.085 ;
      LAYER met4 ;
        RECT 459.730 5046.235 639.270 5050.685 ;
      LAYER met4 ;
        RECT 639.670 5045.835 716.330 5051.085 ;
      LAYER met4 ;
        RECT 716.730 5046.235 896.270 5050.685 ;
      LAYER met4 ;
        RECT 896.670 5045.835 973.330 5051.085 ;
      LAYER met4 ;
        RECT 973.730 5046.235 1153.270 5050.685 ;
      LAYER met4 ;
        RECT 1153.670 5045.835 1230.330 5051.085 ;
      LAYER met4 ;
        RECT 1230.730 5046.235 1411.270 5050.685 ;
      LAYER met4 ;
        RECT 1411.670 5045.835 1488.330 5051.085 ;
      LAYER met4 ;
        RECT 1488.730 5046.235 1668.270 5050.685 ;
      LAYER met4 ;
        RECT 1668.670 5045.835 1740.330 5051.085 ;
      LAYER met4 ;
        RECT 1740.730 5046.235 1920.270 5050.685 ;
      LAYER met4 ;
        RECT 1920.670 5045.835 1997.330 5051.085 ;
      LAYER met4 ;
        RECT 1997.730 5046.235 2365.270 5050.685 ;
      LAYER met4 ;
        RECT 2365.670 5045.835 2442.330 5051.085 ;
      LAYER met4 ;
        RECT 2442.730 5046.235 2622.270 5050.685 ;
      LAYER met4 ;
        RECT 2622.670 5045.835 2699.330 5051.085 ;
      LAYER met4 ;
        RECT 2699.730 5046.235 2879.270 5050.685 ;
      LAYER met4 ;
        RECT 2879.670 5045.835 2951.330 5051.085 ;
      LAYER met4 ;
        RECT 2951.730 5046.235 3131.270 5050.685 ;
      LAYER met4 ;
        RECT 3131.670 5045.835 3208.330 5051.085 ;
      LAYER met4 ;
        RECT 3208.730 5046.235 3389.625 5050.685 ;
      LAYER met4 ;
        RECT 3390.025 5045.835 3588.000 5051.085 ;
        RECT 0.000 5045.135 202.745 5045.835 ;
        RECT 204.000 5045.135 381.000 5045.835 ;
        RECT 381.965 5045.135 459.970 5045.835 ;
        RECT 461.000 5045.135 638.000 5045.835 ;
        RECT 638.965 5045.135 716.970 5045.835 ;
        RECT 718.000 5045.135 895.000 5045.835 ;
        RECT 895.965 5045.135 973.970 5045.835 ;
        RECT 975.000 5045.135 1152.000 5045.835 ;
        RECT 1152.965 5045.135 1230.970 5045.835 ;
        RECT 1232.000 5045.135 1410.000 5045.835 ;
        RECT 1410.965 5045.135 1488.970 5045.835 ;
        RECT 1490.000 5045.135 1667.000 5045.835 ;
        RECT 1667.965 5045.135 1741.035 5045.835 ;
        RECT 1742.000 5045.135 1919.000 5045.835 ;
        RECT 1919.965 5045.135 1997.970 5045.835 ;
        RECT 1999.000 5045.135 2176.000 5045.835 ;
        RECT 2186.000 5045.135 2364.000 5045.835 ;
        RECT 2364.965 5045.135 2442.970 5045.835 ;
        RECT 2444.000 5045.135 2621.000 5045.835 ;
        RECT 2621.965 5045.135 2699.970 5045.835 ;
        RECT 2701.000 5045.135 2878.000 5045.835 ;
        RECT 2878.965 5045.135 2952.035 5045.835 ;
        RECT 2953.000 5045.135 3130.000 5045.835 ;
        RECT 3130.965 5045.135 3208.970 5045.835 ;
        RECT 3210.000 5045.135 3588.000 5045.835 ;
        RECT 0.000 5044.005 176.425 5045.135 ;
      LAYER met4 ;
        RECT 176.825 5044.405 383.610 5044.735 ;
      LAYER met4 ;
        RECT 384.010 5044.505 427.690 5045.135 ;
        RECT 0.000 5040.725 176.690 5044.005 ;
      LAYER met4 ;
        RECT 177.090 5041.125 417.440 5044.105 ;
      LAYER met4 ;
        RECT 0.000 5039.245 182.045 5040.725 ;
      LAYER met4 ;
        RECT 182.445 5039.645 204.000 5040.825 ;
      LAYER met4 ;
        RECT 204.000 5039.745 381.000 5040.725 ;
      LAYER met4 ;
        RECT 381.000 5039.645 382.270 5040.825 ;
      LAYER met4 ;
        RECT 417.840 5040.725 419.360 5044.505 ;
      LAYER met4 ;
        RECT 428.090 5044.405 640.610 5044.735 ;
      LAYER met4 ;
        RECT 641.010 5044.505 684.690 5045.135 ;
      LAYER met4 ;
        RECT 419.760 5041.125 674.440 5044.105 ;
      LAYER met4 ;
        RECT 382.670 5039.745 459.330 5040.725 ;
        RECT 0.000 5036.465 182.725 5039.245 ;
        RECT 0.000 5035.335 180.025 5036.465 ;
      LAYER met4 ;
        RECT 183.125 5036.365 433.145 5039.345 ;
      LAYER met4 ;
        RECT 433.545 5036.465 435.065 5039.745 ;
      LAYER met4 ;
        RECT 459.730 5039.645 461.000 5040.825 ;
      LAYER met4 ;
        RECT 461.000 5039.745 638.000 5040.725 ;
      LAYER met4 ;
        RECT 638.000 5039.645 639.270 5040.825 ;
      LAYER met4 ;
        RECT 674.840 5040.725 676.360 5044.505 ;
      LAYER met4 ;
        RECT 685.090 5044.405 897.610 5044.735 ;
      LAYER met4 ;
        RECT 898.010 5044.505 941.690 5045.135 ;
      LAYER met4 ;
        RECT 676.760 5041.125 931.440 5044.105 ;
      LAYER met4 ;
        RECT 639.670 5039.745 716.330 5040.725 ;
      LAYER met4 ;
        RECT 435.465 5036.365 690.145 5039.345 ;
      LAYER met4 ;
        RECT 690.545 5036.465 692.065 5039.745 ;
      LAYER met4 ;
        RECT 716.730 5039.645 718.000 5040.825 ;
      LAYER met4 ;
        RECT 718.000 5039.745 895.000 5040.725 ;
      LAYER met4 ;
        RECT 895.000 5039.645 896.270 5040.825 ;
      LAYER met4 ;
        RECT 931.840 5040.725 933.360 5044.505 ;
      LAYER met4 ;
        RECT 942.090 5044.405 1154.610 5044.735 ;
      LAYER met4 ;
        RECT 1155.010 5044.505 1198.690 5045.135 ;
      LAYER met4 ;
        RECT 933.760 5041.125 1188.440 5044.105 ;
      LAYER met4 ;
        RECT 896.670 5039.745 973.330 5040.725 ;
      LAYER met4 ;
        RECT 692.465 5036.365 947.145 5039.345 ;
      LAYER met4 ;
        RECT 947.545 5036.465 949.065 5039.745 ;
      LAYER met4 ;
        RECT 973.730 5039.645 975.000 5040.825 ;
      LAYER met4 ;
        RECT 975.000 5039.745 1152.000 5040.725 ;
      LAYER met4 ;
        RECT 1152.000 5039.645 1153.270 5040.825 ;
      LAYER met4 ;
        RECT 1188.840 5040.725 1190.360 5044.505 ;
      LAYER met4 ;
        RECT 1199.090 5044.405 1412.610 5044.735 ;
      LAYER met4 ;
        RECT 1413.010 5044.505 1456.690 5045.135 ;
      LAYER met4 ;
        RECT 1190.760 5041.125 1446.440 5044.105 ;
      LAYER met4 ;
        RECT 1153.670 5039.745 1230.330 5040.725 ;
      LAYER met4 ;
        RECT 949.465 5036.365 1204.145 5039.345 ;
      LAYER met4 ;
        RECT 1204.545 5036.465 1206.065 5039.745 ;
      LAYER met4 ;
        RECT 1230.730 5039.645 1232.000 5040.825 ;
      LAYER met4 ;
        RECT 1232.000 5039.745 1410.000 5040.725 ;
      LAYER met4 ;
        RECT 1410.000 5039.645 1411.270 5040.825 ;
      LAYER met4 ;
        RECT 1446.840 5040.725 1448.360 5044.505 ;
      LAYER met4 ;
        RECT 1457.090 5044.405 1921.610 5044.735 ;
      LAYER met4 ;
        RECT 1922.010 5044.505 1965.690 5045.135 ;
      LAYER met4 ;
        RECT 1448.760 5041.125 1955.440 5044.105 ;
      LAYER met4 ;
        RECT 1411.670 5039.745 1488.330 5040.725 ;
      LAYER met4 ;
        RECT 1206.465 5036.365 1462.145 5039.345 ;
      LAYER met4 ;
        RECT 1462.545 5036.465 1464.065 5039.745 ;
      LAYER met4 ;
        RECT 1488.730 5039.645 1490.000 5040.825 ;
      LAYER met4 ;
        RECT 1490.000 5039.745 1667.000 5040.725 ;
      LAYER met4 ;
        RECT 1667.000 5039.645 1668.270 5040.825 ;
      LAYER met4 ;
        RECT 1668.670 5039.745 1740.330 5040.725 ;
      LAYER met4 ;
        RECT 1740.730 5039.645 1742.000 5040.825 ;
      LAYER met4 ;
        RECT 1742.000 5039.745 1919.000 5040.725 ;
      LAYER met4 ;
        RECT 1919.000 5039.645 1920.270 5040.825 ;
      LAYER met4 ;
        RECT 1955.840 5040.725 1957.360 5044.505 ;
      LAYER met4 ;
        RECT 1966.090 5044.405 2176.000 5044.735 ;
        RECT 2181.000 5044.405 2366.610 5044.735 ;
      LAYER met4 ;
        RECT 2367.010 5044.505 2410.690 5045.135 ;
      LAYER met4 ;
        RECT 1957.760 5041.125 2400.440 5044.105 ;
      LAYER met4 ;
        RECT 1920.670 5039.745 1997.330 5040.725 ;
      LAYER met4 ;
        RECT 1464.465 5036.365 1971.145 5039.345 ;
      LAYER met4 ;
        RECT 1971.545 5036.465 1973.065 5039.745 ;
      LAYER met4 ;
        RECT 1997.730 5039.645 1999.000 5040.825 ;
      LAYER met4 ;
        RECT 2181.000 5040.725 2186.000 5040.825 ;
        RECT 1999.000 5039.745 2176.000 5040.725 ;
        RECT 2181.000 5039.745 2364.000 5040.725 ;
        RECT 2181.000 5039.645 2186.000 5039.745 ;
      LAYER met4 ;
        RECT 2364.000 5039.645 2365.270 5040.825 ;
      LAYER met4 ;
        RECT 2400.840 5040.725 2402.360 5044.505 ;
      LAYER met4 ;
        RECT 2411.090 5044.405 2623.610 5044.735 ;
      LAYER met4 ;
        RECT 2624.010 5044.505 2667.690 5045.135 ;
        RECT 2879.670 5044.505 2951.330 5045.135 ;
        RECT 3133.010 5044.505 3176.690 5045.135 ;
      LAYER met4 ;
        RECT 2402.760 5041.125 2657.440 5044.105 ;
      LAYER met4 ;
        RECT 2365.670 5039.745 2442.330 5040.725 ;
      LAYER met4 ;
        RECT 1973.465 5036.365 2416.145 5039.345 ;
      LAYER met4 ;
        RECT 2416.545 5036.465 2418.065 5039.745 ;
      LAYER met4 ;
        RECT 2442.730 5039.645 2444.000 5040.825 ;
      LAYER met4 ;
        RECT 2444.000 5039.745 2621.000 5040.725 ;
      LAYER met4 ;
        RECT 2621.000 5039.645 2622.270 5040.825 ;
      LAYER met4 ;
        RECT 2657.840 5040.725 2659.360 5044.505 ;
      LAYER met4 ;
        RECT 2659.760 5041.125 3166.440 5044.105 ;
      LAYER met4 ;
        RECT 2622.670 5039.745 2699.330 5040.725 ;
      LAYER met4 ;
        RECT 2418.465 5036.365 2673.145 5039.345 ;
      LAYER met4 ;
        RECT 2673.545 5036.465 2675.065 5039.745 ;
      LAYER met4 ;
        RECT 2699.730 5039.645 2701.000 5040.825 ;
      LAYER met4 ;
        RECT 2701.000 5039.745 2878.000 5040.725 ;
        RECT 2879.670 5039.745 2951.330 5040.725 ;
        RECT 2953.000 5039.745 3130.000 5040.725 ;
      LAYER met4 ;
        RECT 3130.000 5039.645 3131.270 5040.825 ;
      LAYER met4 ;
        RECT 3166.840 5040.725 3168.360 5044.505 ;
      LAYER met4 ;
        RECT 3177.090 5044.405 3411.175 5044.735 ;
        RECT 3168.760 5041.125 3410.910 5044.105 ;
      LAYER met4 ;
        RECT 3411.575 5044.005 3588.000 5045.135 ;
        RECT 3131.670 5039.745 3208.330 5040.725 ;
      LAYER met4 ;
        RECT 2675.465 5036.365 3182.145 5039.345 ;
      LAYER met4 ;
        RECT 3182.545 5036.465 3184.065 5039.745 ;
      LAYER met4 ;
        RECT 3208.730 5039.645 3210.000 5040.825 ;
      LAYER met4 ;
        RECT 3210.000 5039.745 3388.000 5040.725 ;
      LAYER met4 ;
        RECT 3388.000 5039.645 3409.550 5040.825 ;
      LAYER met4 ;
        RECT 3411.310 5040.725 3588.000 5044.005 ;
      LAYER met4 ;
        RECT 3184.465 5036.365 3408.935 5039.345 ;
      LAYER met4 ;
        RECT 3409.950 5039.245 3588.000 5040.725 ;
      LAYER met4 ;
        RECT 180.425 5035.735 383.610 5036.065 ;
      LAYER met4 ;
        RECT 384.010 5035.335 427.690 5035.965 ;
      LAYER met4 ;
        RECT 428.090 5035.735 640.610 5036.065 ;
      LAYER met4 ;
        RECT 641.010 5035.335 684.690 5035.965 ;
      LAYER met4 ;
        RECT 685.090 5035.735 897.610 5036.065 ;
      LAYER met4 ;
        RECT 898.010 5035.335 941.690 5035.965 ;
      LAYER met4 ;
        RECT 942.090 5035.735 1154.610 5036.065 ;
      LAYER met4 ;
        RECT 1155.010 5035.335 1198.690 5035.965 ;
      LAYER met4 ;
        RECT 1199.090 5035.735 1412.610 5036.065 ;
      LAYER met4 ;
        RECT 1413.010 5035.335 1456.690 5035.965 ;
      LAYER met4 ;
        RECT 1457.090 5035.735 1921.610 5036.065 ;
      LAYER met4 ;
        RECT 1922.010 5035.335 1965.690 5035.965 ;
      LAYER met4 ;
        RECT 1966.090 5035.735 2176.000 5036.065 ;
        RECT 2181.000 5035.735 2366.610 5036.065 ;
      LAYER met4 ;
        RECT 2367.010 5035.335 2410.690 5035.965 ;
      LAYER met4 ;
        RECT 2411.090 5035.735 2623.610 5036.065 ;
      LAYER met4 ;
        RECT 2624.010 5035.335 2667.690 5035.965 ;
        RECT 2879.670 5035.335 2951.330 5035.965 ;
        RECT 3133.010 5035.335 3176.690 5035.965 ;
      LAYER met4 ;
        RECT 3177.090 5035.735 3407.575 5036.065 ;
      LAYER met4 ;
        RECT 3409.335 5035.965 3588.000 5039.245 ;
        RECT 3407.975 5035.335 3588.000 5035.965 ;
        RECT 0.000 5034.635 202.745 5035.335 ;
        RECT 381.965 5034.635 459.970 5035.335 ;
        RECT 638.965 5034.635 716.970 5035.335 ;
        RECT 895.965 5034.635 973.970 5035.335 ;
        RECT 1152.965 5034.635 1230.970 5035.335 ;
        RECT 1410.965 5034.635 1488.970 5035.335 ;
        RECT 1667.965 5034.635 1741.035 5035.335 ;
        RECT 1919.965 5034.635 1997.970 5035.335 ;
        RECT 2364.965 5034.635 2442.970 5035.335 ;
        RECT 2621.965 5034.635 2699.970 5035.335 ;
        RECT 2878.965 5034.635 2952.035 5035.335 ;
        RECT 3130.965 5034.635 3208.970 5035.335 ;
        RECT 3388.000 5034.635 3588.000 5035.335 ;
        RECT 0.000 5029.185 202.330 5034.635 ;
      LAYER met4 ;
        RECT 202.730 5029.585 382.270 5034.235 ;
      LAYER met4 ;
        RECT 382.670 5029.185 459.330 5034.635 ;
      LAYER met4 ;
        RECT 459.730 5029.585 639.270 5034.235 ;
      LAYER met4 ;
        RECT 639.670 5029.185 716.330 5034.635 ;
      LAYER met4 ;
        RECT 716.730 5029.585 896.270 5034.235 ;
      LAYER met4 ;
        RECT 896.670 5029.185 973.330 5034.635 ;
      LAYER met4 ;
        RECT 973.730 5029.585 1153.270 5034.235 ;
      LAYER met4 ;
        RECT 1153.670 5029.185 1230.330 5034.635 ;
      LAYER met4 ;
        RECT 1230.730 5029.585 1411.270 5034.235 ;
      LAYER met4 ;
        RECT 1411.670 5029.185 1488.330 5034.635 ;
      LAYER met4 ;
        RECT 1488.730 5029.585 1668.270 5034.235 ;
      LAYER met4 ;
        RECT 1668.670 5029.185 1740.330 5034.635 ;
      LAYER met4 ;
        RECT 1740.730 5029.585 1920.270 5034.235 ;
      LAYER met4 ;
        RECT 1920.670 5029.185 1997.330 5034.635 ;
      LAYER met4 ;
        RECT 1997.730 5029.585 2181.000 5034.235 ;
        RECT 2186.000 5029.585 2365.270 5034.235 ;
      LAYER met4 ;
        RECT 2365.670 5029.185 2442.330 5034.635 ;
      LAYER met4 ;
        RECT 2442.730 5029.585 2622.270 5034.235 ;
      LAYER met4 ;
        RECT 2622.670 5029.185 2699.330 5034.635 ;
      LAYER met4 ;
        RECT 2699.730 5029.585 2879.270 5034.235 ;
      LAYER met4 ;
        RECT 2879.670 5029.185 2951.330 5034.635 ;
      LAYER met4 ;
        RECT 2951.730 5029.585 3131.270 5034.235 ;
      LAYER met4 ;
        RECT 3131.670 5029.185 3208.330 5034.635 ;
      LAYER met4 ;
        RECT 3208.730 5029.585 3389.475 5034.235 ;
      LAYER met4 ;
        RECT 3389.875 5029.185 3588.000 5034.635 ;
        RECT 0.000 5028.585 202.745 5029.185 ;
        RECT 381.965 5028.585 459.970 5029.185 ;
        RECT 638.965 5028.585 716.970 5029.185 ;
        RECT 895.965 5028.585 973.970 5029.185 ;
        RECT 1152.965 5028.585 1230.970 5029.185 ;
        RECT 1410.965 5028.585 1488.970 5029.185 ;
        RECT 1667.965 5028.585 1741.035 5029.185 ;
        RECT 1919.965 5028.585 1997.970 5029.185 ;
        RECT 2364.965 5028.585 2442.970 5029.185 ;
        RECT 2621.965 5028.585 2699.970 5029.185 ;
        RECT 2878.965 5028.585 2952.035 5029.185 ;
        RECT 3130.965 5028.585 3208.970 5029.185 ;
        RECT 3388.000 5028.585 3588.000 5029.185 ;
        RECT 0.000 5024.335 202.330 5028.585 ;
      LAYER met4 ;
        RECT 202.730 5024.735 382.270 5028.185 ;
      LAYER met4 ;
        RECT 382.670 5024.335 459.330 5028.585 ;
      LAYER met4 ;
        RECT 459.730 5024.735 639.270 5028.185 ;
      LAYER met4 ;
        RECT 639.670 5024.335 716.330 5028.585 ;
      LAYER met4 ;
        RECT 716.730 5024.735 896.270 5028.185 ;
      LAYER met4 ;
        RECT 896.670 5024.335 973.330 5028.585 ;
      LAYER met4 ;
        RECT 973.730 5024.735 1153.270 5028.185 ;
      LAYER met4 ;
        RECT 1153.670 5024.335 1230.330 5028.585 ;
      LAYER met4 ;
        RECT 1230.730 5024.735 1411.270 5028.185 ;
      LAYER met4 ;
        RECT 1411.670 5024.335 1488.330 5028.585 ;
      LAYER met4 ;
        RECT 1488.730 5024.735 1668.270 5028.185 ;
      LAYER met4 ;
        RECT 1668.670 5024.335 1740.330 5028.585 ;
      LAYER met4 ;
        RECT 1740.730 5024.735 1920.270 5028.185 ;
      LAYER met4 ;
        RECT 1920.670 5024.335 1997.330 5028.585 ;
      LAYER met4 ;
        RECT 1997.730 5024.735 2176.000 5028.185 ;
        RECT 2181.000 5024.735 2365.270 5028.185 ;
      LAYER met4 ;
        RECT 2365.670 5024.335 2442.330 5028.585 ;
      LAYER met4 ;
        RECT 2442.730 5024.735 2622.270 5028.185 ;
      LAYER met4 ;
        RECT 2622.670 5024.335 2699.330 5028.585 ;
        RECT 2879.670 5024.335 2951.330 5028.585 ;
        RECT 3131.670 5024.335 3208.330 5028.585 ;
      LAYER met4 ;
        RECT 3208.730 5024.735 3389.335 5028.185 ;
      LAYER met4 ;
        RECT 3389.735 5024.335 3588.000 5028.585 ;
        RECT 0.000 5023.735 202.745 5024.335 ;
        RECT 381.965 5023.735 459.970 5024.335 ;
        RECT 638.965 5023.735 716.970 5024.335 ;
        RECT 895.965 5023.735 973.970 5024.335 ;
        RECT 1152.965 5023.735 1230.970 5024.335 ;
        RECT 1410.965 5023.735 1488.970 5024.335 ;
        RECT 1667.965 5023.735 1741.035 5024.335 ;
        RECT 1919.965 5023.735 1997.970 5024.335 ;
        RECT 2364.965 5023.735 2442.970 5024.335 ;
        RECT 2621.965 5023.735 2699.970 5024.335 ;
        RECT 2878.965 5023.735 2952.035 5024.335 ;
        RECT 3130.965 5023.735 3208.970 5024.335 ;
        RECT 3388.000 5023.735 3588.000 5024.335 ;
        RECT 0.000 5019.485 202.330 5023.735 ;
      LAYER met4 ;
        RECT 202.730 5019.885 382.270 5023.335 ;
      LAYER met4 ;
        RECT 382.670 5019.485 459.330 5023.735 ;
      LAYER met4 ;
        RECT 459.730 5019.885 639.270 5023.335 ;
      LAYER met4 ;
        RECT 639.670 5019.485 716.330 5023.735 ;
      LAYER met4 ;
        RECT 716.730 5019.885 896.270 5023.335 ;
      LAYER met4 ;
        RECT 896.670 5019.485 973.330 5023.735 ;
      LAYER met4 ;
        RECT 973.730 5019.885 1153.270 5023.335 ;
      LAYER met4 ;
        RECT 1153.670 5019.485 1230.330 5023.735 ;
      LAYER met4 ;
        RECT 1230.730 5019.885 1411.270 5023.335 ;
      LAYER met4 ;
        RECT 1411.670 5019.485 1488.330 5023.735 ;
      LAYER met4 ;
        RECT 1488.730 5019.885 1668.270 5023.335 ;
      LAYER met4 ;
        RECT 1668.670 5019.485 1740.330 5023.735 ;
      LAYER met4 ;
        RECT 1740.730 5019.885 1920.270 5023.335 ;
      LAYER met4 ;
        RECT 1920.670 5019.485 1997.330 5023.735 ;
      LAYER met4 ;
        RECT 1997.730 5019.885 2365.270 5023.335 ;
      LAYER met4 ;
        RECT 2365.670 5019.485 2442.330 5023.735 ;
      LAYER met4 ;
        RECT 2442.730 5019.885 2622.270 5023.335 ;
      LAYER met4 ;
        RECT 2622.670 5019.485 2699.330 5023.735 ;
      LAYER met4 ;
        RECT 2699.730 5019.885 2879.270 5023.335 ;
      LAYER met4 ;
        RECT 2879.670 5019.485 2951.330 5023.735 ;
      LAYER met4 ;
        RECT 2951.730 5019.885 3131.270 5023.335 ;
      LAYER met4 ;
        RECT 3131.670 5019.485 3208.330 5023.735 ;
      LAYER met4 ;
        RECT 3208.730 5019.885 3389.385 5023.335 ;
      LAYER met4 ;
        RECT 3389.785 5019.485 3588.000 5023.735 ;
        RECT 0.000 5018.885 202.745 5019.485 ;
        RECT 381.965 5018.885 459.970 5019.485 ;
        RECT 638.965 5018.885 716.970 5019.485 ;
        RECT 895.965 5018.885 973.970 5019.485 ;
        RECT 1152.965 5018.885 1230.970 5019.485 ;
        RECT 1410.965 5018.885 1488.970 5019.485 ;
        RECT 1667.965 5018.885 1741.035 5019.485 ;
        RECT 1919.965 5018.885 1997.970 5019.485 ;
        RECT 2364.965 5018.885 2442.970 5019.485 ;
        RECT 2621.965 5018.885 2699.970 5019.485 ;
        RECT 2878.965 5018.885 2952.035 5019.485 ;
        RECT 3130.965 5018.885 3208.970 5019.485 ;
        RECT 3388.000 5018.885 3588.000 5019.485 ;
        RECT 0.000 5013.435 202.330 5018.885 ;
      LAYER met4 ;
        RECT 202.730 5013.835 382.270 5018.485 ;
      LAYER met4 ;
        RECT 382.670 5013.435 459.330 5018.885 ;
      LAYER met4 ;
        RECT 459.730 5013.835 639.270 5018.485 ;
      LAYER met4 ;
        RECT 639.670 5013.435 716.330 5018.885 ;
      LAYER met4 ;
        RECT 716.730 5013.835 896.270 5018.485 ;
      LAYER met4 ;
        RECT 896.670 5013.435 973.330 5018.885 ;
      LAYER met4 ;
        RECT 973.730 5013.835 1153.270 5018.485 ;
      LAYER met4 ;
        RECT 1153.670 5013.435 1230.330 5018.885 ;
      LAYER met4 ;
        RECT 1230.730 5013.835 1411.270 5018.485 ;
      LAYER met4 ;
        RECT 1411.670 5013.435 1488.330 5018.885 ;
        RECT 1668.670 5013.435 1740.330 5018.885 ;
        RECT 1920.670 5013.435 1997.330 5018.885 ;
      LAYER met4 ;
        RECT 1997.730 5013.835 2365.270 5018.485 ;
      LAYER met4 ;
        RECT 2365.670 5013.435 2442.330 5018.885 ;
      LAYER met4 ;
        RECT 2442.730 5013.835 2622.270 5018.485 ;
      LAYER met4 ;
        RECT 2622.670 5013.435 2699.330 5018.885 ;
      LAYER met4 ;
        RECT 2699.730 5013.835 2879.270 5018.485 ;
      LAYER met4 ;
        RECT 2879.670 5013.435 2951.330 5018.885 ;
      LAYER met4 ;
        RECT 2951.730 5013.835 3131.270 5018.485 ;
      LAYER met4 ;
        RECT 3131.670 5013.435 3208.330 5018.885 ;
      LAYER met4 ;
        RECT 3208.730 5013.835 3389.600 5018.485 ;
      LAYER met4 ;
        RECT 3390.000 5013.435 3588.000 5018.885 ;
        RECT 0.000 5012.835 202.745 5013.435 ;
        RECT 381.965 5012.835 459.970 5013.435 ;
        RECT 638.965 5012.835 716.970 5013.435 ;
        RECT 895.965 5012.835 973.970 5013.435 ;
        RECT 1152.965 5012.835 1230.970 5013.435 ;
        RECT 1410.965 5012.835 1488.970 5013.435 ;
        RECT 1667.965 5012.835 1741.035 5013.435 ;
        RECT 1919.965 5012.835 1997.970 5013.435 ;
        RECT 2364.965 5012.835 2442.970 5013.435 ;
        RECT 2621.965 5012.835 2699.970 5013.435 ;
        RECT 2878.965 5012.835 2952.035 5013.435 ;
        RECT 3130.965 5012.835 3208.970 5013.435 ;
        RECT 3388.000 5012.835 3588.000 5013.435 ;
        RECT 0.000 5011.575 202.330 5012.835 ;
        RECT 0.000 4991.045 142.865 5011.575 ;
        RECT 143.995 5011.310 202.330 5011.575 ;
        RECT 0.000 4989.835 104.600 4991.045 ;
      LAYER met4 ;
        RECT 0.000 4988.000 24.215 4989.435 ;
      LAYER met4 ;
        RECT 24.615 4988.000 104.600 4989.835 ;
        RECT 0.000 4851.000 25.965 4988.000 ;
        RECT 102.965 4985.000 105.000 4988.000 ;
      LAYER met4 ;
        RECT 105.000 4985.000 129.965 4990.645 ;
      LAYER met4 ;
        RECT 130.365 4990.025 142.865 4991.045 ;
        RECT 130.365 4989.880 136.915 4990.025 ;
        RECT 130.365 4988.000 131.065 4989.880 ;
        RECT 129.965 4985.000 131.065 4988.000 ;
        RECT 102.965 4982.000 131.065 4985.000 ;
        RECT 102.965 4980.000 105.000 4982.000 ;
      LAYER met4 ;
        RECT 105.000 4980.000 129.965 4982.000 ;
      LAYER met4 ;
        RECT 129.965 4980.000 131.065 4982.000 ;
        RECT 102.965 4972.000 131.065 4980.000 ;
        RECT 102.965 4970.000 105.000 4972.000 ;
      LAYER met4 ;
        RECT 105.000 4970.000 129.965 4972.000 ;
      LAYER met4 ;
        RECT 129.965 4970.000 131.065 4972.000 ;
        RECT 102.965 4952.000 131.065 4970.000 ;
        RECT 102.965 4950.000 105.000 4952.000 ;
      LAYER met4 ;
        RECT 105.000 4950.000 129.965 4952.000 ;
      LAYER met4 ;
        RECT 129.965 4950.000 131.065 4952.000 ;
        RECT 102.965 4932.000 131.065 4950.000 ;
        RECT 102.965 4930.000 105.000 4932.000 ;
      LAYER met4 ;
        RECT 105.000 4930.000 129.965 4932.000 ;
      LAYER met4 ;
        RECT 129.965 4930.000 131.065 4932.000 ;
        RECT 102.965 4912.000 131.065 4930.000 ;
        RECT 102.965 4910.000 105.000 4912.000 ;
      LAYER met4 ;
        RECT 105.000 4910.000 129.965 4912.000 ;
      LAYER met4 ;
        RECT 129.965 4910.000 131.065 4912.000 ;
        RECT 102.965 4892.000 131.065 4910.000 ;
        RECT 102.965 4890.000 105.000 4892.000 ;
      LAYER met4 ;
        RECT 105.000 4890.000 129.965 4892.000 ;
      LAYER met4 ;
        RECT 129.965 4890.000 131.065 4892.000 ;
        RECT 102.965 4872.000 131.065 4890.000 ;
        RECT 102.965 4870.000 105.000 4872.000 ;
      LAYER met4 ;
        RECT 105.000 4870.000 129.965 4872.000 ;
      LAYER met4 ;
        RECT 129.965 4870.000 131.065 4872.000 ;
        RECT 102.965 4852.000 131.065 4870.000 ;
        RECT 102.965 4851.000 105.000 4852.000 ;
      LAYER met4 ;
        RECT 0.000 4849.730 24.215 4851.000 ;
      LAYER met4 ;
        RECT 24.615 4849.330 104.600 4849.970 ;
      LAYER met4 ;
        RECT 105.000 4849.730 129.965 4852.000 ;
      LAYER met4 ;
        RECT 129.965 4851.000 131.065 4852.000 ;
        RECT 130.365 4849.330 131.065 4849.970 ;
      LAYER met4 ;
        RECT 131.465 4849.730 135.915 4989.480 ;
      LAYER met4 ;
        RECT 136.315 4988.000 136.915 4989.880 ;
        RECT 136.315 4851.000 136.915 4986.000 ;
        RECT 136.315 4849.330 136.915 4849.970 ;
      LAYER met4 ;
        RECT 137.315 4849.730 141.765 4989.625 ;
      LAYER met4 ;
        RECT 142.165 4851.000 142.865 4990.025 ;
        RECT 142.165 4849.330 142.865 4849.970 ;
        RECT 0.000 4817.690 142.865 4849.330 ;
      LAYER met4 ;
        RECT 143.265 4818.090 143.595 5011.175 ;
      LAYER met4 ;
        RECT 0.000 4809.360 143.495 4817.690 ;
      LAYER met4 ;
        RECT 143.895 4809.760 146.875 5010.910 ;
      LAYER met4 ;
        RECT 147.275 5009.950 202.330 5011.310 ;
      LAYER met4 ;
        RECT 147.175 4988.000 148.355 5009.550 ;
      LAYER met4 ;
        RECT 148.755 5009.335 202.330 5009.950 ;
        RECT 147.275 4851.000 148.255 4988.000 ;
      LAYER met4 ;
        RECT 147.175 4849.730 148.355 4851.000 ;
      LAYER met4 ;
        RECT 147.275 4825.065 148.255 4849.330 ;
      LAYER met4 ;
        RECT 148.655 4825.465 151.635 5008.935 ;
      LAYER met4 ;
        RECT 152.035 5007.975 202.330 5009.335 ;
        RECT 147.275 4823.545 151.535 4825.065 ;
        RECT 147.275 4809.360 148.255 4823.545 ;
        RECT 0.000 4807.840 148.255 4809.360 ;
        RECT 0.000 4774.010 143.495 4807.840 ;
        RECT 0.000 4772.670 142.865 4774.010 ;
      LAYER met4 ;
        RECT 0.000 4771.000 24.215 4772.270 ;
      LAYER met4 ;
        RECT 24.615 4771.965 104.600 4772.670 ;
        RECT 0.000 4635.000 25.965 4771.000 ;
        RECT 102.965 4769.000 105.000 4771.000 ;
      LAYER met4 ;
        RECT 105.000 4769.000 129.965 4772.270 ;
      LAYER met4 ;
        RECT 130.365 4771.965 131.065 4772.670 ;
        RECT 129.965 4769.000 131.065 4771.000 ;
        RECT 102.965 4766.000 131.065 4769.000 ;
        RECT 102.965 4764.000 105.000 4766.000 ;
      LAYER met4 ;
        RECT 105.000 4764.000 129.965 4766.000 ;
      LAYER met4 ;
        RECT 129.965 4764.000 131.065 4766.000 ;
        RECT 102.965 4756.000 131.065 4764.000 ;
        RECT 102.965 4754.000 105.000 4756.000 ;
      LAYER met4 ;
        RECT 105.000 4754.000 129.965 4756.000 ;
      LAYER met4 ;
        RECT 129.965 4754.000 131.065 4756.000 ;
        RECT 102.965 4736.000 131.065 4754.000 ;
        RECT 102.965 4734.000 105.000 4736.000 ;
      LAYER met4 ;
        RECT 105.000 4734.000 129.965 4736.000 ;
      LAYER met4 ;
        RECT 129.965 4734.000 131.065 4736.000 ;
        RECT 102.965 4716.000 131.065 4734.000 ;
        RECT 102.965 4714.000 105.000 4716.000 ;
      LAYER met4 ;
        RECT 105.000 4714.000 129.965 4716.000 ;
      LAYER met4 ;
        RECT 129.965 4714.000 131.065 4716.000 ;
        RECT 102.965 4696.000 131.065 4714.000 ;
        RECT 102.965 4694.000 105.000 4696.000 ;
      LAYER met4 ;
        RECT 105.000 4694.000 129.965 4696.000 ;
      LAYER met4 ;
        RECT 129.965 4694.000 131.065 4696.000 ;
        RECT 102.965 4676.000 131.065 4694.000 ;
        RECT 102.965 4674.000 105.000 4676.000 ;
      LAYER met4 ;
        RECT 105.000 4674.000 129.965 4676.000 ;
      LAYER met4 ;
        RECT 129.965 4674.000 131.065 4676.000 ;
        RECT 102.965 4656.000 131.065 4674.000 ;
        RECT 102.965 4654.000 105.000 4656.000 ;
      LAYER met4 ;
        RECT 105.000 4654.000 129.965 4656.000 ;
      LAYER met4 ;
        RECT 129.965 4654.000 131.065 4656.000 ;
        RECT 102.965 4636.000 131.065 4654.000 ;
        RECT 102.965 4635.000 105.000 4636.000 ;
      LAYER met4 ;
        RECT 0.000 4633.730 24.215 4635.000 ;
      LAYER met4 ;
        RECT 24.615 4633.330 104.600 4635.000 ;
      LAYER met4 ;
        RECT 105.000 4633.730 129.965 4636.000 ;
      LAYER met4 ;
        RECT 129.965 4635.000 131.065 4636.000 ;
        RECT 130.365 4633.330 131.065 4635.000 ;
      LAYER met4 ;
        RECT 131.465 4633.730 135.915 4772.270 ;
      LAYER met4 ;
        RECT 136.315 4771.965 136.915 4772.670 ;
        RECT 136.315 4633.330 136.915 4770.000 ;
      LAYER met4 ;
        RECT 137.315 4633.730 141.765 4772.270 ;
      LAYER met4 ;
        RECT 142.165 4771.965 142.865 4772.670 ;
        RECT 142.165 4633.330 142.865 4771.000 ;
        RECT 0.000 4561.670 142.865 4633.330 ;
      LAYER met4 ;
        RECT 0.000 4560.000 24.215 4561.270 ;
      LAYER met4 ;
        RECT 24.615 4560.965 104.600 4561.670 ;
        RECT 0.000 4424.000 25.965 4560.000 ;
        RECT 102.965 4558.000 105.000 4560.000 ;
      LAYER met4 ;
        RECT 105.000 4558.000 129.965 4561.270 ;
      LAYER met4 ;
        RECT 130.365 4560.965 131.065 4561.670 ;
        RECT 129.965 4558.000 131.065 4560.000 ;
        RECT 102.965 4555.000 131.065 4558.000 ;
        RECT 102.965 4553.000 105.000 4555.000 ;
      LAYER met4 ;
        RECT 105.000 4553.000 129.965 4555.000 ;
      LAYER met4 ;
        RECT 129.965 4553.000 131.065 4555.000 ;
        RECT 102.965 4545.000 131.065 4553.000 ;
        RECT 102.965 4543.000 105.000 4545.000 ;
      LAYER met4 ;
        RECT 105.000 4543.000 129.965 4545.000 ;
      LAYER met4 ;
        RECT 129.965 4543.000 131.065 4545.000 ;
        RECT 102.965 4525.000 131.065 4543.000 ;
        RECT 102.965 4523.000 105.000 4525.000 ;
      LAYER met4 ;
        RECT 105.000 4523.000 129.965 4525.000 ;
      LAYER met4 ;
        RECT 129.965 4523.000 131.065 4525.000 ;
        RECT 102.965 4505.000 131.065 4523.000 ;
        RECT 102.965 4503.000 105.000 4505.000 ;
      LAYER met4 ;
        RECT 105.000 4503.000 129.965 4505.000 ;
      LAYER met4 ;
        RECT 129.965 4503.000 131.065 4505.000 ;
        RECT 102.965 4485.000 131.065 4503.000 ;
        RECT 102.965 4483.000 105.000 4485.000 ;
      LAYER met4 ;
        RECT 105.000 4483.000 129.965 4485.000 ;
      LAYER met4 ;
        RECT 129.965 4483.000 131.065 4485.000 ;
        RECT 102.965 4465.000 131.065 4483.000 ;
        RECT 102.965 4463.000 105.000 4465.000 ;
      LAYER met4 ;
        RECT 105.000 4463.000 129.965 4465.000 ;
      LAYER met4 ;
        RECT 129.965 4463.000 131.065 4465.000 ;
        RECT 102.965 4445.000 131.065 4463.000 ;
        RECT 102.965 4443.000 105.000 4445.000 ;
      LAYER met4 ;
        RECT 105.000 4443.000 129.965 4445.000 ;
      LAYER met4 ;
        RECT 129.965 4443.000 131.065 4445.000 ;
        RECT 102.965 4425.000 131.065 4443.000 ;
        RECT 102.965 4424.000 105.000 4425.000 ;
      LAYER met4 ;
        RECT 0.000 4422.730 24.215 4424.000 ;
      LAYER met4 ;
        RECT 24.615 4422.330 104.600 4423.035 ;
      LAYER met4 ;
        RECT 105.000 4422.730 129.965 4425.000 ;
      LAYER met4 ;
        RECT 129.965 4424.000 131.065 4425.000 ;
        RECT 130.365 4422.330 131.065 4423.035 ;
      LAYER met4 ;
        RECT 131.465 4422.730 135.915 4561.270 ;
      LAYER met4 ;
        RECT 136.315 4560.965 136.915 4561.670 ;
        RECT 136.315 4424.000 136.915 4559.000 ;
        RECT 136.315 4422.330 136.915 4423.035 ;
      LAYER met4 ;
        RECT 137.315 4422.730 141.765 4561.270 ;
      LAYER met4 ;
        RECT 142.165 4560.965 142.865 4561.670 ;
        RECT 142.165 4424.000 142.865 4560.000 ;
        RECT 142.165 4422.330 142.865 4423.035 ;
        RECT 0.000 4350.670 142.865 4422.330 ;
      LAYER met4 ;
        RECT 0.000 4349.000 24.215 4350.270 ;
      LAYER met4 ;
        RECT 24.615 4349.965 104.600 4350.670 ;
        RECT 0.000 4213.000 25.965 4349.000 ;
        RECT 102.965 4347.000 105.000 4349.000 ;
      LAYER met4 ;
        RECT 105.000 4347.000 129.965 4350.270 ;
      LAYER met4 ;
        RECT 130.365 4349.965 131.065 4350.670 ;
        RECT 129.965 4347.000 131.065 4349.000 ;
        RECT 102.965 4344.000 131.065 4347.000 ;
        RECT 102.965 4342.000 105.000 4344.000 ;
      LAYER met4 ;
        RECT 105.000 4342.000 129.965 4344.000 ;
      LAYER met4 ;
        RECT 129.965 4342.000 131.065 4344.000 ;
        RECT 102.965 4334.000 131.065 4342.000 ;
        RECT 102.965 4332.000 105.000 4334.000 ;
      LAYER met4 ;
        RECT 105.000 4332.000 129.965 4334.000 ;
      LAYER met4 ;
        RECT 129.965 4332.000 131.065 4334.000 ;
        RECT 102.965 4314.000 131.065 4332.000 ;
        RECT 102.965 4312.000 105.000 4314.000 ;
      LAYER met4 ;
        RECT 105.000 4312.000 129.965 4314.000 ;
      LAYER met4 ;
        RECT 129.965 4312.000 131.065 4314.000 ;
        RECT 102.965 4294.000 131.065 4312.000 ;
        RECT 102.965 4292.000 105.000 4294.000 ;
      LAYER met4 ;
        RECT 105.000 4292.000 129.965 4294.000 ;
      LAYER met4 ;
        RECT 129.965 4292.000 131.065 4294.000 ;
        RECT 102.965 4274.000 131.065 4292.000 ;
        RECT 102.965 4272.000 105.000 4274.000 ;
      LAYER met4 ;
        RECT 105.000 4272.000 129.965 4274.000 ;
      LAYER met4 ;
        RECT 129.965 4272.000 131.065 4274.000 ;
        RECT 102.965 4254.000 131.065 4272.000 ;
        RECT 102.965 4252.000 105.000 4254.000 ;
      LAYER met4 ;
        RECT 105.000 4252.000 129.965 4254.000 ;
      LAYER met4 ;
        RECT 129.965 4252.000 131.065 4254.000 ;
        RECT 102.965 4234.000 131.065 4252.000 ;
        RECT 102.965 4232.000 105.000 4234.000 ;
      LAYER met4 ;
        RECT 105.000 4232.000 129.965 4234.000 ;
      LAYER met4 ;
        RECT 129.965 4232.000 131.065 4234.000 ;
        RECT 102.965 4214.000 131.065 4232.000 ;
        RECT 102.965 4213.000 105.000 4214.000 ;
      LAYER met4 ;
        RECT 0.000 4211.730 24.215 4213.000 ;
      LAYER met4 ;
        RECT 24.615 4211.330 104.600 4212.035 ;
      LAYER met4 ;
        RECT 105.000 4211.730 129.965 4214.000 ;
      LAYER met4 ;
        RECT 129.965 4213.000 131.065 4214.000 ;
        RECT 130.365 4211.330 131.065 4212.035 ;
      LAYER met4 ;
        RECT 131.465 4211.730 135.915 4350.270 ;
      LAYER met4 ;
        RECT 136.315 4349.965 136.915 4350.670 ;
        RECT 136.315 4213.000 136.915 4348.000 ;
        RECT 136.315 4211.330 136.915 4212.035 ;
      LAYER met4 ;
        RECT 137.315 4211.730 141.765 4350.270 ;
      LAYER met4 ;
        RECT 142.165 4349.965 142.865 4350.670 ;
        RECT 142.165 4213.000 142.865 4349.000 ;
        RECT 142.165 4211.330 142.865 4212.035 ;
        RECT 0.000 4139.670 143.495 4211.330 ;
      LAYER met4 ;
        RECT 0.000 4138.000 24.215 4139.270 ;
      LAYER met4 ;
        RECT 24.615 4138.965 104.600 4139.670 ;
        RECT 0.000 4002.000 25.965 4138.000 ;
        RECT 102.965 4136.000 105.000 4138.000 ;
      LAYER met4 ;
        RECT 105.000 4136.000 129.965 4139.270 ;
      LAYER met4 ;
        RECT 130.365 4138.965 131.065 4139.670 ;
        RECT 129.965 4136.000 131.065 4138.000 ;
        RECT 102.965 4133.000 131.065 4136.000 ;
        RECT 102.965 4131.000 105.000 4133.000 ;
      LAYER met4 ;
        RECT 105.000 4131.000 129.965 4133.000 ;
      LAYER met4 ;
        RECT 129.965 4131.000 131.065 4133.000 ;
        RECT 102.965 4123.000 131.065 4131.000 ;
        RECT 102.965 4121.000 105.000 4123.000 ;
      LAYER met4 ;
        RECT 105.000 4121.000 129.965 4123.000 ;
      LAYER met4 ;
        RECT 129.965 4121.000 131.065 4123.000 ;
        RECT 102.965 4103.000 131.065 4121.000 ;
        RECT 102.965 4101.000 105.000 4103.000 ;
      LAYER met4 ;
        RECT 105.000 4101.000 129.965 4103.000 ;
      LAYER met4 ;
        RECT 129.965 4101.000 131.065 4103.000 ;
        RECT 102.965 4083.000 131.065 4101.000 ;
        RECT 102.965 4081.000 105.000 4083.000 ;
      LAYER met4 ;
        RECT 105.000 4081.000 129.965 4083.000 ;
      LAYER met4 ;
        RECT 129.965 4081.000 131.065 4083.000 ;
        RECT 102.965 4063.000 131.065 4081.000 ;
        RECT 102.965 4061.000 105.000 4063.000 ;
      LAYER met4 ;
        RECT 105.000 4061.000 129.965 4063.000 ;
      LAYER met4 ;
        RECT 129.965 4061.000 131.065 4063.000 ;
        RECT 102.965 4043.000 131.065 4061.000 ;
        RECT 102.965 4041.000 105.000 4043.000 ;
      LAYER met4 ;
        RECT 105.000 4041.000 129.965 4043.000 ;
      LAYER met4 ;
        RECT 129.965 4041.000 131.065 4043.000 ;
        RECT 102.965 4023.000 131.065 4041.000 ;
        RECT 102.965 4021.000 105.000 4023.000 ;
      LAYER met4 ;
        RECT 105.000 4021.000 129.965 4023.000 ;
      LAYER met4 ;
        RECT 129.965 4021.000 131.065 4023.000 ;
        RECT 102.965 4003.000 131.065 4021.000 ;
        RECT 102.965 4002.000 105.000 4003.000 ;
      LAYER met4 ;
        RECT 0.000 4000.730 24.215 4002.000 ;
      LAYER met4 ;
        RECT 24.615 4000.330 104.600 4000.970 ;
      LAYER met4 ;
        RECT 105.000 4000.730 129.965 4003.000 ;
      LAYER met4 ;
        RECT 129.965 4002.000 131.065 4003.000 ;
        RECT 130.365 4000.330 131.065 4000.970 ;
      LAYER met4 ;
        RECT 131.465 4000.730 135.915 4139.270 ;
      LAYER met4 ;
        RECT 136.315 4138.965 136.915 4139.670 ;
        RECT 136.315 4002.000 136.915 4137.000 ;
        RECT 136.315 4000.330 136.915 4000.970 ;
      LAYER met4 ;
        RECT 137.315 4000.730 141.765 4139.270 ;
      LAYER met4 ;
        RECT 142.165 4138.965 142.865 4139.670 ;
        RECT 142.165 4002.000 142.865 4138.000 ;
        RECT 142.165 4000.330 142.865 4000.970 ;
        RECT 0.000 3968.690 142.865 4000.330 ;
        RECT 0.000 3960.360 143.495 3968.690 ;
      LAYER met4 ;
        RECT 143.895 3960.760 146.875 4807.440 ;
      LAYER met4 ;
        RECT 147.275 4772.670 148.255 4807.840 ;
      LAYER met4 ;
        RECT 147.175 4771.000 148.355 4772.270 ;
      LAYER met4 ;
        RECT 147.275 4635.000 148.255 4771.000 ;
      LAYER met4 ;
        RECT 147.175 4633.730 148.355 4635.000 ;
      LAYER met4 ;
        RECT 147.275 4561.670 148.255 4633.330 ;
      LAYER met4 ;
        RECT 147.175 4560.000 148.355 4561.270 ;
      LAYER met4 ;
        RECT 147.275 4424.000 148.255 4560.000 ;
      LAYER met4 ;
        RECT 147.175 4422.730 148.355 4424.000 ;
      LAYER met4 ;
        RECT 147.275 4350.670 148.255 4422.330 ;
      LAYER met4 ;
        RECT 147.175 4349.000 148.355 4350.270 ;
      LAYER met4 ;
        RECT 147.275 4213.000 148.255 4349.000 ;
        RECT 147.275 4139.670 148.255 4211.330 ;
        RECT 147.275 4002.000 148.255 4138.000 ;
      LAYER met4 ;
        RECT 147.175 4000.730 148.355 4002.000 ;
      LAYER met4 ;
        RECT 147.275 3976.065 148.255 4000.330 ;
      LAYER met4 ;
        RECT 148.655 3976.465 151.635 4823.145 ;
        RECT 151.935 4818.090 152.265 5007.575 ;
      LAYER met4 ;
        RECT 152.665 5007.385 202.330 5007.975 ;
      LAYER met4 ;
        RECT 202.730 5007.785 382.270 5012.435 ;
      LAYER met4 ;
        RECT 382.670 5007.385 459.330 5012.835 ;
      LAYER met4 ;
        RECT 459.730 5007.785 639.270 5012.435 ;
      LAYER met4 ;
        RECT 639.670 5007.385 716.330 5012.835 ;
      LAYER met4 ;
        RECT 716.730 5007.785 896.270 5012.435 ;
      LAYER met4 ;
        RECT 896.670 5007.385 973.330 5012.835 ;
      LAYER met4 ;
        RECT 973.730 5007.785 1153.270 5012.435 ;
      LAYER met4 ;
        RECT 1153.670 5007.385 1230.330 5012.835 ;
      LAYER met4 ;
        RECT 1230.730 5007.785 1411.270 5012.435 ;
      LAYER met4 ;
        RECT 1411.670 5007.385 1488.330 5012.835 ;
      LAYER met4 ;
        RECT 1488.730 5007.785 1668.270 5012.435 ;
      LAYER met4 ;
        RECT 1668.670 5007.385 1740.330 5012.835 ;
      LAYER met4 ;
        RECT 1740.730 5007.785 1920.270 5012.435 ;
      LAYER met4 ;
        RECT 1920.670 5007.385 1997.330 5012.835 ;
      LAYER met4 ;
        RECT 1997.730 5007.785 2365.270 5012.435 ;
      LAYER met4 ;
        RECT 2365.670 5007.385 2442.330 5012.835 ;
      LAYER met4 ;
        RECT 2442.730 5007.785 2622.270 5012.435 ;
      LAYER met4 ;
        RECT 2622.670 5007.385 2699.330 5012.835 ;
      LAYER met4 ;
        RECT 2699.730 5007.785 2879.270 5012.435 ;
      LAYER met4 ;
        RECT 2879.670 5007.385 2951.330 5012.835 ;
      LAYER met4 ;
        RECT 2951.730 5007.785 3131.270 5012.435 ;
      LAYER met4 ;
        RECT 3131.670 5007.385 3208.330 5012.835 ;
      LAYER met4 ;
        RECT 3208.730 5007.785 3389.525 5012.435 ;
      LAYER met4 ;
        RECT 3389.925 5011.575 3588.000 5012.835 ;
        RECT 3389.925 5011.310 3444.005 5011.575 ;
        RECT 3389.925 5007.975 3440.725 5011.310 ;
        RECT 3389.925 5007.385 3435.335 5007.975 ;
        RECT 152.665 5006.785 202.745 5007.385 ;
        RECT 381.965 5006.785 459.970 5007.385 ;
        RECT 638.965 5006.785 716.970 5007.385 ;
        RECT 895.965 5006.785 973.970 5007.385 ;
        RECT 1152.965 5006.785 1230.970 5007.385 ;
        RECT 1410.965 5006.785 1488.970 5007.385 ;
        RECT 1667.965 5006.785 1741.035 5007.385 ;
        RECT 1919.965 5006.785 1997.970 5007.385 ;
        RECT 2364.965 5006.785 2442.970 5007.385 ;
        RECT 2621.965 5006.785 2699.970 5007.385 ;
        RECT 2878.965 5006.785 2952.035 5007.385 ;
        RECT 3130.965 5006.785 3208.970 5007.385 ;
        RECT 3388.000 5006.785 3435.335 5007.385 ;
        RECT 152.665 5002.535 202.345 5006.785 ;
      LAYER met4 ;
        RECT 202.745 5002.935 381.965 5006.385 ;
      LAYER met4 ;
        RECT 382.365 5002.535 459.570 5006.785 ;
      LAYER met4 ;
        RECT 459.970 5002.935 638.965 5006.385 ;
      LAYER met4 ;
        RECT 639.365 5002.535 716.570 5006.785 ;
      LAYER met4 ;
        RECT 716.970 5002.935 895.965 5006.385 ;
      LAYER met4 ;
        RECT 896.365 5002.535 973.570 5006.785 ;
      LAYER met4 ;
        RECT 973.970 5002.935 1152.965 5006.385 ;
      LAYER met4 ;
        RECT 1153.365 5002.535 1230.570 5006.785 ;
      LAYER met4 ;
        RECT 1230.970 5002.935 1410.965 5006.385 ;
      LAYER met4 ;
        RECT 1411.365 5002.535 1488.570 5006.785 ;
      LAYER met4 ;
        RECT 1488.970 5002.935 1667.965 5006.385 ;
      LAYER met4 ;
        RECT 1668.365 5002.535 1740.635 5006.785 ;
      LAYER met4 ;
        RECT 1741.035 5002.935 1919.965 5006.385 ;
      LAYER met4 ;
        RECT 1920.365 5002.535 1997.570 5006.785 ;
      LAYER met4 ;
        RECT 1997.970 5002.935 2176.000 5006.385 ;
        RECT 2181.000 5002.935 2364.965 5006.385 ;
      LAYER met4 ;
        RECT 2365.365 5002.535 2442.570 5006.785 ;
      LAYER met4 ;
        RECT 2442.970 5002.935 2621.965 5006.385 ;
      LAYER met4 ;
        RECT 2622.365 5002.535 2699.570 5006.785 ;
      LAYER met4 ;
        RECT 2699.970 5002.935 2878.965 5006.385 ;
      LAYER met4 ;
        RECT 2879.365 5002.535 2951.635 5006.785 ;
      LAYER met4 ;
        RECT 2952.035 5002.935 3130.965 5006.385 ;
      LAYER met4 ;
        RECT 3131.365 5002.535 3208.570 5006.785 ;
      LAYER met4 ;
        RECT 3208.970 5002.935 3389.470 5006.385 ;
      LAYER met4 ;
        RECT 3389.870 5002.535 3435.335 5006.785 ;
        RECT 152.665 5001.935 202.745 5002.535 ;
        RECT 381.965 5001.935 459.970 5002.535 ;
        RECT 638.965 5001.935 716.970 5002.535 ;
        RECT 895.965 5001.935 973.970 5002.535 ;
        RECT 1152.965 5001.935 1230.970 5002.535 ;
        RECT 1410.965 5001.935 1488.970 5002.535 ;
        RECT 1667.965 5001.935 1741.035 5002.535 ;
        RECT 1919.965 5001.935 1997.970 5002.535 ;
        RECT 2364.965 5001.935 2442.970 5002.535 ;
        RECT 2621.965 5001.935 2699.970 5002.535 ;
        RECT 2878.965 5001.935 2952.035 5002.535 ;
        RECT 3130.965 5001.935 3208.970 5002.535 ;
        RECT 3388.000 5001.935 3435.335 5002.535 ;
        RECT 152.665 4996.485 202.330 5001.935 ;
      LAYER met4 ;
        RECT 202.730 4996.885 382.270 5001.535 ;
      LAYER met4 ;
        RECT 382.670 4996.485 459.330 5001.935 ;
      LAYER met4 ;
        RECT 459.730 4996.885 639.270 5001.535 ;
      LAYER met4 ;
        RECT 639.670 4996.485 716.330 5001.935 ;
      LAYER met4 ;
        RECT 716.730 4996.885 896.270 5001.535 ;
      LAYER met4 ;
        RECT 896.670 4996.485 973.330 5001.935 ;
      LAYER met4 ;
        RECT 973.730 4996.885 1153.270 5001.535 ;
      LAYER met4 ;
        RECT 1153.670 4996.485 1230.330 5001.935 ;
      LAYER met4 ;
        RECT 1230.730 4996.885 1411.270 5001.535 ;
      LAYER met4 ;
        RECT 1411.670 4996.485 1488.330 5001.935 ;
      LAYER met4 ;
        RECT 1488.730 4996.885 1668.270 5001.535 ;
      LAYER met4 ;
        RECT 1668.670 4996.485 1740.330 5001.935 ;
      LAYER met4 ;
        RECT 1740.730 4996.885 1920.270 5001.535 ;
      LAYER met4 ;
        RECT 1920.670 4996.485 1997.330 5001.935 ;
      LAYER met4 ;
        RECT 1997.730 4996.885 2181.000 5001.535 ;
        RECT 2186.000 4996.885 2365.270 5001.535 ;
      LAYER met4 ;
        RECT 2365.670 4996.485 2442.330 5001.935 ;
      LAYER met4 ;
        RECT 2442.730 4996.885 2622.270 5001.535 ;
      LAYER met4 ;
        RECT 2622.670 4996.485 2699.330 5001.935 ;
      LAYER met4 ;
        RECT 2699.730 4996.885 2879.270 5001.535 ;
      LAYER met4 ;
        RECT 2879.670 4996.485 2951.330 5001.935 ;
      LAYER met4 ;
        RECT 2951.730 4996.885 3131.270 5001.535 ;
      LAYER met4 ;
        RECT 3131.670 4996.485 3208.330 5001.935 ;
      LAYER met4 ;
        RECT 3208.730 4996.885 3391.785 5001.535 ;
      LAYER met4 ;
        RECT 3392.185 4996.485 3435.335 5001.935 ;
        RECT 152.665 4995.885 202.745 4996.485 ;
        RECT 381.965 4995.885 459.970 4996.485 ;
        RECT 638.965 4995.885 716.970 4996.485 ;
        RECT 895.965 4995.885 973.970 4996.485 ;
        RECT 1152.965 4995.885 1230.970 4996.485 ;
        RECT 1410.965 4995.885 1488.970 4996.485 ;
        RECT 1667.965 4995.885 1741.035 4996.485 ;
        RECT 1919.965 4995.885 1997.970 4996.485 ;
        RECT 2364.965 4995.885 2442.970 4996.485 ;
        RECT 2621.965 4995.885 2699.970 4996.485 ;
        RECT 2878.965 4995.885 2952.035 4996.485 ;
        RECT 3130.965 4995.885 3208.970 4996.485 ;
        RECT 3388.000 4995.885 3435.335 4996.485 ;
        RECT 152.665 4992.185 202.330 4995.885 ;
        RECT 152.665 4990.000 186.065 4992.185 ;
        RECT 152.665 4989.875 169.115 4990.000 ;
        RECT 152.665 4988.000 153.365 4989.875 ;
        RECT 158.815 4989.785 169.115 4989.875 ;
        RECT 158.815 4989.735 164.265 4989.785 ;
        RECT 152.665 4849.330 153.365 4849.970 ;
      LAYER met4 ;
        RECT 153.765 4849.730 158.415 4989.475 ;
      LAYER met4 ;
        RECT 158.815 4988.000 159.415 4989.735 ;
        RECT 158.815 4849.330 159.415 4849.970 ;
      LAYER met4 ;
        RECT 159.815 4849.730 163.265 4989.335 ;
      LAYER met4 ;
        RECT 163.665 4988.000 164.265 4989.735 ;
        RECT 163.665 4849.330 164.265 4849.970 ;
      LAYER met4 ;
        RECT 164.665 4849.730 168.115 4989.385 ;
      LAYER met4 ;
        RECT 168.515 4988.000 169.115 4989.785 ;
        RECT 174.565 4989.925 186.065 4990.000 ;
        RECT 168.515 4849.330 169.115 4849.970 ;
      LAYER met4 ;
        RECT 169.515 4849.730 174.165 4989.600 ;
      LAYER met4 ;
        RECT 174.565 4988.000 175.165 4989.925 ;
        RECT 180.615 4989.870 186.065 4989.925 ;
        RECT 174.565 4849.330 175.165 4849.970 ;
      LAYER met4 ;
        RECT 175.565 4849.730 180.215 4989.525 ;
      LAYER met4 ;
        RECT 180.615 4988.000 181.215 4989.870 ;
      LAYER met4 ;
        RECT 181.615 4849.970 185.065 4989.470 ;
      LAYER met4 ;
        RECT 185.465 4988.000 186.065 4989.870 ;
        RECT 180.615 4849.570 181.215 4849.970 ;
        RECT 185.465 4849.570 186.065 4849.970 ;
      LAYER met4 ;
        RECT 186.465 4849.730 191.115 4991.785 ;
      LAYER met4 ;
        RECT 191.515 4990.750 202.330 4992.185 ;
        RECT 191.515 4988.000 192.115 4990.750 ;
        RECT 180.615 4849.330 186.065 4849.570 ;
        RECT 191.515 4849.330 192.115 4849.970 ;
      LAYER met4 ;
        RECT 192.515 4849.730 197.965 4990.350 ;
      LAYER met4 ;
        RECT 198.365 4990.035 202.330 4990.750 ;
      LAYER met4 ;
        RECT 202.730 4990.035 382.270 4995.485 ;
      LAYER met4 ;
        RECT 197.965 4989.635 202.330 4990.035 ;
        RECT 382.670 4989.635 459.330 4995.885 ;
      LAYER met4 ;
        RECT 459.730 4990.035 639.270 4995.485 ;
      LAYER met4 ;
        RECT 639.670 4989.635 716.330 4995.885 ;
      LAYER met4 ;
        RECT 716.730 4990.035 896.270 4995.485 ;
      LAYER met4 ;
        RECT 896.670 4989.635 973.330 4995.885 ;
      LAYER met4 ;
        RECT 973.730 4990.035 1153.270 4995.485 ;
      LAYER met4 ;
        RECT 1153.670 4989.635 1230.330 4995.885 ;
      LAYER met4 ;
        RECT 1230.730 4990.035 1411.270 4995.485 ;
      LAYER met4 ;
        RECT 1411.670 4989.635 1488.330 4995.885 ;
      LAYER met4 ;
        RECT 1488.730 4990.035 1668.270 4995.485 ;
      LAYER met4 ;
        RECT 1668.670 4990.035 1740.330 4995.885 ;
      LAYER met4 ;
        RECT 1740.730 4990.035 1920.270 4995.485 ;
      LAYER met4 ;
        RECT 1920.670 4989.635 1997.330 4995.885 ;
      LAYER met4 ;
        RECT 1997.730 4990.035 2365.270 4995.485 ;
      LAYER met4 ;
        RECT 2365.670 4989.635 2442.330 4995.885 ;
      LAYER met4 ;
        RECT 2442.730 4990.035 2622.270 4995.485 ;
      LAYER met4 ;
        RECT 2622.670 4989.635 2699.330 4995.885 ;
      LAYER met4 ;
        RECT 2699.730 4990.035 2879.270 4995.485 ;
      LAYER met4 ;
        RECT 2879.670 4990.035 2951.330 4995.885 ;
      LAYER met4 ;
        RECT 2951.730 4990.035 3131.270 4995.485 ;
      LAYER met4 ;
        RECT 3131.670 4989.635 3208.330 4995.885 ;
      LAYER met4 ;
        RECT 3208.730 4990.035 3390.350 4995.485 ;
      LAYER met4 ;
        POLYGON 3388.000 4990.035 3388.400 4990.035 3388.400 4989.635 ;
        RECT 3388.400 4989.635 3390.035 4990.035 ;
        RECT 3390.750 4989.635 3435.335 4995.885 ;
        RECT 197.965 4988.400 202.745 4989.635 ;
        RECT 381.965 4988.535 459.970 4989.635 ;
        RECT 638.965 4988.535 716.970 4989.635 ;
        RECT 895.965 4988.535 973.970 4989.635 ;
        RECT 1152.965 4988.535 1230.970 4989.635 ;
        RECT 1410.965 4988.535 1488.970 4989.635 ;
        RECT 1919.965 4988.535 1997.970 4989.635 ;
        RECT 2364.965 4988.535 2442.970 4989.635 ;
        RECT 2621.965 4988.535 2699.970 4989.635 ;
        RECT 3130.965 4988.535 3208.970 4989.635 ;
        POLYGON 197.965 4988.400 198.365 4988.400 197.965 4988.000 ;
        RECT 198.365 4988.000 202.745 4988.400 ;
        RECT 3388.000 4985.670 3435.335 4989.635 ;
        RECT 3388.000 4985.255 3389.635 4985.670 ;
        RECT 198.365 4849.330 199.465 4849.970 ;
        RECT 152.665 4817.690 199.465 4849.330 ;
        RECT 152.035 4774.010 199.465 4817.690 ;
        RECT 152.665 4772.670 199.465 4774.010 ;
        RECT 152.665 4771.965 153.365 4772.670 ;
        RECT 152.665 4633.330 153.365 4635.000 ;
      LAYER met4 ;
        RECT 153.765 4633.730 158.415 4772.270 ;
      LAYER met4 ;
        RECT 158.815 4771.965 159.415 4772.670 ;
        RECT 158.815 4633.330 159.415 4635.000 ;
      LAYER met4 ;
        RECT 159.815 4633.730 163.265 4772.270 ;
      LAYER met4 ;
        RECT 163.665 4771.965 164.265 4772.670 ;
        RECT 163.665 4633.330 164.265 4635.000 ;
      LAYER met4 ;
        RECT 164.665 4633.730 168.115 4772.270 ;
      LAYER met4 ;
        RECT 168.515 4771.965 169.115 4772.670 ;
        RECT 168.515 4633.330 169.115 4635.000 ;
      LAYER met4 ;
        RECT 169.515 4633.730 174.165 4772.270 ;
      LAYER met4 ;
        RECT 174.565 4771.965 175.165 4772.670 ;
        RECT 180.615 4772.365 186.065 4772.670 ;
        RECT 174.565 4633.330 175.165 4635.000 ;
      LAYER met4 ;
        RECT 175.565 4633.730 180.215 4772.270 ;
      LAYER met4 ;
        RECT 180.615 4771.965 181.215 4772.365 ;
        RECT 185.465 4771.965 186.065 4772.365 ;
        RECT 191.515 4771.965 192.115 4772.670 ;
        RECT 180.615 4633.635 181.215 4635.000 ;
      LAYER met4 ;
        RECT 181.615 4634.035 185.065 4771.965 ;
      LAYER met4 ;
        RECT 185.465 4633.635 186.065 4635.000 ;
        RECT 180.615 4633.330 186.065 4633.635 ;
        RECT 191.515 4633.330 192.115 4635.000 ;
      LAYER met4 ;
        RECT 192.515 4633.730 197.965 4772.270 ;
      LAYER met4 ;
        RECT 198.365 4771.965 199.465 4772.670 ;
        RECT 3388.535 4836.330 3389.635 4837.035 ;
      LAYER met4 ;
        RECT 3390.035 4836.730 3395.485 4985.270 ;
      LAYER met4 ;
        RECT 3395.885 4985.255 3396.485 4985.670 ;
        RECT 3401.935 4985.655 3407.385 4985.670 ;
        RECT 3395.885 4836.330 3396.485 4837.035 ;
      LAYER met4 ;
        RECT 3396.885 4836.730 3401.535 4985.270 ;
      LAYER met4 ;
        RECT 3401.935 4985.255 3402.535 4985.655 ;
        RECT 3406.785 4985.255 3407.385 4985.655 ;
      LAYER met4 ;
        RECT 3402.935 4837.035 3406.385 4985.255 ;
      LAYER met4 ;
        RECT 3401.935 4836.635 3402.535 4837.035 ;
        RECT 3406.785 4836.635 3407.385 4837.035 ;
      LAYER met4 ;
        RECT 3407.785 4836.730 3412.435 4985.270 ;
      LAYER met4 ;
        RECT 3412.835 4985.255 3413.435 4985.670 ;
        RECT 3401.935 4836.330 3407.385 4836.635 ;
        RECT 3412.835 4836.330 3413.435 4837.035 ;
      LAYER met4 ;
        RECT 3413.835 4836.730 3418.485 4985.270 ;
      LAYER met4 ;
        RECT 3418.885 4985.255 3419.485 4985.670 ;
        RECT 3418.885 4836.330 3419.485 4837.035 ;
      LAYER met4 ;
        RECT 3419.885 4836.730 3423.335 4985.270 ;
      LAYER met4 ;
        RECT 3423.735 4985.255 3424.335 4985.670 ;
        RECT 3423.735 4836.330 3424.335 4837.035 ;
      LAYER met4 ;
        RECT 3424.735 4836.730 3428.185 4985.270 ;
      LAYER met4 ;
        RECT 3428.585 4985.255 3429.185 4985.670 ;
        RECT 3428.585 4836.330 3429.185 4837.035 ;
      LAYER met4 ;
        RECT 3429.585 4836.730 3434.235 4985.270 ;
      LAYER met4 ;
        RECT 3434.635 4985.255 3435.335 4985.670 ;
        RECT 3434.635 4836.330 3435.335 4837.035 ;
        RECT 3388.535 4834.990 3435.335 4836.330 ;
      LAYER met4 ;
        RECT 3435.735 4835.390 3436.065 5007.575 ;
      LAYER met4 ;
        RECT 3436.465 5005.955 3440.725 5007.975 ;
        RECT 3436.465 5005.275 3439.245 5005.955 ;
        RECT 3388.535 4791.310 3435.965 4834.990 ;
        RECT 3388.535 4759.670 3435.335 4791.310 ;
        RECT 3388.535 4759.030 3389.635 4759.670 ;
        RECT 152.665 4561.670 197.965 4633.330 ;
      LAYER met4 ;
        RECT 3390.035 4611.730 3395.485 4759.270 ;
      LAYER met4 ;
        RECT 3395.885 4759.030 3396.485 4759.670 ;
        RECT 3401.935 4759.430 3407.385 4759.670 ;
        RECT 3401.935 4759.030 3402.535 4759.430 ;
        RECT 3406.785 4759.030 3407.385 4759.430 ;
      LAYER met4 ;
        RECT 3402.935 4612.035 3406.385 4759.030 ;
      LAYER met4 ;
        RECT 3395.885 4611.330 3396.485 4612.035 ;
        RECT 3401.935 4611.635 3402.535 4612.035 ;
        RECT 3406.785 4611.635 3407.385 4612.035 ;
      LAYER met4 ;
        RECT 3407.785 4611.730 3412.435 4759.270 ;
      LAYER met4 ;
        RECT 3412.835 4759.030 3413.435 4759.670 ;
        RECT 3401.935 4611.330 3407.385 4611.635 ;
        RECT 3412.835 4611.330 3413.435 4612.035 ;
      LAYER met4 ;
        RECT 3413.835 4611.730 3418.485 4759.270 ;
      LAYER met4 ;
        RECT 3418.885 4759.030 3419.485 4759.670 ;
        RECT 3418.885 4611.330 3419.485 4612.035 ;
      LAYER met4 ;
        RECT 3419.885 4611.730 3423.335 4759.270 ;
      LAYER met4 ;
        RECT 3423.735 4759.030 3424.335 4759.670 ;
        RECT 3423.735 4611.330 3424.335 4612.035 ;
      LAYER met4 ;
        RECT 3424.735 4611.730 3428.185 4759.270 ;
      LAYER met4 ;
        RECT 3428.585 4759.030 3429.185 4759.670 ;
        RECT 3428.585 4611.330 3429.185 4612.035 ;
      LAYER met4 ;
        RECT 3429.585 4611.730 3434.235 4759.270 ;
      LAYER met4 ;
        RECT 3434.635 4759.030 3435.335 4759.670 ;
        RECT 3434.635 4611.330 3435.335 4612.035 ;
        RECT 152.665 4560.965 153.365 4561.670 ;
        RECT 152.665 4422.330 153.365 4423.035 ;
      LAYER met4 ;
        RECT 153.765 4422.730 158.415 4561.270 ;
      LAYER met4 ;
        RECT 158.815 4560.965 159.415 4561.670 ;
        RECT 158.815 4422.330 159.415 4423.035 ;
      LAYER met4 ;
        RECT 159.815 4422.730 163.265 4561.270 ;
      LAYER met4 ;
        RECT 163.665 4560.965 164.265 4561.670 ;
        RECT 163.665 4422.330 164.265 4423.035 ;
      LAYER met4 ;
        RECT 164.665 4422.730 168.115 4561.270 ;
      LAYER met4 ;
        RECT 168.515 4560.965 169.115 4561.670 ;
        RECT 168.515 4422.330 169.115 4423.035 ;
      LAYER met4 ;
        RECT 169.515 4422.730 174.165 4561.270 ;
      LAYER met4 ;
        RECT 174.565 4560.965 175.165 4561.670 ;
        RECT 180.615 4561.365 186.065 4561.670 ;
        RECT 174.565 4422.330 175.165 4423.035 ;
      LAYER met4 ;
        RECT 175.565 4422.730 180.215 4561.270 ;
      LAYER met4 ;
        RECT 180.615 4560.965 181.215 4561.365 ;
        RECT 185.465 4560.965 186.065 4561.365 ;
        RECT 191.515 4560.965 192.115 4561.670 ;
      LAYER met4 ;
        RECT 181.615 4423.035 185.065 4560.965 ;
      LAYER met4 ;
        RECT 180.615 4422.635 181.215 4423.035 ;
        RECT 185.465 4422.635 186.065 4423.035 ;
        RECT 180.615 4422.330 186.065 4422.635 ;
        RECT 191.515 4422.330 192.115 4423.035 ;
      LAYER met4 ;
        RECT 192.515 4422.730 197.965 4561.270 ;
      LAYER met4 ;
        RECT 3390.035 4539.670 3435.335 4611.330 ;
        RECT 152.665 4350.670 197.965 4422.330 ;
        RECT 3388.535 4390.330 3389.635 4391.035 ;
      LAYER met4 ;
        RECT 3390.035 4390.730 3395.485 4539.270 ;
      LAYER met4 ;
        RECT 3395.885 4538.000 3396.485 4539.670 ;
        RECT 3401.935 4539.365 3407.385 4539.670 ;
        RECT 3401.935 4538.000 3402.535 4539.365 ;
      LAYER met4 ;
        RECT 3402.935 4391.035 3406.385 4538.965 ;
      LAYER met4 ;
        RECT 3406.785 4538.000 3407.385 4539.365 ;
        RECT 3395.885 4390.330 3396.485 4391.035 ;
        RECT 3401.935 4390.635 3402.535 4391.035 ;
        RECT 3406.785 4390.635 3407.385 4391.035 ;
      LAYER met4 ;
        RECT 3407.785 4390.730 3412.435 4539.270 ;
      LAYER met4 ;
        RECT 3412.835 4538.000 3413.435 4539.670 ;
        RECT 3401.935 4390.330 3407.385 4390.635 ;
        RECT 3412.835 4390.330 3413.435 4391.035 ;
      LAYER met4 ;
        RECT 3413.835 4390.730 3418.485 4539.270 ;
      LAYER met4 ;
        RECT 3418.885 4538.000 3419.485 4539.670 ;
        RECT 3418.885 4390.330 3419.485 4391.035 ;
      LAYER met4 ;
        RECT 3419.885 4390.730 3423.335 4539.270 ;
      LAYER met4 ;
        RECT 3423.735 4538.000 3424.335 4539.670 ;
        RECT 3423.735 4390.330 3424.335 4391.035 ;
      LAYER met4 ;
        RECT 3424.735 4390.730 3428.185 4539.270 ;
      LAYER met4 ;
        RECT 3428.585 4538.000 3429.185 4539.670 ;
        RECT 3428.585 4390.330 3429.185 4391.035 ;
      LAYER met4 ;
        RECT 3429.585 4390.730 3434.235 4539.270 ;
      LAYER met4 ;
        RECT 3434.635 4538.000 3435.335 4539.670 ;
        RECT 3434.635 4390.330 3435.335 4391.035 ;
        RECT 3388.535 4388.990 3435.335 4390.330 ;
      LAYER met4 ;
        RECT 3435.735 4389.390 3436.065 4790.910 ;
        RECT 3436.365 4785.855 3439.345 5004.875 ;
        RECT 3439.645 4984.000 3440.825 5005.555 ;
      LAYER met4 ;
        RECT 3439.745 4838.000 3440.725 4984.000 ;
      LAYER met4 ;
        RECT 3439.645 4836.730 3440.825 4838.000 ;
      LAYER met4 ;
        RECT 3439.745 4801.160 3440.725 4836.330 ;
      LAYER met4 ;
        RECT 3441.125 4801.560 3444.105 5010.910 ;
        RECT 3444.405 4835.390 3444.735 5011.175 ;
      LAYER met4 ;
        RECT 3445.135 4986.255 3588.000 5011.575 ;
        RECT 3445.135 4985.670 3457.635 4986.255 ;
        RECT 3445.135 4985.255 3445.835 4985.670 ;
        RECT 3445.135 4838.000 3445.835 4984.000 ;
        RECT 3445.135 4836.330 3445.835 4837.035 ;
      LAYER met4 ;
        RECT 3446.235 4836.730 3450.685 4985.270 ;
      LAYER met4 ;
        RECT 3451.085 4985.255 3451.685 4985.670 ;
        RECT 3451.085 4838.000 3451.685 4983.000 ;
        RECT 3451.085 4836.330 3451.685 4837.035 ;
      LAYER met4 ;
        RECT 3452.085 4836.730 3456.535 4985.270 ;
      LAYER met4 ;
        RECT 3456.935 4985.255 3457.635 4985.670 ;
        RECT 3456.935 4982.000 3458.035 4984.000 ;
      LAYER met4 ;
        RECT 3458.035 4982.000 3483.000 4985.855 ;
      LAYER met4 ;
        RECT 3483.400 4985.670 3588.000 4986.255 ;
        RECT 3483.400 4985.255 3563.385 4985.670 ;
      LAYER met4 ;
        RECT 3563.785 4984.000 3588.000 4985.270 ;
      LAYER met4 ;
        RECT 3483.000 4982.000 3485.035 4984.000 ;
        RECT 3456.935 4979.000 3485.035 4982.000 ;
        RECT 3456.935 4977.000 3458.035 4979.000 ;
      LAYER met4 ;
        RECT 3458.035 4977.000 3483.000 4979.000 ;
      LAYER met4 ;
        RECT 3483.000 4977.000 3485.035 4979.000 ;
        RECT 3456.935 4959.000 3485.035 4977.000 ;
        RECT 3456.935 4957.000 3458.035 4959.000 ;
      LAYER met4 ;
        RECT 3458.035 4957.000 3483.000 4959.000 ;
      LAYER met4 ;
        RECT 3483.000 4957.000 3485.035 4959.000 ;
        RECT 3456.935 4939.000 3485.035 4957.000 ;
        RECT 3456.935 4937.000 3458.035 4939.000 ;
      LAYER met4 ;
        RECT 3458.035 4937.000 3483.000 4939.000 ;
      LAYER met4 ;
        RECT 3483.000 4937.000 3485.035 4939.000 ;
        RECT 3456.935 4919.000 3485.035 4937.000 ;
        RECT 3456.935 4917.000 3458.035 4919.000 ;
      LAYER met4 ;
        RECT 3458.035 4917.000 3483.000 4919.000 ;
      LAYER met4 ;
        RECT 3483.000 4917.000 3485.035 4919.000 ;
        RECT 3456.935 4899.000 3485.035 4917.000 ;
        RECT 3456.935 4897.000 3458.035 4899.000 ;
      LAYER met4 ;
        RECT 3458.035 4897.000 3483.000 4899.000 ;
      LAYER met4 ;
        RECT 3483.000 4897.000 3485.035 4899.000 ;
        RECT 3456.935 4879.000 3485.035 4897.000 ;
        RECT 3456.935 4877.000 3458.035 4879.000 ;
      LAYER met4 ;
        RECT 3458.035 4877.000 3483.000 4879.000 ;
      LAYER met4 ;
        RECT 3483.000 4877.000 3485.035 4879.000 ;
        RECT 3456.935 4859.000 3485.035 4877.000 ;
        RECT 3456.935 4857.000 3458.035 4859.000 ;
      LAYER met4 ;
        RECT 3458.035 4857.000 3483.000 4859.000 ;
      LAYER met4 ;
        RECT 3483.000 4857.000 3485.035 4859.000 ;
        RECT 3456.935 4839.000 3485.035 4857.000 ;
        RECT 3456.935 4838.000 3458.035 4839.000 ;
        RECT 3456.935 4836.330 3457.635 4837.035 ;
      LAYER met4 ;
        RECT 3458.035 4836.730 3483.000 4839.000 ;
      LAYER met4 ;
        RECT 3483.000 4838.000 3485.035 4839.000 ;
        RECT 3562.035 4838.000 3588.000 4984.000 ;
        RECT 3483.400 4836.330 3563.385 4837.035 ;
      LAYER met4 ;
        RECT 3563.785 4836.730 3588.000 4838.000 ;
      LAYER met4 ;
        RECT 3445.135 4834.990 3588.000 4836.330 ;
        RECT 3444.505 4801.160 3588.000 4834.990 ;
        RECT 3439.745 4799.640 3588.000 4801.160 ;
        RECT 3439.745 4785.455 3440.725 4799.640 ;
        RECT 3436.465 4783.935 3440.725 4785.455 ;
        RECT 152.665 4349.965 153.365 4350.670 ;
        RECT 152.665 4211.330 153.365 4212.035 ;
      LAYER met4 ;
        RECT 153.765 4211.730 158.415 4350.270 ;
      LAYER met4 ;
        RECT 158.815 4349.965 159.415 4350.670 ;
        RECT 163.665 4349.965 164.265 4350.670 ;
        RECT 158.815 4211.330 159.415 4212.035 ;
        RECT 163.665 4211.330 164.265 4212.035 ;
      LAYER met4 ;
        RECT 164.665 4211.730 168.115 4350.270 ;
      LAYER met4 ;
        RECT 168.515 4349.965 169.115 4350.670 ;
        RECT 168.515 4211.330 169.115 4212.035 ;
      LAYER met4 ;
        RECT 169.515 4211.730 174.165 4350.270 ;
      LAYER met4 ;
        RECT 174.565 4349.965 175.165 4350.670 ;
        RECT 180.615 4350.365 186.065 4350.670 ;
        RECT 174.565 4211.330 175.165 4212.035 ;
      LAYER met4 ;
        RECT 175.565 4211.730 180.215 4350.270 ;
      LAYER met4 ;
        RECT 180.615 4349.965 181.215 4350.365 ;
        RECT 185.465 4349.965 186.065 4350.365 ;
      LAYER met4 ;
        RECT 181.615 4212.035 185.065 4349.965 ;
      LAYER met4 ;
        RECT 180.615 4211.635 181.215 4212.035 ;
        RECT 185.465 4211.635 186.065 4212.035 ;
      LAYER met4 ;
        RECT 186.465 4211.730 191.115 4350.270 ;
      LAYER met4 ;
        RECT 191.515 4349.965 192.115 4350.670 ;
        RECT 180.615 4211.330 186.065 4211.635 ;
        RECT 191.515 4211.330 192.115 4212.035 ;
      LAYER met4 ;
        RECT 192.515 4211.730 197.965 4350.270 ;
      LAYER met4 ;
        RECT 3388.535 4345.310 3435.965 4388.990 ;
        RECT 3388.535 4313.670 3435.335 4345.310 ;
        RECT 3388.535 4313.030 3389.635 4313.670 ;
        RECT 152.035 4139.670 197.965 4211.330 ;
      LAYER met4 ;
        RECT 3390.035 4165.730 3395.485 4313.270 ;
      LAYER met4 ;
        RECT 3395.885 4313.030 3396.485 4313.670 ;
        RECT 3401.935 4313.430 3407.385 4313.670 ;
        RECT 3395.885 4165.330 3396.485 4166.035 ;
      LAYER met4 ;
        RECT 3396.885 4165.730 3401.535 4313.270 ;
      LAYER met4 ;
        RECT 3401.935 4313.030 3402.535 4313.430 ;
        RECT 3406.785 4313.030 3407.385 4313.430 ;
        RECT 3401.935 4165.635 3402.535 4166.035 ;
        RECT 3406.785 4165.635 3407.385 4166.035 ;
      LAYER met4 ;
        RECT 3407.785 4165.730 3412.435 4313.270 ;
      LAYER met4 ;
        RECT 3412.835 4313.030 3413.435 4313.670 ;
        RECT 3401.935 4165.330 3407.385 4165.635 ;
        RECT 3412.835 4165.330 3413.435 4166.035 ;
      LAYER met4 ;
        RECT 3413.835 4165.730 3418.485 4313.270 ;
      LAYER met4 ;
        RECT 3418.885 4313.030 3419.485 4313.670 ;
        RECT 3418.885 4165.330 3419.485 4166.035 ;
      LAYER met4 ;
        RECT 3419.885 4165.730 3423.335 4313.270 ;
      LAYER met4 ;
        RECT 3423.735 4313.030 3424.335 4313.670 ;
        RECT 3423.735 4165.330 3424.335 4166.035 ;
      LAYER met4 ;
        RECT 3424.735 4165.730 3428.185 4313.270 ;
      LAYER met4 ;
        RECT 3428.585 4313.030 3429.185 4313.670 ;
        RECT 3428.585 4165.330 3429.185 4166.035 ;
      LAYER met4 ;
        RECT 3429.585 4165.730 3434.235 4313.270 ;
      LAYER met4 ;
        RECT 3434.635 4313.030 3435.335 4313.670 ;
        RECT 3434.635 4165.330 3435.335 4166.035 ;
        RECT 152.665 4138.965 153.365 4139.670 ;
        RECT 152.665 4000.330 153.365 4000.970 ;
      LAYER met4 ;
        RECT 153.765 4000.730 158.415 4139.270 ;
      LAYER met4 ;
        RECT 158.815 4138.965 159.415 4139.670 ;
        RECT 163.665 4138.965 164.265 4139.670 ;
        RECT 158.815 4000.330 159.415 4000.970 ;
        RECT 163.665 4000.330 164.265 4000.970 ;
      LAYER met4 ;
        RECT 164.665 4000.730 168.115 4139.270 ;
      LAYER met4 ;
        RECT 168.515 4138.965 169.115 4139.670 ;
        RECT 168.515 4000.330 169.115 4000.970 ;
      LAYER met4 ;
        RECT 169.515 4000.730 174.165 4139.270 ;
      LAYER met4 ;
        RECT 174.565 4138.965 175.165 4139.670 ;
        RECT 180.615 4139.365 186.065 4139.670 ;
        RECT 174.565 4000.330 175.165 4000.970 ;
      LAYER met4 ;
        RECT 175.565 4000.730 180.215 4139.270 ;
      LAYER met4 ;
        RECT 180.615 4138.965 181.215 4139.365 ;
        RECT 185.465 4138.965 186.065 4139.365 ;
      LAYER met4 ;
        RECT 181.615 4000.970 185.065 4138.965 ;
      LAYER met4 ;
        RECT 180.615 4000.570 181.215 4000.970 ;
        RECT 185.465 4000.570 186.065 4000.970 ;
      LAYER met4 ;
        RECT 186.465 4000.730 191.115 4139.270 ;
      LAYER met4 ;
        RECT 191.515 4138.965 192.115 4139.670 ;
        RECT 180.615 4000.330 186.065 4000.570 ;
        RECT 191.515 4000.330 192.115 4000.970 ;
      LAYER met4 ;
        RECT 192.515 4000.730 197.965 4139.270 ;
      LAYER met4 ;
        RECT 3390.035 4093.670 3435.335 4165.330 ;
        RECT 198.365 4000.330 199.465 4000.970 ;
        RECT 147.275 3974.545 151.535 3976.065 ;
        RECT 147.275 3960.360 148.255 3974.545 ;
        RECT 0.000 3958.840 148.255 3960.360 ;
        RECT 0.000 3925.010 143.495 3958.840 ;
        RECT 0.000 3923.670 142.865 3925.010 ;
      LAYER met4 ;
        RECT 0.000 3922.000 24.215 3923.270 ;
      LAYER met4 ;
        RECT 24.615 3922.965 104.600 3923.670 ;
        RECT 0.000 3786.000 25.965 3922.000 ;
        RECT 102.965 3920.000 105.000 3922.000 ;
      LAYER met4 ;
        RECT 105.000 3920.000 129.965 3923.270 ;
      LAYER met4 ;
        RECT 130.365 3922.965 131.065 3923.670 ;
        RECT 129.965 3920.000 131.065 3922.000 ;
        RECT 102.965 3917.000 131.065 3920.000 ;
        RECT 102.965 3915.000 105.000 3917.000 ;
      LAYER met4 ;
        RECT 105.000 3915.000 129.965 3917.000 ;
      LAYER met4 ;
        RECT 129.965 3915.000 131.065 3917.000 ;
        RECT 102.965 3907.000 131.065 3915.000 ;
        RECT 102.965 3905.000 105.000 3907.000 ;
      LAYER met4 ;
        RECT 105.000 3905.000 129.965 3907.000 ;
      LAYER met4 ;
        RECT 129.965 3905.000 131.065 3907.000 ;
        RECT 102.965 3887.000 131.065 3905.000 ;
        RECT 102.965 3885.000 105.000 3887.000 ;
      LAYER met4 ;
        RECT 105.000 3885.000 129.965 3887.000 ;
      LAYER met4 ;
        RECT 129.965 3885.000 131.065 3887.000 ;
        RECT 102.965 3867.000 131.065 3885.000 ;
        RECT 102.965 3865.000 105.000 3867.000 ;
      LAYER met4 ;
        RECT 105.000 3865.000 129.965 3867.000 ;
      LAYER met4 ;
        RECT 129.965 3865.000 131.065 3867.000 ;
        RECT 102.965 3847.000 131.065 3865.000 ;
        RECT 102.965 3845.000 105.000 3847.000 ;
      LAYER met4 ;
        RECT 105.000 3845.000 129.965 3847.000 ;
      LAYER met4 ;
        RECT 129.965 3845.000 131.065 3847.000 ;
        RECT 102.965 3827.000 131.065 3845.000 ;
        RECT 102.965 3825.000 105.000 3827.000 ;
      LAYER met4 ;
        RECT 105.000 3825.000 129.965 3827.000 ;
      LAYER met4 ;
        RECT 129.965 3825.000 131.065 3827.000 ;
        RECT 102.965 3807.000 131.065 3825.000 ;
        RECT 102.965 3805.000 105.000 3807.000 ;
      LAYER met4 ;
        RECT 105.000 3805.000 129.965 3807.000 ;
      LAYER met4 ;
        RECT 129.965 3805.000 131.065 3807.000 ;
        RECT 102.965 3787.000 131.065 3805.000 ;
        RECT 102.965 3786.000 105.000 3787.000 ;
      LAYER met4 ;
        RECT 0.000 3784.730 24.215 3786.000 ;
      LAYER met4 ;
        RECT 24.615 3784.330 104.600 3784.970 ;
      LAYER met4 ;
        RECT 105.000 3784.730 129.965 3787.000 ;
      LAYER met4 ;
        RECT 129.965 3786.000 131.065 3787.000 ;
        RECT 130.365 3784.330 131.065 3784.970 ;
      LAYER met4 ;
        RECT 131.465 3784.730 135.915 3923.270 ;
      LAYER met4 ;
        RECT 136.315 3922.965 136.915 3923.670 ;
        RECT 136.315 3786.000 136.915 3921.000 ;
        RECT 136.315 3784.330 136.915 3784.970 ;
      LAYER met4 ;
        RECT 137.315 3784.730 141.765 3923.270 ;
      LAYER met4 ;
        RECT 142.165 3922.965 142.865 3923.670 ;
        RECT 142.165 3786.000 142.865 3922.000 ;
        RECT 142.165 3784.330 142.865 3784.970 ;
        RECT 0.000 3752.690 142.865 3784.330 ;
      LAYER met4 ;
        RECT 143.265 3753.090 143.595 3924.610 ;
      LAYER met4 ;
        RECT 0.000 3744.360 143.495 3752.690 ;
      LAYER met4 ;
        RECT 143.895 3744.760 146.875 3958.440 ;
      LAYER met4 ;
        RECT 147.275 3923.670 148.255 3958.840 ;
      LAYER met4 ;
        RECT 147.175 3922.000 148.355 3923.270 ;
      LAYER met4 ;
        RECT 147.275 3786.000 148.255 3922.000 ;
      LAYER met4 ;
        RECT 147.175 3784.730 148.355 3786.000 ;
      LAYER met4 ;
        RECT 147.275 3760.065 148.255 3784.330 ;
      LAYER met4 ;
        RECT 148.655 3760.465 151.635 3974.145 ;
      LAYER met4 ;
        RECT 152.665 3968.690 199.465 4000.330 ;
        RECT 152.035 3925.010 199.465 3968.690 ;
        RECT 147.275 3758.545 151.535 3760.065 ;
        RECT 147.275 3744.360 148.255 3758.545 ;
        RECT 0.000 3742.840 148.255 3744.360 ;
        RECT 0.000 3709.010 143.495 3742.840 ;
        RECT 0.000 3707.670 142.865 3709.010 ;
      LAYER met4 ;
        RECT 0.000 3706.000 24.215 3707.270 ;
      LAYER met4 ;
        RECT 24.615 3706.965 104.600 3707.670 ;
        RECT 0.000 3570.000 25.965 3706.000 ;
        RECT 102.965 3704.000 105.000 3706.000 ;
      LAYER met4 ;
        RECT 105.000 3704.000 129.965 3707.270 ;
      LAYER met4 ;
        RECT 130.365 3706.965 131.065 3707.670 ;
        RECT 129.965 3704.000 131.065 3706.000 ;
        RECT 102.965 3701.000 131.065 3704.000 ;
        RECT 102.965 3699.000 105.000 3701.000 ;
      LAYER met4 ;
        RECT 105.000 3699.000 129.965 3701.000 ;
      LAYER met4 ;
        RECT 129.965 3699.000 131.065 3701.000 ;
        RECT 102.965 3691.000 131.065 3699.000 ;
        RECT 102.965 3689.000 105.000 3691.000 ;
      LAYER met4 ;
        RECT 105.000 3689.000 129.965 3691.000 ;
      LAYER met4 ;
        RECT 129.965 3689.000 131.065 3691.000 ;
        RECT 102.965 3671.000 131.065 3689.000 ;
        RECT 102.965 3669.000 105.000 3671.000 ;
      LAYER met4 ;
        RECT 105.000 3669.000 129.965 3671.000 ;
      LAYER met4 ;
        RECT 129.965 3669.000 131.065 3671.000 ;
        RECT 102.965 3651.000 131.065 3669.000 ;
        RECT 102.965 3649.000 105.000 3651.000 ;
      LAYER met4 ;
        RECT 105.000 3649.000 129.965 3651.000 ;
      LAYER met4 ;
        RECT 129.965 3649.000 131.065 3651.000 ;
        RECT 102.965 3631.000 131.065 3649.000 ;
        RECT 102.965 3629.000 105.000 3631.000 ;
      LAYER met4 ;
        RECT 105.000 3629.000 129.965 3631.000 ;
      LAYER met4 ;
        RECT 129.965 3629.000 131.065 3631.000 ;
        RECT 102.965 3611.000 131.065 3629.000 ;
        RECT 102.965 3609.000 105.000 3611.000 ;
      LAYER met4 ;
        RECT 105.000 3609.000 129.965 3611.000 ;
      LAYER met4 ;
        RECT 129.965 3609.000 131.065 3611.000 ;
        RECT 102.965 3591.000 131.065 3609.000 ;
        RECT 102.965 3589.000 105.000 3591.000 ;
      LAYER met4 ;
        RECT 105.000 3589.000 129.965 3591.000 ;
      LAYER met4 ;
        RECT 129.965 3589.000 131.065 3591.000 ;
        RECT 102.965 3571.000 131.065 3589.000 ;
        RECT 102.965 3570.000 105.000 3571.000 ;
      LAYER met4 ;
        RECT 0.000 3568.730 24.215 3570.000 ;
      LAYER met4 ;
        RECT 24.615 3568.330 104.600 3568.970 ;
      LAYER met4 ;
        RECT 105.000 3568.730 129.965 3571.000 ;
      LAYER met4 ;
        RECT 129.965 3570.000 131.065 3571.000 ;
        RECT 130.365 3568.330 131.065 3568.970 ;
      LAYER met4 ;
        RECT 131.465 3568.730 135.915 3707.270 ;
      LAYER met4 ;
        RECT 136.315 3706.965 136.915 3707.670 ;
        RECT 136.315 3570.000 136.915 3705.000 ;
        RECT 136.315 3568.330 136.915 3568.970 ;
      LAYER met4 ;
        RECT 137.315 3568.730 141.765 3707.270 ;
      LAYER met4 ;
        RECT 142.165 3706.965 142.865 3707.670 ;
        RECT 142.165 3570.000 142.865 3706.000 ;
        RECT 142.165 3568.330 142.865 3568.970 ;
        RECT 0.000 3536.690 142.865 3568.330 ;
      LAYER met4 ;
        RECT 143.265 3537.090 143.595 3708.610 ;
      LAYER met4 ;
        RECT 0.000 3528.360 143.495 3536.690 ;
      LAYER met4 ;
        RECT 143.895 3528.760 146.875 3742.440 ;
      LAYER met4 ;
        RECT 147.275 3707.670 148.255 3742.840 ;
      LAYER met4 ;
        RECT 147.175 3706.000 148.355 3707.270 ;
      LAYER met4 ;
        RECT 147.275 3570.000 148.255 3706.000 ;
      LAYER met4 ;
        RECT 147.175 3568.730 148.355 3570.000 ;
      LAYER met4 ;
        RECT 147.275 3544.065 148.255 3568.330 ;
      LAYER met4 ;
        RECT 148.655 3544.465 151.635 3758.145 ;
        RECT 151.935 3753.090 152.265 3924.610 ;
      LAYER met4 ;
        RECT 152.665 3923.670 199.465 3925.010 ;
        RECT 152.665 3922.965 153.365 3923.670 ;
        RECT 152.665 3784.330 153.365 3784.970 ;
      LAYER met4 ;
        RECT 153.765 3784.730 158.415 3923.270 ;
      LAYER met4 ;
        RECT 158.815 3922.965 159.415 3923.670 ;
        RECT 158.815 3784.330 159.415 3784.970 ;
      LAYER met4 ;
        RECT 159.815 3784.730 163.265 3923.270 ;
      LAYER met4 ;
        RECT 163.665 3922.965 164.265 3923.670 ;
        RECT 163.665 3784.330 164.265 3784.970 ;
      LAYER met4 ;
        RECT 164.665 3784.730 168.115 3923.270 ;
      LAYER met4 ;
        RECT 168.515 3922.965 169.115 3923.670 ;
        RECT 168.515 3784.330 169.115 3784.970 ;
      LAYER met4 ;
        RECT 169.515 3784.730 174.165 3923.270 ;
      LAYER met4 ;
        RECT 174.565 3922.965 175.165 3923.670 ;
        RECT 180.615 3923.365 186.065 3923.670 ;
        RECT 174.565 3784.330 175.165 3784.970 ;
      LAYER met4 ;
        RECT 175.565 3784.730 180.215 3923.270 ;
      LAYER met4 ;
        RECT 180.615 3922.965 181.215 3923.365 ;
        RECT 185.465 3922.965 186.065 3923.365 ;
      LAYER met4 ;
        RECT 181.615 3784.970 185.065 3922.965 ;
      LAYER met4 ;
        RECT 180.615 3784.570 181.215 3784.970 ;
        RECT 185.465 3784.570 186.065 3784.970 ;
      LAYER met4 ;
        RECT 186.465 3784.730 191.115 3923.270 ;
      LAYER met4 ;
        RECT 191.515 3922.965 192.115 3923.670 ;
        RECT 180.615 3784.330 186.065 3784.570 ;
        RECT 191.515 3784.330 192.115 3784.970 ;
      LAYER met4 ;
        RECT 192.515 3784.730 197.965 3923.270 ;
      LAYER met4 ;
        RECT 198.365 3922.965 199.465 3923.670 ;
        RECT 3388.535 3944.330 3389.635 3945.035 ;
      LAYER met4 ;
        RECT 3390.035 3944.730 3395.485 4093.270 ;
      LAYER met4 ;
        RECT 3395.885 4092.965 3396.485 4093.670 ;
        RECT 3401.935 4093.365 3407.385 4093.670 ;
        RECT 3395.885 3944.330 3396.485 3945.035 ;
      LAYER met4 ;
        RECT 3396.885 3944.730 3401.535 4093.270 ;
      LAYER met4 ;
        RECT 3401.935 4092.965 3402.535 4093.365 ;
        RECT 3406.785 4092.965 3407.385 4093.365 ;
        RECT 3401.935 3944.635 3402.535 3945.035 ;
        RECT 3406.785 3944.635 3407.385 3945.035 ;
      LAYER met4 ;
        RECT 3407.785 3944.730 3412.435 4093.270 ;
      LAYER met4 ;
        RECT 3412.835 4092.965 3413.435 4093.670 ;
        RECT 3401.935 3944.330 3407.385 3944.635 ;
        RECT 3412.835 3944.330 3413.435 3945.035 ;
      LAYER met4 ;
        RECT 3413.835 3944.730 3418.485 4093.270 ;
      LAYER met4 ;
        RECT 3418.885 4092.965 3419.485 4093.670 ;
        RECT 3418.885 3944.330 3419.485 3945.035 ;
      LAYER met4 ;
        RECT 3419.885 3944.730 3423.335 4093.270 ;
      LAYER met4 ;
        RECT 3423.735 4092.965 3424.335 4093.670 ;
        RECT 3423.735 3944.330 3424.335 3945.035 ;
      LAYER met4 ;
        RECT 3424.735 3944.730 3428.185 4093.270 ;
      LAYER met4 ;
        RECT 3428.585 4092.965 3429.185 4093.670 ;
        RECT 3428.585 3944.330 3429.185 3945.035 ;
      LAYER met4 ;
        RECT 3429.585 3944.730 3434.235 4093.270 ;
      LAYER met4 ;
        RECT 3434.635 4092.965 3435.335 4093.670 ;
        RECT 3434.635 3944.330 3435.335 3945.035 ;
        RECT 3388.535 3942.990 3435.335 3944.330 ;
      LAYER met4 ;
        RECT 3435.735 3943.390 3436.065 4344.910 ;
        RECT 3436.365 4339.855 3439.345 4783.535 ;
      LAYER met4 ;
        RECT 3439.745 4759.670 3440.725 4783.935 ;
      LAYER met4 ;
        RECT 3439.645 4758.000 3440.825 4759.270 ;
      LAYER met4 ;
        RECT 3439.745 4613.000 3440.725 4758.000 ;
      LAYER met4 ;
        RECT 3439.645 4611.730 3440.825 4613.000 ;
      LAYER met4 ;
        RECT 3439.745 4539.670 3440.725 4611.330 ;
      LAYER met4 ;
        RECT 3439.645 4538.000 3440.825 4539.270 ;
      LAYER met4 ;
        RECT 3439.745 4392.000 3440.725 4538.000 ;
      LAYER met4 ;
        RECT 3439.645 4390.730 3440.825 4392.000 ;
      LAYER met4 ;
        RECT 3439.745 4355.160 3440.725 4390.330 ;
      LAYER met4 ;
        RECT 3441.125 4355.560 3444.105 4799.240 ;
      LAYER met4 ;
        RECT 3444.505 4791.310 3588.000 4799.640 ;
      LAYER met4 ;
        RECT 3444.405 4389.390 3444.735 4790.910 ;
      LAYER met4 ;
        RECT 3445.135 4759.670 3588.000 4791.310 ;
        RECT 3445.135 4759.030 3445.835 4759.670 ;
        RECT 3445.135 4613.000 3445.835 4758.000 ;
        RECT 3445.135 4611.330 3445.835 4612.035 ;
      LAYER met4 ;
        RECT 3446.235 4611.730 3450.685 4759.270 ;
      LAYER met4 ;
        RECT 3451.085 4759.030 3451.685 4759.670 ;
        RECT 3451.085 4613.000 3451.685 4758.000 ;
        RECT 3451.085 4611.330 3451.685 4612.035 ;
      LAYER met4 ;
        RECT 3452.085 4611.730 3456.535 4759.270 ;
      LAYER met4 ;
        RECT 3456.935 4759.030 3457.635 4759.670 ;
        RECT 3456.935 4757.000 3458.035 4758.000 ;
      LAYER met4 ;
        RECT 3458.035 4757.000 3483.000 4759.270 ;
      LAYER met4 ;
        RECT 3483.400 4759.030 3563.385 4759.670 ;
      LAYER met4 ;
        RECT 3563.785 4758.000 3588.000 4759.270 ;
      LAYER met4 ;
        RECT 3483.000 4757.000 3485.035 4758.000 ;
        RECT 3456.935 4754.000 3485.035 4757.000 ;
        RECT 3456.935 4752.000 3458.035 4754.000 ;
      LAYER met4 ;
        RECT 3458.035 4752.000 3483.000 4754.000 ;
      LAYER met4 ;
        RECT 3483.000 4752.000 3485.035 4754.000 ;
        RECT 3456.935 4734.000 3485.035 4752.000 ;
        RECT 3456.935 4732.000 3458.035 4734.000 ;
      LAYER met4 ;
        RECT 3458.035 4732.000 3483.000 4734.000 ;
      LAYER met4 ;
        RECT 3483.000 4732.000 3485.035 4734.000 ;
        RECT 3456.935 4714.000 3485.035 4732.000 ;
        RECT 3456.935 4712.000 3458.035 4714.000 ;
      LAYER met4 ;
        RECT 3458.035 4712.000 3483.000 4714.000 ;
      LAYER met4 ;
        RECT 3483.000 4712.000 3485.035 4714.000 ;
        RECT 3456.935 4694.000 3485.035 4712.000 ;
        RECT 3456.935 4692.000 3458.035 4694.000 ;
      LAYER met4 ;
        RECT 3458.035 4692.000 3483.000 4694.000 ;
      LAYER met4 ;
        RECT 3483.000 4692.000 3485.035 4694.000 ;
        RECT 3456.935 4674.000 3485.035 4692.000 ;
        RECT 3456.935 4672.000 3458.035 4674.000 ;
      LAYER met4 ;
        RECT 3458.035 4672.000 3483.000 4674.000 ;
      LAYER met4 ;
        RECT 3483.000 4672.000 3485.035 4674.000 ;
        RECT 3456.935 4654.000 3485.035 4672.000 ;
        RECT 3456.935 4652.000 3458.035 4654.000 ;
      LAYER met4 ;
        RECT 3458.035 4652.000 3483.000 4654.000 ;
      LAYER met4 ;
        RECT 3483.000 4652.000 3485.035 4654.000 ;
        RECT 3456.935 4634.000 3485.035 4652.000 ;
        RECT 3456.935 4632.000 3458.035 4634.000 ;
      LAYER met4 ;
        RECT 3458.035 4632.000 3483.000 4634.000 ;
      LAYER met4 ;
        RECT 3483.000 4632.000 3485.035 4634.000 ;
        RECT 3456.935 4614.000 3485.035 4632.000 ;
        RECT 3456.935 4613.000 3458.035 4614.000 ;
        RECT 3456.935 4611.330 3457.635 4612.035 ;
      LAYER met4 ;
        RECT 3458.035 4611.730 3483.000 4614.000 ;
      LAYER met4 ;
        RECT 3483.000 4613.000 3485.035 4614.000 ;
        RECT 3562.035 4613.000 3588.000 4758.000 ;
        RECT 3483.400 4611.330 3563.385 4612.035 ;
      LAYER met4 ;
        RECT 3563.785 4611.730 3588.000 4613.000 ;
      LAYER met4 ;
        RECT 3445.135 4539.670 3588.000 4611.330 ;
        RECT 3445.135 4392.000 3445.835 4539.670 ;
        RECT 3445.135 4390.330 3445.835 4391.035 ;
      LAYER met4 ;
        RECT 3446.235 4390.730 3450.685 4539.270 ;
      LAYER met4 ;
        RECT 3451.085 4538.000 3451.685 4539.670 ;
        RECT 3451.085 4392.000 3451.685 4537.000 ;
        RECT 3451.085 4390.330 3451.685 4391.035 ;
      LAYER met4 ;
        RECT 3452.085 4390.730 3456.535 4539.270 ;
      LAYER met4 ;
        RECT 3456.935 4538.000 3457.635 4539.670 ;
        RECT 3456.935 4536.000 3458.035 4538.000 ;
      LAYER met4 ;
        RECT 3458.035 4536.000 3483.000 4539.270 ;
      LAYER met4 ;
        RECT 3483.400 4538.000 3563.385 4539.670 ;
      LAYER met4 ;
        RECT 3563.785 4538.000 3588.000 4539.270 ;
      LAYER met4 ;
        RECT 3483.000 4536.000 3485.035 4538.000 ;
        RECT 3456.935 4533.000 3485.035 4536.000 ;
        RECT 3456.935 4531.000 3458.035 4533.000 ;
      LAYER met4 ;
        RECT 3458.035 4531.000 3483.000 4533.000 ;
      LAYER met4 ;
        RECT 3483.000 4531.000 3485.035 4533.000 ;
        RECT 3456.935 4513.000 3485.035 4531.000 ;
        RECT 3456.935 4511.000 3458.035 4513.000 ;
      LAYER met4 ;
        RECT 3458.035 4511.000 3483.000 4513.000 ;
      LAYER met4 ;
        RECT 3483.000 4511.000 3485.035 4513.000 ;
        RECT 3456.935 4493.000 3485.035 4511.000 ;
        RECT 3456.935 4491.000 3458.035 4493.000 ;
      LAYER met4 ;
        RECT 3458.035 4491.000 3483.000 4493.000 ;
      LAYER met4 ;
        RECT 3483.000 4491.000 3485.035 4493.000 ;
        RECT 3456.935 4473.000 3485.035 4491.000 ;
        RECT 3456.935 4471.000 3458.035 4473.000 ;
      LAYER met4 ;
        RECT 3458.035 4471.000 3483.000 4473.000 ;
      LAYER met4 ;
        RECT 3483.000 4471.000 3485.035 4473.000 ;
        RECT 3456.935 4453.000 3485.035 4471.000 ;
        RECT 3456.935 4451.000 3458.035 4453.000 ;
      LAYER met4 ;
        RECT 3458.035 4451.000 3483.000 4453.000 ;
      LAYER met4 ;
        RECT 3483.000 4451.000 3485.035 4453.000 ;
        RECT 3456.935 4433.000 3485.035 4451.000 ;
        RECT 3456.935 4431.000 3458.035 4433.000 ;
      LAYER met4 ;
        RECT 3458.035 4431.000 3483.000 4433.000 ;
      LAYER met4 ;
        RECT 3483.000 4431.000 3485.035 4433.000 ;
        RECT 3456.935 4413.000 3485.035 4431.000 ;
        RECT 3456.935 4411.000 3458.035 4413.000 ;
      LAYER met4 ;
        RECT 3458.035 4411.000 3483.000 4413.000 ;
      LAYER met4 ;
        RECT 3483.000 4411.000 3485.035 4413.000 ;
        RECT 3456.935 4393.000 3485.035 4411.000 ;
        RECT 3456.935 4392.000 3458.035 4393.000 ;
        RECT 3456.935 4390.330 3457.635 4391.035 ;
      LAYER met4 ;
        RECT 3458.035 4390.730 3483.000 4393.000 ;
      LAYER met4 ;
        RECT 3483.000 4392.000 3485.035 4393.000 ;
        RECT 3562.035 4392.000 3588.000 4538.000 ;
        RECT 3483.400 4390.330 3563.385 4391.035 ;
      LAYER met4 ;
        RECT 3563.785 4390.730 3588.000 4392.000 ;
      LAYER met4 ;
        RECT 3445.135 4388.990 3588.000 4390.330 ;
        RECT 3444.505 4355.160 3588.000 4388.990 ;
        RECT 3439.745 4353.640 3588.000 4355.160 ;
        RECT 3439.745 4339.455 3440.725 4353.640 ;
        RECT 3436.465 4337.935 3440.725 4339.455 ;
        RECT 3388.535 3899.310 3435.965 3942.990 ;
        RECT 3388.535 3867.670 3435.335 3899.310 ;
        RECT 3388.535 3867.030 3389.635 3867.670 ;
        RECT 198.365 3784.330 199.465 3784.970 ;
        RECT 152.665 3752.690 199.465 3784.330 ;
        RECT 152.035 3709.010 199.465 3752.690 ;
        RECT 147.275 3542.545 151.535 3544.065 ;
        RECT 147.275 3528.360 148.255 3542.545 ;
        RECT 0.000 3526.840 148.255 3528.360 ;
        RECT 0.000 3493.010 143.495 3526.840 ;
        RECT 0.000 3491.670 142.865 3493.010 ;
      LAYER met4 ;
        RECT 0.000 3490.000 24.215 3491.270 ;
      LAYER met4 ;
        RECT 24.615 3490.965 104.600 3491.670 ;
        RECT 0.000 3354.000 25.965 3490.000 ;
        RECT 102.965 3488.000 105.000 3490.000 ;
      LAYER met4 ;
        RECT 105.000 3488.000 129.965 3491.270 ;
      LAYER met4 ;
        RECT 130.365 3490.965 131.065 3491.670 ;
        RECT 129.965 3488.000 131.065 3490.000 ;
        RECT 102.965 3485.000 131.065 3488.000 ;
        RECT 102.965 3483.000 105.000 3485.000 ;
      LAYER met4 ;
        RECT 105.000 3483.000 129.965 3485.000 ;
      LAYER met4 ;
        RECT 129.965 3483.000 131.065 3485.000 ;
        RECT 102.965 3475.000 131.065 3483.000 ;
        RECT 102.965 3473.000 105.000 3475.000 ;
      LAYER met4 ;
        RECT 105.000 3473.000 129.965 3475.000 ;
      LAYER met4 ;
        RECT 129.965 3473.000 131.065 3475.000 ;
        RECT 102.965 3455.000 131.065 3473.000 ;
        RECT 102.965 3453.000 105.000 3455.000 ;
      LAYER met4 ;
        RECT 105.000 3453.000 129.965 3455.000 ;
      LAYER met4 ;
        RECT 129.965 3453.000 131.065 3455.000 ;
        RECT 102.965 3435.000 131.065 3453.000 ;
        RECT 102.965 3433.000 105.000 3435.000 ;
      LAYER met4 ;
        RECT 105.000 3433.000 129.965 3435.000 ;
      LAYER met4 ;
        RECT 129.965 3433.000 131.065 3435.000 ;
        RECT 102.965 3415.000 131.065 3433.000 ;
        RECT 102.965 3413.000 105.000 3415.000 ;
      LAYER met4 ;
        RECT 105.000 3413.000 129.965 3415.000 ;
      LAYER met4 ;
        RECT 129.965 3413.000 131.065 3415.000 ;
        RECT 102.965 3395.000 131.065 3413.000 ;
        RECT 102.965 3393.000 105.000 3395.000 ;
      LAYER met4 ;
        RECT 105.000 3393.000 129.965 3395.000 ;
      LAYER met4 ;
        RECT 129.965 3393.000 131.065 3395.000 ;
        RECT 102.965 3375.000 131.065 3393.000 ;
        RECT 102.965 3373.000 105.000 3375.000 ;
      LAYER met4 ;
        RECT 105.000 3373.000 129.965 3375.000 ;
      LAYER met4 ;
        RECT 129.965 3373.000 131.065 3375.000 ;
        RECT 102.965 3355.000 131.065 3373.000 ;
        RECT 102.965 3354.000 105.000 3355.000 ;
      LAYER met4 ;
        RECT 0.000 3352.730 24.215 3354.000 ;
      LAYER met4 ;
        RECT 24.615 3352.330 104.600 3352.970 ;
      LAYER met4 ;
        RECT 105.000 3352.730 129.965 3355.000 ;
      LAYER met4 ;
        RECT 129.965 3354.000 131.065 3355.000 ;
        RECT 130.365 3352.330 131.065 3352.970 ;
      LAYER met4 ;
        RECT 131.465 3352.730 135.915 3491.270 ;
      LAYER met4 ;
        RECT 136.315 3490.965 136.915 3491.670 ;
        RECT 136.315 3354.000 136.915 3489.000 ;
        RECT 136.315 3352.330 136.915 3352.970 ;
      LAYER met4 ;
        RECT 137.315 3352.730 141.765 3491.270 ;
      LAYER met4 ;
        RECT 142.165 3490.965 142.865 3491.670 ;
        RECT 142.165 3354.000 142.865 3490.000 ;
        RECT 142.165 3352.330 142.865 3352.970 ;
        RECT 0.000 3320.690 142.865 3352.330 ;
      LAYER met4 ;
        RECT 143.265 3321.090 143.595 3492.610 ;
      LAYER met4 ;
        RECT 0.000 3312.360 143.495 3320.690 ;
      LAYER met4 ;
        RECT 143.895 3312.760 146.875 3526.440 ;
      LAYER met4 ;
        RECT 147.275 3491.670 148.255 3526.840 ;
      LAYER met4 ;
        RECT 147.175 3490.000 148.355 3491.270 ;
      LAYER met4 ;
        RECT 147.275 3354.000 148.255 3490.000 ;
      LAYER met4 ;
        RECT 147.175 3352.730 148.355 3354.000 ;
      LAYER met4 ;
        RECT 147.275 3328.065 148.255 3352.330 ;
      LAYER met4 ;
        RECT 148.655 3328.465 151.635 3542.145 ;
        RECT 151.935 3537.090 152.265 3708.610 ;
      LAYER met4 ;
        RECT 152.665 3707.670 199.465 3709.010 ;
        RECT 152.665 3706.965 153.365 3707.670 ;
        RECT 152.665 3568.330 153.365 3568.970 ;
      LAYER met4 ;
        RECT 153.765 3568.730 158.415 3707.270 ;
      LAYER met4 ;
        RECT 158.815 3706.965 159.415 3707.670 ;
        RECT 158.815 3568.330 159.415 3568.970 ;
      LAYER met4 ;
        RECT 159.815 3568.730 163.265 3707.270 ;
      LAYER met4 ;
        RECT 163.665 3706.965 164.265 3707.670 ;
        RECT 163.665 3568.330 164.265 3568.970 ;
      LAYER met4 ;
        RECT 164.665 3568.730 168.115 3707.270 ;
      LAYER met4 ;
        RECT 168.515 3706.965 169.115 3707.670 ;
        RECT 168.515 3568.330 169.115 3568.970 ;
      LAYER met4 ;
        RECT 169.515 3568.730 174.165 3707.270 ;
      LAYER met4 ;
        RECT 174.565 3706.965 175.165 3707.670 ;
        RECT 180.615 3707.365 186.065 3707.670 ;
        RECT 174.565 3568.330 175.165 3568.970 ;
      LAYER met4 ;
        RECT 175.565 3568.730 180.215 3707.270 ;
      LAYER met4 ;
        RECT 180.615 3706.965 181.215 3707.365 ;
        RECT 185.465 3706.965 186.065 3707.365 ;
      LAYER met4 ;
        RECT 181.615 3568.970 185.065 3706.965 ;
      LAYER met4 ;
        RECT 180.615 3568.570 181.215 3568.970 ;
        RECT 185.465 3568.570 186.065 3568.970 ;
      LAYER met4 ;
        RECT 186.465 3568.730 191.115 3707.270 ;
      LAYER met4 ;
        RECT 191.515 3706.965 192.115 3707.670 ;
        RECT 180.615 3568.330 186.065 3568.570 ;
        RECT 191.515 3568.330 192.115 3568.970 ;
      LAYER met4 ;
        RECT 192.515 3568.730 197.965 3707.270 ;
      LAYER met4 ;
        RECT 198.365 3706.965 199.465 3707.670 ;
        RECT 3388.535 3719.330 3389.635 3720.035 ;
      LAYER met4 ;
        RECT 3390.035 3719.730 3395.485 3867.270 ;
      LAYER met4 ;
        RECT 3395.885 3867.030 3396.485 3867.670 ;
        RECT 3401.935 3867.430 3407.385 3867.670 ;
        RECT 3395.885 3719.330 3396.485 3720.035 ;
      LAYER met4 ;
        RECT 3396.885 3719.730 3401.535 3867.270 ;
      LAYER met4 ;
        RECT 3401.935 3867.030 3402.535 3867.430 ;
        RECT 3406.785 3867.030 3407.385 3867.430 ;
      LAYER met4 ;
        RECT 3402.935 3720.035 3406.385 3867.030 ;
      LAYER met4 ;
        RECT 3401.935 3719.635 3402.535 3720.035 ;
        RECT 3406.785 3719.635 3407.385 3720.035 ;
      LAYER met4 ;
        RECT 3407.785 3719.730 3412.435 3867.270 ;
      LAYER met4 ;
        RECT 3412.835 3867.030 3413.435 3867.670 ;
        RECT 3401.935 3719.330 3407.385 3719.635 ;
        RECT 3412.835 3719.330 3413.435 3720.035 ;
      LAYER met4 ;
        RECT 3413.835 3719.730 3418.485 3867.270 ;
      LAYER met4 ;
        RECT 3418.885 3867.030 3419.485 3867.670 ;
        RECT 3418.885 3719.330 3419.485 3720.035 ;
      LAYER met4 ;
        RECT 3419.885 3719.730 3423.335 3867.270 ;
      LAYER met4 ;
        RECT 3423.735 3867.030 3424.335 3867.670 ;
        RECT 3423.735 3719.330 3424.335 3720.035 ;
      LAYER met4 ;
        RECT 3424.735 3719.730 3428.185 3867.270 ;
      LAYER met4 ;
        RECT 3428.585 3867.030 3429.185 3867.670 ;
        RECT 3428.585 3719.330 3429.185 3720.035 ;
      LAYER met4 ;
        RECT 3429.585 3719.730 3434.235 3867.270 ;
      LAYER met4 ;
        RECT 3434.635 3867.030 3435.335 3867.670 ;
        RECT 3434.635 3719.330 3435.335 3720.035 ;
        RECT 3388.535 3717.990 3435.335 3719.330 ;
      LAYER met4 ;
        RECT 3435.735 3718.390 3436.065 3898.910 ;
        RECT 3436.365 3893.855 3439.345 4337.535 ;
      LAYER met4 ;
        RECT 3439.745 4313.670 3440.725 4337.935 ;
      LAYER met4 ;
        RECT 3439.645 4312.000 3440.825 4313.270 ;
      LAYER met4 ;
        RECT 3439.745 4167.000 3440.725 4312.000 ;
      LAYER met4 ;
        RECT 3439.645 4165.730 3440.825 4167.000 ;
      LAYER met4 ;
        RECT 3439.745 4093.670 3440.725 4165.330 ;
      LAYER met4 ;
        RECT 3439.645 4092.000 3440.825 4093.270 ;
      LAYER met4 ;
        RECT 3439.745 3946.000 3440.725 4092.000 ;
      LAYER met4 ;
        RECT 3439.645 3944.730 3440.825 3946.000 ;
      LAYER met4 ;
        RECT 3439.745 3909.160 3440.725 3944.330 ;
      LAYER met4 ;
        RECT 3441.125 3909.560 3444.105 4353.240 ;
      LAYER met4 ;
        RECT 3444.505 4345.310 3588.000 4353.640 ;
      LAYER met4 ;
        RECT 3444.405 3943.390 3444.735 4344.910 ;
      LAYER met4 ;
        RECT 3445.135 4313.670 3588.000 4345.310 ;
        RECT 3445.135 4313.030 3445.835 4313.670 ;
        RECT 3445.135 4167.000 3445.835 4312.000 ;
        RECT 3445.135 4165.330 3445.835 4166.035 ;
      LAYER met4 ;
        RECT 3446.235 4165.730 3450.685 4313.270 ;
      LAYER met4 ;
        RECT 3451.085 4313.030 3451.685 4313.670 ;
        RECT 3451.085 4167.000 3451.685 4312.000 ;
        RECT 3451.085 4165.330 3451.685 4166.035 ;
      LAYER met4 ;
        RECT 3452.085 4165.730 3456.535 4313.270 ;
      LAYER met4 ;
        RECT 3456.935 4313.030 3457.635 4313.670 ;
        RECT 3456.935 4311.000 3458.035 4312.000 ;
      LAYER met4 ;
        RECT 3458.035 4311.000 3483.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4313.030 3563.385 4313.670 ;
      LAYER met4 ;
        RECT 3563.785 4312.000 3588.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.000 4311.000 3485.035 4312.000 ;
        RECT 3456.935 4308.000 3485.035 4311.000 ;
        RECT 3456.935 4306.000 3458.035 4308.000 ;
      LAYER met4 ;
        RECT 3458.035 4306.000 3483.000 4308.000 ;
      LAYER met4 ;
        RECT 3483.000 4306.000 3485.035 4308.000 ;
        RECT 3456.935 4288.000 3485.035 4306.000 ;
        RECT 3456.935 4286.000 3458.035 4288.000 ;
      LAYER met4 ;
        RECT 3458.035 4286.000 3483.000 4288.000 ;
      LAYER met4 ;
        RECT 3483.000 4286.000 3485.035 4288.000 ;
        RECT 3456.935 4268.000 3485.035 4286.000 ;
        RECT 3456.935 4266.000 3458.035 4268.000 ;
      LAYER met4 ;
        RECT 3458.035 4266.000 3483.000 4268.000 ;
      LAYER met4 ;
        RECT 3483.000 4266.000 3485.035 4268.000 ;
        RECT 3456.935 4248.000 3485.035 4266.000 ;
        RECT 3456.935 4246.000 3458.035 4248.000 ;
      LAYER met4 ;
        RECT 3458.035 4246.000 3483.000 4248.000 ;
      LAYER met4 ;
        RECT 3483.000 4246.000 3485.035 4248.000 ;
        RECT 3456.935 4228.000 3485.035 4246.000 ;
        RECT 3456.935 4226.000 3458.035 4228.000 ;
      LAYER met4 ;
        RECT 3458.035 4226.000 3483.000 4228.000 ;
      LAYER met4 ;
        RECT 3483.000 4226.000 3485.035 4228.000 ;
        RECT 3456.935 4208.000 3485.035 4226.000 ;
        RECT 3456.935 4206.000 3458.035 4208.000 ;
      LAYER met4 ;
        RECT 3458.035 4206.000 3483.000 4208.000 ;
      LAYER met4 ;
        RECT 3483.000 4206.000 3485.035 4208.000 ;
        RECT 3456.935 4188.000 3485.035 4206.000 ;
        RECT 3456.935 4186.000 3458.035 4188.000 ;
      LAYER met4 ;
        RECT 3458.035 4186.000 3483.000 4188.000 ;
      LAYER met4 ;
        RECT 3483.000 4186.000 3485.035 4188.000 ;
        RECT 3456.935 4168.000 3485.035 4186.000 ;
        RECT 3456.935 4167.000 3458.035 4168.000 ;
        RECT 3456.935 4165.330 3457.635 4166.035 ;
      LAYER met4 ;
        RECT 3458.035 4165.730 3483.000 4168.000 ;
      LAYER met4 ;
        RECT 3483.000 4167.000 3485.035 4168.000 ;
        RECT 3562.035 4167.000 3588.000 4312.000 ;
        RECT 3483.400 4165.330 3563.385 4166.035 ;
      LAYER met4 ;
        RECT 3563.785 4165.730 3588.000 4167.000 ;
      LAYER met4 ;
        RECT 3445.135 4093.670 3588.000 4165.330 ;
        RECT 3445.135 4092.965 3445.835 4093.670 ;
        RECT 3445.135 3946.000 3445.835 4092.000 ;
        RECT 3445.135 3944.330 3445.835 3945.035 ;
      LAYER met4 ;
        RECT 3446.235 3944.730 3450.685 4093.270 ;
      LAYER met4 ;
        RECT 3451.085 4092.965 3451.685 4093.670 ;
        RECT 3451.085 3946.000 3451.685 4091.000 ;
        RECT 3451.085 3944.330 3451.685 3945.035 ;
      LAYER met4 ;
        RECT 3452.085 3944.730 3456.535 4093.270 ;
      LAYER met4 ;
        RECT 3456.935 4092.965 3457.635 4093.670 ;
        RECT 3456.935 4090.000 3458.035 4092.000 ;
      LAYER met4 ;
        RECT 3458.035 4090.000 3483.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 4092.965 3563.385 4093.670 ;
      LAYER met4 ;
        RECT 3563.785 4092.000 3588.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.000 4090.000 3485.035 4092.000 ;
        RECT 3456.935 4087.000 3485.035 4090.000 ;
        RECT 3456.935 4085.000 3458.035 4087.000 ;
      LAYER met4 ;
        RECT 3458.035 4085.000 3483.000 4087.000 ;
      LAYER met4 ;
        RECT 3483.000 4085.000 3485.035 4087.000 ;
        RECT 3456.935 4067.000 3485.035 4085.000 ;
        RECT 3456.935 4065.000 3458.035 4067.000 ;
      LAYER met4 ;
        RECT 3458.035 4065.000 3483.000 4067.000 ;
      LAYER met4 ;
        RECT 3483.000 4065.000 3485.035 4067.000 ;
        RECT 3456.935 4047.000 3485.035 4065.000 ;
        RECT 3456.935 4045.000 3458.035 4047.000 ;
      LAYER met4 ;
        RECT 3458.035 4045.000 3483.000 4047.000 ;
      LAYER met4 ;
        RECT 3483.000 4045.000 3485.035 4047.000 ;
        RECT 3456.935 4027.000 3485.035 4045.000 ;
        RECT 3456.935 4025.000 3458.035 4027.000 ;
      LAYER met4 ;
        RECT 3458.035 4025.000 3483.000 4027.000 ;
      LAYER met4 ;
        RECT 3483.000 4025.000 3485.035 4027.000 ;
        RECT 3456.935 4007.000 3485.035 4025.000 ;
        RECT 3456.935 4005.000 3458.035 4007.000 ;
      LAYER met4 ;
        RECT 3458.035 4005.000 3483.000 4007.000 ;
      LAYER met4 ;
        RECT 3483.000 4005.000 3485.035 4007.000 ;
        RECT 3456.935 3987.000 3485.035 4005.000 ;
        RECT 3456.935 3985.000 3458.035 3987.000 ;
      LAYER met4 ;
        RECT 3458.035 3985.000 3483.000 3987.000 ;
      LAYER met4 ;
        RECT 3483.000 3985.000 3485.035 3987.000 ;
        RECT 3456.935 3967.000 3485.035 3985.000 ;
        RECT 3456.935 3965.000 3458.035 3967.000 ;
      LAYER met4 ;
        RECT 3458.035 3965.000 3483.000 3967.000 ;
      LAYER met4 ;
        RECT 3483.000 3965.000 3485.035 3967.000 ;
        RECT 3456.935 3947.000 3485.035 3965.000 ;
        RECT 3456.935 3946.000 3458.035 3947.000 ;
        RECT 3456.935 3944.330 3457.635 3945.035 ;
      LAYER met4 ;
        RECT 3458.035 3944.730 3483.000 3947.000 ;
      LAYER met4 ;
        RECT 3483.000 3946.000 3485.035 3947.000 ;
        RECT 3562.035 3946.000 3588.000 4092.000 ;
        RECT 3483.400 3944.330 3563.385 3945.035 ;
      LAYER met4 ;
        RECT 3563.785 3944.730 3588.000 3946.000 ;
      LAYER met4 ;
        RECT 3445.135 3942.990 3588.000 3944.330 ;
        RECT 3444.505 3909.160 3588.000 3942.990 ;
        RECT 3439.745 3907.640 3588.000 3909.160 ;
        RECT 3439.745 3893.455 3440.725 3907.640 ;
        RECT 3436.465 3891.935 3440.725 3893.455 ;
        RECT 3388.535 3674.310 3435.965 3717.990 ;
        RECT 3388.535 3642.670 3435.335 3674.310 ;
        RECT 3388.535 3642.030 3389.635 3642.670 ;
        RECT 198.365 3568.330 199.465 3568.970 ;
        RECT 152.665 3536.690 199.465 3568.330 ;
        RECT 152.035 3493.010 199.465 3536.690 ;
        RECT 147.275 3326.545 151.535 3328.065 ;
        RECT 147.275 3312.360 148.255 3326.545 ;
        RECT 0.000 3310.840 148.255 3312.360 ;
        RECT 0.000 3277.010 143.495 3310.840 ;
        RECT 0.000 3275.670 142.865 3277.010 ;
      LAYER met4 ;
        RECT 0.000 3274.000 24.215 3275.270 ;
      LAYER met4 ;
        RECT 24.615 3274.965 104.600 3275.670 ;
        RECT 0.000 3138.000 25.965 3274.000 ;
        RECT 102.965 3272.000 105.000 3274.000 ;
      LAYER met4 ;
        RECT 105.000 3272.000 129.965 3275.270 ;
      LAYER met4 ;
        RECT 130.365 3274.965 131.065 3275.670 ;
        RECT 129.965 3272.000 131.065 3274.000 ;
        RECT 102.965 3269.000 131.065 3272.000 ;
        RECT 102.965 3267.000 105.000 3269.000 ;
      LAYER met4 ;
        RECT 105.000 3267.000 129.965 3269.000 ;
      LAYER met4 ;
        RECT 129.965 3267.000 131.065 3269.000 ;
        RECT 102.965 3259.000 131.065 3267.000 ;
        RECT 102.965 3257.000 105.000 3259.000 ;
      LAYER met4 ;
        RECT 105.000 3257.000 129.965 3259.000 ;
      LAYER met4 ;
        RECT 129.965 3257.000 131.065 3259.000 ;
        RECT 102.965 3239.000 131.065 3257.000 ;
        RECT 102.965 3237.000 105.000 3239.000 ;
      LAYER met4 ;
        RECT 105.000 3237.000 129.965 3239.000 ;
      LAYER met4 ;
        RECT 129.965 3237.000 131.065 3239.000 ;
        RECT 102.965 3219.000 131.065 3237.000 ;
        RECT 102.965 3217.000 105.000 3219.000 ;
      LAYER met4 ;
        RECT 105.000 3217.000 129.965 3219.000 ;
      LAYER met4 ;
        RECT 129.965 3217.000 131.065 3219.000 ;
        RECT 102.965 3199.000 131.065 3217.000 ;
        RECT 102.965 3197.000 105.000 3199.000 ;
      LAYER met4 ;
        RECT 105.000 3197.000 129.965 3199.000 ;
      LAYER met4 ;
        RECT 129.965 3197.000 131.065 3199.000 ;
        RECT 102.965 3179.000 131.065 3197.000 ;
        RECT 102.965 3177.000 105.000 3179.000 ;
      LAYER met4 ;
        RECT 105.000 3177.000 129.965 3179.000 ;
      LAYER met4 ;
        RECT 129.965 3177.000 131.065 3179.000 ;
        RECT 102.965 3159.000 131.065 3177.000 ;
        RECT 102.965 3157.000 105.000 3159.000 ;
      LAYER met4 ;
        RECT 105.000 3157.000 129.965 3159.000 ;
      LAYER met4 ;
        RECT 129.965 3157.000 131.065 3159.000 ;
        RECT 102.965 3139.000 131.065 3157.000 ;
        RECT 102.965 3138.000 105.000 3139.000 ;
      LAYER met4 ;
        RECT 0.000 3136.730 24.215 3138.000 ;
      LAYER met4 ;
        RECT 24.615 3136.330 104.600 3136.970 ;
      LAYER met4 ;
        RECT 105.000 3136.730 129.965 3139.000 ;
      LAYER met4 ;
        RECT 129.965 3138.000 131.065 3139.000 ;
        RECT 130.365 3136.330 131.065 3136.970 ;
      LAYER met4 ;
        RECT 131.465 3136.730 135.915 3275.270 ;
      LAYER met4 ;
        RECT 136.315 3274.965 136.915 3275.670 ;
        RECT 136.315 3138.000 136.915 3273.000 ;
        RECT 136.315 3136.330 136.915 3136.970 ;
      LAYER met4 ;
        RECT 137.315 3136.730 141.765 3275.270 ;
      LAYER met4 ;
        RECT 142.165 3274.965 142.865 3275.670 ;
        RECT 142.165 3138.000 142.865 3274.000 ;
        RECT 142.165 3136.330 142.865 3136.970 ;
        RECT 0.000 3104.690 142.865 3136.330 ;
      LAYER met4 ;
        RECT 143.265 3105.090 143.595 3276.610 ;
      LAYER met4 ;
        RECT 0.000 3096.360 143.495 3104.690 ;
      LAYER met4 ;
        RECT 143.895 3096.760 146.875 3310.440 ;
      LAYER met4 ;
        RECT 147.275 3275.670 148.255 3310.840 ;
      LAYER met4 ;
        RECT 147.175 3274.000 148.355 3275.270 ;
      LAYER met4 ;
        RECT 147.275 3138.000 148.255 3274.000 ;
      LAYER met4 ;
        RECT 147.175 3136.730 148.355 3138.000 ;
      LAYER met4 ;
        RECT 147.275 3112.065 148.255 3136.330 ;
      LAYER met4 ;
        RECT 148.655 3112.465 151.635 3326.145 ;
        RECT 151.935 3321.090 152.265 3492.610 ;
      LAYER met4 ;
        RECT 152.665 3491.670 199.465 3493.010 ;
        RECT 152.665 3490.965 153.365 3491.670 ;
        RECT 152.665 3352.330 153.365 3352.970 ;
      LAYER met4 ;
        RECT 153.765 3352.730 158.415 3491.270 ;
      LAYER met4 ;
        RECT 158.815 3490.965 159.415 3491.670 ;
        RECT 158.815 3352.330 159.415 3352.970 ;
      LAYER met4 ;
        RECT 159.815 3352.730 163.265 3491.270 ;
      LAYER met4 ;
        RECT 163.665 3490.965 164.265 3491.670 ;
        RECT 163.665 3352.330 164.265 3352.970 ;
      LAYER met4 ;
        RECT 164.665 3352.730 168.115 3491.270 ;
      LAYER met4 ;
        RECT 168.515 3490.965 169.115 3491.670 ;
        RECT 168.515 3352.330 169.115 3352.970 ;
      LAYER met4 ;
        RECT 169.515 3352.730 174.165 3491.270 ;
      LAYER met4 ;
        RECT 174.565 3490.965 175.165 3491.670 ;
        RECT 180.615 3491.365 186.065 3491.670 ;
        RECT 174.565 3352.330 175.165 3352.970 ;
      LAYER met4 ;
        RECT 175.565 3352.730 180.215 3491.270 ;
      LAYER met4 ;
        RECT 180.615 3490.965 181.215 3491.365 ;
        RECT 185.465 3490.965 186.065 3491.365 ;
      LAYER met4 ;
        RECT 181.615 3352.970 185.065 3490.965 ;
      LAYER met4 ;
        RECT 180.615 3352.570 181.215 3352.970 ;
        RECT 185.465 3352.570 186.065 3352.970 ;
      LAYER met4 ;
        RECT 186.465 3352.730 191.115 3491.270 ;
      LAYER met4 ;
        RECT 191.515 3490.965 192.115 3491.670 ;
        RECT 180.615 3352.330 186.065 3352.570 ;
        RECT 191.515 3352.330 192.115 3352.970 ;
      LAYER met4 ;
        RECT 192.515 3352.730 197.965 3491.270 ;
      LAYER met4 ;
        RECT 198.365 3490.965 199.465 3491.670 ;
        RECT 3388.535 3494.330 3389.635 3495.035 ;
      LAYER met4 ;
        RECT 3390.035 3494.730 3395.485 3642.270 ;
      LAYER met4 ;
        RECT 3395.885 3642.030 3396.485 3642.670 ;
        RECT 3401.935 3642.430 3407.385 3642.670 ;
        RECT 3395.885 3494.330 3396.485 3495.035 ;
      LAYER met4 ;
        RECT 3396.885 3494.730 3401.535 3642.270 ;
      LAYER met4 ;
        RECT 3401.935 3642.030 3402.535 3642.430 ;
        RECT 3406.785 3642.030 3407.385 3642.430 ;
      LAYER met4 ;
        RECT 3402.935 3495.035 3406.385 3642.030 ;
      LAYER met4 ;
        RECT 3401.935 3494.635 3402.535 3495.035 ;
        RECT 3406.785 3494.635 3407.385 3495.035 ;
      LAYER met4 ;
        RECT 3407.785 3494.730 3412.435 3642.270 ;
      LAYER met4 ;
        RECT 3412.835 3642.030 3413.435 3642.670 ;
        RECT 3401.935 3494.330 3407.385 3494.635 ;
        RECT 3412.835 3494.330 3413.435 3495.035 ;
      LAYER met4 ;
        RECT 3413.835 3494.730 3418.485 3642.270 ;
      LAYER met4 ;
        RECT 3418.885 3642.030 3419.485 3642.670 ;
        RECT 3418.885 3494.330 3419.485 3495.035 ;
      LAYER met4 ;
        RECT 3419.885 3494.730 3423.335 3642.270 ;
      LAYER met4 ;
        RECT 3423.735 3642.030 3424.335 3642.670 ;
        RECT 3423.735 3494.330 3424.335 3495.035 ;
      LAYER met4 ;
        RECT 3424.735 3494.730 3428.185 3642.270 ;
      LAYER met4 ;
        RECT 3428.585 3642.030 3429.185 3642.670 ;
        RECT 3428.585 3494.330 3429.185 3495.035 ;
      LAYER met4 ;
        RECT 3429.585 3494.730 3434.235 3642.270 ;
      LAYER met4 ;
        RECT 3434.635 3642.030 3435.335 3642.670 ;
        RECT 3434.635 3494.330 3435.335 3495.035 ;
        RECT 3388.535 3492.990 3435.335 3494.330 ;
      LAYER met4 ;
        RECT 3435.735 3493.390 3436.065 3673.910 ;
        RECT 3436.365 3668.855 3439.345 3891.535 ;
      LAYER met4 ;
        RECT 3439.745 3867.670 3440.725 3891.935 ;
      LAYER met4 ;
        RECT 3439.645 3866.000 3440.825 3867.270 ;
      LAYER met4 ;
        RECT 3439.745 3721.000 3440.725 3866.000 ;
      LAYER met4 ;
        RECT 3439.645 3719.730 3440.825 3721.000 ;
      LAYER met4 ;
        RECT 3439.745 3684.160 3440.725 3719.330 ;
      LAYER met4 ;
        RECT 3441.125 3684.560 3444.105 3907.240 ;
      LAYER met4 ;
        RECT 3444.505 3899.310 3588.000 3907.640 ;
      LAYER met4 ;
        RECT 3444.405 3718.390 3444.735 3898.910 ;
      LAYER met4 ;
        RECT 3445.135 3867.670 3588.000 3899.310 ;
        RECT 3445.135 3867.030 3445.835 3867.670 ;
        RECT 3445.135 3721.000 3445.835 3866.000 ;
        RECT 3445.135 3719.330 3445.835 3720.035 ;
      LAYER met4 ;
        RECT 3446.235 3719.730 3450.685 3867.270 ;
      LAYER met4 ;
        RECT 3451.085 3867.030 3451.685 3867.670 ;
        RECT 3451.085 3721.000 3451.685 3866.000 ;
        RECT 3451.085 3719.330 3451.685 3720.035 ;
      LAYER met4 ;
        RECT 3452.085 3719.730 3456.535 3867.270 ;
      LAYER met4 ;
        RECT 3456.935 3867.030 3457.635 3867.670 ;
        RECT 3456.935 3865.000 3458.035 3866.000 ;
      LAYER met4 ;
        RECT 3458.035 3865.000 3483.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3867.030 3563.385 3867.670 ;
      LAYER met4 ;
        RECT 3563.785 3866.000 3588.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.000 3865.000 3485.035 3866.000 ;
        RECT 3456.935 3862.000 3485.035 3865.000 ;
        RECT 3456.935 3860.000 3458.035 3862.000 ;
      LAYER met4 ;
        RECT 3458.035 3860.000 3483.000 3862.000 ;
      LAYER met4 ;
        RECT 3483.000 3860.000 3485.035 3862.000 ;
        RECT 3456.935 3842.000 3485.035 3860.000 ;
        RECT 3456.935 3840.000 3458.035 3842.000 ;
      LAYER met4 ;
        RECT 3458.035 3840.000 3483.000 3842.000 ;
      LAYER met4 ;
        RECT 3483.000 3840.000 3485.035 3842.000 ;
        RECT 3456.935 3822.000 3485.035 3840.000 ;
        RECT 3456.935 3820.000 3458.035 3822.000 ;
      LAYER met4 ;
        RECT 3458.035 3820.000 3483.000 3822.000 ;
      LAYER met4 ;
        RECT 3483.000 3820.000 3485.035 3822.000 ;
        RECT 3456.935 3802.000 3485.035 3820.000 ;
        RECT 3456.935 3800.000 3458.035 3802.000 ;
      LAYER met4 ;
        RECT 3458.035 3800.000 3483.000 3802.000 ;
      LAYER met4 ;
        RECT 3483.000 3800.000 3485.035 3802.000 ;
        RECT 3456.935 3782.000 3485.035 3800.000 ;
        RECT 3456.935 3780.000 3458.035 3782.000 ;
      LAYER met4 ;
        RECT 3458.035 3780.000 3483.000 3782.000 ;
      LAYER met4 ;
        RECT 3483.000 3780.000 3485.035 3782.000 ;
        RECT 3456.935 3762.000 3485.035 3780.000 ;
        RECT 3456.935 3760.000 3458.035 3762.000 ;
      LAYER met4 ;
        RECT 3458.035 3760.000 3483.000 3762.000 ;
      LAYER met4 ;
        RECT 3483.000 3760.000 3485.035 3762.000 ;
        RECT 3456.935 3742.000 3485.035 3760.000 ;
        RECT 3456.935 3740.000 3458.035 3742.000 ;
      LAYER met4 ;
        RECT 3458.035 3740.000 3483.000 3742.000 ;
      LAYER met4 ;
        RECT 3483.000 3740.000 3485.035 3742.000 ;
        RECT 3456.935 3722.000 3485.035 3740.000 ;
        RECT 3456.935 3721.000 3458.035 3722.000 ;
        RECT 3456.935 3719.330 3457.635 3720.035 ;
      LAYER met4 ;
        RECT 3458.035 3719.730 3483.000 3722.000 ;
      LAYER met4 ;
        RECT 3483.000 3721.000 3485.035 3722.000 ;
        RECT 3562.035 3721.000 3588.000 3866.000 ;
        RECT 3483.400 3719.330 3563.385 3720.035 ;
      LAYER met4 ;
        RECT 3563.785 3719.730 3588.000 3721.000 ;
      LAYER met4 ;
        RECT 3445.135 3717.990 3588.000 3719.330 ;
        RECT 3444.505 3684.160 3588.000 3717.990 ;
        RECT 3439.745 3682.640 3588.000 3684.160 ;
        RECT 3439.745 3668.455 3440.725 3682.640 ;
        RECT 3436.465 3666.935 3440.725 3668.455 ;
        RECT 3388.535 3449.310 3435.965 3492.990 ;
        RECT 3388.535 3417.670 3435.335 3449.310 ;
        RECT 3388.535 3417.030 3389.635 3417.670 ;
        RECT 198.365 3352.330 199.465 3352.970 ;
        RECT 152.665 3320.690 199.465 3352.330 ;
        RECT 152.035 3277.010 199.465 3320.690 ;
        RECT 147.275 3110.545 151.535 3112.065 ;
        RECT 147.275 3096.360 148.255 3110.545 ;
        RECT 0.000 3094.840 148.255 3096.360 ;
        RECT 0.000 3061.010 143.495 3094.840 ;
        RECT 0.000 3059.670 142.865 3061.010 ;
      LAYER met4 ;
        RECT 0.000 3058.000 24.215 3059.270 ;
      LAYER met4 ;
        RECT 24.615 3058.965 104.600 3059.670 ;
        RECT 0.000 2922.000 25.965 3058.000 ;
        RECT 102.965 3056.000 105.000 3058.000 ;
      LAYER met4 ;
        RECT 105.000 3056.000 129.965 3059.270 ;
      LAYER met4 ;
        RECT 130.365 3058.965 131.065 3059.670 ;
        RECT 129.965 3056.000 131.065 3058.000 ;
        RECT 102.965 3053.000 131.065 3056.000 ;
        RECT 102.965 3051.000 105.000 3053.000 ;
      LAYER met4 ;
        RECT 105.000 3051.000 129.965 3053.000 ;
      LAYER met4 ;
        RECT 129.965 3051.000 131.065 3053.000 ;
        RECT 102.965 3043.000 131.065 3051.000 ;
        RECT 102.965 3041.000 105.000 3043.000 ;
      LAYER met4 ;
        RECT 105.000 3041.000 129.965 3043.000 ;
      LAYER met4 ;
        RECT 129.965 3041.000 131.065 3043.000 ;
        RECT 102.965 3023.000 131.065 3041.000 ;
        RECT 102.965 3021.000 105.000 3023.000 ;
      LAYER met4 ;
        RECT 105.000 3021.000 129.965 3023.000 ;
      LAYER met4 ;
        RECT 129.965 3021.000 131.065 3023.000 ;
        RECT 102.965 3003.000 131.065 3021.000 ;
        RECT 102.965 3001.000 105.000 3003.000 ;
      LAYER met4 ;
        RECT 105.000 3001.000 129.965 3003.000 ;
      LAYER met4 ;
        RECT 129.965 3001.000 131.065 3003.000 ;
        RECT 102.965 2983.000 131.065 3001.000 ;
        RECT 102.965 2981.000 105.000 2983.000 ;
      LAYER met4 ;
        RECT 105.000 2981.000 129.965 2983.000 ;
      LAYER met4 ;
        RECT 129.965 2981.000 131.065 2983.000 ;
        RECT 102.965 2963.000 131.065 2981.000 ;
        RECT 102.965 2961.000 105.000 2963.000 ;
      LAYER met4 ;
        RECT 105.000 2961.000 129.965 2963.000 ;
      LAYER met4 ;
        RECT 129.965 2961.000 131.065 2963.000 ;
        RECT 102.965 2943.000 131.065 2961.000 ;
        RECT 102.965 2941.000 105.000 2943.000 ;
      LAYER met4 ;
        RECT 105.000 2941.000 129.965 2943.000 ;
      LAYER met4 ;
        RECT 129.965 2941.000 131.065 2943.000 ;
        RECT 102.965 2923.000 131.065 2941.000 ;
        RECT 102.965 2922.000 105.000 2923.000 ;
      LAYER met4 ;
        RECT 0.000 2920.730 24.215 2922.000 ;
      LAYER met4 ;
        RECT 24.615 2920.330 104.600 2920.970 ;
      LAYER met4 ;
        RECT 105.000 2920.730 129.965 2923.000 ;
      LAYER met4 ;
        RECT 129.965 2922.000 131.065 2923.000 ;
        RECT 130.365 2920.330 131.065 2920.970 ;
      LAYER met4 ;
        RECT 131.465 2920.730 135.915 3059.270 ;
      LAYER met4 ;
        RECT 136.315 3058.965 136.915 3059.670 ;
        RECT 136.315 2922.000 136.915 3057.000 ;
        RECT 136.315 2920.330 136.915 2920.970 ;
      LAYER met4 ;
        RECT 137.315 2920.730 141.765 3059.270 ;
      LAYER met4 ;
        RECT 142.165 3058.965 142.865 3059.670 ;
        RECT 142.165 2922.000 142.865 3058.000 ;
        RECT 142.165 2920.330 142.865 2920.970 ;
        RECT 0.000 2888.690 142.865 2920.330 ;
      LAYER met4 ;
        RECT 143.265 2889.090 143.595 3060.610 ;
      LAYER met4 ;
        RECT 0.000 2880.360 143.495 2888.690 ;
      LAYER met4 ;
        RECT 143.895 2880.760 146.875 3094.440 ;
      LAYER met4 ;
        RECT 147.275 3059.670 148.255 3094.840 ;
      LAYER met4 ;
        RECT 147.175 3058.000 148.355 3059.270 ;
      LAYER met4 ;
        RECT 147.275 2922.000 148.255 3058.000 ;
      LAYER met4 ;
        RECT 147.175 2920.730 148.355 2922.000 ;
      LAYER met4 ;
        RECT 147.275 2896.065 148.255 2920.330 ;
      LAYER met4 ;
        RECT 148.655 2896.465 151.635 3110.145 ;
        RECT 151.935 3105.090 152.265 3276.610 ;
      LAYER met4 ;
        RECT 152.665 3275.670 199.465 3277.010 ;
        RECT 152.665 3274.965 153.365 3275.670 ;
        RECT 152.665 3136.330 153.365 3136.970 ;
      LAYER met4 ;
        RECT 153.765 3136.730 158.415 3275.270 ;
      LAYER met4 ;
        RECT 158.815 3274.965 159.415 3275.670 ;
        RECT 158.815 3136.330 159.415 3136.970 ;
      LAYER met4 ;
        RECT 159.815 3136.730 163.265 3275.270 ;
      LAYER met4 ;
        RECT 163.665 3274.965 164.265 3275.670 ;
        RECT 163.665 3136.330 164.265 3136.970 ;
      LAYER met4 ;
        RECT 164.665 3136.730 168.115 3275.270 ;
      LAYER met4 ;
        RECT 168.515 3274.965 169.115 3275.670 ;
        RECT 168.515 3136.330 169.115 3136.970 ;
      LAYER met4 ;
        RECT 169.515 3136.730 174.165 3275.270 ;
      LAYER met4 ;
        RECT 174.565 3274.965 175.165 3275.670 ;
        RECT 180.615 3275.365 186.065 3275.670 ;
        RECT 174.565 3136.330 175.165 3136.970 ;
      LAYER met4 ;
        RECT 175.565 3136.730 180.215 3275.270 ;
      LAYER met4 ;
        RECT 180.615 3274.965 181.215 3275.365 ;
        RECT 185.465 3274.965 186.065 3275.365 ;
      LAYER met4 ;
        RECT 181.615 3136.970 185.065 3274.965 ;
      LAYER met4 ;
        RECT 180.615 3136.570 181.215 3136.970 ;
        RECT 185.465 3136.570 186.065 3136.970 ;
      LAYER met4 ;
        RECT 186.465 3136.730 191.115 3275.270 ;
      LAYER met4 ;
        RECT 191.515 3274.965 192.115 3275.670 ;
        RECT 180.615 3136.330 186.065 3136.570 ;
        RECT 191.515 3136.330 192.115 3136.970 ;
      LAYER met4 ;
        RECT 192.515 3136.730 197.965 3275.270 ;
      LAYER met4 ;
        RECT 198.365 3274.965 199.465 3275.670 ;
        RECT 3388.535 3268.330 3389.635 3269.035 ;
      LAYER met4 ;
        RECT 3390.035 3268.730 3395.485 3417.270 ;
      LAYER met4 ;
        RECT 3395.885 3417.030 3396.485 3417.670 ;
        RECT 3401.935 3417.430 3407.385 3417.670 ;
        RECT 3395.885 3268.330 3396.485 3269.035 ;
      LAYER met4 ;
        RECT 3396.885 3268.730 3401.535 3417.270 ;
      LAYER met4 ;
        RECT 3401.935 3417.030 3402.535 3417.430 ;
        RECT 3406.785 3417.030 3407.385 3417.430 ;
      LAYER met4 ;
        RECT 3402.935 3269.035 3406.385 3417.030 ;
      LAYER met4 ;
        RECT 3401.935 3268.635 3402.535 3269.035 ;
        RECT 3406.785 3268.635 3407.385 3269.035 ;
      LAYER met4 ;
        RECT 3407.785 3268.730 3412.435 3417.270 ;
      LAYER met4 ;
        RECT 3412.835 3417.030 3413.435 3417.670 ;
        RECT 3401.935 3268.330 3407.385 3268.635 ;
        RECT 3412.835 3268.330 3413.435 3269.035 ;
      LAYER met4 ;
        RECT 3413.835 3268.730 3418.485 3417.270 ;
      LAYER met4 ;
        RECT 3418.885 3417.030 3419.485 3417.670 ;
        RECT 3418.885 3268.330 3419.485 3269.035 ;
      LAYER met4 ;
        RECT 3419.885 3268.730 3423.335 3417.270 ;
      LAYER met4 ;
        RECT 3423.735 3417.030 3424.335 3417.670 ;
        RECT 3423.735 3268.330 3424.335 3269.035 ;
      LAYER met4 ;
        RECT 3424.735 3268.730 3428.185 3417.270 ;
      LAYER met4 ;
        RECT 3428.585 3417.030 3429.185 3417.670 ;
        RECT 3428.585 3268.330 3429.185 3269.035 ;
      LAYER met4 ;
        RECT 3429.585 3268.730 3434.235 3417.270 ;
      LAYER met4 ;
        RECT 3434.635 3417.030 3435.335 3417.670 ;
        RECT 3434.635 3268.330 3435.335 3269.035 ;
        RECT 3388.535 3266.990 3435.335 3268.330 ;
      LAYER met4 ;
        RECT 3435.735 3267.390 3436.065 3448.910 ;
        RECT 3436.365 3443.855 3439.345 3666.535 ;
      LAYER met4 ;
        RECT 3439.745 3642.670 3440.725 3666.935 ;
      LAYER met4 ;
        RECT 3439.645 3641.000 3440.825 3642.270 ;
      LAYER met4 ;
        RECT 3439.745 3496.000 3440.725 3641.000 ;
      LAYER met4 ;
        RECT 3439.645 3494.730 3440.825 3496.000 ;
      LAYER met4 ;
        RECT 3439.745 3459.160 3440.725 3494.330 ;
      LAYER met4 ;
        RECT 3441.125 3459.560 3444.105 3682.240 ;
      LAYER met4 ;
        RECT 3444.505 3674.310 3588.000 3682.640 ;
      LAYER met4 ;
        RECT 3444.405 3493.390 3444.735 3673.910 ;
      LAYER met4 ;
        RECT 3445.135 3642.670 3588.000 3674.310 ;
        RECT 3445.135 3642.030 3445.835 3642.670 ;
        RECT 3445.135 3496.000 3445.835 3641.000 ;
        RECT 3445.135 3494.330 3445.835 3495.035 ;
      LAYER met4 ;
        RECT 3446.235 3494.730 3450.685 3642.270 ;
      LAYER met4 ;
        RECT 3451.085 3642.030 3451.685 3642.670 ;
        RECT 3451.085 3496.000 3451.685 3641.000 ;
        RECT 3451.085 3494.330 3451.685 3495.035 ;
      LAYER met4 ;
        RECT 3452.085 3494.730 3456.535 3642.270 ;
      LAYER met4 ;
        RECT 3456.935 3642.030 3457.635 3642.670 ;
        RECT 3456.935 3640.000 3458.035 3641.000 ;
      LAYER met4 ;
        RECT 3458.035 3640.000 3483.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3642.030 3563.385 3642.670 ;
      LAYER met4 ;
        RECT 3563.785 3641.000 3588.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.000 3640.000 3485.035 3641.000 ;
        RECT 3456.935 3637.000 3485.035 3640.000 ;
        RECT 3456.935 3635.000 3458.035 3637.000 ;
      LAYER met4 ;
        RECT 3458.035 3635.000 3483.000 3637.000 ;
      LAYER met4 ;
        RECT 3483.000 3635.000 3485.035 3637.000 ;
        RECT 3456.935 3617.000 3485.035 3635.000 ;
        RECT 3456.935 3615.000 3458.035 3617.000 ;
      LAYER met4 ;
        RECT 3458.035 3615.000 3483.000 3617.000 ;
      LAYER met4 ;
        RECT 3483.000 3615.000 3485.035 3617.000 ;
        RECT 3456.935 3597.000 3485.035 3615.000 ;
        RECT 3456.935 3595.000 3458.035 3597.000 ;
      LAYER met4 ;
        RECT 3458.035 3595.000 3483.000 3597.000 ;
      LAYER met4 ;
        RECT 3483.000 3595.000 3485.035 3597.000 ;
        RECT 3456.935 3577.000 3485.035 3595.000 ;
        RECT 3456.935 3575.000 3458.035 3577.000 ;
      LAYER met4 ;
        RECT 3458.035 3575.000 3483.000 3577.000 ;
      LAYER met4 ;
        RECT 3483.000 3575.000 3485.035 3577.000 ;
        RECT 3456.935 3557.000 3485.035 3575.000 ;
        RECT 3456.935 3555.000 3458.035 3557.000 ;
      LAYER met4 ;
        RECT 3458.035 3555.000 3483.000 3557.000 ;
      LAYER met4 ;
        RECT 3483.000 3555.000 3485.035 3557.000 ;
        RECT 3456.935 3537.000 3485.035 3555.000 ;
        RECT 3456.935 3535.000 3458.035 3537.000 ;
      LAYER met4 ;
        RECT 3458.035 3535.000 3483.000 3537.000 ;
      LAYER met4 ;
        RECT 3483.000 3535.000 3485.035 3537.000 ;
        RECT 3456.935 3517.000 3485.035 3535.000 ;
        RECT 3456.935 3515.000 3458.035 3517.000 ;
      LAYER met4 ;
        RECT 3458.035 3515.000 3483.000 3517.000 ;
      LAYER met4 ;
        RECT 3483.000 3515.000 3485.035 3517.000 ;
        RECT 3456.935 3497.000 3485.035 3515.000 ;
        RECT 3456.935 3496.000 3458.035 3497.000 ;
        RECT 3456.935 3494.330 3457.635 3495.035 ;
      LAYER met4 ;
        RECT 3458.035 3494.730 3483.000 3497.000 ;
      LAYER met4 ;
        RECT 3483.000 3496.000 3485.035 3497.000 ;
        RECT 3562.035 3496.000 3588.000 3641.000 ;
        RECT 3483.400 3494.330 3563.385 3495.035 ;
      LAYER met4 ;
        RECT 3563.785 3494.730 3588.000 3496.000 ;
      LAYER met4 ;
        RECT 3445.135 3492.990 3588.000 3494.330 ;
        RECT 3444.505 3459.160 3588.000 3492.990 ;
        RECT 3439.745 3457.640 3588.000 3459.160 ;
        RECT 3439.745 3443.455 3440.725 3457.640 ;
        RECT 3436.465 3441.935 3440.725 3443.455 ;
        RECT 3388.535 3223.310 3435.965 3266.990 ;
        RECT 3388.535 3191.670 3435.335 3223.310 ;
        RECT 3388.535 3191.030 3389.635 3191.670 ;
        RECT 198.365 3136.330 199.465 3136.970 ;
        RECT 152.665 3104.690 199.465 3136.330 ;
        RECT 152.035 3061.010 199.465 3104.690 ;
        RECT 147.275 2894.545 151.535 2896.065 ;
        RECT 147.275 2880.360 148.255 2894.545 ;
        RECT 0.000 2878.840 148.255 2880.360 ;
        RECT 0.000 2845.010 143.495 2878.840 ;
        RECT 0.000 2843.670 142.865 2845.010 ;
      LAYER met4 ;
        RECT 0.000 2842.000 24.215 2843.270 ;
      LAYER met4 ;
        RECT 24.615 2842.965 104.600 2843.670 ;
        RECT 0.000 2706.000 25.965 2842.000 ;
        RECT 102.965 2840.000 105.000 2842.000 ;
      LAYER met4 ;
        RECT 105.000 2840.000 129.965 2843.270 ;
      LAYER met4 ;
        RECT 130.365 2842.965 131.065 2843.670 ;
        RECT 129.965 2840.000 131.065 2842.000 ;
        RECT 102.965 2837.000 131.065 2840.000 ;
        RECT 102.965 2835.000 105.000 2837.000 ;
      LAYER met4 ;
        RECT 105.000 2835.000 129.965 2837.000 ;
      LAYER met4 ;
        RECT 129.965 2835.000 131.065 2837.000 ;
        RECT 102.965 2827.000 131.065 2835.000 ;
        RECT 102.965 2825.000 105.000 2827.000 ;
      LAYER met4 ;
        RECT 105.000 2825.000 129.965 2827.000 ;
      LAYER met4 ;
        RECT 129.965 2825.000 131.065 2827.000 ;
        RECT 102.965 2807.000 131.065 2825.000 ;
        RECT 102.965 2805.000 105.000 2807.000 ;
      LAYER met4 ;
        RECT 105.000 2805.000 129.965 2807.000 ;
      LAYER met4 ;
        RECT 129.965 2805.000 131.065 2807.000 ;
        RECT 102.965 2787.000 131.065 2805.000 ;
        RECT 102.965 2785.000 105.000 2787.000 ;
      LAYER met4 ;
        RECT 105.000 2785.000 129.965 2787.000 ;
      LAYER met4 ;
        RECT 129.965 2785.000 131.065 2787.000 ;
        RECT 102.965 2767.000 131.065 2785.000 ;
        RECT 102.965 2765.000 105.000 2767.000 ;
      LAYER met4 ;
        RECT 105.000 2765.000 129.965 2767.000 ;
      LAYER met4 ;
        RECT 129.965 2765.000 131.065 2767.000 ;
        RECT 102.965 2747.000 131.065 2765.000 ;
        RECT 102.965 2745.000 105.000 2747.000 ;
      LAYER met4 ;
        RECT 105.000 2745.000 129.965 2747.000 ;
      LAYER met4 ;
        RECT 129.965 2745.000 131.065 2747.000 ;
        RECT 102.965 2727.000 131.065 2745.000 ;
        RECT 102.965 2725.000 105.000 2727.000 ;
      LAYER met4 ;
        RECT 105.000 2725.000 129.965 2727.000 ;
      LAYER met4 ;
        RECT 129.965 2725.000 131.065 2727.000 ;
        RECT 102.965 2707.000 131.065 2725.000 ;
        RECT 102.965 2706.000 105.000 2707.000 ;
      LAYER met4 ;
        RECT 0.000 2704.730 24.215 2706.000 ;
      LAYER met4 ;
        RECT 24.615 2704.330 104.600 2704.970 ;
      LAYER met4 ;
        RECT 105.000 2704.730 129.965 2707.000 ;
      LAYER met4 ;
        RECT 129.965 2706.000 131.065 2707.000 ;
        RECT 130.365 2704.330 131.065 2704.970 ;
      LAYER met4 ;
        RECT 131.465 2704.730 135.915 2843.270 ;
      LAYER met4 ;
        RECT 136.315 2842.965 136.915 2843.670 ;
        RECT 136.315 2706.000 136.915 2841.000 ;
        RECT 136.315 2704.330 136.915 2704.970 ;
      LAYER met4 ;
        RECT 137.315 2704.730 141.765 2843.270 ;
      LAYER met4 ;
        RECT 142.165 2842.965 142.865 2843.670 ;
        RECT 142.165 2706.000 142.865 2842.000 ;
        RECT 142.165 2704.330 142.865 2704.970 ;
        RECT 0.000 2672.690 142.865 2704.330 ;
      LAYER met4 ;
        RECT 143.265 2673.090 143.595 2844.610 ;
      LAYER met4 ;
        RECT 0.000 2664.360 143.495 2672.690 ;
      LAYER met4 ;
        RECT 143.895 2664.760 146.875 2878.440 ;
      LAYER met4 ;
        RECT 147.275 2843.670 148.255 2878.840 ;
      LAYER met4 ;
        RECT 147.175 2842.000 148.355 2843.270 ;
      LAYER met4 ;
        RECT 147.275 2706.000 148.255 2842.000 ;
      LAYER met4 ;
        RECT 147.175 2704.730 148.355 2706.000 ;
      LAYER met4 ;
        RECT 147.275 2680.065 148.255 2704.330 ;
      LAYER met4 ;
        RECT 148.655 2680.465 151.635 2894.145 ;
        RECT 151.935 2889.090 152.265 3060.610 ;
      LAYER met4 ;
        RECT 152.665 3059.670 199.465 3061.010 ;
        RECT 152.665 3058.965 153.365 3059.670 ;
        RECT 152.665 2920.330 153.365 2920.970 ;
      LAYER met4 ;
        RECT 153.765 2920.730 158.415 3059.270 ;
      LAYER met4 ;
        RECT 158.815 3058.965 159.415 3059.670 ;
        RECT 158.815 2920.330 159.415 2920.970 ;
      LAYER met4 ;
        RECT 159.815 2920.730 163.265 3059.270 ;
      LAYER met4 ;
        RECT 163.665 3058.965 164.265 3059.670 ;
        RECT 163.665 2920.330 164.265 2920.970 ;
      LAYER met4 ;
        RECT 164.665 2920.730 168.115 3059.270 ;
      LAYER met4 ;
        RECT 168.515 3058.965 169.115 3059.670 ;
        RECT 168.515 2920.330 169.115 2920.970 ;
      LAYER met4 ;
        RECT 169.515 2920.730 174.165 3059.270 ;
      LAYER met4 ;
        RECT 174.565 3058.965 175.165 3059.670 ;
        RECT 180.615 3059.365 186.065 3059.670 ;
        RECT 174.565 2920.330 175.165 2920.970 ;
      LAYER met4 ;
        RECT 175.565 2920.730 180.215 3059.270 ;
      LAYER met4 ;
        RECT 180.615 3058.965 181.215 3059.365 ;
        RECT 185.465 3058.965 186.065 3059.365 ;
      LAYER met4 ;
        RECT 181.615 2920.970 185.065 3058.965 ;
      LAYER met4 ;
        RECT 180.615 2920.570 181.215 2920.970 ;
        RECT 185.465 2920.570 186.065 2920.970 ;
      LAYER met4 ;
        RECT 186.465 2920.730 191.115 3059.270 ;
      LAYER met4 ;
        RECT 191.515 3058.965 192.115 3059.670 ;
        RECT 180.615 2920.330 186.065 2920.570 ;
        RECT 191.515 2920.330 192.115 2920.970 ;
      LAYER met4 ;
        RECT 192.515 2920.730 197.965 3059.270 ;
      LAYER met4 ;
        RECT 198.365 3058.965 199.465 3059.670 ;
        RECT 3388.535 3043.330 3389.635 3044.035 ;
      LAYER met4 ;
        RECT 3390.035 3043.730 3395.485 3191.270 ;
      LAYER met4 ;
        RECT 3395.885 3191.030 3396.485 3191.670 ;
        RECT 3401.935 3191.430 3407.385 3191.670 ;
        RECT 3395.885 3043.330 3396.485 3044.035 ;
      LAYER met4 ;
        RECT 3396.885 3043.730 3401.535 3191.270 ;
      LAYER met4 ;
        RECT 3401.935 3191.030 3402.535 3191.430 ;
        RECT 3406.785 3191.030 3407.385 3191.430 ;
      LAYER met4 ;
        RECT 3402.935 3044.035 3406.385 3191.030 ;
      LAYER met4 ;
        RECT 3401.935 3043.635 3402.535 3044.035 ;
        RECT 3406.785 3043.635 3407.385 3044.035 ;
      LAYER met4 ;
        RECT 3407.785 3043.730 3412.435 3191.270 ;
      LAYER met4 ;
        RECT 3412.835 3191.030 3413.435 3191.670 ;
        RECT 3401.935 3043.330 3407.385 3043.635 ;
        RECT 3412.835 3043.330 3413.435 3044.035 ;
      LAYER met4 ;
        RECT 3413.835 3043.730 3418.485 3191.270 ;
      LAYER met4 ;
        RECT 3418.885 3191.030 3419.485 3191.670 ;
        RECT 3418.885 3043.330 3419.485 3044.035 ;
      LAYER met4 ;
        RECT 3419.885 3043.730 3423.335 3191.270 ;
      LAYER met4 ;
        RECT 3423.735 3191.030 3424.335 3191.670 ;
        RECT 3423.735 3043.330 3424.335 3044.035 ;
      LAYER met4 ;
        RECT 3424.735 3043.730 3428.185 3191.270 ;
      LAYER met4 ;
        RECT 3428.585 3191.030 3429.185 3191.670 ;
        RECT 3428.585 3043.330 3429.185 3044.035 ;
      LAYER met4 ;
        RECT 3429.585 3043.730 3434.235 3191.270 ;
      LAYER met4 ;
        RECT 3434.635 3191.030 3435.335 3191.670 ;
        RECT 3434.635 3043.330 3435.335 3044.035 ;
        RECT 3388.535 3041.990 3435.335 3043.330 ;
      LAYER met4 ;
        RECT 3435.735 3042.390 3436.065 3222.910 ;
        RECT 3436.365 3217.855 3439.345 3441.535 ;
      LAYER met4 ;
        RECT 3439.745 3417.670 3440.725 3441.935 ;
      LAYER met4 ;
        RECT 3439.645 3416.000 3440.825 3417.270 ;
      LAYER met4 ;
        RECT 3439.745 3270.000 3440.725 3416.000 ;
      LAYER met4 ;
        RECT 3439.645 3268.730 3440.825 3270.000 ;
      LAYER met4 ;
        RECT 3439.745 3233.160 3440.725 3268.330 ;
      LAYER met4 ;
        RECT 3441.125 3233.560 3444.105 3457.240 ;
      LAYER met4 ;
        RECT 3444.505 3449.310 3588.000 3457.640 ;
      LAYER met4 ;
        RECT 3444.405 3267.390 3444.735 3448.910 ;
      LAYER met4 ;
        RECT 3445.135 3417.670 3588.000 3449.310 ;
        RECT 3445.135 3417.030 3445.835 3417.670 ;
        RECT 3445.135 3270.000 3445.835 3416.000 ;
        RECT 3445.135 3268.330 3445.835 3269.035 ;
      LAYER met4 ;
        RECT 3446.235 3268.730 3450.685 3417.270 ;
      LAYER met4 ;
        RECT 3451.085 3417.030 3451.685 3417.670 ;
        RECT 3451.085 3270.000 3451.685 3415.000 ;
        RECT 3451.085 3268.330 3451.685 3269.035 ;
      LAYER met4 ;
        RECT 3452.085 3268.730 3456.535 3417.270 ;
      LAYER met4 ;
        RECT 3456.935 3417.030 3457.635 3417.670 ;
        RECT 3456.935 3414.000 3458.035 3416.000 ;
      LAYER met4 ;
        RECT 3458.035 3414.000 3483.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3417.030 3563.385 3417.670 ;
      LAYER met4 ;
        RECT 3563.785 3416.000 3588.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.000 3414.000 3485.035 3416.000 ;
        RECT 3456.935 3411.000 3485.035 3414.000 ;
        RECT 3456.935 3409.000 3458.035 3411.000 ;
      LAYER met4 ;
        RECT 3458.035 3409.000 3483.000 3411.000 ;
      LAYER met4 ;
        RECT 3483.000 3409.000 3485.035 3411.000 ;
        RECT 3456.935 3391.000 3485.035 3409.000 ;
        RECT 3456.935 3389.000 3458.035 3391.000 ;
      LAYER met4 ;
        RECT 3458.035 3389.000 3483.000 3391.000 ;
      LAYER met4 ;
        RECT 3483.000 3389.000 3485.035 3391.000 ;
        RECT 3456.935 3371.000 3485.035 3389.000 ;
        RECT 3456.935 3369.000 3458.035 3371.000 ;
      LAYER met4 ;
        RECT 3458.035 3369.000 3483.000 3371.000 ;
      LAYER met4 ;
        RECT 3483.000 3369.000 3485.035 3371.000 ;
        RECT 3456.935 3351.000 3485.035 3369.000 ;
        RECT 3456.935 3349.000 3458.035 3351.000 ;
      LAYER met4 ;
        RECT 3458.035 3349.000 3483.000 3351.000 ;
      LAYER met4 ;
        RECT 3483.000 3349.000 3485.035 3351.000 ;
        RECT 3456.935 3331.000 3485.035 3349.000 ;
        RECT 3456.935 3329.000 3458.035 3331.000 ;
      LAYER met4 ;
        RECT 3458.035 3329.000 3483.000 3331.000 ;
      LAYER met4 ;
        RECT 3483.000 3329.000 3485.035 3331.000 ;
        RECT 3456.935 3311.000 3485.035 3329.000 ;
        RECT 3456.935 3309.000 3458.035 3311.000 ;
      LAYER met4 ;
        RECT 3458.035 3309.000 3483.000 3311.000 ;
      LAYER met4 ;
        RECT 3483.000 3309.000 3485.035 3311.000 ;
        RECT 3456.935 3291.000 3485.035 3309.000 ;
        RECT 3456.935 3289.000 3458.035 3291.000 ;
      LAYER met4 ;
        RECT 3458.035 3289.000 3483.000 3291.000 ;
      LAYER met4 ;
        RECT 3483.000 3289.000 3485.035 3291.000 ;
        RECT 3456.935 3271.000 3485.035 3289.000 ;
        RECT 3456.935 3270.000 3458.035 3271.000 ;
        RECT 3456.935 3268.330 3457.635 3269.035 ;
      LAYER met4 ;
        RECT 3458.035 3268.730 3483.000 3271.000 ;
      LAYER met4 ;
        RECT 3483.000 3270.000 3485.035 3271.000 ;
        RECT 3562.035 3270.000 3588.000 3416.000 ;
        RECT 3483.400 3268.330 3563.385 3269.035 ;
      LAYER met4 ;
        RECT 3563.785 3268.730 3588.000 3270.000 ;
      LAYER met4 ;
        RECT 3445.135 3266.990 3588.000 3268.330 ;
        RECT 3444.505 3233.160 3588.000 3266.990 ;
        RECT 3439.745 3231.640 3588.000 3233.160 ;
        RECT 3439.745 3217.455 3440.725 3231.640 ;
        RECT 3436.465 3215.935 3440.725 3217.455 ;
        RECT 3388.535 2998.310 3435.965 3041.990 ;
        RECT 3388.535 2966.670 3435.335 2998.310 ;
        RECT 3388.535 2966.030 3389.635 2966.670 ;
        RECT 198.365 2920.330 199.465 2920.970 ;
        RECT 152.665 2888.690 199.465 2920.330 ;
        RECT 152.035 2845.010 199.465 2888.690 ;
        RECT 147.275 2678.545 151.535 2680.065 ;
        RECT 147.275 2664.360 148.255 2678.545 ;
        RECT 0.000 2662.840 148.255 2664.360 ;
        RECT 0.000 2629.010 143.495 2662.840 ;
        RECT 0.000 2627.670 142.865 2629.010 ;
      LAYER met4 ;
        RECT 0.000 2626.000 24.215 2627.270 ;
      LAYER met4 ;
        RECT 24.615 2626.965 104.600 2627.670 ;
        RECT 0.000 2490.000 25.965 2626.000 ;
        RECT 102.965 2624.000 105.000 2626.000 ;
      LAYER met4 ;
        RECT 105.000 2624.000 129.965 2627.270 ;
      LAYER met4 ;
        RECT 130.365 2626.965 131.065 2627.670 ;
        RECT 129.965 2624.000 131.065 2626.000 ;
        RECT 102.965 2621.000 131.065 2624.000 ;
        RECT 102.965 2619.000 105.000 2621.000 ;
      LAYER met4 ;
        RECT 105.000 2619.000 129.965 2621.000 ;
      LAYER met4 ;
        RECT 129.965 2619.000 131.065 2621.000 ;
        RECT 102.965 2611.000 131.065 2619.000 ;
        RECT 102.965 2609.000 105.000 2611.000 ;
      LAYER met4 ;
        RECT 105.000 2609.000 129.965 2611.000 ;
      LAYER met4 ;
        RECT 129.965 2609.000 131.065 2611.000 ;
        RECT 102.965 2591.000 131.065 2609.000 ;
        RECT 102.965 2589.000 105.000 2591.000 ;
      LAYER met4 ;
        RECT 105.000 2589.000 129.965 2591.000 ;
      LAYER met4 ;
        RECT 129.965 2589.000 131.065 2591.000 ;
        RECT 102.965 2571.000 131.065 2589.000 ;
        RECT 102.965 2569.000 105.000 2571.000 ;
      LAYER met4 ;
        RECT 105.000 2569.000 129.965 2571.000 ;
      LAYER met4 ;
        RECT 129.965 2569.000 131.065 2571.000 ;
        RECT 102.965 2551.000 131.065 2569.000 ;
        RECT 102.965 2549.000 105.000 2551.000 ;
      LAYER met4 ;
        RECT 105.000 2549.000 129.965 2551.000 ;
      LAYER met4 ;
        RECT 129.965 2549.000 131.065 2551.000 ;
        RECT 102.965 2531.000 131.065 2549.000 ;
        RECT 102.965 2529.000 105.000 2531.000 ;
      LAYER met4 ;
        RECT 105.000 2529.000 129.965 2531.000 ;
      LAYER met4 ;
        RECT 129.965 2529.000 131.065 2531.000 ;
        RECT 102.965 2511.000 131.065 2529.000 ;
        RECT 102.965 2509.000 105.000 2511.000 ;
      LAYER met4 ;
        RECT 105.000 2509.000 129.965 2511.000 ;
      LAYER met4 ;
        RECT 129.965 2509.000 131.065 2511.000 ;
        RECT 102.965 2491.000 131.065 2509.000 ;
        RECT 102.965 2490.000 105.000 2491.000 ;
      LAYER met4 ;
        RECT 0.000 2488.730 24.215 2490.000 ;
      LAYER met4 ;
        RECT 24.615 2488.330 104.600 2489.035 ;
      LAYER met4 ;
        RECT 105.000 2488.730 129.965 2491.000 ;
      LAYER met4 ;
        RECT 129.965 2490.000 131.065 2491.000 ;
        RECT 130.365 2488.330 131.065 2489.035 ;
      LAYER met4 ;
        RECT 131.465 2488.730 135.915 2627.270 ;
      LAYER met4 ;
        RECT 136.315 2626.965 136.915 2627.670 ;
        RECT 136.315 2490.000 136.915 2625.000 ;
        RECT 136.315 2488.330 136.915 2489.035 ;
      LAYER met4 ;
        RECT 137.315 2488.730 141.765 2627.270 ;
      LAYER met4 ;
        RECT 142.165 2626.965 142.865 2627.670 ;
        RECT 142.165 2490.000 142.865 2626.000 ;
        RECT 142.165 2488.330 142.865 2489.035 ;
        RECT 0.000 2416.670 142.865 2488.330 ;
      LAYER met4 ;
        RECT 0.000 2415.000 24.215 2416.270 ;
      LAYER met4 ;
        RECT 24.615 2415.965 104.600 2416.670 ;
        RECT 0.000 2279.000 25.965 2415.000 ;
        RECT 102.965 2413.000 105.000 2415.000 ;
      LAYER met4 ;
        RECT 105.000 2413.000 129.965 2416.270 ;
      LAYER met4 ;
        RECT 130.365 2415.965 131.065 2416.670 ;
        RECT 129.965 2413.000 131.065 2415.000 ;
        RECT 102.965 2410.000 131.065 2413.000 ;
        RECT 102.965 2408.000 105.000 2410.000 ;
      LAYER met4 ;
        RECT 105.000 2408.000 129.965 2410.000 ;
      LAYER met4 ;
        RECT 129.965 2408.000 131.065 2410.000 ;
        RECT 102.965 2400.000 131.065 2408.000 ;
        RECT 102.965 2398.000 105.000 2400.000 ;
      LAYER met4 ;
        RECT 105.000 2398.000 129.965 2400.000 ;
      LAYER met4 ;
        RECT 129.965 2398.000 131.065 2400.000 ;
        RECT 102.965 2380.000 131.065 2398.000 ;
        RECT 102.965 2378.000 105.000 2380.000 ;
      LAYER met4 ;
        RECT 105.000 2378.000 129.965 2380.000 ;
      LAYER met4 ;
        RECT 129.965 2378.000 131.065 2380.000 ;
        RECT 102.965 2360.000 131.065 2378.000 ;
        RECT 102.965 2358.000 105.000 2360.000 ;
      LAYER met4 ;
        RECT 105.000 2358.000 129.965 2360.000 ;
      LAYER met4 ;
        RECT 129.965 2358.000 131.065 2360.000 ;
        RECT 102.965 2340.000 131.065 2358.000 ;
        RECT 102.965 2338.000 105.000 2340.000 ;
      LAYER met4 ;
        RECT 105.000 2338.000 129.965 2340.000 ;
      LAYER met4 ;
        RECT 129.965 2338.000 131.065 2340.000 ;
        RECT 102.965 2320.000 131.065 2338.000 ;
        RECT 102.965 2318.000 105.000 2320.000 ;
      LAYER met4 ;
        RECT 105.000 2318.000 129.965 2320.000 ;
      LAYER met4 ;
        RECT 129.965 2318.000 131.065 2320.000 ;
        RECT 102.965 2300.000 131.065 2318.000 ;
        RECT 102.965 2298.000 105.000 2300.000 ;
      LAYER met4 ;
        RECT 105.000 2298.000 129.965 2300.000 ;
      LAYER met4 ;
        RECT 129.965 2298.000 131.065 2300.000 ;
        RECT 102.965 2280.000 131.065 2298.000 ;
        RECT 102.965 2279.000 105.000 2280.000 ;
      LAYER met4 ;
        RECT 0.000 2277.730 24.215 2279.000 ;
      LAYER met4 ;
        RECT 24.615 2277.330 104.600 2279.000 ;
      LAYER met4 ;
        RECT 105.000 2277.730 129.965 2280.000 ;
      LAYER met4 ;
        RECT 129.965 2279.000 131.065 2280.000 ;
        RECT 130.365 2277.330 131.065 2279.000 ;
      LAYER met4 ;
        RECT 131.465 2277.730 135.915 2416.270 ;
      LAYER met4 ;
        RECT 136.315 2415.965 136.915 2416.670 ;
        RECT 136.315 2277.330 136.915 2414.000 ;
      LAYER met4 ;
        RECT 137.315 2277.730 141.765 2416.270 ;
      LAYER met4 ;
        RECT 142.165 2415.965 142.865 2416.670 ;
        RECT 142.165 2277.330 142.865 2415.000 ;
        RECT 0.000 2205.670 142.865 2277.330 ;
      LAYER met4 ;
        RECT 0.000 2204.000 24.215 2205.270 ;
      LAYER met4 ;
        RECT 24.615 2204.965 104.600 2205.670 ;
        RECT 0.000 2068.000 25.965 2204.000 ;
        RECT 102.965 2202.000 105.000 2204.000 ;
      LAYER met4 ;
        RECT 105.000 2202.000 129.965 2205.270 ;
      LAYER met4 ;
        RECT 130.365 2204.965 131.065 2205.670 ;
        RECT 129.965 2202.000 131.065 2204.000 ;
        RECT 102.965 2199.000 131.065 2202.000 ;
        RECT 102.965 2197.000 105.000 2199.000 ;
      LAYER met4 ;
        RECT 105.000 2197.000 129.965 2199.000 ;
      LAYER met4 ;
        RECT 129.965 2197.000 131.065 2199.000 ;
        RECT 102.965 2189.000 131.065 2197.000 ;
        RECT 102.965 2187.000 105.000 2189.000 ;
      LAYER met4 ;
        RECT 105.000 2187.000 129.965 2189.000 ;
      LAYER met4 ;
        RECT 129.965 2187.000 131.065 2189.000 ;
        RECT 102.965 2169.000 131.065 2187.000 ;
        RECT 102.965 2167.000 105.000 2169.000 ;
      LAYER met4 ;
        RECT 105.000 2167.000 129.965 2169.000 ;
      LAYER met4 ;
        RECT 129.965 2167.000 131.065 2169.000 ;
        RECT 102.965 2149.000 131.065 2167.000 ;
        RECT 102.965 2147.000 105.000 2149.000 ;
      LAYER met4 ;
        RECT 105.000 2147.000 129.965 2149.000 ;
      LAYER met4 ;
        RECT 129.965 2147.000 131.065 2149.000 ;
        RECT 102.965 2129.000 131.065 2147.000 ;
        RECT 102.965 2127.000 105.000 2129.000 ;
      LAYER met4 ;
        RECT 105.000 2127.000 129.965 2129.000 ;
      LAYER met4 ;
        RECT 129.965 2127.000 131.065 2129.000 ;
        RECT 102.965 2109.000 131.065 2127.000 ;
        RECT 102.965 2107.000 105.000 2109.000 ;
      LAYER met4 ;
        RECT 105.000 2107.000 129.965 2109.000 ;
      LAYER met4 ;
        RECT 129.965 2107.000 131.065 2109.000 ;
        RECT 102.965 2089.000 131.065 2107.000 ;
        RECT 102.965 2087.000 105.000 2089.000 ;
      LAYER met4 ;
        RECT 105.000 2087.000 129.965 2089.000 ;
      LAYER met4 ;
        RECT 129.965 2087.000 131.065 2089.000 ;
        RECT 102.965 2069.000 131.065 2087.000 ;
        RECT 102.965 2068.000 105.000 2069.000 ;
      LAYER met4 ;
        RECT 0.000 2066.730 24.215 2068.000 ;
      LAYER met4 ;
        RECT 24.615 2066.330 104.600 2066.970 ;
      LAYER met4 ;
        RECT 105.000 2066.730 129.965 2069.000 ;
      LAYER met4 ;
        RECT 129.965 2068.000 131.065 2069.000 ;
        RECT 130.365 2066.330 131.065 2066.970 ;
      LAYER met4 ;
        RECT 131.465 2066.730 135.915 2205.270 ;
      LAYER met4 ;
        RECT 136.315 2204.965 136.915 2205.670 ;
        RECT 136.315 2068.000 136.915 2203.000 ;
        RECT 136.315 2066.330 136.915 2066.970 ;
      LAYER met4 ;
        RECT 137.315 2066.730 141.765 2205.270 ;
      LAYER met4 ;
        RECT 142.165 2204.965 142.865 2205.670 ;
        RECT 142.165 2068.000 142.865 2204.000 ;
        RECT 142.165 2066.330 142.865 2066.970 ;
        RECT 0.000 2034.690 142.865 2066.330 ;
      LAYER met4 ;
        RECT 143.265 2035.090 143.595 2628.610 ;
      LAYER met4 ;
        RECT 0.000 2026.360 143.495 2034.690 ;
      LAYER met4 ;
        RECT 143.895 2026.760 146.875 2662.440 ;
      LAYER met4 ;
        RECT 147.275 2627.670 148.255 2662.840 ;
      LAYER met4 ;
        RECT 147.175 2626.000 148.355 2627.270 ;
      LAYER met4 ;
        RECT 147.275 2490.000 148.255 2626.000 ;
      LAYER met4 ;
        RECT 147.175 2488.730 148.355 2490.000 ;
      LAYER met4 ;
        RECT 147.275 2416.670 148.255 2488.330 ;
      LAYER met4 ;
        RECT 147.175 2415.000 148.355 2416.270 ;
      LAYER met4 ;
        RECT 147.275 2279.000 148.255 2415.000 ;
      LAYER met4 ;
        RECT 147.175 2277.730 148.355 2279.000 ;
      LAYER met4 ;
        RECT 147.275 2205.670 148.255 2277.330 ;
      LAYER met4 ;
        RECT 147.175 2204.000 148.355 2205.270 ;
      LAYER met4 ;
        RECT 147.275 2068.000 148.255 2204.000 ;
      LAYER met4 ;
        RECT 147.175 2066.730 148.355 2068.000 ;
      LAYER met4 ;
        RECT 147.275 2042.065 148.255 2066.330 ;
      LAYER met4 ;
        RECT 148.655 2042.465 151.635 2678.145 ;
        RECT 151.935 2673.090 152.265 2844.610 ;
      LAYER met4 ;
        RECT 152.665 2843.670 199.465 2845.010 ;
        RECT 152.665 2842.965 153.365 2843.670 ;
        RECT 152.665 2704.330 153.365 2704.970 ;
      LAYER met4 ;
        RECT 153.765 2704.730 158.415 2843.270 ;
      LAYER met4 ;
        RECT 158.815 2842.965 159.415 2843.670 ;
        RECT 158.815 2704.330 159.415 2704.970 ;
      LAYER met4 ;
        RECT 159.815 2704.730 163.265 2843.270 ;
      LAYER met4 ;
        RECT 163.665 2842.965 164.265 2843.670 ;
        RECT 163.665 2704.330 164.265 2704.970 ;
      LAYER met4 ;
        RECT 164.665 2704.730 168.115 2843.270 ;
      LAYER met4 ;
        RECT 168.515 2842.965 169.115 2843.670 ;
        RECT 168.515 2704.330 169.115 2704.970 ;
      LAYER met4 ;
        RECT 169.515 2704.730 174.165 2843.270 ;
      LAYER met4 ;
        RECT 174.565 2842.965 175.165 2843.670 ;
        RECT 180.615 2843.365 186.065 2843.670 ;
        RECT 174.565 2704.330 175.165 2704.970 ;
      LAYER met4 ;
        RECT 175.565 2704.730 180.215 2843.270 ;
      LAYER met4 ;
        RECT 180.615 2842.965 181.215 2843.365 ;
        RECT 185.465 2842.965 186.065 2843.365 ;
      LAYER met4 ;
        RECT 181.615 2704.970 185.065 2842.965 ;
      LAYER met4 ;
        RECT 180.615 2704.570 181.215 2704.970 ;
        RECT 185.465 2704.570 186.065 2704.970 ;
      LAYER met4 ;
        RECT 186.465 2704.730 191.115 2843.270 ;
      LAYER met4 ;
        RECT 191.515 2842.965 192.115 2843.670 ;
        RECT 180.615 2704.330 186.065 2704.570 ;
        RECT 191.515 2704.330 192.115 2704.970 ;
      LAYER met4 ;
        RECT 192.515 2704.730 197.965 2843.270 ;
      LAYER met4 ;
        RECT 198.365 2842.965 199.465 2843.670 ;
        RECT 3388.535 2817.330 3389.635 2818.035 ;
      LAYER met4 ;
        RECT 3390.035 2817.730 3395.485 2966.270 ;
      LAYER met4 ;
        RECT 3395.885 2966.030 3396.485 2966.670 ;
        RECT 3401.935 2966.430 3407.385 2966.670 ;
        RECT 3395.885 2817.330 3396.485 2818.035 ;
      LAYER met4 ;
        RECT 3396.885 2817.730 3401.535 2966.270 ;
      LAYER met4 ;
        RECT 3401.935 2966.030 3402.535 2966.430 ;
        RECT 3406.785 2966.030 3407.385 2966.430 ;
      LAYER met4 ;
        RECT 3402.935 2818.035 3406.385 2966.030 ;
      LAYER met4 ;
        RECT 3401.935 2817.635 3402.535 2818.035 ;
        RECT 3406.785 2817.635 3407.385 2818.035 ;
      LAYER met4 ;
        RECT 3407.785 2817.730 3412.435 2966.270 ;
      LAYER met4 ;
        RECT 3412.835 2966.030 3413.435 2966.670 ;
        RECT 3401.935 2817.330 3407.385 2817.635 ;
        RECT 3412.835 2817.330 3413.435 2818.035 ;
      LAYER met4 ;
        RECT 3413.835 2817.730 3418.485 2966.270 ;
      LAYER met4 ;
        RECT 3418.885 2966.030 3419.485 2966.670 ;
        RECT 3418.885 2817.330 3419.485 2818.035 ;
      LAYER met4 ;
        RECT 3419.885 2817.730 3423.335 2966.270 ;
      LAYER met4 ;
        RECT 3423.735 2966.030 3424.335 2966.670 ;
        RECT 3423.735 2817.330 3424.335 2818.035 ;
      LAYER met4 ;
        RECT 3424.735 2817.730 3428.185 2966.270 ;
      LAYER met4 ;
        RECT 3428.585 2966.030 3429.185 2966.670 ;
        RECT 3428.585 2817.330 3429.185 2818.035 ;
      LAYER met4 ;
        RECT 3429.585 2817.730 3434.235 2966.270 ;
      LAYER met4 ;
        RECT 3434.635 2966.030 3435.335 2966.670 ;
        RECT 3434.635 2817.330 3435.335 2818.035 ;
        RECT 3388.535 2815.990 3435.335 2817.330 ;
      LAYER met4 ;
        RECT 3435.735 2816.390 3436.065 2997.910 ;
        RECT 3436.365 2992.855 3439.345 3215.535 ;
      LAYER met4 ;
        RECT 3439.745 3191.670 3440.725 3215.935 ;
      LAYER met4 ;
        RECT 3439.645 3190.000 3440.825 3191.270 ;
      LAYER met4 ;
        RECT 3439.745 3045.000 3440.725 3190.000 ;
      LAYER met4 ;
        RECT 3439.645 3043.730 3440.825 3045.000 ;
      LAYER met4 ;
        RECT 3439.745 3008.160 3440.725 3043.330 ;
      LAYER met4 ;
        RECT 3441.125 3008.560 3444.105 3231.240 ;
      LAYER met4 ;
        RECT 3444.505 3223.310 3588.000 3231.640 ;
      LAYER met4 ;
        RECT 3444.405 3042.390 3444.735 3222.910 ;
      LAYER met4 ;
        RECT 3445.135 3191.670 3588.000 3223.310 ;
        RECT 3445.135 3191.030 3445.835 3191.670 ;
        RECT 3445.135 3045.000 3445.835 3190.000 ;
        RECT 3445.135 3043.330 3445.835 3044.035 ;
      LAYER met4 ;
        RECT 3446.235 3043.730 3450.685 3191.270 ;
      LAYER met4 ;
        RECT 3451.085 3191.030 3451.685 3191.670 ;
        RECT 3451.085 3045.000 3451.685 3190.000 ;
        RECT 3451.085 3043.330 3451.685 3044.035 ;
      LAYER met4 ;
        RECT 3452.085 3043.730 3456.535 3191.270 ;
      LAYER met4 ;
        RECT 3456.935 3191.030 3457.635 3191.670 ;
        RECT 3456.935 3189.000 3458.035 3190.000 ;
      LAYER met4 ;
        RECT 3458.035 3189.000 3483.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3191.030 3563.385 3191.670 ;
      LAYER met4 ;
        RECT 3563.785 3190.000 3588.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.000 3189.000 3485.035 3190.000 ;
        RECT 3456.935 3186.000 3485.035 3189.000 ;
        RECT 3456.935 3184.000 3458.035 3186.000 ;
      LAYER met4 ;
        RECT 3458.035 3184.000 3483.000 3186.000 ;
      LAYER met4 ;
        RECT 3483.000 3184.000 3485.035 3186.000 ;
        RECT 3456.935 3166.000 3485.035 3184.000 ;
        RECT 3456.935 3164.000 3458.035 3166.000 ;
      LAYER met4 ;
        RECT 3458.035 3164.000 3483.000 3166.000 ;
      LAYER met4 ;
        RECT 3483.000 3164.000 3485.035 3166.000 ;
        RECT 3456.935 3146.000 3485.035 3164.000 ;
        RECT 3456.935 3144.000 3458.035 3146.000 ;
      LAYER met4 ;
        RECT 3458.035 3144.000 3483.000 3146.000 ;
      LAYER met4 ;
        RECT 3483.000 3144.000 3485.035 3146.000 ;
        RECT 3456.935 3126.000 3485.035 3144.000 ;
        RECT 3456.935 3124.000 3458.035 3126.000 ;
      LAYER met4 ;
        RECT 3458.035 3124.000 3483.000 3126.000 ;
      LAYER met4 ;
        RECT 3483.000 3124.000 3485.035 3126.000 ;
        RECT 3456.935 3106.000 3485.035 3124.000 ;
        RECT 3456.935 3104.000 3458.035 3106.000 ;
      LAYER met4 ;
        RECT 3458.035 3104.000 3483.000 3106.000 ;
      LAYER met4 ;
        RECT 3483.000 3104.000 3485.035 3106.000 ;
        RECT 3456.935 3086.000 3485.035 3104.000 ;
        RECT 3456.935 3084.000 3458.035 3086.000 ;
      LAYER met4 ;
        RECT 3458.035 3084.000 3483.000 3086.000 ;
      LAYER met4 ;
        RECT 3483.000 3084.000 3485.035 3086.000 ;
        RECT 3456.935 3066.000 3485.035 3084.000 ;
        RECT 3456.935 3064.000 3458.035 3066.000 ;
      LAYER met4 ;
        RECT 3458.035 3064.000 3483.000 3066.000 ;
      LAYER met4 ;
        RECT 3483.000 3064.000 3485.035 3066.000 ;
        RECT 3456.935 3046.000 3485.035 3064.000 ;
        RECT 3456.935 3045.000 3458.035 3046.000 ;
        RECT 3456.935 3043.330 3457.635 3044.035 ;
      LAYER met4 ;
        RECT 3458.035 3043.730 3483.000 3046.000 ;
      LAYER met4 ;
        RECT 3483.000 3045.000 3485.035 3046.000 ;
        RECT 3562.035 3045.000 3588.000 3190.000 ;
        RECT 3483.400 3043.330 3563.385 3044.035 ;
      LAYER met4 ;
        RECT 3563.785 3043.730 3588.000 3045.000 ;
      LAYER met4 ;
        RECT 3445.135 3041.990 3588.000 3043.330 ;
        RECT 3444.505 3008.160 3588.000 3041.990 ;
        RECT 3439.745 3006.640 3588.000 3008.160 ;
        RECT 3439.745 2992.455 3440.725 3006.640 ;
        RECT 3436.465 2990.935 3440.725 2992.455 ;
        RECT 3388.535 2772.310 3435.965 2815.990 ;
        RECT 3388.535 2740.670 3435.335 2772.310 ;
        RECT 3388.535 2740.030 3389.635 2740.670 ;
        RECT 198.365 2704.330 199.465 2704.970 ;
        RECT 152.665 2672.690 199.465 2704.330 ;
        RECT 152.035 2629.010 199.465 2672.690 ;
        RECT 147.275 2040.545 151.535 2042.065 ;
        RECT 147.275 2026.360 148.255 2040.545 ;
        RECT 0.000 2024.840 148.255 2026.360 ;
        RECT 0.000 1991.010 143.495 2024.840 ;
        RECT 0.000 1989.670 142.865 1991.010 ;
      LAYER met4 ;
        RECT 0.000 1988.000 24.215 1989.270 ;
      LAYER met4 ;
        RECT 24.615 1988.965 104.600 1989.670 ;
        RECT 0.000 1852.000 25.965 1988.000 ;
        RECT 102.965 1986.000 105.000 1988.000 ;
      LAYER met4 ;
        RECT 105.000 1986.000 129.965 1989.270 ;
      LAYER met4 ;
        RECT 130.365 1988.965 131.065 1989.670 ;
        RECT 129.965 1986.000 131.065 1988.000 ;
        RECT 102.965 1983.000 131.065 1986.000 ;
        RECT 102.965 1981.000 105.000 1983.000 ;
      LAYER met4 ;
        RECT 105.000 1981.000 129.965 1983.000 ;
      LAYER met4 ;
        RECT 129.965 1981.000 131.065 1983.000 ;
        RECT 102.965 1973.000 131.065 1981.000 ;
        RECT 102.965 1971.000 105.000 1973.000 ;
      LAYER met4 ;
        RECT 105.000 1971.000 129.965 1973.000 ;
      LAYER met4 ;
        RECT 129.965 1971.000 131.065 1973.000 ;
        RECT 102.965 1953.000 131.065 1971.000 ;
        RECT 102.965 1951.000 105.000 1953.000 ;
      LAYER met4 ;
        RECT 105.000 1951.000 129.965 1953.000 ;
      LAYER met4 ;
        RECT 129.965 1951.000 131.065 1953.000 ;
        RECT 102.965 1933.000 131.065 1951.000 ;
        RECT 102.965 1931.000 105.000 1933.000 ;
      LAYER met4 ;
        RECT 105.000 1931.000 129.965 1933.000 ;
      LAYER met4 ;
        RECT 129.965 1931.000 131.065 1933.000 ;
        RECT 102.965 1913.000 131.065 1931.000 ;
        RECT 102.965 1911.000 105.000 1913.000 ;
      LAYER met4 ;
        RECT 105.000 1911.000 129.965 1913.000 ;
      LAYER met4 ;
        RECT 129.965 1911.000 131.065 1913.000 ;
        RECT 102.965 1893.000 131.065 1911.000 ;
        RECT 102.965 1891.000 105.000 1893.000 ;
      LAYER met4 ;
        RECT 105.000 1891.000 129.965 1893.000 ;
      LAYER met4 ;
        RECT 129.965 1891.000 131.065 1893.000 ;
        RECT 102.965 1873.000 131.065 1891.000 ;
        RECT 102.965 1871.000 105.000 1873.000 ;
      LAYER met4 ;
        RECT 105.000 1871.000 129.965 1873.000 ;
      LAYER met4 ;
        RECT 129.965 1871.000 131.065 1873.000 ;
        RECT 102.965 1853.000 131.065 1871.000 ;
        RECT 102.965 1852.000 105.000 1853.000 ;
      LAYER met4 ;
        RECT 0.000 1850.730 24.215 1852.000 ;
      LAYER met4 ;
        RECT 24.615 1850.330 104.600 1850.970 ;
      LAYER met4 ;
        RECT 105.000 1850.730 129.965 1853.000 ;
      LAYER met4 ;
        RECT 129.965 1852.000 131.065 1853.000 ;
        RECT 130.365 1850.330 131.065 1850.970 ;
      LAYER met4 ;
        RECT 131.465 1850.730 135.915 1989.270 ;
      LAYER met4 ;
        RECT 136.315 1988.965 136.915 1989.670 ;
        RECT 136.315 1852.000 136.915 1987.000 ;
        RECT 136.315 1850.330 136.915 1850.970 ;
      LAYER met4 ;
        RECT 137.315 1850.730 141.765 1989.270 ;
      LAYER met4 ;
        RECT 142.165 1988.965 142.865 1989.670 ;
        RECT 142.165 1852.000 142.865 1988.000 ;
        RECT 142.165 1850.330 142.865 1850.970 ;
        RECT 0.000 1818.690 142.865 1850.330 ;
      LAYER met4 ;
        RECT 143.265 1819.090 143.595 1990.610 ;
      LAYER met4 ;
        RECT 0.000 1810.360 143.495 1818.690 ;
      LAYER met4 ;
        RECT 143.895 1810.760 146.875 2024.440 ;
      LAYER met4 ;
        RECT 147.275 1989.670 148.255 2024.840 ;
      LAYER met4 ;
        RECT 147.175 1988.000 148.355 1989.270 ;
      LAYER met4 ;
        RECT 147.275 1852.000 148.255 1988.000 ;
      LAYER met4 ;
        RECT 147.175 1850.730 148.355 1852.000 ;
      LAYER met4 ;
        RECT 147.275 1826.065 148.255 1850.330 ;
      LAYER met4 ;
        RECT 148.655 1826.465 151.635 2040.145 ;
        RECT 151.935 2035.090 152.265 2628.610 ;
      LAYER met4 ;
        RECT 152.665 2627.670 199.465 2629.010 ;
        RECT 152.665 2626.965 153.365 2627.670 ;
        RECT 152.665 2488.330 153.365 2489.035 ;
      LAYER met4 ;
        RECT 153.765 2488.730 158.415 2627.270 ;
      LAYER met4 ;
        RECT 158.815 2626.965 159.415 2627.670 ;
        RECT 158.815 2488.330 159.415 2489.035 ;
      LAYER met4 ;
        RECT 159.815 2488.730 163.265 2627.270 ;
      LAYER met4 ;
        RECT 163.665 2626.965 164.265 2627.670 ;
        RECT 163.665 2488.330 164.265 2489.035 ;
      LAYER met4 ;
        RECT 164.665 2488.730 168.115 2627.270 ;
      LAYER met4 ;
        RECT 168.515 2626.965 169.115 2627.670 ;
        RECT 168.515 2488.330 169.115 2489.035 ;
      LAYER met4 ;
        RECT 169.515 2488.730 174.165 2627.270 ;
      LAYER met4 ;
        RECT 174.565 2626.965 175.165 2627.670 ;
        RECT 180.615 2627.365 186.065 2627.670 ;
        RECT 174.565 2488.330 175.165 2489.035 ;
      LAYER met4 ;
        RECT 175.565 2488.730 180.215 2627.270 ;
      LAYER met4 ;
        RECT 180.615 2626.965 181.215 2627.365 ;
        RECT 185.465 2626.965 186.065 2627.365 ;
        RECT 180.615 2488.635 181.215 2489.035 ;
        RECT 185.465 2488.635 186.065 2489.035 ;
      LAYER met4 ;
        RECT 186.465 2488.730 191.115 2627.270 ;
      LAYER met4 ;
        RECT 191.515 2626.965 192.115 2627.670 ;
        RECT 180.615 2488.330 186.065 2488.635 ;
        RECT 191.515 2488.330 192.115 2489.035 ;
      LAYER met4 ;
        RECT 192.515 2488.730 197.965 2627.270 ;
      LAYER met4 ;
        RECT 198.365 2626.965 199.465 2627.670 ;
      LAYER met4 ;
        RECT 3390.035 2592.730 3395.485 2740.270 ;
      LAYER met4 ;
        RECT 3395.885 2740.030 3396.485 2740.670 ;
        RECT 3401.935 2740.430 3407.385 2740.670 ;
        RECT 3395.885 2592.330 3396.485 2593.035 ;
      LAYER met4 ;
        RECT 3396.885 2592.730 3401.535 2740.270 ;
      LAYER met4 ;
        RECT 3401.935 2740.030 3402.535 2740.430 ;
        RECT 3406.785 2740.030 3407.385 2740.430 ;
      LAYER met4 ;
        RECT 3402.935 2593.035 3406.385 2740.030 ;
      LAYER met4 ;
        RECT 3401.935 2592.635 3402.535 2593.035 ;
        RECT 3406.785 2592.635 3407.385 2593.035 ;
      LAYER met4 ;
        RECT 3407.785 2592.730 3412.435 2740.270 ;
      LAYER met4 ;
        RECT 3412.835 2740.030 3413.435 2740.670 ;
        RECT 3401.935 2592.330 3407.385 2592.635 ;
        RECT 3412.835 2592.330 3413.435 2593.035 ;
      LAYER met4 ;
        RECT 3413.835 2592.730 3418.485 2740.270 ;
      LAYER met4 ;
        RECT 3418.885 2740.030 3419.485 2740.670 ;
        RECT 3418.885 2592.330 3419.485 2593.035 ;
      LAYER met4 ;
        RECT 3419.885 2592.730 3423.335 2740.270 ;
      LAYER met4 ;
        RECT 3423.735 2740.030 3424.335 2740.670 ;
        RECT 3423.735 2592.330 3424.335 2593.035 ;
      LAYER met4 ;
        RECT 3424.735 2592.730 3428.185 2740.270 ;
      LAYER met4 ;
        RECT 3428.585 2740.030 3429.185 2740.670 ;
        RECT 3428.585 2592.330 3429.185 2593.035 ;
      LAYER met4 ;
        RECT 3429.585 2592.730 3434.235 2740.270 ;
      LAYER met4 ;
        RECT 3434.635 2740.030 3435.335 2740.670 ;
        RECT 3434.635 2592.330 3435.335 2593.035 ;
        RECT 3390.035 2520.670 3435.335 2592.330 ;
        RECT 152.665 2416.670 197.965 2488.330 ;
        RECT 152.665 2415.965 153.365 2416.670 ;
        RECT 158.815 2415.965 159.415 2416.670 ;
        RECT 152.665 2277.330 153.365 2279.000 ;
        RECT 158.815 2277.330 159.415 2279.000 ;
      LAYER met4 ;
        RECT 159.815 2277.730 163.265 2416.270 ;
      LAYER met4 ;
        RECT 163.665 2415.965 164.265 2416.670 ;
        RECT 163.665 2277.330 164.265 2279.000 ;
      LAYER met4 ;
        RECT 164.665 2277.730 168.115 2416.270 ;
      LAYER met4 ;
        RECT 168.515 2415.965 169.115 2416.670 ;
        RECT 168.515 2277.330 169.115 2279.000 ;
      LAYER met4 ;
        RECT 169.515 2277.730 174.165 2416.270 ;
      LAYER met4 ;
        RECT 174.565 2415.965 175.165 2416.670 ;
        RECT 180.615 2416.365 186.065 2416.670 ;
        RECT 174.565 2277.330 175.165 2279.000 ;
      LAYER met4 ;
        RECT 175.565 2277.730 180.215 2416.270 ;
      LAYER met4 ;
        RECT 180.615 2415.965 181.215 2416.365 ;
        RECT 185.465 2415.965 186.065 2416.365 ;
        RECT 180.615 2277.635 181.215 2279.000 ;
        RECT 185.465 2277.635 186.065 2279.000 ;
      LAYER met4 ;
        RECT 186.465 2277.730 191.115 2416.270 ;
      LAYER met4 ;
        RECT 191.515 2415.965 192.115 2416.670 ;
        RECT 180.615 2277.330 186.065 2277.635 ;
        RECT 191.515 2277.330 192.115 2279.000 ;
      LAYER met4 ;
        RECT 192.515 2277.730 197.965 2416.270 ;
        RECT 3390.035 2372.730 3395.485 2520.270 ;
      LAYER met4 ;
        RECT 3395.885 2519.965 3396.485 2520.670 ;
        RECT 3401.935 2520.365 3407.385 2520.670 ;
        RECT 3395.885 2372.330 3396.485 2373.035 ;
      LAYER met4 ;
        RECT 3396.885 2372.730 3401.535 2520.270 ;
      LAYER met4 ;
        RECT 3401.935 2519.965 3402.535 2520.365 ;
        RECT 3406.785 2519.965 3407.385 2520.365 ;
      LAYER met4 ;
        RECT 3402.935 2373.035 3406.385 2519.965 ;
      LAYER met4 ;
        RECT 3401.935 2372.635 3402.535 2373.035 ;
        RECT 3406.785 2372.635 3407.385 2373.035 ;
      LAYER met4 ;
        RECT 3407.785 2372.730 3412.435 2520.270 ;
      LAYER met4 ;
        RECT 3412.835 2519.965 3413.435 2520.670 ;
        RECT 3401.935 2372.330 3407.385 2372.635 ;
        RECT 3412.835 2372.330 3413.435 2373.035 ;
      LAYER met4 ;
        RECT 3413.835 2372.730 3418.485 2520.270 ;
      LAYER met4 ;
        RECT 3418.885 2519.965 3419.485 2520.670 ;
        RECT 3418.885 2372.330 3419.485 2373.035 ;
      LAYER met4 ;
        RECT 3419.885 2372.730 3423.335 2520.270 ;
      LAYER met4 ;
        RECT 3423.735 2519.965 3424.335 2520.670 ;
        RECT 3423.735 2372.330 3424.335 2373.035 ;
      LAYER met4 ;
        RECT 3424.735 2372.730 3428.185 2520.270 ;
      LAYER met4 ;
        RECT 3428.585 2519.965 3429.185 2520.670 ;
        RECT 3434.635 2519.965 3435.335 2520.670 ;
        RECT 3428.585 2372.330 3429.185 2373.035 ;
        RECT 3434.635 2372.330 3435.335 2373.035 ;
        RECT 3390.035 2300.670 3435.335 2372.330 ;
        RECT 152.665 2205.670 197.965 2277.330 ;
        RECT 152.665 2204.965 153.365 2205.670 ;
        RECT 158.815 2204.965 159.415 2205.670 ;
        RECT 152.665 2066.330 153.365 2066.970 ;
        RECT 158.815 2066.330 159.415 2066.970 ;
      LAYER met4 ;
        RECT 159.815 2066.730 163.265 2205.270 ;
      LAYER met4 ;
        RECT 163.665 2204.965 164.265 2205.670 ;
        RECT 163.665 2066.330 164.265 2066.970 ;
      LAYER met4 ;
        RECT 164.665 2066.730 168.115 2205.270 ;
      LAYER met4 ;
        RECT 168.515 2204.965 169.115 2205.670 ;
        RECT 168.515 2066.330 169.115 2066.970 ;
      LAYER met4 ;
        RECT 169.515 2066.730 174.165 2205.270 ;
      LAYER met4 ;
        RECT 174.565 2204.965 175.165 2205.670 ;
        RECT 180.615 2205.365 186.065 2205.670 ;
        RECT 174.565 2066.330 175.165 2066.970 ;
      LAYER met4 ;
        RECT 175.565 2066.730 180.215 2205.270 ;
      LAYER met4 ;
        RECT 180.615 2204.965 181.215 2205.365 ;
        RECT 185.465 2204.965 186.065 2205.365 ;
      LAYER met4 ;
        RECT 181.615 2066.970 185.065 2204.965 ;
      LAYER met4 ;
        RECT 180.615 2066.570 181.215 2066.970 ;
        RECT 185.465 2066.570 186.065 2066.970 ;
      LAYER met4 ;
        RECT 186.465 2066.730 191.115 2205.270 ;
      LAYER met4 ;
        RECT 191.515 2204.965 192.115 2205.670 ;
        RECT 180.615 2066.330 186.065 2066.570 ;
        RECT 191.515 2066.330 192.115 2066.970 ;
      LAYER met4 ;
        RECT 192.515 2066.730 197.965 2205.270 ;
        RECT 3390.035 2151.730 3395.485 2300.270 ;
      LAYER met4 ;
        RECT 3395.885 2299.000 3396.485 2300.670 ;
        RECT 3401.935 2300.365 3407.385 2300.670 ;
        RECT 3395.885 2151.330 3396.485 2152.035 ;
      LAYER met4 ;
        RECT 3396.885 2151.730 3401.535 2300.270 ;
      LAYER met4 ;
        RECT 3401.935 2299.000 3402.535 2300.365 ;
      LAYER met4 ;
        RECT 3402.935 2152.035 3406.385 2299.965 ;
      LAYER met4 ;
        RECT 3406.785 2299.000 3407.385 2300.365 ;
        RECT 3401.935 2151.635 3402.535 2152.035 ;
        RECT 3406.785 2151.635 3407.385 2152.035 ;
      LAYER met4 ;
        RECT 3407.785 2151.730 3412.435 2300.270 ;
      LAYER met4 ;
        RECT 3412.835 2299.000 3413.435 2300.670 ;
        RECT 3401.935 2151.330 3407.385 2151.635 ;
        RECT 3412.835 2151.330 3413.435 2152.035 ;
      LAYER met4 ;
        RECT 3413.835 2151.730 3418.485 2300.270 ;
      LAYER met4 ;
        RECT 3418.885 2299.000 3419.485 2300.670 ;
        RECT 3418.885 2151.330 3419.485 2152.035 ;
      LAYER met4 ;
        RECT 3419.885 2151.730 3423.335 2300.270 ;
      LAYER met4 ;
        RECT 3423.735 2299.000 3424.335 2300.670 ;
        RECT 3423.735 2151.330 3424.335 2152.035 ;
      LAYER met4 ;
        RECT 3424.735 2151.730 3428.185 2300.270 ;
      LAYER met4 ;
        RECT 3428.585 2299.000 3429.185 2300.670 ;
        RECT 3434.635 2299.000 3435.335 2300.670 ;
        RECT 3428.585 2151.330 3429.185 2152.035 ;
        RECT 3434.635 2151.330 3435.335 2152.035 ;
      LAYER met4 ;
        RECT 3435.735 2151.730 3436.065 2771.910 ;
        RECT 3436.365 2766.855 3439.345 2990.535 ;
      LAYER met4 ;
        RECT 3439.745 2966.670 3440.725 2990.935 ;
      LAYER met4 ;
        RECT 3439.645 2965.000 3440.825 2966.270 ;
      LAYER met4 ;
        RECT 3439.745 2819.000 3440.725 2965.000 ;
      LAYER met4 ;
        RECT 3439.645 2817.730 3440.825 2819.000 ;
      LAYER met4 ;
        RECT 3439.745 2782.160 3440.725 2817.330 ;
      LAYER met4 ;
        RECT 3441.125 2782.560 3444.105 3006.240 ;
      LAYER met4 ;
        RECT 3444.505 2998.310 3588.000 3006.640 ;
      LAYER met4 ;
        RECT 3444.405 2816.390 3444.735 2997.910 ;
      LAYER met4 ;
        RECT 3445.135 2966.670 3588.000 2998.310 ;
        RECT 3445.135 2966.030 3445.835 2966.670 ;
        RECT 3445.135 2819.000 3445.835 2965.000 ;
        RECT 3445.135 2817.330 3445.835 2818.035 ;
      LAYER met4 ;
        RECT 3446.235 2817.730 3450.685 2966.270 ;
      LAYER met4 ;
        RECT 3451.085 2966.030 3451.685 2966.670 ;
        RECT 3451.085 2819.000 3451.685 2964.000 ;
        RECT 3451.085 2817.330 3451.685 2818.035 ;
      LAYER met4 ;
        RECT 3452.085 2817.730 3456.535 2966.270 ;
      LAYER met4 ;
        RECT 3456.935 2966.030 3457.635 2966.670 ;
        RECT 3456.935 2963.000 3458.035 2965.000 ;
      LAYER met4 ;
        RECT 3458.035 2963.000 3483.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2966.030 3563.385 2966.670 ;
      LAYER met4 ;
        RECT 3563.785 2965.000 3588.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.000 2963.000 3485.035 2965.000 ;
        RECT 3456.935 2960.000 3485.035 2963.000 ;
        RECT 3456.935 2958.000 3458.035 2960.000 ;
      LAYER met4 ;
        RECT 3458.035 2958.000 3483.000 2960.000 ;
      LAYER met4 ;
        RECT 3483.000 2958.000 3485.035 2960.000 ;
        RECT 3456.935 2940.000 3485.035 2958.000 ;
        RECT 3456.935 2938.000 3458.035 2940.000 ;
      LAYER met4 ;
        RECT 3458.035 2938.000 3483.000 2940.000 ;
      LAYER met4 ;
        RECT 3483.000 2938.000 3485.035 2940.000 ;
        RECT 3456.935 2920.000 3485.035 2938.000 ;
        RECT 3456.935 2918.000 3458.035 2920.000 ;
      LAYER met4 ;
        RECT 3458.035 2918.000 3483.000 2920.000 ;
      LAYER met4 ;
        RECT 3483.000 2918.000 3485.035 2920.000 ;
        RECT 3456.935 2900.000 3485.035 2918.000 ;
        RECT 3456.935 2898.000 3458.035 2900.000 ;
      LAYER met4 ;
        RECT 3458.035 2898.000 3483.000 2900.000 ;
      LAYER met4 ;
        RECT 3483.000 2898.000 3485.035 2900.000 ;
        RECT 3456.935 2880.000 3485.035 2898.000 ;
        RECT 3456.935 2878.000 3458.035 2880.000 ;
      LAYER met4 ;
        RECT 3458.035 2878.000 3483.000 2880.000 ;
      LAYER met4 ;
        RECT 3483.000 2878.000 3485.035 2880.000 ;
        RECT 3456.935 2860.000 3485.035 2878.000 ;
        RECT 3456.935 2858.000 3458.035 2860.000 ;
      LAYER met4 ;
        RECT 3458.035 2858.000 3483.000 2860.000 ;
      LAYER met4 ;
        RECT 3483.000 2858.000 3485.035 2860.000 ;
        RECT 3456.935 2840.000 3485.035 2858.000 ;
        RECT 3456.935 2838.000 3458.035 2840.000 ;
      LAYER met4 ;
        RECT 3458.035 2838.000 3483.000 2840.000 ;
      LAYER met4 ;
        RECT 3483.000 2838.000 3485.035 2840.000 ;
        RECT 3456.935 2820.000 3485.035 2838.000 ;
        RECT 3456.935 2819.000 3458.035 2820.000 ;
        RECT 3456.935 2817.330 3457.635 2818.035 ;
      LAYER met4 ;
        RECT 3458.035 2817.730 3483.000 2820.000 ;
      LAYER met4 ;
        RECT 3483.000 2819.000 3485.035 2820.000 ;
        RECT 3562.035 2819.000 3588.000 2965.000 ;
        RECT 3483.400 2817.330 3563.385 2818.035 ;
      LAYER met4 ;
        RECT 3563.785 2817.730 3588.000 2819.000 ;
      LAYER met4 ;
        RECT 3445.135 2815.990 3588.000 2817.330 ;
        RECT 3444.505 2782.160 3588.000 2815.990 ;
        RECT 3439.745 2780.640 3588.000 2782.160 ;
        RECT 3439.745 2766.455 3440.725 2780.640 ;
        RECT 3436.465 2764.935 3440.725 2766.455 ;
        RECT 3390.035 2079.670 3435.965 2151.330 ;
        RECT 198.365 2066.330 199.465 2066.970 ;
        RECT 152.665 2034.690 199.465 2066.330 ;
        RECT 152.035 1991.010 199.465 2034.690 ;
        RECT 147.275 1824.545 151.535 1826.065 ;
        RECT 147.275 1810.360 148.255 1824.545 ;
        RECT 0.000 1808.840 148.255 1810.360 ;
        RECT 0.000 1775.010 143.495 1808.840 ;
        RECT 0.000 1773.670 142.865 1775.010 ;
      LAYER met4 ;
        RECT 0.000 1772.000 24.215 1773.270 ;
      LAYER met4 ;
        RECT 24.615 1772.965 104.600 1773.670 ;
        RECT 0.000 1636.000 25.965 1772.000 ;
        RECT 102.965 1770.000 105.000 1772.000 ;
      LAYER met4 ;
        RECT 105.000 1770.000 129.965 1773.270 ;
      LAYER met4 ;
        RECT 130.365 1772.965 131.065 1773.670 ;
        RECT 129.965 1770.000 131.065 1772.000 ;
        RECT 102.965 1767.000 131.065 1770.000 ;
        RECT 102.965 1765.000 105.000 1767.000 ;
      LAYER met4 ;
        RECT 105.000 1765.000 129.965 1767.000 ;
      LAYER met4 ;
        RECT 129.965 1765.000 131.065 1767.000 ;
        RECT 102.965 1757.000 131.065 1765.000 ;
        RECT 102.965 1755.000 105.000 1757.000 ;
      LAYER met4 ;
        RECT 105.000 1755.000 129.965 1757.000 ;
      LAYER met4 ;
        RECT 129.965 1755.000 131.065 1757.000 ;
        RECT 102.965 1737.000 131.065 1755.000 ;
        RECT 102.965 1735.000 105.000 1737.000 ;
      LAYER met4 ;
        RECT 105.000 1735.000 129.965 1737.000 ;
      LAYER met4 ;
        RECT 129.965 1735.000 131.065 1737.000 ;
        RECT 102.965 1717.000 131.065 1735.000 ;
        RECT 102.965 1715.000 105.000 1717.000 ;
      LAYER met4 ;
        RECT 105.000 1715.000 129.965 1717.000 ;
      LAYER met4 ;
        RECT 129.965 1715.000 131.065 1717.000 ;
        RECT 102.965 1697.000 131.065 1715.000 ;
        RECT 102.965 1695.000 105.000 1697.000 ;
      LAYER met4 ;
        RECT 105.000 1695.000 129.965 1697.000 ;
      LAYER met4 ;
        RECT 129.965 1695.000 131.065 1697.000 ;
        RECT 102.965 1677.000 131.065 1695.000 ;
        RECT 102.965 1675.000 105.000 1677.000 ;
      LAYER met4 ;
        RECT 105.000 1675.000 129.965 1677.000 ;
      LAYER met4 ;
        RECT 129.965 1675.000 131.065 1677.000 ;
        RECT 102.965 1657.000 131.065 1675.000 ;
        RECT 102.965 1655.000 105.000 1657.000 ;
      LAYER met4 ;
        RECT 105.000 1655.000 129.965 1657.000 ;
      LAYER met4 ;
        RECT 129.965 1655.000 131.065 1657.000 ;
        RECT 102.965 1637.000 131.065 1655.000 ;
        RECT 102.965 1636.000 105.000 1637.000 ;
      LAYER met4 ;
        RECT 0.000 1634.730 24.215 1636.000 ;
      LAYER met4 ;
        RECT 24.615 1634.330 104.600 1634.970 ;
      LAYER met4 ;
        RECT 105.000 1634.730 129.965 1637.000 ;
      LAYER met4 ;
        RECT 129.965 1636.000 131.065 1637.000 ;
        RECT 130.365 1634.330 131.065 1634.970 ;
      LAYER met4 ;
        RECT 131.465 1634.730 135.915 1773.270 ;
      LAYER met4 ;
        RECT 136.315 1772.965 136.915 1773.670 ;
        RECT 136.315 1636.000 136.915 1771.000 ;
        RECT 136.315 1634.330 136.915 1634.970 ;
      LAYER met4 ;
        RECT 137.315 1634.730 141.765 1773.270 ;
      LAYER met4 ;
        RECT 142.165 1772.965 142.865 1773.670 ;
        RECT 142.165 1636.000 142.865 1772.000 ;
        RECT 142.165 1634.330 142.865 1634.970 ;
        RECT 0.000 1602.690 142.865 1634.330 ;
      LAYER met4 ;
        RECT 143.265 1603.090 143.595 1774.610 ;
      LAYER met4 ;
        RECT 0.000 1594.360 143.495 1602.690 ;
      LAYER met4 ;
        RECT 143.895 1594.760 146.875 1808.440 ;
      LAYER met4 ;
        RECT 147.275 1773.670 148.255 1808.840 ;
      LAYER met4 ;
        RECT 147.175 1772.000 148.355 1773.270 ;
      LAYER met4 ;
        RECT 147.275 1636.000 148.255 1772.000 ;
      LAYER met4 ;
        RECT 147.175 1634.730 148.355 1636.000 ;
      LAYER met4 ;
        RECT 147.275 1610.065 148.255 1634.330 ;
      LAYER met4 ;
        RECT 148.655 1610.465 151.635 1824.145 ;
        RECT 151.935 1819.090 152.265 1990.610 ;
      LAYER met4 ;
        RECT 152.665 1989.670 199.465 1991.010 ;
        RECT 152.665 1988.965 153.365 1989.670 ;
        RECT 152.665 1850.330 153.365 1850.970 ;
      LAYER met4 ;
        RECT 153.765 1850.730 158.415 1989.270 ;
      LAYER met4 ;
        RECT 158.815 1988.965 159.415 1989.670 ;
        RECT 158.815 1850.330 159.415 1850.970 ;
      LAYER met4 ;
        RECT 159.815 1850.730 163.265 1989.270 ;
      LAYER met4 ;
        RECT 163.665 1988.965 164.265 1989.670 ;
        RECT 163.665 1850.330 164.265 1850.970 ;
      LAYER met4 ;
        RECT 164.665 1850.730 168.115 1989.270 ;
      LAYER met4 ;
        RECT 168.515 1988.965 169.115 1989.670 ;
        RECT 168.515 1850.330 169.115 1850.970 ;
      LAYER met4 ;
        RECT 169.515 1850.730 174.165 1989.270 ;
      LAYER met4 ;
        RECT 174.565 1988.965 175.165 1989.670 ;
        RECT 180.615 1989.365 186.065 1989.670 ;
        RECT 174.565 1850.330 175.165 1850.970 ;
      LAYER met4 ;
        RECT 175.565 1850.730 180.215 1989.270 ;
      LAYER met4 ;
        RECT 180.615 1988.965 181.215 1989.365 ;
        RECT 185.465 1988.965 186.065 1989.365 ;
      LAYER met4 ;
        RECT 181.615 1850.970 185.065 1988.965 ;
      LAYER met4 ;
        RECT 180.615 1850.570 181.215 1850.970 ;
        RECT 185.465 1850.570 186.065 1850.970 ;
      LAYER met4 ;
        RECT 186.465 1850.730 191.115 1989.270 ;
      LAYER met4 ;
        RECT 191.515 1988.965 192.115 1989.670 ;
        RECT 180.615 1850.330 186.065 1850.570 ;
        RECT 191.515 1850.330 192.115 1850.970 ;
      LAYER met4 ;
        RECT 192.515 1850.730 197.965 1989.270 ;
      LAYER met4 ;
        RECT 198.365 1988.965 199.465 1989.670 ;
        RECT 3388.535 1931.330 3389.635 1932.035 ;
      LAYER met4 ;
        RECT 3390.035 1931.730 3395.485 2079.270 ;
      LAYER met4 ;
        RECT 3395.885 2078.965 3396.485 2079.670 ;
        RECT 3401.935 2079.365 3407.385 2079.670 ;
        RECT 3395.885 1931.330 3396.485 1932.035 ;
      LAYER met4 ;
        RECT 3396.885 1931.730 3401.535 2079.270 ;
      LAYER met4 ;
        RECT 3401.935 2078.965 3402.535 2079.365 ;
        RECT 3406.785 2078.965 3407.385 2079.365 ;
      LAYER met4 ;
        RECT 3402.935 1932.035 3406.385 2078.965 ;
      LAYER met4 ;
        RECT 3401.935 1931.635 3402.535 1932.035 ;
        RECT 3406.785 1931.635 3407.385 1932.035 ;
      LAYER met4 ;
        RECT 3407.785 1931.730 3412.435 2079.270 ;
      LAYER met4 ;
        RECT 3412.835 2078.965 3413.435 2079.670 ;
        RECT 3401.935 1931.330 3407.385 1931.635 ;
        RECT 3412.835 1931.330 3413.435 1932.035 ;
      LAYER met4 ;
        RECT 3413.835 1931.730 3418.485 2079.270 ;
      LAYER met4 ;
        RECT 3418.885 2078.965 3419.485 2079.670 ;
        RECT 3418.885 1931.330 3419.485 1932.035 ;
      LAYER met4 ;
        RECT 3419.885 1931.730 3423.335 2079.270 ;
      LAYER met4 ;
        RECT 3423.735 2078.965 3424.335 2079.670 ;
        RECT 3423.735 1931.330 3424.335 1932.035 ;
      LAYER met4 ;
        RECT 3424.735 1931.730 3428.185 2079.270 ;
      LAYER met4 ;
        RECT 3428.585 2078.965 3429.185 2079.670 ;
        RECT 3428.585 1931.330 3429.185 1932.035 ;
      LAYER met4 ;
        RECT 3429.585 1931.730 3434.235 2079.270 ;
      LAYER met4 ;
        RECT 3434.635 2078.965 3435.335 2079.670 ;
        RECT 3434.635 1931.330 3435.335 1932.035 ;
        RECT 3388.535 1929.990 3435.335 1931.330 ;
      LAYER met4 ;
        RECT 3435.735 1930.390 3436.065 2079.270 ;
      LAYER met4 ;
        RECT 3388.535 1886.310 3435.965 1929.990 ;
        RECT 3388.535 1854.670 3435.335 1886.310 ;
        RECT 3388.535 1854.030 3389.635 1854.670 ;
        RECT 198.365 1850.330 199.465 1850.970 ;
        RECT 152.665 1818.690 199.465 1850.330 ;
        RECT 152.035 1775.010 199.465 1818.690 ;
        RECT 147.275 1608.545 151.535 1610.065 ;
        RECT 147.275 1594.360 148.255 1608.545 ;
        RECT 0.000 1592.840 148.255 1594.360 ;
        RECT 0.000 1559.010 143.495 1592.840 ;
        RECT 0.000 1557.670 142.865 1559.010 ;
      LAYER met4 ;
        RECT 0.000 1556.000 24.215 1557.270 ;
      LAYER met4 ;
        RECT 24.615 1556.965 104.600 1557.670 ;
        RECT 0.000 1420.000 25.965 1556.000 ;
        RECT 102.965 1554.000 105.000 1556.000 ;
      LAYER met4 ;
        RECT 105.000 1554.000 129.965 1557.270 ;
      LAYER met4 ;
        RECT 130.365 1556.965 131.065 1557.670 ;
        RECT 129.965 1554.000 131.065 1556.000 ;
        RECT 102.965 1551.000 131.065 1554.000 ;
        RECT 102.965 1549.000 105.000 1551.000 ;
      LAYER met4 ;
        RECT 105.000 1549.000 129.965 1551.000 ;
      LAYER met4 ;
        RECT 129.965 1549.000 131.065 1551.000 ;
        RECT 102.965 1541.000 131.065 1549.000 ;
        RECT 102.965 1539.000 105.000 1541.000 ;
      LAYER met4 ;
        RECT 105.000 1539.000 129.965 1541.000 ;
      LAYER met4 ;
        RECT 129.965 1539.000 131.065 1541.000 ;
        RECT 102.965 1521.000 131.065 1539.000 ;
        RECT 102.965 1519.000 105.000 1521.000 ;
      LAYER met4 ;
        RECT 105.000 1519.000 129.965 1521.000 ;
      LAYER met4 ;
        RECT 129.965 1519.000 131.065 1521.000 ;
        RECT 102.965 1501.000 131.065 1519.000 ;
        RECT 102.965 1499.000 105.000 1501.000 ;
      LAYER met4 ;
        RECT 105.000 1499.000 129.965 1501.000 ;
      LAYER met4 ;
        RECT 129.965 1499.000 131.065 1501.000 ;
        RECT 102.965 1481.000 131.065 1499.000 ;
        RECT 102.965 1479.000 105.000 1481.000 ;
      LAYER met4 ;
        RECT 105.000 1479.000 129.965 1481.000 ;
      LAYER met4 ;
        RECT 129.965 1479.000 131.065 1481.000 ;
        RECT 102.965 1461.000 131.065 1479.000 ;
        RECT 102.965 1459.000 105.000 1461.000 ;
      LAYER met4 ;
        RECT 105.000 1459.000 129.965 1461.000 ;
      LAYER met4 ;
        RECT 129.965 1459.000 131.065 1461.000 ;
        RECT 102.965 1441.000 131.065 1459.000 ;
        RECT 102.965 1439.000 105.000 1441.000 ;
      LAYER met4 ;
        RECT 105.000 1439.000 129.965 1441.000 ;
      LAYER met4 ;
        RECT 129.965 1439.000 131.065 1441.000 ;
        RECT 102.965 1421.000 131.065 1439.000 ;
        RECT 102.965 1420.000 105.000 1421.000 ;
      LAYER met4 ;
        RECT 0.000 1418.730 24.215 1420.000 ;
      LAYER met4 ;
        RECT 24.615 1418.330 104.600 1418.970 ;
      LAYER met4 ;
        RECT 105.000 1418.730 129.965 1421.000 ;
      LAYER met4 ;
        RECT 129.965 1420.000 131.065 1421.000 ;
        RECT 130.365 1418.330 131.065 1418.970 ;
      LAYER met4 ;
        RECT 131.465 1418.730 135.915 1557.270 ;
      LAYER met4 ;
        RECT 136.315 1556.965 136.915 1557.670 ;
        RECT 136.315 1420.000 136.915 1555.000 ;
        RECT 136.315 1418.330 136.915 1418.970 ;
      LAYER met4 ;
        RECT 137.315 1418.730 141.765 1557.270 ;
      LAYER met4 ;
        RECT 142.165 1556.965 142.865 1557.670 ;
        RECT 142.165 1420.000 142.865 1556.000 ;
        RECT 142.165 1418.330 142.865 1418.970 ;
        RECT 0.000 1386.690 142.865 1418.330 ;
      LAYER met4 ;
        RECT 143.265 1387.090 143.595 1558.610 ;
      LAYER met4 ;
        RECT 0.000 1378.360 143.495 1386.690 ;
      LAYER met4 ;
        RECT 143.895 1378.760 146.875 1592.440 ;
      LAYER met4 ;
        RECT 147.275 1557.670 148.255 1592.840 ;
      LAYER met4 ;
        RECT 147.175 1556.000 148.355 1557.270 ;
      LAYER met4 ;
        RECT 147.275 1420.000 148.255 1556.000 ;
      LAYER met4 ;
        RECT 147.175 1418.730 148.355 1420.000 ;
      LAYER met4 ;
        RECT 147.275 1394.065 148.255 1418.330 ;
      LAYER met4 ;
        RECT 148.655 1394.465 151.635 1608.145 ;
        RECT 151.935 1603.090 152.265 1774.610 ;
      LAYER met4 ;
        RECT 152.665 1773.670 199.465 1775.010 ;
        RECT 152.665 1772.965 153.365 1773.670 ;
        RECT 152.665 1634.330 153.365 1634.970 ;
      LAYER met4 ;
        RECT 153.765 1634.730 158.415 1773.270 ;
      LAYER met4 ;
        RECT 158.815 1772.965 159.415 1773.670 ;
        RECT 158.815 1634.330 159.415 1634.970 ;
      LAYER met4 ;
        RECT 159.815 1634.730 163.265 1773.270 ;
      LAYER met4 ;
        RECT 163.665 1772.965 164.265 1773.670 ;
        RECT 163.665 1634.330 164.265 1634.970 ;
      LAYER met4 ;
        RECT 164.665 1634.730 168.115 1773.270 ;
      LAYER met4 ;
        RECT 168.515 1772.965 169.115 1773.670 ;
        RECT 168.515 1634.330 169.115 1634.970 ;
      LAYER met4 ;
        RECT 169.515 1634.730 174.165 1773.270 ;
      LAYER met4 ;
        RECT 174.565 1772.965 175.165 1773.670 ;
        RECT 180.615 1773.365 186.065 1773.670 ;
        RECT 174.565 1634.330 175.165 1634.970 ;
      LAYER met4 ;
        RECT 175.565 1634.730 180.215 1773.270 ;
      LAYER met4 ;
        RECT 180.615 1772.965 181.215 1773.365 ;
        RECT 185.465 1772.965 186.065 1773.365 ;
      LAYER met4 ;
        RECT 181.615 1634.970 185.065 1772.965 ;
      LAYER met4 ;
        RECT 180.615 1634.570 181.215 1634.970 ;
        RECT 185.465 1634.570 186.065 1634.970 ;
      LAYER met4 ;
        RECT 186.465 1634.730 191.115 1773.270 ;
      LAYER met4 ;
        RECT 191.515 1772.965 192.115 1773.670 ;
        RECT 180.615 1634.330 186.065 1634.570 ;
        RECT 191.515 1634.330 192.115 1634.970 ;
      LAYER met4 ;
        RECT 192.515 1634.730 197.965 1773.270 ;
      LAYER met4 ;
        RECT 198.365 1772.965 199.465 1773.670 ;
        RECT 3388.535 1705.330 3389.635 1706.035 ;
      LAYER met4 ;
        RECT 3390.035 1705.730 3395.485 1854.270 ;
      LAYER met4 ;
        RECT 3395.885 1854.030 3396.485 1854.670 ;
        RECT 3401.935 1854.430 3407.385 1854.670 ;
        RECT 3395.885 1705.330 3396.485 1706.035 ;
      LAYER met4 ;
        RECT 3396.885 1705.730 3401.535 1854.270 ;
      LAYER met4 ;
        RECT 3401.935 1854.030 3402.535 1854.430 ;
        RECT 3406.785 1854.030 3407.385 1854.430 ;
      LAYER met4 ;
        RECT 3402.935 1706.035 3406.385 1854.030 ;
      LAYER met4 ;
        RECT 3401.935 1705.635 3402.535 1706.035 ;
        RECT 3406.785 1705.635 3407.385 1706.035 ;
      LAYER met4 ;
        RECT 3407.785 1705.730 3412.435 1854.270 ;
      LAYER met4 ;
        RECT 3412.835 1854.030 3413.435 1854.670 ;
        RECT 3401.935 1705.330 3407.385 1705.635 ;
        RECT 3412.835 1705.330 3413.435 1706.035 ;
      LAYER met4 ;
        RECT 3413.835 1705.730 3418.485 1854.270 ;
      LAYER met4 ;
        RECT 3418.885 1854.030 3419.485 1854.670 ;
        RECT 3418.885 1705.330 3419.485 1706.035 ;
      LAYER met4 ;
        RECT 3419.885 1705.730 3423.335 1854.270 ;
      LAYER met4 ;
        RECT 3423.735 1854.030 3424.335 1854.670 ;
        RECT 3423.735 1705.330 3424.335 1706.035 ;
      LAYER met4 ;
        RECT 3424.735 1705.730 3428.185 1854.270 ;
      LAYER met4 ;
        RECT 3428.585 1854.030 3429.185 1854.670 ;
        RECT 3428.585 1705.330 3429.185 1706.035 ;
      LAYER met4 ;
        RECT 3429.585 1705.730 3434.235 1854.270 ;
      LAYER met4 ;
        RECT 3434.635 1854.030 3435.335 1854.670 ;
        RECT 3434.635 1705.330 3435.335 1706.035 ;
        RECT 3388.535 1703.990 3435.335 1705.330 ;
      LAYER met4 ;
        RECT 3435.735 1704.390 3436.065 1885.910 ;
        RECT 3436.365 1880.855 3439.345 2764.535 ;
      LAYER met4 ;
        RECT 3439.745 2740.670 3440.725 2764.935 ;
      LAYER met4 ;
        RECT 3439.645 2739.000 3440.825 2740.270 ;
      LAYER met4 ;
        RECT 3439.745 2594.000 3440.725 2739.000 ;
      LAYER met4 ;
        RECT 3439.645 2592.730 3440.825 2594.000 ;
      LAYER met4 ;
        RECT 3439.745 2520.670 3440.725 2592.330 ;
      LAYER met4 ;
        RECT 3439.645 2519.000 3440.825 2520.270 ;
      LAYER met4 ;
        RECT 3439.745 2374.000 3440.725 2519.000 ;
      LAYER met4 ;
        RECT 3439.645 2372.730 3440.825 2374.000 ;
      LAYER met4 ;
        RECT 3439.745 2300.670 3440.725 2372.330 ;
      LAYER met4 ;
        RECT 3439.645 2299.000 3440.825 2300.270 ;
      LAYER met4 ;
        RECT 3439.745 2153.000 3440.725 2299.000 ;
      LAYER met4 ;
        RECT 3439.645 2151.730 3440.825 2153.000 ;
      LAYER met4 ;
        RECT 3439.745 2079.670 3440.725 2151.330 ;
      LAYER met4 ;
        RECT 3439.645 2078.000 3440.825 2079.270 ;
      LAYER met4 ;
        RECT 3439.745 1933.000 3440.725 2078.000 ;
      LAYER met4 ;
        RECT 3439.645 1931.730 3440.825 1933.000 ;
      LAYER met4 ;
        RECT 3439.745 1896.160 3440.725 1931.330 ;
      LAYER met4 ;
        RECT 3441.125 1896.560 3444.105 2780.240 ;
      LAYER met4 ;
        RECT 3444.505 2772.310 3588.000 2780.640 ;
      LAYER met4 ;
        RECT 3444.405 2151.730 3444.735 2771.910 ;
      LAYER met4 ;
        RECT 3445.135 2740.670 3588.000 2772.310 ;
        RECT 3445.135 2740.030 3445.835 2740.670 ;
        RECT 3445.135 2594.000 3445.835 2739.000 ;
        RECT 3445.135 2592.330 3445.835 2593.035 ;
      LAYER met4 ;
        RECT 3446.235 2592.730 3450.685 2740.270 ;
      LAYER met4 ;
        RECT 3451.085 2740.030 3451.685 2740.670 ;
        RECT 3451.085 2594.000 3451.685 2739.000 ;
        RECT 3451.085 2592.330 3451.685 2593.035 ;
      LAYER met4 ;
        RECT 3452.085 2592.730 3456.535 2740.270 ;
      LAYER met4 ;
        RECT 3456.935 2740.030 3457.635 2740.670 ;
        RECT 3456.935 2738.000 3458.035 2739.000 ;
      LAYER met4 ;
        RECT 3458.035 2738.000 3483.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2740.030 3563.385 2740.670 ;
      LAYER met4 ;
        RECT 3563.785 2739.000 3588.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.000 2738.000 3485.035 2739.000 ;
        RECT 3456.935 2735.000 3485.035 2738.000 ;
        RECT 3456.935 2733.000 3458.035 2735.000 ;
      LAYER met4 ;
        RECT 3458.035 2733.000 3483.000 2735.000 ;
      LAYER met4 ;
        RECT 3483.000 2733.000 3485.035 2735.000 ;
        RECT 3456.935 2715.000 3485.035 2733.000 ;
        RECT 3456.935 2713.000 3458.035 2715.000 ;
      LAYER met4 ;
        RECT 3458.035 2713.000 3483.000 2715.000 ;
      LAYER met4 ;
        RECT 3483.000 2713.000 3485.035 2715.000 ;
        RECT 3456.935 2695.000 3485.035 2713.000 ;
        RECT 3456.935 2693.000 3458.035 2695.000 ;
      LAYER met4 ;
        RECT 3458.035 2693.000 3483.000 2695.000 ;
      LAYER met4 ;
        RECT 3483.000 2693.000 3485.035 2695.000 ;
        RECT 3456.935 2675.000 3485.035 2693.000 ;
        RECT 3456.935 2673.000 3458.035 2675.000 ;
      LAYER met4 ;
        RECT 3458.035 2673.000 3483.000 2675.000 ;
      LAYER met4 ;
        RECT 3483.000 2673.000 3485.035 2675.000 ;
        RECT 3456.935 2655.000 3485.035 2673.000 ;
        RECT 3456.935 2653.000 3458.035 2655.000 ;
      LAYER met4 ;
        RECT 3458.035 2653.000 3483.000 2655.000 ;
      LAYER met4 ;
        RECT 3483.000 2653.000 3485.035 2655.000 ;
        RECT 3456.935 2635.000 3485.035 2653.000 ;
        RECT 3456.935 2633.000 3458.035 2635.000 ;
      LAYER met4 ;
        RECT 3458.035 2633.000 3483.000 2635.000 ;
      LAYER met4 ;
        RECT 3483.000 2633.000 3485.035 2635.000 ;
        RECT 3456.935 2615.000 3485.035 2633.000 ;
        RECT 3456.935 2613.000 3458.035 2615.000 ;
      LAYER met4 ;
        RECT 3458.035 2613.000 3483.000 2615.000 ;
      LAYER met4 ;
        RECT 3483.000 2613.000 3485.035 2615.000 ;
        RECT 3456.935 2595.000 3485.035 2613.000 ;
        RECT 3456.935 2594.000 3458.035 2595.000 ;
        RECT 3456.935 2592.330 3457.635 2593.035 ;
      LAYER met4 ;
        RECT 3458.035 2592.730 3483.000 2595.000 ;
      LAYER met4 ;
        RECT 3483.000 2594.000 3485.035 2595.000 ;
        RECT 3562.035 2594.000 3588.000 2739.000 ;
        RECT 3483.400 2592.330 3563.385 2593.035 ;
      LAYER met4 ;
        RECT 3563.785 2592.730 3588.000 2594.000 ;
      LAYER met4 ;
        RECT 3445.135 2520.670 3588.000 2592.330 ;
        RECT 3445.135 2519.965 3445.835 2520.670 ;
        RECT 3445.135 2374.000 3445.835 2519.000 ;
        RECT 3445.135 2372.330 3445.835 2373.035 ;
      LAYER met4 ;
        RECT 3446.235 2372.730 3450.685 2520.270 ;
      LAYER met4 ;
        RECT 3451.085 2519.965 3451.685 2520.670 ;
        RECT 3451.085 2374.000 3451.685 2519.000 ;
        RECT 3451.085 2372.330 3451.685 2373.035 ;
      LAYER met4 ;
        RECT 3452.085 2372.730 3456.535 2520.270 ;
      LAYER met4 ;
        RECT 3456.935 2519.965 3457.635 2520.670 ;
        RECT 3456.935 2518.000 3458.035 2519.000 ;
      LAYER met4 ;
        RECT 3458.035 2518.000 3483.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2519.965 3563.385 2520.670 ;
      LAYER met4 ;
        RECT 3563.785 2519.000 3588.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.000 2518.000 3485.035 2519.000 ;
        RECT 3456.935 2515.000 3485.035 2518.000 ;
        RECT 3456.935 2513.000 3458.035 2515.000 ;
      LAYER met4 ;
        RECT 3458.035 2513.000 3483.000 2515.000 ;
      LAYER met4 ;
        RECT 3483.000 2513.000 3485.035 2515.000 ;
        RECT 3456.935 2495.000 3485.035 2513.000 ;
        RECT 3456.935 2493.000 3458.035 2495.000 ;
      LAYER met4 ;
        RECT 3458.035 2493.000 3483.000 2495.000 ;
      LAYER met4 ;
        RECT 3483.000 2493.000 3485.035 2495.000 ;
        RECT 3456.935 2475.000 3485.035 2493.000 ;
        RECT 3456.935 2473.000 3458.035 2475.000 ;
      LAYER met4 ;
        RECT 3458.035 2473.000 3483.000 2475.000 ;
      LAYER met4 ;
        RECT 3483.000 2473.000 3485.035 2475.000 ;
        RECT 3456.935 2455.000 3485.035 2473.000 ;
        RECT 3456.935 2453.000 3458.035 2455.000 ;
      LAYER met4 ;
        RECT 3458.035 2453.000 3483.000 2455.000 ;
      LAYER met4 ;
        RECT 3483.000 2453.000 3485.035 2455.000 ;
        RECT 3456.935 2435.000 3485.035 2453.000 ;
        RECT 3456.935 2433.000 3458.035 2435.000 ;
      LAYER met4 ;
        RECT 3458.035 2433.000 3483.000 2435.000 ;
      LAYER met4 ;
        RECT 3483.000 2433.000 3485.035 2435.000 ;
        RECT 3456.935 2415.000 3485.035 2433.000 ;
        RECT 3456.935 2413.000 3458.035 2415.000 ;
      LAYER met4 ;
        RECT 3458.035 2413.000 3483.000 2415.000 ;
      LAYER met4 ;
        RECT 3483.000 2413.000 3485.035 2415.000 ;
        RECT 3456.935 2395.000 3485.035 2413.000 ;
        RECT 3456.935 2393.000 3458.035 2395.000 ;
      LAYER met4 ;
        RECT 3458.035 2393.000 3483.000 2395.000 ;
      LAYER met4 ;
        RECT 3483.000 2393.000 3485.035 2395.000 ;
        RECT 3456.935 2375.000 3485.035 2393.000 ;
        RECT 3456.935 2374.000 3458.035 2375.000 ;
        RECT 3456.935 2372.330 3457.635 2373.035 ;
      LAYER met4 ;
        RECT 3458.035 2372.730 3483.000 2375.000 ;
      LAYER met4 ;
        RECT 3483.000 2374.000 3485.035 2375.000 ;
        RECT 3562.035 2374.000 3588.000 2519.000 ;
        RECT 3483.400 2372.330 3563.385 2373.035 ;
      LAYER met4 ;
        RECT 3563.785 2372.730 3588.000 2374.000 ;
      LAYER met4 ;
        RECT 3445.135 2300.670 3588.000 2372.330 ;
        RECT 3445.135 2153.000 3445.835 2300.670 ;
        RECT 3445.135 2151.330 3445.835 2152.035 ;
      LAYER met4 ;
        RECT 3446.235 2151.730 3450.685 2300.270 ;
      LAYER met4 ;
        RECT 3451.085 2299.000 3451.685 2300.670 ;
        RECT 3451.085 2153.000 3451.685 2298.000 ;
        RECT 3451.085 2151.330 3451.685 2152.035 ;
      LAYER met4 ;
        RECT 3452.085 2151.730 3456.535 2300.270 ;
      LAYER met4 ;
        RECT 3456.935 2299.000 3457.635 2300.670 ;
        RECT 3456.935 2297.000 3458.035 2299.000 ;
      LAYER met4 ;
        RECT 3458.035 2297.000 3483.000 2300.270 ;
      LAYER met4 ;
        RECT 3483.400 2299.000 3563.385 2300.670 ;
      LAYER met4 ;
        RECT 3563.785 2299.000 3588.000 2300.270 ;
      LAYER met4 ;
        RECT 3483.000 2297.000 3485.035 2299.000 ;
        RECT 3456.935 2294.000 3485.035 2297.000 ;
        RECT 3456.935 2292.000 3458.035 2294.000 ;
      LAYER met4 ;
        RECT 3458.035 2292.000 3483.000 2294.000 ;
      LAYER met4 ;
        RECT 3483.000 2292.000 3485.035 2294.000 ;
        RECT 3456.935 2274.000 3485.035 2292.000 ;
        RECT 3456.935 2272.000 3458.035 2274.000 ;
      LAYER met4 ;
        RECT 3458.035 2272.000 3483.000 2274.000 ;
      LAYER met4 ;
        RECT 3483.000 2272.000 3485.035 2274.000 ;
        RECT 3456.935 2254.000 3485.035 2272.000 ;
        RECT 3456.935 2252.000 3458.035 2254.000 ;
      LAYER met4 ;
        RECT 3458.035 2252.000 3483.000 2254.000 ;
      LAYER met4 ;
        RECT 3483.000 2252.000 3485.035 2254.000 ;
        RECT 3456.935 2234.000 3485.035 2252.000 ;
        RECT 3456.935 2232.000 3458.035 2234.000 ;
      LAYER met4 ;
        RECT 3458.035 2232.000 3483.000 2234.000 ;
      LAYER met4 ;
        RECT 3483.000 2232.000 3485.035 2234.000 ;
        RECT 3456.935 2214.000 3485.035 2232.000 ;
        RECT 3456.935 2212.000 3458.035 2214.000 ;
      LAYER met4 ;
        RECT 3458.035 2212.000 3483.000 2214.000 ;
      LAYER met4 ;
        RECT 3483.000 2212.000 3485.035 2214.000 ;
        RECT 3456.935 2194.000 3485.035 2212.000 ;
        RECT 3456.935 2192.000 3458.035 2194.000 ;
      LAYER met4 ;
        RECT 3458.035 2192.000 3483.000 2194.000 ;
      LAYER met4 ;
        RECT 3483.000 2192.000 3485.035 2194.000 ;
        RECT 3456.935 2174.000 3485.035 2192.000 ;
        RECT 3456.935 2172.000 3458.035 2174.000 ;
      LAYER met4 ;
        RECT 3458.035 2172.000 3483.000 2174.000 ;
      LAYER met4 ;
        RECT 3483.000 2172.000 3485.035 2174.000 ;
        RECT 3456.935 2154.000 3485.035 2172.000 ;
        RECT 3456.935 2153.000 3458.035 2154.000 ;
        RECT 3456.935 2151.330 3457.635 2152.035 ;
      LAYER met4 ;
        RECT 3458.035 2151.730 3483.000 2154.000 ;
      LAYER met4 ;
        RECT 3483.000 2153.000 3485.035 2154.000 ;
        RECT 3562.035 2153.000 3588.000 2299.000 ;
        RECT 3483.400 2151.330 3563.385 2152.035 ;
      LAYER met4 ;
        RECT 3563.785 2151.730 3588.000 2153.000 ;
      LAYER met4 ;
        RECT 3444.505 2079.670 3588.000 2151.330 ;
      LAYER met4 ;
        RECT 3444.405 1930.390 3444.735 2079.270 ;
      LAYER met4 ;
        RECT 3445.135 2078.965 3445.835 2079.670 ;
        RECT 3445.135 1933.000 3445.835 2078.000 ;
        RECT 3445.135 1931.330 3445.835 1932.035 ;
      LAYER met4 ;
        RECT 3446.235 1931.730 3450.685 2079.270 ;
      LAYER met4 ;
        RECT 3451.085 2078.965 3451.685 2079.670 ;
        RECT 3451.085 1933.000 3451.685 2078.000 ;
        RECT 3451.085 1931.330 3451.685 1932.035 ;
      LAYER met4 ;
        RECT 3452.085 1931.730 3456.535 2079.270 ;
      LAYER met4 ;
        RECT 3456.935 2078.965 3457.635 2079.670 ;
        RECT 3456.935 2077.000 3458.035 2078.000 ;
      LAYER met4 ;
        RECT 3458.035 2077.000 3483.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 2078.965 3563.385 2079.670 ;
      LAYER met4 ;
        RECT 3563.785 2078.000 3588.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.000 2077.000 3485.035 2078.000 ;
        RECT 3456.935 2074.000 3485.035 2077.000 ;
        RECT 3456.935 2072.000 3458.035 2074.000 ;
      LAYER met4 ;
        RECT 3458.035 2072.000 3483.000 2074.000 ;
      LAYER met4 ;
        RECT 3483.000 2072.000 3485.035 2074.000 ;
        RECT 3456.935 2054.000 3485.035 2072.000 ;
        RECT 3456.935 2052.000 3458.035 2054.000 ;
      LAYER met4 ;
        RECT 3458.035 2052.000 3483.000 2054.000 ;
      LAYER met4 ;
        RECT 3483.000 2052.000 3485.035 2054.000 ;
        RECT 3456.935 2034.000 3485.035 2052.000 ;
        RECT 3456.935 2032.000 3458.035 2034.000 ;
      LAYER met4 ;
        RECT 3458.035 2032.000 3483.000 2034.000 ;
      LAYER met4 ;
        RECT 3483.000 2032.000 3485.035 2034.000 ;
        RECT 3456.935 2014.000 3485.035 2032.000 ;
        RECT 3456.935 2012.000 3458.035 2014.000 ;
      LAYER met4 ;
        RECT 3458.035 2012.000 3483.000 2014.000 ;
      LAYER met4 ;
        RECT 3483.000 2012.000 3485.035 2014.000 ;
        RECT 3456.935 1994.000 3485.035 2012.000 ;
        RECT 3456.935 1992.000 3458.035 1994.000 ;
      LAYER met4 ;
        RECT 3458.035 1992.000 3483.000 1994.000 ;
      LAYER met4 ;
        RECT 3483.000 1992.000 3485.035 1994.000 ;
        RECT 3456.935 1974.000 3485.035 1992.000 ;
        RECT 3456.935 1972.000 3458.035 1974.000 ;
      LAYER met4 ;
        RECT 3458.035 1972.000 3483.000 1974.000 ;
      LAYER met4 ;
        RECT 3483.000 1972.000 3485.035 1974.000 ;
        RECT 3456.935 1954.000 3485.035 1972.000 ;
        RECT 3456.935 1952.000 3458.035 1954.000 ;
      LAYER met4 ;
        RECT 3458.035 1952.000 3483.000 1954.000 ;
      LAYER met4 ;
        RECT 3483.000 1952.000 3485.035 1954.000 ;
        RECT 3456.935 1934.000 3485.035 1952.000 ;
        RECT 3456.935 1933.000 3458.035 1934.000 ;
        RECT 3456.935 1931.330 3457.635 1932.035 ;
      LAYER met4 ;
        RECT 3458.035 1931.730 3483.000 1934.000 ;
      LAYER met4 ;
        RECT 3483.000 1933.000 3485.035 1934.000 ;
        RECT 3562.035 1933.000 3588.000 2078.000 ;
        RECT 3483.400 1931.330 3563.385 1932.035 ;
      LAYER met4 ;
        RECT 3563.785 1931.730 3588.000 1933.000 ;
      LAYER met4 ;
        RECT 3445.135 1929.990 3588.000 1931.330 ;
        RECT 3444.505 1896.160 3588.000 1929.990 ;
        RECT 3439.745 1894.640 3588.000 1896.160 ;
        RECT 3439.745 1880.455 3440.725 1894.640 ;
        RECT 3436.465 1878.935 3440.725 1880.455 ;
        RECT 3388.535 1660.310 3435.965 1703.990 ;
        RECT 198.365 1634.330 199.465 1634.970 ;
        RECT 152.665 1602.690 199.465 1634.330 ;
        RECT 3388.535 1628.670 3435.335 1660.310 ;
        RECT 3388.535 1628.030 3389.635 1628.670 ;
        RECT 152.035 1559.010 199.465 1602.690 ;
        RECT 147.275 1392.545 151.535 1394.065 ;
        RECT 147.275 1378.360 148.255 1392.545 ;
        RECT 0.000 1376.840 148.255 1378.360 ;
        RECT 0.000 1343.010 143.495 1376.840 ;
        RECT 0.000 1341.670 142.865 1343.010 ;
      LAYER met4 ;
        RECT 0.000 1340.000 24.215 1341.270 ;
      LAYER met4 ;
        RECT 24.615 1340.965 104.600 1341.670 ;
        RECT 0.000 1204.000 25.965 1340.000 ;
        RECT 102.965 1338.000 105.000 1340.000 ;
      LAYER met4 ;
        RECT 105.000 1338.000 129.965 1341.270 ;
      LAYER met4 ;
        RECT 130.365 1340.965 131.065 1341.670 ;
        RECT 129.965 1338.000 131.065 1340.000 ;
        RECT 102.965 1335.000 131.065 1338.000 ;
        RECT 102.965 1333.000 105.000 1335.000 ;
      LAYER met4 ;
        RECT 105.000 1333.000 129.965 1335.000 ;
      LAYER met4 ;
        RECT 129.965 1333.000 131.065 1335.000 ;
        RECT 102.965 1325.000 131.065 1333.000 ;
        RECT 102.965 1323.000 105.000 1325.000 ;
      LAYER met4 ;
        RECT 105.000 1323.000 129.965 1325.000 ;
      LAYER met4 ;
        RECT 129.965 1323.000 131.065 1325.000 ;
        RECT 102.965 1305.000 131.065 1323.000 ;
        RECT 102.965 1303.000 105.000 1305.000 ;
      LAYER met4 ;
        RECT 105.000 1303.000 129.965 1305.000 ;
      LAYER met4 ;
        RECT 129.965 1303.000 131.065 1305.000 ;
        RECT 102.965 1285.000 131.065 1303.000 ;
        RECT 102.965 1283.000 105.000 1285.000 ;
      LAYER met4 ;
        RECT 105.000 1283.000 129.965 1285.000 ;
      LAYER met4 ;
        RECT 129.965 1283.000 131.065 1285.000 ;
        RECT 102.965 1265.000 131.065 1283.000 ;
        RECT 102.965 1263.000 105.000 1265.000 ;
      LAYER met4 ;
        RECT 105.000 1263.000 129.965 1265.000 ;
      LAYER met4 ;
        RECT 129.965 1263.000 131.065 1265.000 ;
        RECT 102.965 1245.000 131.065 1263.000 ;
        RECT 102.965 1243.000 105.000 1245.000 ;
      LAYER met4 ;
        RECT 105.000 1243.000 129.965 1245.000 ;
      LAYER met4 ;
        RECT 129.965 1243.000 131.065 1245.000 ;
        RECT 102.965 1225.000 131.065 1243.000 ;
        RECT 102.965 1223.000 105.000 1225.000 ;
      LAYER met4 ;
        RECT 105.000 1223.000 129.965 1225.000 ;
      LAYER met4 ;
        RECT 129.965 1223.000 131.065 1225.000 ;
        RECT 102.965 1205.000 131.065 1223.000 ;
        RECT 102.965 1204.000 105.000 1205.000 ;
      LAYER met4 ;
        RECT 0.000 1202.730 24.215 1204.000 ;
      LAYER met4 ;
        RECT 24.615 1202.330 104.600 1202.970 ;
      LAYER met4 ;
        RECT 105.000 1202.730 129.965 1205.000 ;
      LAYER met4 ;
        RECT 129.965 1204.000 131.065 1205.000 ;
        RECT 130.365 1202.330 131.065 1202.970 ;
      LAYER met4 ;
        RECT 131.465 1202.730 135.915 1341.270 ;
      LAYER met4 ;
        RECT 136.315 1340.965 136.915 1341.670 ;
        RECT 136.315 1204.000 136.915 1339.000 ;
        RECT 136.315 1202.330 136.915 1202.970 ;
      LAYER met4 ;
        RECT 137.315 1202.730 141.765 1341.270 ;
      LAYER met4 ;
        RECT 142.165 1340.965 142.865 1341.670 ;
        RECT 142.165 1204.000 142.865 1340.000 ;
        RECT 142.165 1202.330 142.865 1202.970 ;
        RECT 0.000 1170.690 142.865 1202.330 ;
      LAYER met4 ;
        RECT 143.265 1171.090 143.595 1342.610 ;
      LAYER met4 ;
        RECT 0.000 1162.360 143.495 1170.690 ;
      LAYER met4 ;
        RECT 143.895 1162.760 146.875 1376.440 ;
      LAYER met4 ;
        RECT 147.275 1341.670 148.255 1376.840 ;
      LAYER met4 ;
        RECT 147.175 1340.000 148.355 1341.270 ;
      LAYER met4 ;
        RECT 147.275 1204.000 148.255 1340.000 ;
      LAYER met4 ;
        RECT 147.175 1202.730 148.355 1204.000 ;
      LAYER met4 ;
        RECT 147.275 1178.065 148.255 1202.330 ;
      LAYER met4 ;
        RECT 148.655 1178.465 151.635 1392.145 ;
        RECT 151.935 1387.090 152.265 1558.610 ;
      LAYER met4 ;
        RECT 152.665 1557.670 199.465 1559.010 ;
        RECT 152.665 1556.965 153.365 1557.670 ;
        RECT 152.665 1418.330 153.365 1418.970 ;
      LAYER met4 ;
        RECT 153.765 1418.730 158.415 1557.270 ;
      LAYER met4 ;
        RECT 158.815 1556.965 159.415 1557.670 ;
        RECT 158.815 1418.330 159.415 1418.970 ;
      LAYER met4 ;
        RECT 159.815 1418.730 163.265 1557.270 ;
      LAYER met4 ;
        RECT 163.665 1556.965 164.265 1557.670 ;
        RECT 163.665 1418.330 164.265 1418.970 ;
      LAYER met4 ;
        RECT 164.665 1418.730 168.115 1557.270 ;
      LAYER met4 ;
        RECT 168.515 1556.965 169.115 1557.670 ;
        RECT 168.515 1418.330 169.115 1418.970 ;
      LAYER met4 ;
        RECT 169.515 1418.730 174.165 1557.270 ;
      LAYER met4 ;
        RECT 174.565 1556.965 175.165 1557.670 ;
        RECT 180.615 1557.365 186.065 1557.670 ;
        RECT 174.565 1418.330 175.165 1418.970 ;
      LAYER met4 ;
        RECT 175.565 1418.730 180.215 1557.270 ;
      LAYER met4 ;
        RECT 180.615 1556.965 181.215 1557.365 ;
        RECT 185.465 1556.965 186.065 1557.365 ;
      LAYER met4 ;
        RECT 181.615 1418.970 185.065 1556.965 ;
      LAYER met4 ;
        RECT 180.615 1418.570 181.215 1418.970 ;
        RECT 185.465 1418.570 186.065 1418.970 ;
      LAYER met4 ;
        RECT 186.465 1418.730 191.115 1557.270 ;
      LAYER met4 ;
        RECT 191.515 1556.965 192.115 1557.670 ;
        RECT 180.615 1418.330 186.065 1418.570 ;
        RECT 191.515 1418.330 192.115 1418.970 ;
      LAYER met4 ;
        RECT 192.515 1418.730 197.965 1557.270 ;
      LAYER met4 ;
        RECT 198.365 1556.965 199.465 1557.670 ;
        RECT 3388.535 1480.330 3389.635 1481.035 ;
      LAYER met4 ;
        RECT 3390.035 1480.730 3395.485 1628.270 ;
      LAYER met4 ;
        RECT 3395.885 1628.030 3396.485 1628.670 ;
        RECT 3401.935 1628.430 3407.385 1628.670 ;
        RECT 3395.885 1480.330 3396.485 1481.035 ;
      LAYER met4 ;
        RECT 3396.885 1480.730 3401.535 1628.270 ;
      LAYER met4 ;
        RECT 3401.935 1628.030 3402.535 1628.430 ;
        RECT 3406.785 1628.030 3407.385 1628.430 ;
      LAYER met4 ;
        RECT 3402.935 1481.035 3406.385 1628.030 ;
      LAYER met4 ;
        RECT 3401.935 1480.635 3402.535 1481.035 ;
        RECT 3406.785 1480.635 3407.385 1481.035 ;
      LAYER met4 ;
        RECT 3407.785 1480.730 3412.435 1628.270 ;
      LAYER met4 ;
        RECT 3412.835 1628.030 3413.435 1628.670 ;
        RECT 3401.935 1480.330 3407.385 1480.635 ;
        RECT 3412.835 1480.330 3413.435 1481.035 ;
      LAYER met4 ;
        RECT 3413.835 1480.730 3418.485 1628.270 ;
      LAYER met4 ;
        RECT 3418.885 1628.030 3419.485 1628.670 ;
        RECT 3418.885 1480.330 3419.485 1481.035 ;
      LAYER met4 ;
        RECT 3419.885 1480.730 3423.335 1628.270 ;
      LAYER met4 ;
        RECT 3423.735 1628.030 3424.335 1628.670 ;
        RECT 3423.735 1480.330 3424.335 1481.035 ;
      LAYER met4 ;
        RECT 3424.735 1480.730 3428.185 1628.270 ;
      LAYER met4 ;
        RECT 3428.585 1628.030 3429.185 1628.670 ;
        RECT 3428.585 1480.330 3429.185 1481.035 ;
      LAYER met4 ;
        RECT 3429.585 1480.730 3434.235 1628.270 ;
      LAYER met4 ;
        RECT 3434.635 1628.030 3435.335 1628.670 ;
        RECT 3434.635 1480.330 3435.335 1481.035 ;
        RECT 3388.535 1478.990 3435.335 1480.330 ;
      LAYER met4 ;
        RECT 3435.735 1479.390 3436.065 1659.910 ;
        RECT 3436.365 1654.855 3439.345 1878.535 ;
      LAYER met4 ;
        RECT 3439.745 1854.670 3440.725 1878.935 ;
      LAYER met4 ;
        RECT 3439.645 1853.000 3440.825 1854.270 ;
      LAYER met4 ;
        RECT 3439.745 1707.000 3440.725 1853.000 ;
      LAYER met4 ;
        RECT 3439.645 1705.730 3440.825 1707.000 ;
      LAYER met4 ;
        RECT 3439.745 1670.160 3440.725 1705.330 ;
      LAYER met4 ;
        RECT 3441.125 1670.560 3444.105 1894.240 ;
      LAYER met4 ;
        RECT 3444.505 1886.310 3588.000 1894.640 ;
      LAYER met4 ;
        RECT 3444.405 1704.390 3444.735 1885.910 ;
      LAYER met4 ;
        RECT 3445.135 1854.670 3588.000 1886.310 ;
        RECT 3445.135 1854.030 3445.835 1854.670 ;
        RECT 3445.135 1707.000 3445.835 1853.000 ;
        RECT 3445.135 1705.330 3445.835 1706.035 ;
      LAYER met4 ;
        RECT 3446.235 1705.730 3450.685 1854.270 ;
      LAYER met4 ;
        RECT 3451.085 1854.030 3451.685 1854.670 ;
        RECT 3451.085 1707.000 3451.685 1852.000 ;
        RECT 3451.085 1705.330 3451.685 1706.035 ;
      LAYER met4 ;
        RECT 3452.085 1705.730 3456.535 1854.270 ;
      LAYER met4 ;
        RECT 3456.935 1854.030 3457.635 1854.670 ;
        RECT 3456.935 1851.000 3458.035 1853.000 ;
      LAYER met4 ;
        RECT 3458.035 1851.000 3483.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1854.030 3563.385 1854.670 ;
      LAYER met4 ;
        RECT 3563.785 1853.000 3588.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.000 1851.000 3485.035 1853.000 ;
        RECT 3456.935 1848.000 3485.035 1851.000 ;
        RECT 3456.935 1846.000 3458.035 1848.000 ;
      LAYER met4 ;
        RECT 3458.035 1846.000 3483.000 1848.000 ;
      LAYER met4 ;
        RECT 3483.000 1846.000 3485.035 1848.000 ;
        RECT 3456.935 1828.000 3485.035 1846.000 ;
        RECT 3456.935 1826.000 3458.035 1828.000 ;
      LAYER met4 ;
        RECT 3458.035 1826.000 3483.000 1828.000 ;
      LAYER met4 ;
        RECT 3483.000 1826.000 3485.035 1828.000 ;
        RECT 3456.935 1808.000 3485.035 1826.000 ;
        RECT 3456.935 1806.000 3458.035 1808.000 ;
      LAYER met4 ;
        RECT 3458.035 1806.000 3483.000 1808.000 ;
      LAYER met4 ;
        RECT 3483.000 1806.000 3485.035 1808.000 ;
        RECT 3456.935 1788.000 3485.035 1806.000 ;
        RECT 3456.935 1786.000 3458.035 1788.000 ;
      LAYER met4 ;
        RECT 3458.035 1786.000 3483.000 1788.000 ;
      LAYER met4 ;
        RECT 3483.000 1786.000 3485.035 1788.000 ;
        RECT 3456.935 1768.000 3485.035 1786.000 ;
        RECT 3456.935 1766.000 3458.035 1768.000 ;
      LAYER met4 ;
        RECT 3458.035 1766.000 3483.000 1768.000 ;
      LAYER met4 ;
        RECT 3483.000 1766.000 3485.035 1768.000 ;
        RECT 3456.935 1748.000 3485.035 1766.000 ;
        RECT 3456.935 1746.000 3458.035 1748.000 ;
      LAYER met4 ;
        RECT 3458.035 1746.000 3483.000 1748.000 ;
      LAYER met4 ;
        RECT 3483.000 1746.000 3485.035 1748.000 ;
        RECT 3456.935 1728.000 3485.035 1746.000 ;
        RECT 3456.935 1726.000 3458.035 1728.000 ;
      LAYER met4 ;
        RECT 3458.035 1726.000 3483.000 1728.000 ;
      LAYER met4 ;
        RECT 3483.000 1726.000 3485.035 1728.000 ;
        RECT 3456.935 1708.000 3485.035 1726.000 ;
        RECT 3456.935 1707.000 3458.035 1708.000 ;
        RECT 3456.935 1705.330 3457.635 1706.035 ;
      LAYER met4 ;
        RECT 3458.035 1705.730 3483.000 1708.000 ;
      LAYER met4 ;
        RECT 3483.000 1707.000 3485.035 1708.000 ;
        RECT 3562.035 1707.000 3588.000 1853.000 ;
        RECT 3483.400 1705.330 3563.385 1706.035 ;
      LAYER met4 ;
        RECT 3563.785 1705.730 3588.000 1707.000 ;
      LAYER met4 ;
        RECT 3445.135 1703.990 3588.000 1705.330 ;
        RECT 3444.505 1670.160 3588.000 1703.990 ;
        RECT 3439.745 1668.640 3588.000 1670.160 ;
        RECT 3439.745 1654.455 3440.725 1668.640 ;
        RECT 3436.465 1652.935 3440.725 1654.455 ;
        RECT 3388.535 1435.310 3435.965 1478.990 ;
        RECT 198.365 1418.330 199.465 1418.970 ;
        RECT 152.665 1386.690 199.465 1418.330 ;
        RECT 3388.535 1403.670 3435.335 1435.310 ;
        RECT 3388.535 1403.030 3389.635 1403.670 ;
        RECT 152.035 1343.010 199.465 1386.690 ;
        RECT 147.275 1176.545 151.535 1178.065 ;
        RECT 147.275 1162.360 148.255 1176.545 ;
        RECT 0.000 1160.840 148.255 1162.360 ;
        RECT 0.000 1127.010 143.495 1160.840 ;
        RECT 0.000 1125.670 142.865 1127.010 ;
      LAYER met4 ;
        RECT 0.000 1124.000 24.215 1125.270 ;
      LAYER met4 ;
        RECT 24.615 1124.965 104.600 1125.670 ;
        RECT 0.000 988.000 25.965 1124.000 ;
        RECT 102.965 1122.000 105.000 1124.000 ;
      LAYER met4 ;
        RECT 105.000 1122.000 129.965 1125.270 ;
      LAYER met4 ;
        RECT 130.365 1124.965 131.065 1125.670 ;
        RECT 129.965 1122.000 131.065 1124.000 ;
        RECT 102.965 1119.000 131.065 1122.000 ;
        RECT 102.965 1117.000 105.000 1119.000 ;
      LAYER met4 ;
        RECT 105.000 1117.000 129.965 1119.000 ;
      LAYER met4 ;
        RECT 129.965 1117.000 131.065 1119.000 ;
        RECT 102.965 1109.000 131.065 1117.000 ;
        RECT 102.965 1107.000 105.000 1109.000 ;
      LAYER met4 ;
        RECT 105.000 1107.000 129.965 1109.000 ;
      LAYER met4 ;
        RECT 129.965 1107.000 131.065 1109.000 ;
        RECT 102.965 1089.000 131.065 1107.000 ;
        RECT 102.965 1087.000 105.000 1089.000 ;
      LAYER met4 ;
        RECT 105.000 1087.000 129.965 1089.000 ;
      LAYER met4 ;
        RECT 129.965 1087.000 131.065 1089.000 ;
        RECT 102.965 1069.000 131.065 1087.000 ;
        RECT 102.965 1067.000 105.000 1069.000 ;
      LAYER met4 ;
        RECT 105.000 1067.000 129.965 1069.000 ;
      LAYER met4 ;
        RECT 129.965 1067.000 131.065 1069.000 ;
        RECT 102.965 1049.000 131.065 1067.000 ;
        RECT 102.965 1047.000 105.000 1049.000 ;
      LAYER met4 ;
        RECT 105.000 1047.000 129.965 1049.000 ;
      LAYER met4 ;
        RECT 129.965 1047.000 131.065 1049.000 ;
        RECT 102.965 1029.000 131.065 1047.000 ;
        RECT 102.965 1027.000 105.000 1029.000 ;
      LAYER met4 ;
        RECT 105.000 1027.000 129.965 1029.000 ;
      LAYER met4 ;
        RECT 129.965 1027.000 131.065 1029.000 ;
        RECT 102.965 1009.000 131.065 1027.000 ;
        RECT 102.965 1007.000 105.000 1009.000 ;
      LAYER met4 ;
        RECT 105.000 1007.000 129.965 1009.000 ;
      LAYER met4 ;
        RECT 129.965 1007.000 131.065 1009.000 ;
        RECT 102.965 989.000 131.065 1007.000 ;
        RECT 102.965 988.000 105.000 989.000 ;
      LAYER met4 ;
        RECT 0.000 986.730 24.215 988.000 ;
      LAYER met4 ;
        RECT 24.615 986.330 104.600 986.970 ;
      LAYER met4 ;
        RECT 105.000 986.730 129.965 989.000 ;
      LAYER met4 ;
        RECT 129.965 988.000 131.065 989.000 ;
        RECT 130.365 986.330 131.065 986.970 ;
      LAYER met4 ;
        RECT 131.465 986.730 135.915 1125.270 ;
      LAYER met4 ;
        RECT 136.315 1124.965 136.915 1125.670 ;
        RECT 136.315 988.000 136.915 1123.000 ;
        RECT 136.315 986.330 136.915 986.970 ;
      LAYER met4 ;
        RECT 137.315 986.730 141.765 1125.270 ;
      LAYER met4 ;
        RECT 142.165 1124.965 142.865 1125.670 ;
        RECT 142.165 988.000 142.865 1124.000 ;
        RECT 142.165 986.330 142.865 986.970 ;
        RECT 0.000 954.690 142.865 986.330 ;
      LAYER met4 ;
        RECT 143.265 955.090 143.595 1126.610 ;
      LAYER met4 ;
        RECT 0.000 946.360 143.495 954.690 ;
      LAYER met4 ;
        RECT 143.895 946.760 146.875 1160.440 ;
      LAYER met4 ;
        RECT 147.275 1125.670 148.255 1160.840 ;
      LAYER met4 ;
        RECT 147.175 1124.000 148.355 1125.270 ;
      LAYER met4 ;
        RECT 147.275 988.000 148.255 1124.000 ;
      LAYER met4 ;
        RECT 147.175 986.730 148.355 988.000 ;
      LAYER met4 ;
        RECT 147.275 962.065 148.255 986.330 ;
      LAYER met4 ;
        RECT 148.655 962.465 151.635 1176.145 ;
        RECT 151.935 1171.090 152.265 1342.610 ;
      LAYER met4 ;
        RECT 152.665 1341.670 199.465 1343.010 ;
        RECT 152.665 1340.965 153.365 1341.670 ;
        RECT 152.665 1202.330 153.365 1202.970 ;
      LAYER met4 ;
        RECT 153.765 1202.730 158.415 1341.270 ;
      LAYER met4 ;
        RECT 158.815 1340.965 159.415 1341.670 ;
        RECT 158.815 1202.330 159.415 1202.970 ;
      LAYER met4 ;
        RECT 159.815 1202.730 163.265 1341.270 ;
      LAYER met4 ;
        RECT 163.665 1340.965 164.265 1341.670 ;
        RECT 163.665 1202.330 164.265 1202.970 ;
      LAYER met4 ;
        RECT 164.665 1202.730 168.115 1341.270 ;
      LAYER met4 ;
        RECT 168.515 1340.965 169.115 1341.670 ;
        RECT 168.515 1202.330 169.115 1202.970 ;
      LAYER met4 ;
        RECT 169.515 1202.730 174.165 1341.270 ;
      LAYER met4 ;
        RECT 174.565 1340.965 175.165 1341.670 ;
        RECT 180.615 1341.365 186.065 1341.670 ;
        RECT 174.565 1202.330 175.165 1202.970 ;
      LAYER met4 ;
        RECT 175.565 1202.730 180.215 1341.270 ;
      LAYER met4 ;
        RECT 180.615 1340.965 181.215 1341.365 ;
        RECT 185.465 1340.965 186.065 1341.365 ;
      LAYER met4 ;
        RECT 181.615 1202.970 185.065 1340.965 ;
      LAYER met4 ;
        RECT 180.615 1202.570 181.215 1202.970 ;
        RECT 185.465 1202.570 186.065 1202.970 ;
      LAYER met4 ;
        RECT 186.465 1202.730 191.115 1341.270 ;
      LAYER met4 ;
        RECT 191.515 1340.965 192.115 1341.670 ;
        RECT 180.615 1202.330 186.065 1202.570 ;
        RECT 191.515 1202.330 192.115 1202.970 ;
      LAYER met4 ;
        RECT 192.515 1202.730 197.965 1341.270 ;
      LAYER met4 ;
        RECT 198.365 1340.965 199.465 1341.670 ;
        RECT 3388.535 1255.330 3389.635 1256.035 ;
      LAYER met4 ;
        RECT 3390.035 1255.730 3395.485 1403.270 ;
      LAYER met4 ;
        RECT 3395.885 1403.030 3396.485 1403.670 ;
        RECT 3401.935 1403.430 3407.385 1403.670 ;
        RECT 3395.885 1255.330 3396.485 1256.035 ;
      LAYER met4 ;
        RECT 3396.885 1255.730 3401.535 1403.270 ;
      LAYER met4 ;
        RECT 3401.935 1403.030 3402.535 1403.430 ;
        RECT 3406.785 1403.030 3407.385 1403.430 ;
      LAYER met4 ;
        RECT 3402.935 1256.035 3406.385 1403.030 ;
      LAYER met4 ;
        RECT 3401.935 1255.635 3402.535 1256.035 ;
        RECT 3406.785 1255.635 3407.385 1256.035 ;
      LAYER met4 ;
        RECT 3407.785 1255.730 3412.435 1403.270 ;
      LAYER met4 ;
        RECT 3412.835 1403.030 3413.435 1403.670 ;
        RECT 3401.935 1255.330 3407.385 1255.635 ;
        RECT 3412.835 1255.330 3413.435 1256.035 ;
      LAYER met4 ;
        RECT 3413.835 1255.730 3418.485 1403.270 ;
      LAYER met4 ;
        RECT 3418.885 1403.030 3419.485 1403.670 ;
        RECT 3418.885 1255.330 3419.485 1256.035 ;
      LAYER met4 ;
        RECT 3419.885 1255.730 3423.335 1403.270 ;
      LAYER met4 ;
        RECT 3423.735 1403.030 3424.335 1403.670 ;
        RECT 3423.735 1255.330 3424.335 1256.035 ;
      LAYER met4 ;
        RECT 3424.735 1255.730 3428.185 1403.270 ;
      LAYER met4 ;
        RECT 3428.585 1403.030 3429.185 1403.670 ;
        RECT 3428.585 1255.330 3429.185 1256.035 ;
      LAYER met4 ;
        RECT 3429.585 1255.730 3434.235 1403.270 ;
      LAYER met4 ;
        RECT 3434.635 1403.030 3435.335 1403.670 ;
        RECT 3434.635 1255.330 3435.335 1256.035 ;
        RECT 3388.535 1253.990 3435.335 1255.330 ;
      LAYER met4 ;
        RECT 3435.735 1254.390 3436.065 1434.910 ;
        RECT 3436.365 1429.855 3439.345 1652.535 ;
      LAYER met4 ;
        RECT 3439.745 1628.670 3440.725 1652.935 ;
      LAYER met4 ;
        RECT 3439.645 1627.000 3440.825 1628.270 ;
      LAYER met4 ;
        RECT 3439.745 1482.000 3440.725 1627.000 ;
      LAYER met4 ;
        RECT 3439.645 1480.730 3440.825 1482.000 ;
      LAYER met4 ;
        RECT 3439.745 1445.160 3440.725 1480.330 ;
      LAYER met4 ;
        RECT 3441.125 1445.560 3444.105 1668.240 ;
      LAYER met4 ;
        RECT 3444.505 1660.310 3588.000 1668.640 ;
      LAYER met4 ;
        RECT 3444.405 1479.390 3444.735 1659.910 ;
      LAYER met4 ;
        RECT 3445.135 1628.670 3588.000 1660.310 ;
        RECT 3445.135 1628.030 3445.835 1628.670 ;
        RECT 3445.135 1482.000 3445.835 1627.000 ;
        RECT 3445.135 1480.330 3445.835 1481.035 ;
      LAYER met4 ;
        RECT 3446.235 1480.730 3450.685 1628.270 ;
      LAYER met4 ;
        RECT 3451.085 1628.030 3451.685 1628.670 ;
        RECT 3451.085 1482.000 3451.685 1627.000 ;
        RECT 3451.085 1480.330 3451.685 1481.035 ;
      LAYER met4 ;
        RECT 3452.085 1480.730 3456.535 1628.270 ;
      LAYER met4 ;
        RECT 3456.935 1628.030 3457.635 1628.670 ;
        RECT 3456.935 1626.000 3458.035 1627.000 ;
      LAYER met4 ;
        RECT 3458.035 1626.000 3483.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1628.030 3563.385 1628.670 ;
      LAYER met4 ;
        RECT 3563.785 1627.000 3588.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.000 1626.000 3485.035 1627.000 ;
        RECT 3456.935 1623.000 3485.035 1626.000 ;
        RECT 3456.935 1621.000 3458.035 1623.000 ;
      LAYER met4 ;
        RECT 3458.035 1621.000 3483.000 1623.000 ;
      LAYER met4 ;
        RECT 3483.000 1621.000 3485.035 1623.000 ;
        RECT 3456.935 1603.000 3485.035 1621.000 ;
        RECT 3456.935 1601.000 3458.035 1603.000 ;
      LAYER met4 ;
        RECT 3458.035 1601.000 3483.000 1603.000 ;
      LAYER met4 ;
        RECT 3483.000 1601.000 3485.035 1603.000 ;
        RECT 3456.935 1583.000 3485.035 1601.000 ;
        RECT 3456.935 1581.000 3458.035 1583.000 ;
      LAYER met4 ;
        RECT 3458.035 1581.000 3483.000 1583.000 ;
      LAYER met4 ;
        RECT 3483.000 1581.000 3485.035 1583.000 ;
        RECT 3456.935 1563.000 3485.035 1581.000 ;
        RECT 3456.935 1561.000 3458.035 1563.000 ;
      LAYER met4 ;
        RECT 3458.035 1561.000 3483.000 1563.000 ;
      LAYER met4 ;
        RECT 3483.000 1561.000 3485.035 1563.000 ;
        RECT 3456.935 1543.000 3485.035 1561.000 ;
        RECT 3456.935 1541.000 3458.035 1543.000 ;
      LAYER met4 ;
        RECT 3458.035 1541.000 3483.000 1543.000 ;
      LAYER met4 ;
        RECT 3483.000 1541.000 3485.035 1543.000 ;
        RECT 3456.935 1523.000 3485.035 1541.000 ;
        RECT 3456.935 1521.000 3458.035 1523.000 ;
      LAYER met4 ;
        RECT 3458.035 1521.000 3483.000 1523.000 ;
      LAYER met4 ;
        RECT 3483.000 1521.000 3485.035 1523.000 ;
        RECT 3456.935 1503.000 3485.035 1521.000 ;
        RECT 3456.935 1501.000 3458.035 1503.000 ;
      LAYER met4 ;
        RECT 3458.035 1501.000 3483.000 1503.000 ;
      LAYER met4 ;
        RECT 3483.000 1501.000 3485.035 1503.000 ;
        RECT 3456.935 1483.000 3485.035 1501.000 ;
        RECT 3456.935 1482.000 3458.035 1483.000 ;
        RECT 3456.935 1480.330 3457.635 1481.035 ;
      LAYER met4 ;
        RECT 3458.035 1480.730 3483.000 1483.000 ;
      LAYER met4 ;
        RECT 3483.000 1482.000 3485.035 1483.000 ;
        RECT 3562.035 1482.000 3588.000 1627.000 ;
        RECT 3483.400 1480.330 3563.385 1481.035 ;
      LAYER met4 ;
        RECT 3563.785 1480.730 3588.000 1482.000 ;
      LAYER met4 ;
        RECT 3445.135 1478.990 3588.000 1480.330 ;
        RECT 3444.505 1445.160 3588.000 1478.990 ;
        RECT 3439.745 1443.640 3588.000 1445.160 ;
        RECT 3439.745 1429.455 3440.725 1443.640 ;
        RECT 3436.465 1427.935 3440.725 1429.455 ;
        RECT 3388.535 1210.310 3435.965 1253.990 ;
        RECT 198.365 1202.330 199.465 1202.970 ;
        RECT 152.665 1170.690 199.465 1202.330 ;
        RECT 3388.535 1178.670 3435.335 1210.310 ;
        RECT 3388.535 1178.030 3389.635 1178.670 ;
        RECT 152.035 1127.010 199.465 1170.690 ;
        RECT 147.275 960.545 151.535 962.065 ;
        RECT 147.275 946.360 148.255 960.545 ;
        RECT 0.000 944.840 148.255 946.360 ;
        RECT 0.000 911.010 143.495 944.840 ;
        RECT 0.000 909.670 142.865 911.010 ;
      LAYER met4 ;
        RECT 0.000 908.000 24.215 909.270 ;
      LAYER met4 ;
        RECT 24.615 908.965 104.600 909.670 ;
        RECT 0.000 772.000 25.965 908.000 ;
        RECT 102.965 906.000 105.000 908.000 ;
      LAYER met4 ;
        RECT 105.000 906.000 129.965 909.270 ;
      LAYER met4 ;
        RECT 130.365 908.965 131.065 909.670 ;
        RECT 129.965 906.000 131.065 908.000 ;
        RECT 102.965 903.000 131.065 906.000 ;
        RECT 102.965 901.000 105.000 903.000 ;
      LAYER met4 ;
        RECT 105.000 901.000 129.965 903.000 ;
      LAYER met4 ;
        RECT 129.965 901.000 131.065 903.000 ;
        RECT 102.965 893.000 131.065 901.000 ;
        RECT 102.965 891.000 105.000 893.000 ;
      LAYER met4 ;
        RECT 105.000 891.000 129.965 893.000 ;
      LAYER met4 ;
        RECT 129.965 891.000 131.065 893.000 ;
        RECT 102.965 873.000 131.065 891.000 ;
        RECT 102.965 871.000 105.000 873.000 ;
      LAYER met4 ;
        RECT 105.000 871.000 129.965 873.000 ;
      LAYER met4 ;
        RECT 129.965 871.000 131.065 873.000 ;
        RECT 102.965 853.000 131.065 871.000 ;
        RECT 102.965 851.000 105.000 853.000 ;
      LAYER met4 ;
        RECT 105.000 851.000 129.965 853.000 ;
      LAYER met4 ;
        RECT 129.965 851.000 131.065 853.000 ;
        RECT 102.965 833.000 131.065 851.000 ;
        RECT 102.965 831.000 105.000 833.000 ;
      LAYER met4 ;
        RECT 105.000 831.000 129.965 833.000 ;
      LAYER met4 ;
        RECT 129.965 831.000 131.065 833.000 ;
        RECT 102.965 813.000 131.065 831.000 ;
        RECT 102.965 811.000 105.000 813.000 ;
      LAYER met4 ;
        RECT 105.000 811.000 129.965 813.000 ;
      LAYER met4 ;
        RECT 129.965 811.000 131.065 813.000 ;
        RECT 102.965 793.000 131.065 811.000 ;
        RECT 102.965 791.000 105.000 793.000 ;
      LAYER met4 ;
        RECT 105.000 791.000 129.965 793.000 ;
      LAYER met4 ;
        RECT 129.965 791.000 131.065 793.000 ;
        RECT 102.965 773.000 131.065 791.000 ;
        RECT 102.965 772.000 105.000 773.000 ;
        RECT 0.000 762.000 24.215 772.000 ;
        RECT 0.000 626.000 25.965 762.000 ;
        RECT 102.965 760.000 105.000 762.000 ;
      LAYER met4 ;
        RECT 105.000 760.000 129.965 773.000 ;
      LAYER met4 ;
        RECT 129.965 772.000 131.065 773.000 ;
        RECT 129.965 760.000 131.065 762.000 ;
        RECT 102.965 757.000 131.065 760.000 ;
        RECT 102.965 755.000 105.000 757.000 ;
      LAYER met4 ;
        RECT 105.000 755.000 129.965 757.000 ;
      LAYER met4 ;
        RECT 129.965 755.000 131.065 757.000 ;
        RECT 102.965 747.000 131.065 755.000 ;
        RECT 102.965 745.000 105.000 747.000 ;
      LAYER met4 ;
        RECT 105.000 745.000 129.965 747.000 ;
      LAYER met4 ;
        RECT 129.965 745.000 131.065 747.000 ;
        RECT 102.965 727.000 131.065 745.000 ;
        RECT 102.965 725.000 105.000 727.000 ;
      LAYER met4 ;
        RECT 105.000 725.000 129.965 727.000 ;
      LAYER met4 ;
        RECT 129.965 725.000 131.065 727.000 ;
        RECT 102.965 707.000 131.065 725.000 ;
        RECT 102.965 705.000 105.000 707.000 ;
      LAYER met4 ;
        RECT 105.000 705.000 129.965 707.000 ;
      LAYER met4 ;
        RECT 129.965 705.000 131.065 707.000 ;
        RECT 102.965 687.000 131.065 705.000 ;
        RECT 102.965 685.000 105.000 687.000 ;
      LAYER met4 ;
        RECT 105.000 685.000 129.965 687.000 ;
      LAYER met4 ;
        RECT 129.965 685.000 131.065 687.000 ;
        RECT 102.965 667.000 131.065 685.000 ;
        RECT 102.965 665.000 105.000 667.000 ;
      LAYER met4 ;
        RECT 105.000 665.000 129.965 667.000 ;
      LAYER met4 ;
        RECT 129.965 665.000 131.065 667.000 ;
        RECT 102.965 647.000 131.065 665.000 ;
        RECT 102.965 645.000 105.000 647.000 ;
      LAYER met4 ;
        RECT 105.000 645.000 129.965 647.000 ;
      LAYER met4 ;
        RECT 129.965 645.000 131.065 647.000 ;
        RECT 102.965 627.000 131.065 645.000 ;
        RECT 102.965 626.000 105.000 627.000 ;
        RECT 129.965 626.000 131.065 627.000 ;
      LAYER met4 ;
        RECT 0.000 624.730 24.215 626.000 ;
      LAYER met4 ;
        RECT 24.615 624.330 104.600 625.035 ;
        RECT 130.365 624.330 131.065 625.035 ;
      LAYER met4 ;
        RECT 131.465 624.730 135.915 909.270 ;
      LAYER met4 ;
        RECT 136.315 908.965 136.915 909.670 ;
        RECT 136.315 772.000 136.915 907.000 ;
        RECT 136.315 626.000 136.915 761.000 ;
        RECT 136.315 624.330 136.915 625.035 ;
      LAYER met4 ;
        RECT 137.315 624.730 141.765 909.270 ;
      LAYER met4 ;
        RECT 142.165 908.965 142.865 909.670 ;
        RECT 142.165 772.000 142.865 908.000 ;
      LAYER met4 ;
        RECT 143.265 767.000 143.595 910.610 ;
      LAYER met4 ;
        RECT 142.165 626.000 142.865 762.000 ;
        RECT 142.165 624.330 142.865 625.035 ;
        RECT 0.000 552.670 142.865 624.330 ;
      LAYER met4 ;
        RECT 0.000 551.000 24.215 552.270 ;
      LAYER met4 ;
        RECT 24.615 551.965 104.600 552.670 ;
        RECT 130.365 551.965 131.065 552.670 ;
        RECT 0.000 416.470 25.965 551.000 ;
        RECT 0.000 415.000 0.035 416.470 ;
      LAYER met4 ;
        RECT 0.035 415.000 24.215 416.470 ;
      LAYER met4 ;
        RECT 24.215 415.000 25.965 416.470 ;
        RECT 102.965 549.000 105.000 551.000 ;
        RECT 129.965 549.000 131.065 551.000 ;
        RECT 102.965 546.000 131.065 549.000 ;
        RECT 102.965 544.000 105.000 546.000 ;
      LAYER met4 ;
        RECT 105.000 544.000 129.965 546.000 ;
      LAYER met4 ;
        RECT 129.965 544.000 131.065 546.000 ;
        RECT 102.965 536.000 131.065 544.000 ;
        RECT 102.965 534.000 105.000 536.000 ;
      LAYER met4 ;
        RECT 105.000 534.000 129.965 536.000 ;
      LAYER met4 ;
        RECT 129.965 534.000 131.065 536.000 ;
        RECT 102.965 516.000 131.065 534.000 ;
        RECT 102.965 514.000 105.000 516.000 ;
      LAYER met4 ;
        RECT 105.000 514.000 129.965 516.000 ;
      LAYER met4 ;
        RECT 129.965 514.000 131.065 516.000 ;
        RECT 102.965 496.000 131.065 514.000 ;
        RECT 102.965 494.000 105.000 496.000 ;
      LAYER met4 ;
        RECT 105.000 494.000 129.965 496.000 ;
      LAYER met4 ;
        RECT 129.965 494.000 131.065 496.000 ;
        RECT 102.965 476.000 131.065 494.000 ;
        RECT 102.965 474.000 105.000 476.000 ;
      LAYER met4 ;
        RECT 105.000 474.000 129.965 476.000 ;
      LAYER met4 ;
        RECT 129.965 474.000 131.065 476.000 ;
        RECT 102.965 456.000 131.065 474.000 ;
        RECT 102.965 454.000 105.000 456.000 ;
      LAYER met4 ;
        RECT 105.000 454.000 129.965 456.000 ;
      LAYER met4 ;
        RECT 129.965 454.000 131.065 456.000 ;
        RECT 102.965 436.000 131.065 454.000 ;
        RECT 102.965 434.000 105.000 436.000 ;
      LAYER met4 ;
        RECT 105.000 434.000 129.965 436.000 ;
      LAYER met4 ;
        RECT 129.965 434.000 131.065 436.000 ;
        RECT 102.965 416.000 131.065 434.000 ;
        RECT 102.965 415.000 105.000 416.000 ;
      LAYER met4 ;
        RECT 0.000 413.730 24.215 415.000 ;
      LAYER met4 ;
        RECT 24.215 414.785 24.250 415.000 ;
        RECT 24.615 413.330 104.600 415.000 ;
      LAYER met4 ;
        RECT 105.000 413.730 129.965 416.000 ;
      LAYER met4 ;
        RECT 129.965 415.000 131.065 416.000 ;
        RECT 130.365 413.330 131.065 415.000 ;
      LAYER met4 ;
        RECT 131.465 413.730 135.915 552.270 ;
      LAYER met4 ;
        RECT 136.315 551.965 136.915 552.670 ;
        RECT 136.315 413.330 136.915 550.000 ;
      LAYER met4 ;
        RECT 137.315 413.730 141.765 552.270 ;
      LAYER met4 ;
        RECT 142.165 551.965 142.865 552.670 ;
        RECT 142.165 413.330 142.865 551.000 ;
        RECT 0.000 341.670 142.865 413.330 ;
      LAYER met4 ;
        RECT 0.000 340.000 24.215 341.270 ;
      LAYER met4 ;
        RECT 24.615 340.000 104.600 341.670 ;
        RECT 0.000 204.000 25.965 340.000 ;
        RECT 102.965 338.000 105.000 340.000 ;
      LAYER met4 ;
        RECT 105.000 338.000 129.965 341.270 ;
      LAYER met4 ;
        RECT 130.365 340.000 131.065 341.670 ;
        RECT 129.965 338.000 131.065 340.000 ;
        RECT 102.965 335.000 131.065 338.000 ;
        RECT 102.965 333.000 105.000 335.000 ;
      LAYER met4 ;
        RECT 105.000 333.000 129.965 335.000 ;
      LAYER met4 ;
        RECT 129.965 333.000 131.065 335.000 ;
        RECT 102.965 325.000 131.065 333.000 ;
        RECT 102.965 323.000 105.000 325.000 ;
      LAYER met4 ;
        RECT 105.000 323.000 129.965 325.000 ;
      LAYER met4 ;
        RECT 129.965 323.000 131.065 325.000 ;
        RECT 102.965 305.000 131.065 323.000 ;
        RECT 102.965 303.000 105.000 305.000 ;
      LAYER met4 ;
        RECT 105.000 303.000 129.965 305.000 ;
      LAYER met4 ;
        RECT 129.965 303.000 131.065 305.000 ;
        RECT 102.965 285.000 131.065 303.000 ;
        RECT 102.965 283.000 105.000 285.000 ;
      LAYER met4 ;
        RECT 105.000 283.000 129.965 285.000 ;
      LAYER met4 ;
        RECT 129.965 283.000 131.065 285.000 ;
        RECT 102.965 265.000 131.065 283.000 ;
        RECT 102.965 263.000 105.000 265.000 ;
      LAYER met4 ;
        RECT 105.000 263.000 129.965 265.000 ;
      LAYER met4 ;
        RECT 129.965 263.000 131.065 265.000 ;
        RECT 102.965 245.000 131.065 263.000 ;
        RECT 102.965 243.000 105.000 245.000 ;
      LAYER met4 ;
        RECT 105.000 243.000 129.965 245.000 ;
      LAYER met4 ;
        RECT 129.965 243.000 131.065 245.000 ;
        RECT 102.965 225.000 131.065 243.000 ;
        RECT 102.965 223.000 105.000 225.000 ;
      LAYER met4 ;
        RECT 105.000 223.000 129.965 225.000 ;
      LAYER met4 ;
        RECT 129.965 223.000 131.065 225.000 ;
        RECT 102.965 205.000 131.065 223.000 ;
        RECT 102.965 204.000 105.000 205.000 ;
      LAYER met4 ;
        RECT 0.000 202.730 24.215 204.000 ;
      LAYER met4 ;
        RECT 24.615 202.330 104.600 202.745 ;
        RECT 0.000 201.745 104.600 202.330 ;
      LAYER met4 ;
        RECT 105.000 202.145 129.965 205.000 ;
      LAYER met4 ;
        RECT 129.965 204.000 131.065 205.000 ;
        RECT 130.365 202.330 131.065 202.745 ;
      LAYER met4 ;
        RECT 131.465 202.730 135.915 341.270 ;
      LAYER met4 ;
        RECT 136.315 340.000 136.915 341.670 ;
        RECT 136.315 204.000 136.915 339.000 ;
        RECT 136.315 202.330 136.915 202.745 ;
      LAYER met4 ;
        RECT 137.315 202.730 141.765 341.270 ;
      LAYER met4 ;
        RECT 142.165 204.000 142.865 341.670 ;
        RECT 142.165 202.330 142.865 202.745 ;
        RECT 130.365 201.745 142.865 202.330 ;
        RECT 0.000 176.425 142.865 201.745 ;
      LAYER met4 ;
        RECT 143.265 176.825 143.595 762.000 ;
        RECT 143.895 177.090 146.875 944.440 ;
      LAYER met4 ;
        RECT 147.275 909.670 148.255 944.840 ;
      LAYER met4 ;
        RECT 147.175 908.000 148.355 909.270 ;
      LAYER met4 ;
        RECT 147.275 772.000 148.255 908.000 ;
        RECT 147.175 767.000 148.355 772.000 ;
        RECT 147.275 626.000 148.255 762.000 ;
      LAYER met4 ;
        RECT 147.175 624.730 148.355 626.000 ;
      LAYER met4 ;
        RECT 147.275 552.670 148.255 624.330 ;
      LAYER met4 ;
        RECT 147.175 551.000 148.355 552.270 ;
      LAYER met4 ;
        RECT 147.275 415.000 148.255 551.000 ;
      LAYER met4 ;
        RECT 147.175 413.730 148.355 415.000 ;
      LAYER met4 ;
        RECT 147.275 341.670 148.255 413.330 ;
      LAYER met4 ;
        RECT 147.175 340.000 148.355 341.270 ;
      LAYER met4 ;
        RECT 147.275 204.000 148.255 340.000 ;
      LAYER met4 ;
        RECT 147.175 182.445 148.355 204.000 ;
        RECT 148.655 183.125 151.635 960.145 ;
        RECT 151.935 955.090 152.265 1126.610 ;
      LAYER met4 ;
        RECT 152.665 1125.670 199.465 1127.010 ;
        RECT 152.665 1124.965 153.365 1125.670 ;
        RECT 152.665 986.330 153.365 986.970 ;
      LAYER met4 ;
        RECT 153.765 986.730 158.415 1125.270 ;
      LAYER met4 ;
        RECT 158.815 1124.965 159.415 1125.670 ;
        RECT 158.815 986.330 159.415 986.970 ;
      LAYER met4 ;
        RECT 159.815 986.730 163.265 1125.270 ;
      LAYER met4 ;
        RECT 163.665 1124.965 164.265 1125.670 ;
        RECT 163.665 986.330 164.265 986.970 ;
      LAYER met4 ;
        RECT 164.665 986.730 168.115 1125.270 ;
      LAYER met4 ;
        RECT 168.515 1124.965 169.115 1125.670 ;
        RECT 168.515 986.330 169.115 986.970 ;
      LAYER met4 ;
        RECT 169.515 986.730 174.165 1125.270 ;
      LAYER met4 ;
        RECT 174.565 1124.965 175.165 1125.670 ;
        RECT 180.615 1125.365 186.065 1125.670 ;
        RECT 174.565 986.330 175.165 986.970 ;
      LAYER met4 ;
        RECT 175.565 986.730 180.215 1125.270 ;
      LAYER met4 ;
        RECT 180.615 1124.965 181.215 1125.365 ;
        RECT 185.465 1124.965 186.065 1125.365 ;
      LAYER met4 ;
        RECT 181.615 986.970 185.065 1124.965 ;
      LAYER met4 ;
        RECT 180.615 986.570 181.215 986.970 ;
        RECT 185.465 986.570 186.065 986.970 ;
      LAYER met4 ;
        RECT 186.465 986.730 191.115 1125.270 ;
      LAYER met4 ;
        RECT 191.515 1124.965 192.115 1125.670 ;
        RECT 180.615 986.330 186.065 986.570 ;
        RECT 191.515 986.330 192.115 986.970 ;
      LAYER met4 ;
        RECT 192.515 986.730 197.965 1125.270 ;
      LAYER met4 ;
        RECT 198.365 1124.965 199.465 1125.670 ;
        RECT 3388.535 1029.330 3389.635 1030.035 ;
      LAYER met4 ;
        RECT 3390.035 1029.730 3395.485 1178.270 ;
      LAYER met4 ;
        RECT 3395.885 1178.030 3396.485 1178.670 ;
        RECT 3401.935 1178.430 3407.385 1178.670 ;
        RECT 3395.885 1029.330 3396.485 1030.035 ;
      LAYER met4 ;
        RECT 3396.885 1029.730 3401.535 1178.270 ;
      LAYER met4 ;
        RECT 3401.935 1178.030 3402.535 1178.430 ;
        RECT 3406.785 1178.030 3407.385 1178.430 ;
      LAYER met4 ;
        RECT 3402.935 1030.035 3406.385 1178.030 ;
      LAYER met4 ;
        RECT 3401.935 1029.635 3402.535 1030.035 ;
        RECT 3406.785 1029.635 3407.385 1030.035 ;
      LAYER met4 ;
        RECT 3407.785 1029.730 3412.435 1178.270 ;
      LAYER met4 ;
        RECT 3412.835 1178.030 3413.435 1178.670 ;
        RECT 3401.935 1029.330 3407.385 1029.635 ;
        RECT 3412.835 1029.330 3413.435 1030.035 ;
      LAYER met4 ;
        RECT 3413.835 1029.730 3418.485 1178.270 ;
      LAYER met4 ;
        RECT 3418.885 1178.030 3419.485 1178.670 ;
        RECT 3418.885 1029.330 3419.485 1030.035 ;
      LAYER met4 ;
        RECT 3419.885 1029.730 3423.335 1178.270 ;
      LAYER met4 ;
        RECT 3423.735 1178.030 3424.335 1178.670 ;
        RECT 3423.735 1029.330 3424.335 1030.035 ;
      LAYER met4 ;
        RECT 3424.735 1029.730 3428.185 1178.270 ;
      LAYER met4 ;
        RECT 3428.585 1178.030 3429.185 1178.670 ;
        RECT 3428.585 1029.330 3429.185 1030.035 ;
      LAYER met4 ;
        RECT 3429.585 1029.730 3434.235 1178.270 ;
      LAYER met4 ;
        RECT 3434.635 1178.030 3435.335 1178.670 ;
        RECT 3434.635 1029.330 3435.335 1030.035 ;
        RECT 3388.535 1027.990 3435.335 1029.330 ;
      LAYER met4 ;
        RECT 3435.735 1028.390 3436.065 1209.910 ;
        RECT 3436.365 1204.855 3439.345 1427.535 ;
      LAYER met4 ;
        RECT 3439.745 1403.670 3440.725 1427.935 ;
      LAYER met4 ;
        RECT 3439.645 1402.000 3440.825 1403.270 ;
      LAYER met4 ;
        RECT 3439.745 1257.000 3440.725 1402.000 ;
      LAYER met4 ;
        RECT 3439.645 1255.730 3440.825 1257.000 ;
      LAYER met4 ;
        RECT 3439.745 1220.160 3440.725 1255.330 ;
      LAYER met4 ;
        RECT 3441.125 1220.560 3444.105 1443.240 ;
      LAYER met4 ;
        RECT 3444.505 1435.310 3588.000 1443.640 ;
      LAYER met4 ;
        RECT 3444.405 1254.390 3444.735 1434.910 ;
      LAYER met4 ;
        RECT 3445.135 1403.670 3588.000 1435.310 ;
        RECT 3445.135 1403.030 3445.835 1403.670 ;
        RECT 3445.135 1257.000 3445.835 1402.000 ;
        RECT 3445.135 1255.330 3445.835 1256.035 ;
      LAYER met4 ;
        RECT 3446.235 1255.730 3450.685 1403.270 ;
      LAYER met4 ;
        RECT 3451.085 1403.030 3451.685 1403.670 ;
        RECT 3451.085 1257.000 3451.685 1402.000 ;
        RECT 3451.085 1255.330 3451.685 1256.035 ;
      LAYER met4 ;
        RECT 3452.085 1255.730 3456.535 1403.270 ;
      LAYER met4 ;
        RECT 3456.935 1403.030 3457.635 1403.670 ;
        RECT 3456.935 1401.000 3458.035 1402.000 ;
      LAYER met4 ;
        RECT 3458.035 1401.000 3483.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1403.030 3563.385 1403.670 ;
      LAYER met4 ;
        RECT 3563.785 1402.000 3588.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.000 1401.000 3485.035 1402.000 ;
        RECT 3456.935 1398.000 3485.035 1401.000 ;
        RECT 3456.935 1396.000 3458.035 1398.000 ;
      LAYER met4 ;
        RECT 3458.035 1396.000 3483.000 1398.000 ;
      LAYER met4 ;
        RECT 3483.000 1396.000 3485.035 1398.000 ;
        RECT 3456.935 1378.000 3485.035 1396.000 ;
        RECT 3456.935 1376.000 3458.035 1378.000 ;
      LAYER met4 ;
        RECT 3458.035 1376.000 3483.000 1378.000 ;
      LAYER met4 ;
        RECT 3483.000 1376.000 3485.035 1378.000 ;
        RECT 3456.935 1358.000 3485.035 1376.000 ;
        RECT 3456.935 1356.000 3458.035 1358.000 ;
      LAYER met4 ;
        RECT 3458.035 1356.000 3483.000 1358.000 ;
      LAYER met4 ;
        RECT 3483.000 1356.000 3485.035 1358.000 ;
        RECT 3456.935 1338.000 3485.035 1356.000 ;
        RECT 3456.935 1336.000 3458.035 1338.000 ;
      LAYER met4 ;
        RECT 3458.035 1336.000 3483.000 1338.000 ;
      LAYER met4 ;
        RECT 3483.000 1336.000 3485.035 1338.000 ;
        RECT 3456.935 1318.000 3485.035 1336.000 ;
        RECT 3456.935 1316.000 3458.035 1318.000 ;
      LAYER met4 ;
        RECT 3458.035 1316.000 3483.000 1318.000 ;
      LAYER met4 ;
        RECT 3483.000 1316.000 3485.035 1318.000 ;
        RECT 3456.935 1298.000 3485.035 1316.000 ;
        RECT 3456.935 1296.000 3458.035 1298.000 ;
      LAYER met4 ;
        RECT 3458.035 1296.000 3483.000 1298.000 ;
      LAYER met4 ;
        RECT 3483.000 1296.000 3485.035 1298.000 ;
        RECT 3456.935 1278.000 3485.035 1296.000 ;
        RECT 3456.935 1276.000 3458.035 1278.000 ;
      LAYER met4 ;
        RECT 3458.035 1276.000 3483.000 1278.000 ;
      LAYER met4 ;
        RECT 3483.000 1276.000 3485.035 1278.000 ;
        RECT 3456.935 1258.000 3485.035 1276.000 ;
        RECT 3456.935 1257.000 3458.035 1258.000 ;
        RECT 3456.935 1255.330 3457.635 1256.035 ;
      LAYER met4 ;
        RECT 3458.035 1255.730 3483.000 1258.000 ;
      LAYER met4 ;
        RECT 3483.000 1257.000 3485.035 1258.000 ;
        RECT 3562.035 1257.000 3588.000 1402.000 ;
        RECT 3483.400 1255.330 3563.385 1256.035 ;
      LAYER met4 ;
        RECT 3563.785 1255.730 3588.000 1257.000 ;
      LAYER met4 ;
        RECT 3445.135 1253.990 3588.000 1255.330 ;
        RECT 3444.505 1220.160 3588.000 1253.990 ;
        RECT 3439.745 1218.640 3588.000 1220.160 ;
        RECT 3439.745 1204.455 3440.725 1218.640 ;
        RECT 3436.465 1202.935 3440.725 1204.455 ;
        RECT 198.365 986.330 199.465 986.970 ;
        RECT 152.665 954.690 199.465 986.330 ;
        RECT 152.035 911.010 199.465 954.690 ;
        RECT 3388.535 984.310 3435.965 1027.990 ;
        RECT 3388.535 952.670 3435.335 984.310 ;
        RECT 3388.535 952.030 3389.635 952.670 ;
      LAYER met4 ;
        RECT 151.935 767.000 152.265 910.610 ;
      LAYER met4 ;
        RECT 152.665 909.670 199.465 911.010 ;
        RECT 152.665 908.965 153.365 909.670 ;
      LAYER met4 ;
        RECT 153.765 772.000 158.415 909.270 ;
      LAYER met4 ;
        RECT 158.815 908.965 159.415 909.670 ;
      LAYER met4 ;
        RECT 159.815 767.000 163.265 909.270 ;
      LAYER met4 ;
        RECT 163.665 908.965 164.265 909.670 ;
        RECT 148.755 182.045 151.535 182.725 ;
        RECT 147.275 180.025 151.535 182.045 ;
      LAYER met4 ;
        RECT 151.935 180.425 152.265 762.000 ;
      LAYER met4 ;
        RECT 152.665 624.330 153.365 625.035 ;
      LAYER met4 ;
        RECT 153.765 624.730 158.415 767.000 ;
      LAYER met4 ;
        RECT 158.815 624.330 159.415 625.035 ;
      LAYER met4 ;
        RECT 159.815 624.730 163.265 762.000 ;
      LAYER met4 ;
        RECT 163.665 624.330 164.265 625.035 ;
      LAYER met4 ;
        RECT 164.665 624.730 168.115 909.270 ;
      LAYER met4 ;
        RECT 168.515 908.965 169.115 909.670 ;
        RECT 168.515 624.330 169.115 625.035 ;
      LAYER met4 ;
        RECT 169.515 624.730 174.165 909.270 ;
      LAYER met4 ;
        RECT 174.565 908.965 175.165 909.670 ;
        RECT 180.615 909.365 186.065 909.670 ;
        RECT 180.615 908.965 181.215 909.365 ;
        RECT 185.465 908.965 186.065 909.365 ;
      LAYER met4 ;
        RECT 181.615 767.000 185.065 908.965 ;
        RECT 186.465 772.000 191.115 909.270 ;
      LAYER met4 ;
        RECT 191.515 908.965 192.115 909.670 ;
      LAYER met4 ;
        RECT 181.615 625.035 185.065 762.000 ;
      LAYER met4 ;
        RECT 174.565 624.330 175.165 625.035 ;
        RECT 180.615 624.635 181.215 625.035 ;
        RECT 185.465 624.635 186.065 625.035 ;
      LAYER met4 ;
        RECT 186.465 624.730 191.115 767.000 ;
      LAYER met4 ;
        RECT 180.615 624.330 186.065 624.635 ;
        RECT 191.515 624.330 192.115 625.035 ;
      LAYER met4 ;
        RECT 192.515 624.730 197.965 909.270 ;
      LAYER met4 ;
        RECT 198.365 908.965 199.465 909.670 ;
        RECT 3388.535 804.330 3389.635 805.035 ;
      LAYER met4 ;
        RECT 3390.035 804.730 3395.485 952.270 ;
      LAYER met4 ;
        RECT 3395.885 952.030 3396.485 952.670 ;
        RECT 3401.935 952.430 3407.385 952.670 ;
        RECT 3395.885 804.330 3396.485 805.035 ;
      LAYER met4 ;
        RECT 3396.885 804.730 3401.535 952.270 ;
      LAYER met4 ;
        RECT 3401.935 952.030 3402.535 952.430 ;
        RECT 3406.785 952.030 3407.385 952.430 ;
      LAYER met4 ;
        RECT 3402.935 805.035 3406.385 952.030 ;
      LAYER met4 ;
        RECT 3401.935 804.635 3402.535 805.035 ;
        RECT 3406.785 804.635 3407.385 805.035 ;
      LAYER met4 ;
        RECT 3407.785 804.730 3412.435 952.270 ;
      LAYER met4 ;
        RECT 3412.835 952.030 3413.435 952.670 ;
        RECT 3401.935 804.330 3407.385 804.635 ;
        RECT 3412.835 804.330 3413.435 805.035 ;
      LAYER met4 ;
        RECT 3413.835 804.730 3418.485 952.270 ;
      LAYER met4 ;
        RECT 3418.885 952.030 3419.485 952.670 ;
        RECT 3418.885 804.330 3419.485 805.035 ;
      LAYER met4 ;
        RECT 3419.885 804.730 3423.335 952.270 ;
      LAYER met4 ;
        RECT 3423.735 952.030 3424.335 952.670 ;
        RECT 3423.735 804.330 3424.335 805.035 ;
      LAYER met4 ;
        RECT 3424.735 804.730 3428.185 952.270 ;
      LAYER met4 ;
        RECT 3428.585 952.030 3429.185 952.670 ;
        RECT 3428.585 804.330 3429.185 805.035 ;
      LAYER met4 ;
        RECT 3429.585 804.730 3434.235 952.270 ;
      LAYER met4 ;
        RECT 3434.635 952.030 3435.335 952.670 ;
        RECT 3434.635 804.330 3435.335 805.035 ;
        RECT 3388.535 802.990 3435.335 804.330 ;
      LAYER met4 ;
        RECT 3435.735 803.390 3436.065 983.910 ;
        RECT 3436.365 978.855 3439.345 1202.535 ;
      LAYER met4 ;
        RECT 3439.745 1178.670 3440.725 1202.935 ;
      LAYER met4 ;
        RECT 3439.645 1177.000 3440.825 1178.270 ;
      LAYER met4 ;
        RECT 3439.745 1031.000 3440.725 1177.000 ;
      LAYER met4 ;
        RECT 3439.645 1029.730 3440.825 1031.000 ;
      LAYER met4 ;
        RECT 3439.745 994.160 3440.725 1029.330 ;
      LAYER met4 ;
        RECT 3441.125 994.560 3444.105 1218.240 ;
      LAYER met4 ;
        RECT 3444.505 1210.310 3588.000 1218.640 ;
      LAYER met4 ;
        RECT 3444.405 1028.390 3444.735 1209.910 ;
      LAYER met4 ;
        RECT 3445.135 1178.670 3588.000 1210.310 ;
        RECT 3445.135 1178.030 3445.835 1178.670 ;
        RECT 3445.135 1031.000 3445.835 1177.000 ;
        RECT 3445.135 1029.330 3445.835 1030.035 ;
      LAYER met4 ;
        RECT 3446.235 1029.730 3450.685 1178.270 ;
      LAYER met4 ;
        RECT 3451.085 1178.030 3451.685 1178.670 ;
        RECT 3451.085 1031.000 3451.685 1176.000 ;
        RECT 3451.085 1029.330 3451.685 1030.035 ;
      LAYER met4 ;
        RECT 3452.085 1029.730 3456.535 1178.270 ;
      LAYER met4 ;
        RECT 3456.935 1178.030 3457.635 1178.670 ;
        RECT 3456.935 1175.000 3458.035 1177.000 ;
      LAYER met4 ;
        RECT 3458.035 1175.000 3483.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1178.030 3563.385 1178.670 ;
      LAYER met4 ;
        RECT 3563.785 1177.000 3588.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.000 1175.000 3485.035 1177.000 ;
        RECT 3456.935 1172.000 3485.035 1175.000 ;
        RECT 3456.935 1170.000 3458.035 1172.000 ;
      LAYER met4 ;
        RECT 3458.035 1170.000 3483.000 1172.000 ;
      LAYER met4 ;
        RECT 3483.000 1170.000 3485.035 1172.000 ;
        RECT 3456.935 1152.000 3485.035 1170.000 ;
        RECT 3456.935 1150.000 3458.035 1152.000 ;
      LAYER met4 ;
        RECT 3458.035 1150.000 3483.000 1152.000 ;
      LAYER met4 ;
        RECT 3483.000 1150.000 3485.035 1152.000 ;
        RECT 3456.935 1132.000 3485.035 1150.000 ;
        RECT 3456.935 1130.000 3458.035 1132.000 ;
      LAYER met4 ;
        RECT 3458.035 1130.000 3483.000 1132.000 ;
      LAYER met4 ;
        RECT 3483.000 1130.000 3485.035 1132.000 ;
        RECT 3456.935 1112.000 3485.035 1130.000 ;
        RECT 3456.935 1110.000 3458.035 1112.000 ;
      LAYER met4 ;
        RECT 3458.035 1110.000 3483.000 1112.000 ;
      LAYER met4 ;
        RECT 3483.000 1110.000 3485.035 1112.000 ;
        RECT 3456.935 1092.000 3485.035 1110.000 ;
        RECT 3456.935 1090.000 3458.035 1092.000 ;
      LAYER met4 ;
        RECT 3458.035 1090.000 3483.000 1092.000 ;
      LAYER met4 ;
        RECT 3483.000 1090.000 3485.035 1092.000 ;
        RECT 3456.935 1072.000 3485.035 1090.000 ;
        RECT 3456.935 1070.000 3458.035 1072.000 ;
      LAYER met4 ;
        RECT 3458.035 1070.000 3483.000 1072.000 ;
      LAYER met4 ;
        RECT 3483.000 1070.000 3485.035 1072.000 ;
        RECT 3456.935 1052.000 3485.035 1070.000 ;
        RECT 3456.935 1050.000 3458.035 1052.000 ;
      LAYER met4 ;
        RECT 3458.035 1050.000 3483.000 1052.000 ;
      LAYER met4 ;
        RECT 3483.000 1050.000 3485.035 1052.000 ;
        RECT 3456.935 1032.000 3485.035 1050.000 ;
        RECT 3456.935 1031.000 3458.035 1032.000 ;
        RECT 3456.935 1029.330 3457.635 1030.035 ;
      LAYER met4 ;
        RECT 3458.035 1029.730 3483.000 1032.000 ;
      LAYER met4 ;
        RECT 3483.000 1031.000 3485.035 1032.000 ;
        RECT 3562.035 1031.000 3588.000 1177.000 ;
        RECT 3483.400 1029.330 3563.385 1030.035 ;
      LAYER met4 ;
        RECT 3563.785 1029.730 3588.000 1031.000 ;
      LAYER met4 ;
        RECT 3445.135 1027.990 3588.000 1029.330 ;
        RECT 3444.505 994.160 3588.000 1027.990 ;
        RECT 3439.745 992.640 3588.000 994.160 ;
        RECT 3439.745 978.455 3440.725 992.640 ;
        RECT 3436.465 976.935 3440.725 978.455 ;
        RECT 3388.535 759.310 3435.965 802.990 ;
        RECT 3388.535 727.670 3435.335 759.310 ;
        RECT 3388.535 727.030 3389.635 727.670 ;
        RECT 152.665 552.670 197.965 624.330 ;
        RECT 3388.535 578.330 3389.635 579.035 ;
      LAYER met4 ;
        RECT 3390.035 578.730 3395.485 727.270 ;
      LAYER met4 ;
        RECT 3395.885 727.030 3396.485 727.670 ;
        RECT 3401.935 727.430 3407.385 727.670 ;
        RECT 3395.885 578.330 3396.485 579.035 ;
      LAYER met4 ;
        RECT 3396.885 578.730 3401.535 727.270 ;
      LAYER met4 ;
        RECT 3401.935 727.030 3402.535 727.430 ;
        RECT 3406.785 727.030 3407.385 727.430 ;
      LAYER met4 ;
        RECT 3402.935 579.035 3406.385 727.030 ;
      LAYER met4 ;
        RECT 3401.935 578.635 3402.535 579.035 ;
        RECT 3406.785 578.635 3407.385 579.035 ;
      LAYER met4 ;
        RECT 3407.785 578.730 3412.435 727.270 ;
      LAYER met4 ;
        RECT 3412.835 727.030 3413.435 727.670 ;
        RECT 3401.935 578.330 3407.385 578.635 ;
        RECT 3412.835 578.330 3413.435 579.035 ;
      LAYER met4 ;
        RECT 3413.835 578.730 3418.485 727.270 ;
      LAYER met4 ;
        RECT 3418.885 727.030 3419.485 727.670 ;
        RECT 3418.885 578.330 3419.485 579.035 ;
      LAYER met4 ;
        RECT 3419.885 578.730 3423.335 727.270 ;
      LAYER met4 ;
        RECT 3423.735 727.030 3424.335 727.670 ;
        RECT 3423.735 578.330 3424.335 579.035 ;
      LAYER met4 ;
        RECT 3424.735 578.730 3428.185 727.270 ;
      LAYER met4 ;
        RECT 3428.585 727.030 3429.185 727.670 ;
        RECT 3428.585 578.330 3429.185 579.035 ;
      LAYER met4 ;
        RECT 3429.585 578.730 3434.235 727.270 ;
      LAYER met4 ;
        RECT 3434.635 727.030 3435.335 727.670 ;
        RECT 3434.635 578.330 3435.335 579.035 ;
        RECT 3388.535 576.990 3435.335 578.330 ;
      LAYER met4 ;
        RECT 3435.735 577.390 3436.065 758.910 ;
        RECT 3436.365 753.855 3439.345 976.535 ;
      LAYER met4 ;
        RECT 3439.745 952.670 3440.725 976.935 ;
      LAYER met4 ;
        RECT 3439.645 951.000 3440.825 952.270 ;
      LAYER met4 ;
        RECT 3439.745 806.000 3440.725 951.000 ;
      LAYER met4 ;
        RECT 3439.645 804.730 3440.825 806.000 ;
      LAYER met4 ;
        RECT 3439.745 769.160 3440.725 804.330 ;
      LAYER met4 ;
        RECT 3441.125 769.560 3444.105 992.240 ;
      LAYER met4 ;
        RECT 3444.505 984.310 3588.000 992.640 ;
      LAYER met4 ;
        RECT 3444.405 803.390 3444.735 983.910 ;
      LAYER met4 ;
        RECT 3445.135 952.670 3588.000 984.310 ;
        RECT 3445.135 952.030 3445.835 952.670 ;
        RECT 3445.135 806.000 3445.835 951.000 ;
        RECT 3445.135 804.330 3445.835 805.035 ;
      LAYER met4 ;
        RECT 3446.235 804.730 3450.685 952.270 ;
      LAYER met4 ;
        RECT 3451.085 952.030 3451.685 952.670 ;
        RECT 3451.085 806.000 3451.685 951.000 ;
        RECT 3451.085 804.330 3451.685 805.035 ;
      LAYER met4 ;
        RECT 3452.085 804.730 3456.535 952.270 ;
      LAYER met4 ;
        RECT 3456.935 952.030 3457.635 952.670 ;
        RECT 3456.935 950.000 3458.035 951.000 ;
      LAYER met4 ;
        RECT 3458.035 950.000 3483.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 952.030 3563.385 952.670 ;
      LAYER met4 ;
        RECT 3563.785 951.000 3588.000 952.270 ;
      LAYER met4 ;
        RECT 3483.000 950.000 3485.035 951.000 ;
        RECT 3456.935 947.000 3485.035 950.000 ;
        RECT 3456.935 945.000 3458.035 947.000 ;
      LAYER met4 ;
        RECT 3458.035 945.000 3483.000 947.000 ;
      LAYER met4 ;
        RECT 3483.000 945.000 3485.035 947.000 ;
        RECT 3456.935 927.000 3485.035 945.000 ;
        RECT 3456.935 925.000 3458.035 927.000 ;
      LAYER met4 ;
        RECT 3458.035 925.000 3483.000 927.000 ;
      LAYER met4 ;
        RECT 3483.000 925.000 3485.035 927.000 ;
        RECT 3456.935 907.000 3485.035 925.000 ;
        RECT 3456.935 905.000 3458.035 907.000 ;
      LAYER met4 ;
        RECT 3458.035 905.000 3483.000 907.000 ;
      LAYER met4 ;
        RECT 3483.000 905.000 3485.035 907.000 ;
        RECT 3456.935 887.000 3485.035 905.000 ;
        RECT 3456.935 885.000 3458.035 887.000 ;
      LAYER met4 ;
        RECT 3458.035 885.000 3483.000 887.000 ;
      LAYER met4 ;
        RECT 3483.000 885.000 3485.035 887.000 ;
        RECT 3456.935 867.000 3485.035 885.000 ;
        RECT 3456.935 865.000 3458.035 867.000 ;
      LAYER met4 ;
        RECT 3458.035 865.000 3483.000 867.000 ;
      LAYER met4 ;
        RECT 3483.000 865.000 3485.035 867.000 ;
        RECT 3456.935 847.000 3485.035 865.000 ;
        RECT 3456.935 845.000 3458.035 847.000 ;
      LAYER met4 ;
        RECT 3458.035 845.000 3483.000 847.000 ;
      LAYER met4 ;
        RECT 3483.000 845.000 3485.035 847.000 ;
        RECT 3456.935 827.000 3485.035 845.000 ;
        RECT 3456.935 825.000 3458.035 827.000 ;
      LAYER met4 ;
        RECT 3458.035 825.000 3483.000 827.000 ;
      LAYER met4 ;
        RECT 3483.000 825.000 3485.035 827.000 ;
        RECT 3456.935 807.000 3485.035 825.000 ;
        RECT 3456.935 806.000 3458.035 807.000 ;
        RECT 3456.935 804.330 3457.635 805.035 ;
      LAYER met4 ;
        RECT 3458.035 804.730 3483.000 807.000 ;
      LAYER met4 ;
        RECT 3483.000 806.000 3485.035 807.000 ;
        RECT 3562.035 806.000 3588.000 951.000 ;
        RECT 3483.400 804.330 3563.385 805.035 ;
      LAYER met4 ;
        RECT 3563.785 804.730 3588.000 806.000 ;
      LAYER met4 ;
        RECT 3445.135 802.990 3588.000 804.330 ;
        RECT 3444.505 769.160 3588.000 802.990 ;
        RECT 3439.745 767.640 3588.000 769.160 ;
        RECT 3439.745 753.455 3440.725 767.640 ;
        RECT 3436.465 751.935 3440.725 753.455 ;
        RECT 152.665 551.965 153.365 552.670 ;
        RECT 152.665 413.330 153.365 415.000 ;
      LAYER met4 ;
        RECT 153.765 413.730 158.415 552.270 ;
      LAYER met4 ;
        RECT 158.815 551.965 159.415 552.670 ;
        RECT 158.815 413.330 159.415 415.000 ;
      LAYER met4 ;
        RECT 159.815 413.730 163.265 552.270 ;
      LAYER met4 ;
        RECT 163.665 551.965 164.265 552.670 ;
        RECT 163.665 413.330 164.265 415.000 ;
      LAYER met4 ;
        RECT 164.665 413.730 168.115 552.270 ;
      LAYER met4 ;
        RECT 168.515 551.965 169.115 552.670 ;
        RECT 168.515 413.330 169.115 415.000 ;
      LAYER met4 ;
        RECT 169.515 413.730 174.165 552.270 ;
      LAYER met4 ;
        RECT 174.565 551.965 175.165 552.670 ;
        RECT 180.615 552.365 186.065 552.670 ;
        RECT 180.615 551.965 181.215 552.365 ;
        RECT 185.465 551.965 186.065 552.365 ;
        RECT 191.515 551.965 192.115 552.670 ;
        RECT 174.165 414.935 174.200 425.935 ;
        RECT 174.565 413.330 175.165 415.000 ;
        RECT 180.615 413.635 181.215 415.000 ;
      LAYER met4 ;
        RECT 181.615 414.035 185.065 551.965 ;
      LAYER met4 ;
        RECT 185.465 413.635 186.065 415.000 ;
        RECT 180.615 413.330 186.065 413.635 ;
        RECT 191.515 413.330 192.115 415.000 ;
      LAYER met4 ;
        RECT 192.515 413.730 197.965 552.270 ;
      LAYER met4 ;
        RECT 3388.535 533.310 3435.965 576.990 ;
        RECT 3388.535 501.670 3435.335 533.310 ;
        RECT 3388.535 501.030 3389.635 501.670 ;
        RECT 152.665 341.670 197.965 413.330 ;
        RECT 152.665 340.000 153.365 341.670 ;
        RECT 152.665 202.330 153.365 202.745 ;
      LAYER met4 ;
        RECT 153.765 202.730 158.415 341.270 ;
      LAYER met4 ;
        RECT 158.415 329.025 158.450 340.070 ;
        RECT 158.815 340.000 159.415 341.670 ;
        RECT 158.815 202.330 159.415 202.745 ;
      LAYER met4 ;
        RECT 159.815 202.730 163.265 341.270 ;
      LAYER met4 ;
        RECT 163.665 340.000 164.265 341.670 ;
        RECT 163.665 202.330 164.265 202.745 ;
      LAYER met4 ;
        RECT 164.665 202.730 168.115 341.270 ;
      LAYER met4 ;
        RECT 168.515 340.000 169.115 341.670 ;
        RECT 168.515 202.330 169.115 202.745 ;
      LAYER met4 ;
        RECT 169.515 202.730 174.165 341.270 ;
      LAYER met4 ;
        RECT 174.565 340.000 175.165 341.670 ;
        RECT 180.615 341.365 186.065 341.670 ;
        RECT 174.565 202.330 175.165 202.745 ;
      LAYER met4 ;
        RECT 175.565 202.730 180.215 341.270 ;
      LAYER met4 ;
        RECT 180.615 340.000 181.215 341.365 ;
      LAYER met4 ;
        RECT 181.615 202.745 185.065 340.965 ;
      LAYER met4 ;
        RECT 185.465 340.000 186.065 341.365 ;
        RECT 191.515 340.000 192.115 341.670 ;
        RECT 180.615 202.345 181.215 202.745 ;
        RECT 185.465 202.345 186.065 202.745 ;
        RECT 180.615 202.330 186.065 202.345 ;
        RECT 191.515 202.330 192.115 202.745 ;
      LAYER met4 ;
        RECT 192.515 202.730 197.965 341.270 ;
      LAYER met4 ;
        RECT 198.365 202.330 200.000 202.745 ;
        RECT 152.665 198.365 200.000 202.330 ;
        RECT 3385.255 199.600 3389.635 200.000 ;
        POLYGON 3390.035 200.000 3390.035 199.600 3389.635 199.600 ;
        RECT 933.030 198.365 1011.035 199.465 ;
        RECT 1476.030 198.365 1554.035 199.465 ;
        RECT 1750.030 198.365 1828.035 199.465 ;
        RECT 2024.030 198.365 2102.035 199.465 ;
        RECT 2298.030 198.365 2376.035 199.465 ;
        RECT 2572.030 198.365 2650.035 199.465 ;
        RECT 3385.255 198.365 3390.035 199.600 ;
        RECT 152.665 192.115 197.250 198.365 ;
        RECT 197.965 197.965 199.600 198.365 ;
        POLYGON 199.600 198.365 200.000 197.965 199.600 197.965 ;
      LAYER met4 ;
        RECT 197.650 192.515 395.270 197.965 ;
      LAYER met4 ;
        RECT 395.670 192.115 467.330 197.965 ;
      LAYER met4 ;
        RECT 467.730 192.515 664.270 197.965 ;
      LAYER met4 ;
        RECT 664.670 192.115 736.330 197.965 ;
      LAYER met4 ;
        RECT 736.730 192.515 933.270 197.965 ;
      LAYER met4 ;
        RECT 933.670 192.115 1010.330 198.365 ;
      LAYER met4 ;
        RECT 1010.730 192.515 1207.270 197.965 ;
      LAYER met4 ;
        RECT 1207.670 192.115 1279.330 197.965 ;
      LAYER met4 ;
        RECT 1279.730 192.515 1476.270 197.965 ;
      LAYER met4 ;
        RECT 1476.670 192.115 1553.330 198.365 ;
      LAYER met4 ;
        RECT 1553.730 192.515 1750.270 197.965 ;
      LAYER met4 ;
        RECT 1750.670 192.115 1827.330 198.365 ;
      LAYER met4 ;
        RECT 1827.730 192.515 2024.270 197.965 ;
      LAYER met4 ;
        RECT 2024.670 192.115 2101.330 198.365 ;
      LAYER met4 ;
        RECT 2101.730 192.515 2298.270 197.965 ;
      LAYER met4 ;
        RECT 2298.670 192.115 2375.330 198.365 ;
      LAYER met4 ;
        RECT 2375.730 192.515 2572.270 197.965 ;
      LAYER met4 ;
        RECT 2572.670 192.115 2649.330 198.365 ;
        RECT 3385.670 197.965 3390.035 198.365 ;
      LAYER met4 ;
        RECT 2649.730 192.515 2846.270 197.965 ;
      LAYER met4 ;
        RECT 2846.670 192.115 2918.330 197.965 ;
      LAYER met4 ;
        RECT 2918.730 192.515 3115.270 197.965 ;
      LAYER met4 ;
        RECT 3115.670 192.115 3187.330 197.965 ;
      LAYER met4 ;
        RECT 3187.730 192.515 3385.270 197.965 ;
      LAYER met4 ;
        RECT 3385.670 197.250 3389.635 197.965 ;
      LAYER met4 ;
        RECT 3390.035 197.650 3395.485 501.270 ;
      LAYER met4 ;
        RECT 3395.885 501.030 3396.485 501.670 ;
        RECT 3401.935 501.430 3407.385 501.670 ;
      LAYER met4 ;
        RECT 3396.885 355.000 3401.535 501.270 ;
      LAYER met4 ;
        RECT 3401.935 501.030 3402.535 501.430 ;
        RECT 3406.785 501.030 3407.385 501.430 ;
      LAYER met4 ;
        RECT 3402.935 350.000 3406.385 501.030 ;
      LAYER met4 ;
        RECT 3395.885 197.250 3396.485 200.000 ;
        RECT 3385.670 195.815 3396.485 197.250 ;
      LAYER met4 ;
        RECT 3396.885 196.215 3401.535 350.000 ;
      LAYER met4 ;
        RECT 3401.935 198.130 3402.535 200.000 ;
      LAYER met4 ;
        RECT 3402.935 198.530 3406.385 345.000 ;
      LAYER met4 ;
        RECT 3406.785 198.130 3407.385 200.000 ;
      LAYER met4 ;
        RECT 3407.785 198.475 3412.435 501.270 ;
      LAYER met4 ;
        RECT 3412.835 501.030 3413.435 501.670 ;
        RECT 3401.935 198.075 3407.385 198.130 ;
        RECT 3412.835 198.075 3413.435 200.000 ;
      LAYER met4 ;
        RECT 3413.835 198.400 3418.485 501.270 ;
      LAYER met4 ;
        RECT 3418.885 501.030 3419.485 501.670 ;
        RECT 3401.935 198.000 3413.435 198.075 ;
        RECT 3418.885 198.215 3419.485 200.000 ;
      LAYER met4 ;
        RECT 3419.885 198.615 3423.335 501.270 ;
      LAYER met4 ;
        RECT 3423.735 501.030 3424.335 501.670 ;
      LAYER met4 ;
        RECT 3424.735 350.000 3428.185 501.270 ;
      LAYER met4 ;
        RECT 3428.585 501.030 3429.185 501.670 ;
      LAYER met4 ;
        RECT 3429.585 355.000 3434.235 501.270 ;
      LAYER met4 ;
        RECT 3434.635 501.030 3435.335 501.670 ;
      LAYER met4 ;
        RECT 3435.735 350.000 3436.065 532.910 ;
        RECT 3436.365 527.855 3439.345 751.535 ;
      LAYER met4 ;
        RECT 3439.745 727.670 3440.725 751.935 ;
      LAYER met4 ;
        RECT 3439.645 726.000 3440.825 727.270 ;
      LAYER met4 ;
        RECT 3439.745 580.000 3440.725 726.000 ;
      LAYER met4 ;
        RECT 3439.645 578.730 3440.825 580.000 ;
      LAYER met4 ;
        RECT 3439.745 543.160 3440.725 578.330 ;
      LAYER met4 ;
        RECT 3441.125 543.560 3444.105 767.240 ;
      LAYER met4 ;
        RECT 3444.505 759.310 3588.000 767.640 ;
      LAYER met4 ;
        RECT 3444.405 577.390 3444.735 758.910 ;
      LAYER met4 ;
        RECT 3445.135 727.670 3588.000 759.310 ;
        RECT 3445.135 727.030 3445.835 727.670 ;
        RECT 3445.135 580.000 3445.835 726.000 ;
        RECT 3445.135 578.330 3445.835 579.035 ;
      LAYER met4 ;
        RECT 3446.235 578.730 3450.685 727.270 ;
      LAYER met4 ;
        RECT 3451.085 727.030 3451.685 727.670 ;
        RECT 3451.085 580.000 3451.685 725.000 ;
        RECT 3451.085 578.330 3451.685 579.035 ;
      LAYER met4 ;
        RECT 3452.085 578.730 3456.535 727.270 ;
      LAYER met4 ;
        RECT 3456.935 727.030 3457.635 727.670 ;
        RECT 3456.935 724.000 3458.035 726.000 ;
      LAYER met4 ;
        RECT 3458.035 724.000 3483.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 727.030 3563.385 727.670 ;
      LAYER met4 ;
        RECT 3563.785 726.000 3588.000 727.270 ;
      LAYER met4 ;
        RECT 3483.000 724.000 3485.035 726.000 ;
        RECT 3456.935 721.000 3485.035 724.000 ;
        RECT 3456.935 719.000 3458.035 721.000 ;
      LAYER met4 ;
        RECT 3458.035 719.000 3483.000 721.000 ;
      LAYER met4 ;
        RECT 3483.000 719.000 3485.035 721.000 ;
        RECT 3456.935 701.000 3485.035 719.000 ;
        RECT 3456.935 699.000 3458.035 701.000 ;
      LAYER met4 ;
        RECT 3458.035 699.000 3483.000 701.000 ;
      LAYER met4 ;
        RECT 3483.000 699.000 3485.035 701.000 ;
        RECT 3456.935 681.000 3485.035 699.000 ;
        RECT 3456.935 679.000 3458.035 681.000 ;
      LAYER met4 ;
        RECT 3458.035 679.000 3483.000 681.000 ;
      LAYER met4 ;
        RECT 3483.000 679.000 3485.035 681.000 ;
        RECT 3456.935 661.000 3485.035 679.000 ;
        RECT 3456.935 659.000 3458.035 661.000 ;
      LAYER met4 ;
        RECT 3458.035 659.000 3483.000 661.000 ;
      LAYER met4 ;
        RECT 3483.000 659.000 3485.035 661.000 ;
        RECT 3456.935 641.000 3485.035 659.000 ;
        RECT 3456.935 639.000 3458.035 641.000 ;
      LAYER met4 ;
        RECT 3458.035 639.000 3483.000 641.000 ;
      LAYER met4 ;
        RECT 3483.000 639.000 3485.035 641.000 ;
        RECT 3456.935 621.000 3485.035 639.000 ;
        RECT 3456.935 619.000 3458.035 621.000 ;
      LAYER met4 ;
        RECT 3458.035 619.000 3483.000 621.000 ;
      LAYER met4 ;
        RECT 3483.000 619.000 3485.035 621.000 ;
        RECT 3456.935 601.000 3485.035 619.000 ;
        RECT 3456.935 599.000 3458.035 601.000 ;
      LAYER met4 ;
        RECT 3458.035 599.000 3483.000 601.000 ;
      LAYER met4 ;
        RECT 3483.000 599.000 3485.035 601.000 ;
        RECT 3456.935 581.000 3485.035 599.000 ;
        RECT 3456.935 580.000 3458.035 581.000 ;
        RECT 3456.935 578.330 3457.635 579.035 ;
      LAYER met4 ;
        RECT 3458.035 578.730 3483.000 581.000 ;
      LAYER met4 ;
        RECT 3483.000 580.000 3485.035 581.000 ;
        RECT 3562.035 580.000 3588.000 726.000 ;
        RECT 3483.400 578.330 3563.385 579.035 ;
      LAYER met4 ;
        RECT 3563.785 578.730 3588.000 580.000 ;
      LAYER met4 ;
        RECT 3445.135 576.990 3588.000 578.330 ;
        RECT 3444.505 543.160 3588.000 576.990 ;
        RECT 3439.745 541.640 3588.000 543.160 ;
        RECT 3439.745 527.455 3440.725 541.640 ;
        RECT 3436.465 525.935 3440.725 527.455 ;
        RECT 3423.735 198.265 3424.335 200.000 ;
      LAYER met4 ;
        RECT 3424.735 198.665 3428.185 345.000 ;
      LAYER met4 ;
        RECT 3428.585 198.265 3429.185 200.000 ;
      LAYER met4 ;
        RECT 3429.585 198.525 3434.235 350.000 ;
      LAYER met4 ;
        RECT 3423.735 198.215 3429.185 198.265 ;
        RECT 3418.885 198.125 3429.185 198.215 ;
        RECT 3434.635 198.125 3435.335 200.000 ;
        RECT 3418.885 198.000 3435.335 198.125 ;
        RECT 3401.935 195.815 3435.335 198.000 ;
        RECT 3385.670 192.115 3435.335 195.815 ;
        RECT 152.665 191.515 200.000 192.115 ;
        RECT 394.965 191.515 468.035 192.115 ;
        RECT 663.965 191.515 737.035 192.115 ;
        RECT 933.030 191.515 1011.035 192.115 ;
        RECT 1206.000 191.515 1281.000 192.115 ;
        RECT 1476.030 191.515 1554.035 192.115 ;
        RECT 1750.030 191.515 1828.035 192.115 ;
        RECT 2024.030 191.515 2102.035 192.115 ;
        RECT 2298.030 191.515 2376.035 192.115 ;
        RECT 2572.030 191.515 2650.035 192.115 ;
        RECT 2845.965 191.515 2919.035 192.115 ;
        RECT 3114.965 191.515 3188.035 192.115 ;
        RECT 3385.255 191.515 3435.335 192.115 ;
        RECT 152.665 186.065 195.815 191.515 ;
      LAYER met4 ;
        RECT 196.215 186.465 395.270 191.115 ;
      LAYER met4 ;
        RECT 395.670 186.065 467.330 191.515 ;
      LAYER met4 ;
        RECT 467.730 186.465 664.270 191.115 ;
      LAYER met4 ;
        RECT 664.670 186.065 736.330 191.515 ;
      LAYER met4 ;
        RECT 736.730 186.465 933.270 191.115 ;
      LAYER met4 ;
        RECT 933.670 186.065 1010.330 191.515 ;
      LAYER met4 ;
        RECT 1010.730 186.465 1207.270 191.115 ;
      LAYER met4 ;
        RECT 1207.670 186.065 1279.330 191.515 ;
      LAYER met4 ;
        RECT 1279.730 186.465 1476.270 191.115 ;
      LAYER met4 ;
        RECT 1476.670 186.065 1553.330 191.515 ;
      LAYER met4 ;
        RECT 1553.730 186.465 1750.270 191.115 ;
      LAYER met4 ;
        RECT 1750.670 186.065 1827.330 191.515 ;
      LAYER met4 ;
        RECT 1827.730 186.465 2024.270 191.115 ;
      LAYER met4 ;
        RECT 2024.670 186.065 2101.330 191.515 ;
      LAYER met4 ;
        RECT 2101.730 186.465 2298.270 191.115 ;
      LAYER met4 ;
        RECT 2298.670 186.065 2375.330 191.515 ;
      LAYER met4 ;
        RECT 2375.730 186.465 2572.270 191.115 ;
      LAYER met4 ;
        RECT 2572.670 186.065 2649.330 191.515 ;
      LAYER met4 ;
        RECT 2649.730 186.465 2846.270 191.115 ;
      LAYER met4 ;
        RECT 2846.670 186.065 2918.330 191.515 ;
      LAYER met4 ;
        RECT 2918.730 186.465 3115.270 191.115 ;
      LAYER met4 ;
        RECT 3115.670 186.065 3187.330 191.515 ;
      LAYER met4 ;
        RECT 3187.730 186.465 3385.270 191.115 ;
      LAYER met4 ;
        RECT 3385.670 186.065 3435.335 191.515 ;
        RECT 152.665 185.465 200.000 186.065 ;
        RECT 394.965 185.465 468.035 186.065 ;
        RECT 663.965 185.465 737.035 186.065 ;
        RECT 933.030 185.465 1011.035 186.065 ;
        RECT 1206.000 185.465 1281.000 186.065 ;
        RECT 1476.030 185.465 1554.035 186.065 ;
        RECT 1750.030 185.465 1828.035 186.065 ;
        RECT 2024.030 185.465 2102.035 186.065 ;
        RECT 2298.030 185.465 2376.035 186.065 ;
        RECT 2572.030 185.465 2650.035 186.065 ;
        RECT 2845.965 185.465 2919.035 186.065 ;
        RECT 3114.965 185.465 3188.035 186.065 ;
        RECT 3385.255 185.465 3435.335 186.065 ;
        RECT 152.665 181.215 198.130 185.465 ;
      LAYER met4 ;
        RECT 198.530 181.615 394.965 185.065 ;
      LAYER met4 ;
        RECT 395.365 181.215 467.635 185.465 ;
      LAYER met4 ;
        RECT 468.035 181.615 663.965 185.065 ;
      LAYER met4 ;
        RECT 664.365 181.215 736.635 185.465 ;
      LAYER met4 ;
        RECT 737.035 181.615 933.030 185.065 ;
      LAYER met4 ;
        RECT 933.430 181.215 1010.635 185.465 ;
      LAYER met4 ;
        RECT 1011.035 181.615 1206.965 185.065 ;
      LAYER met4 ;
        RECT 1207.365 181.215 1279.635 185.465 ;
      LAYER met4 ;
        RECT 1280.035 181.615 1476.030 185.065 ;
      LAYER met4 ;
        RECT 1476.430 181.215 1553.635 185.465 ;
      LAYER met4 ;
        RECT 1554.035 181.615 1750.030 185.065 ;
      LAYER met4 ;
        RECT 1750.430 181.215 1827.635 185.465 ;
      LAYER met4 ;
        RECT 1828.035 181.615 2024.030 185.065 ;
      LAYER met4 ;
        RECT 2024.430 181.215 2101.635 185.465 ;
      LAYER met4 ;
        RECT 2102.035 181.615 2298.030 185.065 ;
      LAYER met4 ;
        RECT 2298.430 181.215 2375.635 185.465 ;
      LAYER met4 ;
        RECT 2376.035 181.615 2572.030 185.065 ;
      LAYER met4 ;
        RECT 2572.430 181.215 2649.635 185.465 ;
      LAYER met4 ;
        RECT 2650.035 181.615 2845.965 185.065 ;
      LAYER met4 ;
        RECT 2846.365 181.215 2918.635 185.465 ;
        RECT 3115.365 181.215 3187.635 185.465 ;
        RECT 3385.655 181.215 3435.335 185.465 ;
        RECT 152.665 180.615 200.000 181.215 ;
        RECT 394.965 180.615 468.035 181.215 ;
        RECT 663.965 180.615 737.035 181.215 ;
        RECT 933.030 180.615 1011.035 181.215 ;
        RECT 1206.000 180.615 1281.000 181.215 ;
        RECT 1476.030 180.615 1554.035 181.215 ;
        RECT 1750.030 180.615 1828.035 181.215 ;
        RECT 2024.030 180.615 2102.035 181.215 ;
        RECT 2298.030 180.615 2376.035 181.215 ;
        RECT 2572.030 180.615 2650.035 181.215 ;
        RECT 2845.965 180.615 2919.035 181.215 ;
        RECT 3114.965 180.615 3188.035 181.215 ;
        RECT 3385.255 180.615 3435.335 181.215 ;
        RECT 152.665 180.025 198.075 180.615 ;
        RECT 147.275 176.690 198.075 180.025 ;
        RECT 143.995 176.425 198.075 176.690 ;
        RECT 0.000 175.165 198.075 176.425 ;
      LAYER met4 ;
        RECT 198.475 175.565 395.270 180.215 ;
      LAYER met4 ;
        RECT 395.670 175.165 467.330 180.615 ;
      LAYER met4 ;
        RECT 467.730 175.565 664.270 180.215 ;
      LAYER met4 ;
        RECT 664.670 175.165 736.330 180.615 ;
      LAYER met4 ;
        RECT 736.730 175.565 933.270 180.215 ;
      LAYER met4 ;
        RECT 933.670 175.165 1010.330 180.615 ;
      LAYER met4 ;
        RECT 1010.730 175.565 1207.270 180.215 ;
      LAYER met4 ;
        RECT 1207.670 175.165 1279.330 180.615 ;
      LAYER met4 ;
        RECT 1279.730 175.565 1476.270 180.215 ;
      LAYER met4 ;
        RECT 1476.670 175.165 1553.330 180.615 ;
      LAYER met4 ;
        RECT 1553.730 175.565 1750.270 180.215 ;
      LAYER met4 ;
        RECT 1750.670 175.165 1827.330 180.615 ;
      LAYER met4 ;
        RECT 1827.730 175.565 2024.270 180.215 ;
      LAYER met4 ;
        RECT 2024.670 175.165 2101.330 180.615 ;
      LAYER met4 ;
        RECT 2101.730 175.565 2298.270 180.215 ;
      LAYER met4 ;
        RECT 2298.670 175.165 2375.330 180.615 ;
      LAYER met4 ;
        RECT 2375.730 175.565 2572.270 180.215 ;
      LAYER met4 ;
        RECT 2572.670 175.165 2649.330 180.615 ;
      LAYER met4 ;
        RECT 2649.730 175.565 2846.270 180.215 ;
      LAYER met4 ;
        RECT 2846.670 175.165 2918.330 180.615 ;
      LAYER met4 ;
        RECT 2918.730 175.565 3115.270 180.215 ;
      LAYER met4 ;
        RECT 3115.670 175.165 3187.330 180.615 ;
      LAYER met4 ;
        RECT 3187.730 175.565 3385.270 180.215 ;
      LAYER met4 ;
        RECT 3385.670 180.025 3435.335 180.615 ;
      LAYER met4 ;
        RECT 3435.735 180.425 3436.065 345.000 ;
      LAYER met4 ;
        RECT 3385.670 178.665 3435.965 180.025 ;
      LAYER met4 ;
        RECT 3436.365 179.065 3439.345 525.535 ;
      LAYER met4 ;
        RECT 3439.745 501.670 3440.725 525.935 ;
      LAYER met4 ;
        RECT 3439.645 500.000 3440.825 501.270 ;
      LAYER met4 ;
        RECT 3439.745 355.000 3440.725 500.000 ;
        RECT 3439.645 350.000 3440.825 355.000 ;
        RECT 3439.745 200.000 3440.725 345.000 ;
        RECT 3385.670 178.050 3439.245 178.665 ;
      LAYER met4 ;
        RECT 3439.645 178.450 3440.825 200.000 ;
      LAYER met4 ;
        RECT 3385.670 176.690 3440.725 178.050 ;
      LAYER met4 ;
        RECT 3441.125 177.090 3444.105 541.240 ;
      LAYER met4 ;
        RECT 3444.505 533.310 3588.000 541.640 ;
      LAYER met4 ;
        RECT 3444.405 350.000 3444.735 532.910 ;
      LAYER met4 ;
        RECT 3445.135 501.670 3588.000 533.310 ;
        RECT 3445.135 501.030 3445.835 501.670 ;
        RECT 3445.135 355.000 3445.835 500.000 ;
      LAYER met4 ;
        RECT 3444.405 176.825 3444.735 345.000 ;
      LAYER met4 ;
        RECT 3445.135 197.975 3445.835 345.000 ;
      LAYER met4 ;
        RECT 3446.235 198.375 3450.685 501.270 ;
      LAYER met4 ;
        RECT 3451.085 501.030 3451.685 501.670 ;
        RECT 3451.085 355.000 3451.685 500.000 ;
        RECT 3451.085 198.120 3451.685 345.000 ;
      LAYER met4 ;
        RECT 3452.085 198.520 3456.535 501.270 ;
      LAYER met4 ;
        RECT 3456.935 501.030 3457.635 501.670 ;
        RECT 3456.935 499.000 3458.035 500.000 ;
      LAYER met4 ;
        RECT 3458.035 499.000 3483.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 501.030 3563.385 501.670 ;
      LAYER met4 ;
        RECT 3563.785 500.000 3588.000 501.270 ;
      LAYER met4 ;
        RECT 3483.000 499.000 3485.035 500.000 ;
        RECT 3456.935 496.000 3485.035 499.000 ;
        RECT 3456.935 494.000 3458.035 496.000 ;
      LAYER met4 ;
        RECT 3458.035 494.000 3483.000 496.000 ;
      LAYER met4 ;
        RECT 3483.000 494.000 3485.035 496.000 ;
        RECT 3456.935 476.000 3485.035 494.000 ;
        RECT 3456.935 474.000 3458.035 476.000 ;
      LAYER met4 ;
        RECT 3458.035 474.000 3483.000 476.000 ;
      LAYER met4 ;
        RECT 3483.000 474.000 3485.035 476.000 ;
        RECT 3456.935 456.000 3485.035 474.000 ;
        RECT 3456.935 454.000 3458.035 456.000 ;
      LAYER met4 ;
        RECT 3458.035 454.000 3483.000 456.000 ;
      LAYER met4 ;
        RECT 3483.000 454.000 3485.035 456.000 ;
        RECT 3456.935 436.000 3485.035 454.000 ;
        RECT 3456.935 434.000 3458.035 436.000 ;
      LAYER met4 ;
        RECT 3458.035 434.000 3483.000 436.000 ;
      LAYER met4 ;
        RECT 3483.000 434.000 3485.035 436.000 ;
        RECT 3456.935 416.000 3485.035 434.000 ;
        RECT 3456.935 414.000 3458.035 416.000 ;
      LAYER met4 ;
        RECT 3458.035 414.000 3483.000 416.000 ;
      LAYER met4 ;
        RECT 3483.000 414.000 3485.035 416.000 ;
        RECT 3456.935 396.000 3485.035 414.000 ;
        RECT 3456.935 394.000 3458.035 396.000 ;
      LAYER met4 ;
        RECT 3458.035 394.000 3483.000 396.000 ;
      LAYER met4 ;
        RECT 3483.000 394.000 3485.035 396.000 ;
        RECT 3456.935 376.000 3485.035 394.000 ;
        RECT 3456.935 374.000 3458.035 376.000 ;
      LAYER met4 ;
        RECT 3458.035 374.000 3483.000 376.000 ;
      LAYER met4 ;
        RECT 3483.000 374.000 3485.035 376.000 ;
        RECT 3456.935 356.000 3485.035 374.000 ;
        RECT 3456.935 355.000 3458.035 356.000 ;
        RECT 3456.935 344.000 3458.035 345.000 ;
      LAYER met4 ;
        RECT 3458.035 344.000 3483.000 356.000 ;
      LAYER met4 ;
        RECT 3483.000 355.000 3485.035 356.000 ;
        RECT 3562.035 355.000 3588.000 500.000 ;
        RECT 3563.785 345.000 3588.000 355.000 ;
        RECT 3483.000 344.000 3485.035 345.000 ;
        RECT 3456.935 341.000 3485.035 344.000 ;
        RECT 3456.935 339.000 3458.035 341.000 ;
      LAYER met4 ;
        RECT 3458.035 339.000 3483.000 341.000 ;
      LAYER met4 ;
        RECT 3483.000 339.000 3485.035 341.000 ;
        RECT 3456.935 321.000 3485.035 339.000 ;
        RECT 3456.935 319.000 3458.035 321.000 ;
      LAYER met4 ;
        RECT 3458.035 319.000 3483.000 321.000 ;
      LAYER met4 ;
        RECT 3483.000 319.000 3485.035 321.000 ;
        RECT 3456.935 301.000 3485.035 319.000 ;
        RECT 3456.935 299.000 3458.035 301.000 ;
      LAYER met4 ;
        RECT 3458.035 299.000 3483.000 301.000 ;
      LAYER met4 ;
        RECT 3483.000 299.000 3485.035 301.000 ;
        RECT 3456.935 281.000 3485.035 299.000 ;
        RECT 3456.935 279.000 3458.035 281.000 ;
      LAYER met4 ;
        RECT 3458.035 279.000 3483.000 281.000 ;
      LAYER met4 ;
        RECT 3483.000 279.000 3485.035 281.000 ;
        RECT 3456.935 261.000 3485.035 279.000 ;
        RECT 3456.935 259.000 3458.035 261.000 ;
      LAYER met4 ;
        RECT 3458.035 259.000 3483.000 261.000 ;
      LAYER met4 ;
        RECT 3483.000 259.000 3485.035 261.000 ;
        RECT 3456.935 241.000 3485.035 259.000 ;
        RECT 3456.935 239.000 3458.035 241.000 ;
      LAYER met4 ;
        RECT 3458.035 239.000 3483.000 241.000 ;
      LAYER met4 ;
        RECT 3483.000 239.000 3485.035 241.000 ;
        RECT 3456.935 221.000 3485.035 239.000 ;
        RECT 3456.935 219.000 3458.035 221.000 ;
      LAYER met4 ;
        RECT 3458.035 219.000 3483.000 221.000 ;
      LAYER met4 ;
        RECT 3483.000 219.000 3485.035 221.000 ;
        RECT 3456.935 201.000 3485.035 219.000 ;
        RECT 3456.935 200.000 3458.035 201.000 ;
        RECT 3456.935 198.120 3457.635 200.000 ;
        RECT 3451.085 197.975 3457.635 198.120 ;
        RECT 3445.135 196.955 3457.635 197.975 ;
      LAYER met4 ;
        RECT 3458.035 197.355 3483.000 201.000 ;
      LAYER met4 ;
        RECT 3483.000 200.000 3485.035 201.000 ;
        RECT 3562.035 200.000 3588.000 345.000 ;
        RECT 3483.400 198.165 3563.385 200.000 ;
      LAYER met4 ;
        RECT 3563.785 198.565 3588.000 200.000 ;
      LAYER met4 ;
        RECT 3483.400 196.955 3588.000 198.165 ;
        RECT 3385.670 176.425 3444.005 176.690 ;
        RECT 3445.135 176.425 3588.000 196.955 ;
        RECT 3385.670 175.165 3588.000 176.425 ;
        RECT 0.000 174.565 200.000 175.165 ;
        RECT 394.965 174.565 468.035 175.165 ;
        RECT 663.965 174.565 737.035 175.165 ;
        RECT 933.030 174.565 1011.035 175.165 ;
        RECT 1206.000 174.565 1281.000 175.165 ;
        RECT 1476.030 174.565 1554.035 175.165 ;
        RECT 1750.030 174.565 1828.035 175.165 ;
        RECT 2024.030 174.565 2102.035 175.165 ;
        RECT 2298.030 174.565 2376.035 175.165 ;
        RECT 2572.030 174.565 2650.035 175.165 ;
        RECT 2845.965 174.565 2919.035 175.165 ;
        RECT 3114.965 174.565 3188.035 175.165 ;
        RECT 3385.255 174.565 3588.000 175.165 ;
        RECT 0.000 169.115 198.000 174.565 ;
      LAYER met4 ;
        RECT 198.400 169.515 395.270 174.165 ;
      LAYER met4 ;
        RECT 395.670 169.115 467.330 174.565 ;
      LAYER met4 ;
        RECT 467.730 169.515 664.270 174.165 ;
      LAYER met4 ;
        RECT 664.670 169.115 736.330 174.565 ;
      LAYER met4 ;
        RECT 736.730 169.515 933.270 174.165 ;
      LAYER met4 ;
        RECT 933.670 169.115 1010.330 174.565 ;
        RECT 1195.065 174.165 1206.065 174.200 ;
      LAYER met4 ;
        RECT 1010.730 169.515 1207.270 174.165 ;
      LAYER met4 ;
        RECT 1207.670 169.115 1279.330 174.565 ;
      LAYER met4 ;
        RECT 1279.730 169.515 1476.270 174.165 ;
      LAYER met4 ;
        RECT 1476.670 169.115 1553.330 174.565 ;
      LAYER met4 ;
        RECT 1553.730 169.515 1750.270 174.165 ;
      LAYER met4 ;
        RECT 1750.670 169.115 1827.330 174.565 ;
      LAYER met4 ;
        RECT 1827.730 169.515 2024.270 174.165 ;
      LAYER met4 ;
        RECT 2024.670 169.115 2101.330 174.565 ;
      LAYER met4 ;
        RECT 2101.730 169.515 2298.270 174.165 ;
      LAYER met4 ;
        RECT 2298.670 169.115 2375.330 174.565 ;
      LAYER met4 ;
        RECT 2375.730 169.515 2572.270 174.165 ;
      LAYER met4 ;
        RECT 2572.670 169.115 2649.330 174.565 ;
      LAYER met4 ;
        RECT 2649.730 169.515 2846.270 174.165 ;
      LAYER met4 ;
        RECT 2846.670 169.115 2918.330 174.565 ;
      LAYER met4 ;
        RECT 2918.730 169.515 3115.270 174.165 ;
      LAYER met4 ;
        RECT 3115.670 169.115 3187.330 174.565 ;
      LAYER met4 ;
        RECT 3187.730 169.515 3385.270 174.165 ;
      LAYER met4 ;
        RECT 3385.670 169.115 3588.000 174.565 ;
        RECT 0.000 168.515 200.000 169.115 ;
        RECT 394.965 168.515 468.035 169.115 ;
        RECT 663.965 168.515 737.035 169.115 ;
        RECT 933.030 168.515 1011.035 169.115 ;
        RECT 1206.000 168.515 1281.000 169.115 ;
        RECT 1476.030 168.515 1554.035 169.115 ;
        RECT 1750.030 168.515 1828.035 169.115 ;
        RECT 2024.030 168.515 2102.035 169.115 ;
        RECT 2298.030 168.515 2376.035 169.115 ;
        RECT 2572.030 168.515 2650.035 169.115 ;
        RECT 2845.965 168.515 2919.035 169.115 ;
        RECT 3114.965 168.515 3188.035 169.115 ;
        RECT 3385.255 168.515 3588.000 169.115 ;
        RECT 0.000 164.265 198.215 168.515 ;
      LAYER met4 ;
        RECT 198.615 164.665 395.270 168.115 ;
      LAYER met4 ;
        RECT 395.670 164.265 467.330 168.515 ;
      LAYER met4 ;
        RECT 467.730 164.665 664.270 168.115 ;
      LAYER met4 ;
        RECT 664.670 164.265 736.330 168.515 ;
      LAYER met4 ;
        RECT 736.730 164.665 933.270 168.115 ;
      LAYER met4 ;
        RECT 933.670 164.265 1010.330 168.515 ;
      LAYER met4 ;
        RECT 1010.730 164.665 1207.270 168.115 ;
      LAYER met4 ;
        RECT 1207.670 164.265 1279.330 168.515 ;
      LAYER met4 ;
        RECT 1279.730 164.665 1476.270 168.115 ;
      LAYER met4 ;
        RECT 1476.670 164.265 1553.330 168.515 ;
      LAYER met4 ;
        RECT 1553.730 164.665 1750.270 168.115 ;
      LAYER met4 ;
        RECT 1750.670 164.265 1827.330 168.515 ;
      LAYER met4 ;
        RECT 1827.730 164.665 2024.270 168.115 ;
      LAYER met4 ;
        RECT 2024.670 164.265 2101.330 168.515 ;
      LAYER met4 ;
        RECT 2101.730 164.665 2298.270 168.115 ;
      LAYER met4 ;
        RECT 2298.670 164.265 2375.330 168.515 ;
      LAYER met4 ;
        RECT 2375.730 164.665 2572.270 168.115 ;
      LAYER met4 ;
        RECT 2572.670 164.265 2649.330 168.515 ;
      LAYER met4 ;
        RECT 2649.730 164.665 2846.270 168.115 ;
      LAYER met4 ;
        RECT 2846.670 164.265 2918.330 168.515 ;
      LAYER met4 ;
        RECT 2918.730 164.665 3115.270 168.115 ;
      LAYER met4 ;
        RECT 3115.670 164.265 3187.330 168.515 ;
      LAYER met4 ;
        RECT 3187.730 164.665 3385.270 168.115 ;
      LAYER met4 ;
        RECT 3385.670 164.265 3588.000 168.515 ;
        RECT 0.000 163.665 200.000 164.265 ;
        RECT 394.965 163.665 468.035 164.265 ;
        RECT 663.965 163.665 737.035 164.265 ;
        RECT 933.030 163.665 1011.035 164.265 ;
        RECT 1206.000 163.665 1281.000 164.265 ;
        RECT 1476.030 163.665 1554.035 164.265 ;
        RECT 1750.030 163.665 1828.035 164.265 ;
        RECT 2024.030 163.665 2102.035 164.265 ;
        RECT 2298.030 163.665 2376.035 164.265 ;
        RECT 2572.030 163.665 2650.035 164.265 ;
        RECT 2845.965 163.665 2919.035 164.265 ;
        RECT 3114.965 163.665 3188.035 164.265 ;
        RECT 3385.255 163.665 3588.000 164.265 ;
        RECT 0.000 159.415 198.265 163.665 ;
        RECT 395.670 159.415 467.330 163.665 ;
        RECT 664.670 159.415 736.330 163.665 ;
      LAYER met4 ;
        RECT 736.730 159.815 933.270 163.265 ;
      LAYER met4 ;
        RECT 933.670 159.415 1010.330 163.665 ;
      LAYER met4 ;
        RECT 1010.730 159.815 1207.270 163.265 ;
      LAYER met4 ;
        RECT 1207.670 159.415 1279.330 163.665 ;
      LAYER met4 ;
        RECT 1279.730 159.815 1476.270 163.265 ;
      LAYER met4 ;
        RECT 1476.670 159.415 1553.330 163.665 ;
      LAYER met4 ;
        RECT 1553.730 159.815 1750.270 163.265 ;
      LAYER met4 ;
        RECT 1750.670 159.415 1827.330 163.665 ;
      LAYER met4 ;
        RECT 1827.730 159.815 2024.270 163.265 ;
      LAYER met4 ;
        RECT 2024.670 159.415 2101.330 163.665 ;
      LAYER met4 ;
        RECT 2101.730 159.815 2298.270 163.265 ;
      LAYER met4 ;
        RECT 2298.670 159.415 2375.330 163.665 ;
      LAYER met4 ;
        RECT 2375.730 159.815 2572.270 163.265 ;
      LAYER met4 ;
        RECT 2572.670 159.415 2649.330 163.665 ;
      LAYER met4 ;
        RECT 2649.730 159.815 2846.270 163.265 ;
      LAYER met4 ;
        RECT 2846.670 159.415 2918.330 163.665 ;
      LAYER met4 ;
        RECT 2918.730 159.815 3115.270 163.265 ;
      LAYER met4 ;
        RECT 3115.670 159.415 3187.330 163.665 ;
      LAYER met4 ;
        RECT 3187.730 159.815 3385.270 163.265 ;
      LAYER met4 ;
        RECT 3385.670 159.415 3588.000 163.665 ;
        RECT 0.000 158.815 200.000 159.415 ;
        RECT 394.965 158.815 468.035 159.415 ;
        RECT 663.965 158.815 737.035 159.415 ;
        RECT 933.030 158.815 1011.035 159.415 ;
        RECT 1206.000 158.815 1281.000 159.415 ;
        RECT 1476.030 158.815 1554.035 159.415 ;
        RECT 1750.030 158.815 1828.035 159.415 ;
        RECT 2024.030 158.815 2102.035 159.415 ;
        RECT 2298.030 158.815 2376.035 159.415 ;
        RECT 2572.030 158.815 2650.035 159.415 ;
        RECT 2845.965 158.815 2919.035 159.415 ;
        RECT 3114.965 158.815 3188.035 159.415 ;
        RECT 3385.255 158.815 3588.000 159.415 ;
        RECT 0.000 153.365 198.125 158.815 ;
      LAYER met4 ;
        RECT 198.525 153.765 395.270 158.415 ;
      LAYER met4 ;
        RECT 395.670 153.365 467.330 158.815 ;
        RECT 664.670 158.770 736.330 158.815 ;
      LAYER met4 ;
        RECT 467.730 158.370 664.270 158.415 ;
        RECT 467.730 153.810 664.345 158.370 ;
        RECT 467.730 153.765 664.270 153.810 ;
      LAYER met4 ;
        RECT 664.745 153.410 736.330 158.770 ;
      LAYER met4 ;
        RECT 736.730 153.765 933.270 158.415 ;
      LAYER met4 ;
        RECT 664.670 153.365 736.330 153.410 ;
        RECT 933.670 153.365 1010.330 158.815 ;
        RECT 1207.670 153.365 1279.330 158.815 ;
        RECT 1280.930 158.415 1291.975 158.450 ;
        RECT 1476.670 153.365 1553.330 158.815 ;
      LAYER met4 ;
        RECT 1553.730 153.765 1750.270 158.415 ;
      LAYER met4 ;
        RECT 1750.670 153.365 1827.330 158.815 ;
      LAYER met4 ;
        RECT 1827.730 153.765 2024.270 158.415 ;
      LAYER met4 ;
        RECT 2024.670 153.365 2101.330 158.815 ;
      LAYER met4 ;
        RECT 2101.730 153.765 2298.270 158.415 ;
      LAYER met4 ;
        RECT 2298.670 153.365 2375.330 158.815 ;
      LAYER met4 ;
        RECT 2375.730 153.765 2572.270 158.415 ;
      LAYER met4 ;
        RECT 2572.670 153.365 2649.330 158.815 ;
      LAYER met4 ;
        RECT 2649.730 153.765 2846.270 158.415 ;
      LAYER met4 ;
        RECT 2846.670 153.365 2918.330 158.815 ;
      LAYER met4 ;
        RECT 2918.730 153.765 3115.270 158.415 ;
      LAYER met4 ;
        RECT 3115.670 153.365 3187.330 158.815 ;
      LAYER met4 ;
        RECT 3187.730 153.765 3385.270 158.415 ;
      LAYER met4 ;
        RECT 3385.670 153.365 3588.000 158.815 ;
        RECT 0.000 152.665 200.000 153.365 ;
        RECT 394.965 152.665 468.035 153.365 ;
        RECT 663.965 152.665 737.035 153.365 ;
        RECT 933.030 152.665 1011.035 153.365 ;
        RECT 1206.000 152.665 1281.000 153.365 ;
        RECT 1476.030 152.665 1554.035 153.365 ;
        RECT 1750.030 152.665 1828.035 153.365 ;
        RECT 2024.030 152.665 2102.035 153.365 ;
        RECT 2298.030 152.665 2376.035 153.365 ;
        RECT 2572.030 152.665 2650.035 153.365 ;
        RECT 2845.965 152.665 2919.035 153.365 ;
        RECT 3114.965 152.665 3188.035 153.365 ;
        RECT 3385.255 152.665 3588.000 153.365 ;
        RECT 0.000 152.035 180.025 152.665 ;
        RECT 395.670 152.035 467.330 152.665 ;
        RECT 965.310 152.035 1008.990 152.665 ;
        RECT 0.000 148.755 178.665 152.035 ;
      LAYER met4 ;
        RECT 1009.390 151.935 1507.910 152.265 ;
      LAYER met4 ;
        RECT 1508.310 152.035 1551.990 152.665 ;
      LAYER met4 ;
        RECT 1552.390 151.935 1781.910 152.265 ;
      LAYER met4 ;
        RECT 1782.310 152.035 1825.990 152.665 ;
      LAYER met4 ;
        RECT 1826.390 151.935 2055.910 152.265 ;
      LAYER met4 ;
        RECT 2056.310 152.035 2099.990 152.665 ;
      LAYER met4 ;
        RECT 2100.390 151.935 2329.910 152.265 ;
      LAYER met4 ;
        RECT 2330.310 152.035 2373.990 152.665 ;
      LAYER met4 ;
        RECT 2374.390 151.935 2603.910 152.265 ;
      LAYER met4 ;
        RECT 2604.310 152.035 2647.990 152.665 ;
      LAYER met4 ;
        RECT 2648.390 151.935 3407.575 152.265 ;
      LAYER met4 ;
        RECT 0.000 147.275 178.050 148.755 ;
      LAYER met4 ;
        RECT 179.065 148.655 957.535 151.635 ;
      LAYER met4 ;
        RECT 0.000 143.995 176.690 147.275 ;
      LAYER met4 ;
        RECT 178.450 147.175 200.000 148.355 ;
      LAYER met4 ;
        RECT 237.000 148.255 357.000 148.355 ;
        RECT 506.000 148.255 626.000 148.355 ;
        RECT 200.000 147.275 394.000 148.255 ;
        RECT 395.670 147.275 467.330 148.255 ;
        RECT 469.000 147.275 663.000 148.255 ;
        RECT 237.000 147.175 357.000 147.275 ;
        RECT 506.000 147.175 626.000 147.275 ;
      LAYER met4 ;
        RECT 663.000 147.175 664.270 148.355 ;
      LAYER met4 ;
        RECT 664.670 147.275 736.330 148.255 ;
      LAYER met4 ;
        RECT 736.730 147.175 738.000 148.355 ;
      LAYER met4 ;
        RECT 775.000 148.255 895.000 148.355 ;
        RECT 738.000 147.275 932.000 148.255 ;
        RECT 775.000 147.175 895.000 147.275 ;
      LAYER met4 ;
        RECT 932.000 147.175 933.270 148.355 ;
      LAYER met4 ;
        RECT 957.935 148.255 959.455 151.535 ;
      LAYER met4 ;
        RECT 959.855 148.655 1500.535 151.635 ;
      LAYER met4 ;
        RECT 933.670 147.275 1010.330 148.255 ;
        RECT 0.000 142.865 176.425 143.995 ;
      LAYER met4 ;
        RECT 177.090 143.895 973.240 146.875 ;
      LAYER met4 ;
        RECT 973.640 143.495 975.160 147.275 ;
      LAYER met4 ;
        RECT 1010.730 147.175 1012.000 148.355 ;
      LAYER met4 ;
        RECT 1049.000 148.255 1169.000 148.355 ;
        RECT 1012.000 147.275 1206.000 148.255 ;
        RECT 1049.000 147.175 1169.000 147.275 ;
      LAYER met4 ;
        RECT 1206.000 147.175 1207.270 148.355 ;
      LAYER met4 ;
        RECT 1207.670 147.275 1279.330 148.255 ;
      LAYER met4 ;
        RECT 1279.730 147.175 1281.000 148.355 ;
      LAYER met4 ;
        RECT 1318.000 148.255 1438.000 148.355 ;
        RECT 1281.000 147.275 1475.000 148.255 ;
        RECT 1318.000 147.175 1438.000 147.275 ;
      LAYER met4 ;
        RECT 1475.000 147.175 1476.270 148.355 ;
      LAYER met4 ;
        RECT 1500.935 148.255 1502.455 151.535 ;
      LAYER met4 ;
        RECT 1502.855 148.655 1774.535 151.635 ;
      LAYER met4 ;
        RECT 1476.670 147.275 1553.330 148.255 ;
      LAYER met4 ;
        RECT 975.560 143.895 1516.240 146.875 ;
      LAYER met4 ;
        RECT 395.670 142.865 467.330 143.495 ;
        RECT 965.310 142.865 1008.990 143.495 ;
      LAYER met4 ;
        RECT 1009.390 143.265 1507.910 143.595 ;
      LAYER met4 ;
        RECT 1516.640 143.495 1518.160 147.275 ;
      LAYER met4 ;
        RECT 1553.730 147.175 1555.000 148.355 ;
      LAYER met4 ;
        RECT 1592.000 148.255 1712.000 148.355 ;
        RECT 1555.000 147.275 1749.000 148.255 ;
        RECT 1592.000 147.175 1712.000 147.275 ;
      LAYER met4 ;
        RECT 1749.000 147.175 1750.270 148.355 ;
      LAYER met4 ;
        RECT 1774.935 148.255 1776.455 151.535 ;
      LAYER met4 ;
        RECT 1776.855 148.655 2048.535 151.635 ;
      LAYER met4 ;
        RECT 1750.670 147.275 1827.330 148.255 ;
      LAYER met4 ;
        RECT 1518.560 143.895 1790.240 146.875 ;
      LAYER met4 ;
        RECT 1508.310 142.865 1551.990 143.495 ;
      LAYER met4 ;
        RECT 1552.390 143.265 1781.910 143.595 ;
      LAYER met4 ;
        RECT 1790.640 143.495 1792.160 147.275 ;
      LAYER met4 ;
        RECT 1827.730 147.175 1829.000 148.355 ;
      LAYER met4 ;
        RECT 1866.000 148.255 1986.000 148.355 ;
        RECT 1829.000 147.275 2023.000 148.255 ;
        RECT 1866.000 147.175 1986.000 147.275 ;
      LAYER met4 ;
        RECT 2023.000 147.175 2024.270 148.355 ;
      LAYER met4 ;
        RECT 2048.935 148.255 2050.455 151.535 ;
      LAYER met4 ;
        RECT 2050.855 148.655 2322.535 151.635 ;
      LAYER met4 ;
        RECT 2024.670 147.275 2101.330 148.255 ;
      LAYER met4 ;
        RECT 1792.560 143.895 2064.240 146.875 ;
      LAYER met4 ;
        RECT 1782.310 142.865 1825.990 143.495 ;
      LAYER met4 ;
        RECT 1826.390 143.265 2055.910 143.595 ;
      LAYER met4 ;
        RECT 2064.640 143.495 2066.160 147.275 ;
      LAYER met4 ;
        RECT 2101.730 147.175 2103.000 148.355 ;
      LAYER met4 ;
        RECT 2140.000 148.255 2260.000 148.355 ;
        RECT 2103.000 147.275 2297.000 148.255 ;
        RECT 2140.000 147.175 2260.000 147.275 ;
      LAYER met4 ;
        RECT 2297.000 147.175 2298.270 148.355 ;
      LAYER met4 ;
        RECT 2322.935 148.255 2324.455 151.535 ;
      LAYER met4 ;
        RECT 2324.855 148.655 2596.535 151.635 ;
      LAYER met4 ;
        RECT 2298.670 147.275 2375.330 148.255 ;
      LAYER met4 ;
        RECT 2066.560 143.895 2338.240 146.875 ;
      LAYER met4 ;
        RECT 2056.310 142.865 2099.990 143.495 ;
      LAYER met4 ;
        RECT 2100.390 143.265 2329.910 143.595 ;
      LAYER met4 ;
        RECT 2338.640 143.495 2340.160 147.275 ;
      LAYER met4 ;
        RECT 2375.730 147.175 2377.000 148.355 ;
      LAYER met4 ;
        RECT 2414.000 148.255 2534.000 148.355 ;
        RECT 2377.000 147.275 2571.000 148.255 ;
        RECT 2414.000 147.175 2534.000 147.275 ;
      LAYER met4 ;
        RECT 2571.000 147.175 2572.270 148.355 ;
      LAYER met4 ;
        RECT 2596.935 148.255 2598.455 151.535 ;
      LAYER met4 ;
        RECT 2598.855 148.655 3404.875 151.635 ;
      LAYER met4 ;
        RECT 3407.975 151.535 3588.000 152.665 ;
        RECT 3405.275 148.755 3588.000 151.535 ;
        RECT 2572.670 147.275 2649.330 148.255 ;
      LAYER met4 ;
        RECT 2340.560 143.895 2612.240 146.875 ;
      LAYER met4 ;
        RECT 2330.310 142.865 2373.990 143.495 ;
      LAYER met4 ;
        RECT 2374.390 143.265 2603.910 143.595 ;
      LAYER met4 ;
        RECT 2612.640 143.495 2614.160 147.275 ;
      LAYER met4 ;
        RECT 2649.730 147.175 2651.000 148.355 ;
      LAYER met4 ;
        RECT 2688.000 148.255 2808.000 148.355 ;
        RECT 2651.000 147.275 2845.000 148.255 ;
        RECT 2688.000 147.175 2808.000 147.275 ;
      LAYER met4 ;
        RECT 2845.000 147.175 2846.270 148.355 ;
      LAYER met4 ;
        RECT 2846.670 147.275 2918.330 148.255 ;
      LAYER met4 ;
        RECT 2918.730 147.175 2920.000 148.355 ;
      LAYER met4 ;
        RECT 2957.000 148.255 3077.000 148.355 ;
        RECT 2920.000 147.275 3114.000 148.255 ;
        RECT 2957.000 147.175 3077.000 147.275 ;
      LAYER met4 ;
        RECT 3114.000 147.175 3115.270 148.355 ;
      LAYER met4 ;
        RECT 3115.670 147.275 3187.330 148.255 ;
      LAYER met4 ;
        RECT 3187.730 147.175 3189.000 148.355 ;
      LAYER met4 ;
        RECT 3226.000 148.255 3346.000 148.355 ;
        RECT 3189.000 147.275 3384.000 148.255 ;
        RECT 3226.000 147.175 3346.000 147.275 ;
      LAYER met4 ;
        RECT 3384.000 147.175 3405.555 148.355 ;
      LAYER met4 ;
        RECT 3405.955 147.275 3588.000 148.755 ;
      LAYER met4 ;
        RECT 2614.560 143.895 3410.910 146.875 ;
      LAYER met4 ;
        RECT 3411.310 143.995 3588.000 147.275 ;
        RECT 2604.310 142.865 2647.990 143.495 ;
      LAYER met4 ;
        RECT 2648.390 143.265 3411.175 143.595 ;
      LAYER met4 ;
        RECT 3411.575 142.865 3588.000 143.995 ;
        RECT 0.000 142.165 237.000 142.865 ;
        RECT 357.000 142.165 394.000 142.865 ;
        RECT 394.965 142.165 468.035 142.865 ;
        RECT 469.000 142.165 506.000 142.865 ;
        RECT 626.000 142.165 663.000 142.865 ;
        RECT 663.965 142.165 737.035 142.865 ;
        RECT 738.000 142.165 775.000 142.865 ;
        RECT 895.000 142.165 932.000 142.865 ;
        RECT 933.030 142.165 1011.035 142.865 ;
        RECT 1012.000 142.165 1049.000 142.865 ;
        RECT 1169.000 142.165 1318.000 142.865 ;
        RECT 1438.000 142.165 1475.000 142.865 ;
        RECT 1476.030 142.165 1554.035 142.865 ;
        RECT 1555.000 142.165 1592.000 142.865 ;
        RECT 1712.000 142.165 1749.000 142.865 ;
        RECT 1750.030 142.165 1828.035 142.865 ;
        RECT 1829.000 142.165 1866.000 142.865 ;
        RECT 1986.000 142.165 2023.000 142.865 ;
        RECT 2024.030 142.165 2102.035 142.865 ;
        RECT 2103.000 142.165 2140.000 142.865 ;
        RECT 2260.000 142.165 2297.000 142.865 ;
        RECT 2298.030 142.165 2376.035 142.865 ;
        RECT 2377.000 142.165 2414.000 142.865 ;
        RECT 2534.000 142.165 2571.000 142.865 ;
        RECT 2572.030 142.165 2650.035 142.865 ;
        RECT 2651.000 142.165 2688.000 142.865 ;
        RECT 2808.000 142.165 2845.000 142.865 ;
        RECT 2845.965 142.165 2919.035 142.865 ;
        RECT 2920.000 142.165 2957.000 142.865 ;
        RECT 3077.000 142.165 3114.000 142.865 ;
        RECT 3114.965 142.165 3188.035 142.865 ;
        RECT 3189.000 142.165 3226.000 142.865 ;
        RECT 3346.000 142.165 3384.000 142.865 ;
        RECT 3385.255 142.165 3588.000 142.865 ;
        RECT 0.000 136.915 197.975 142.165 ;
      LAYER met4 ;
        RECT 198.375 137.315 395.270 141.765 ;
      LAYER met4 ;
        RECT 395.670 136.915 467.330 142.165 ;
      LAYER met4 ;
        RECT 467.730 137.315 664.270 141.765 ;
      LAYER met4 ;
        RECT 664.670 136.915 736.330 142.165 ;
      LAYER met4 ;
        RECT 736.730 137.315 933.270 141.765 ;
      LAYER met4 ;
        RECT 933.670 136.915 1010.330 142.165 ;
      LAYER met4 ;
        RECT 1010.730 137.315 1207.270 141.765 ;
      LAYER met4 ;
        RECT 1207.670 136.915 1279.330 142.165 ;
      LAYER met4 ;
        RECT 1279.730 137.315 1476.270 141.765 ;
      LAYER met4 ;
        RECT 1476.670 136.915 1553.330 142.165 ;
      LAYER met4 ;
        RECT 1553.730 137.315 1750.270 141.765 ;
      LAYER met4 ;
        RECT 1750.670 136.915 1827.330 142.165 ;
      LAYER met4 ;
        RECT 1827.730 137.315 2024.270 141.765 ;
      LAYER met4 ;
        RECT 2024.670 136.915 2101.330 142.165 ;
      LAYER met4 ;
        RECT 2101.730 137.315 2298.270 141.765 ;
      LAYER met4 ;
        RECT 2298.670 136.915 2375.330 142.165 ;
      LAYER met4 ;
        RECT 2375.730 137.315 2572.270 141.765 ;
      LAYER met4 ;
        RECT 2572.670 136.915 2649.330 142.165 ;
      LAYER met4 ;
        RECT 2649.730 137.315 2846.270 141.765 ;
      LAYER met4 ;
        RECT 2846.670 136.915 2918.330 142.165 ;
      LAYER met4 ;
        RECT 2918.730 137.315 3115.270 141.765 ;
      LAYER met4 ;
        RECT 3115.670 136.915 3187.330 142.165 ;
      LAYER met4 ;
        RECT 3187.730 137.315 3385.270 141.765 ;
      LAYER met4 ;
        RECT 3385.670 136.915 3588.000 142.165 ;
        RECT 0.000 136.315 235.000 136.915 ;
        RECT 357.000 136.315 392.000 136.915 ;
        RECT 394.965 136.315 468.035 136.915 ;
        RECT 469.000 136.315 504.000 136.915 ;
        RECT 626.000 136.315 661.000 136.915 ;
        RECT 663.965 136.315 737.035 136.915 ;
        RECT 738.000 136.315 773.000 136.915 ;
        RECT 895.000 136.315 930.000 136.915 ;
        RECT 933.030 136.315 1011.035 136.915 ;
        RECT 1012.000 136.315 1047.000 136.915 ;
        RECT 1169.000 136.315 1204.000 136.915 ;
        RECT 1206.000 136.315 1316.000 136.915 ;
        RECT 1438.000 136.315 1473.000 136.915 ;
        RECT 1476.030 136.315 1554.035 136.915 ;
        RECT 1555.000 136.315 1590.000 136.915 ;
        RECT 1712.000 136.315 1747.000 136.915 ;
        RECT 1750.030 136.315 1828.035 136.915 ;
        RECT 1829.000 136.315 1864.000 136.915 ;
        RECT 1986.000 136.315 2021.000 136.915 ;
        RECT 2024.030 136.315 2102.035 136.915 ;
        RECT 2103.000 136.315 2138.000 136.915 ;
        RECT 2260.000 136.315 2295.000 136.915 ;
        RECT 2298.030 136.315 2376.035 136.915 ;
        RECT 2377.000 136.315 2412.000 136.915 ;
        RECT 2534.000 136.315 2569.000 136.915 ;
        RECT 2572.030 136.315 2650.035 136.915 ;
        RECT 2651.000 136.315 2686.000 136.915 ;
        RECT 2808.000 136.315 2843.000 136.915 ;
        RECT 2845.965 136.315 2919.035 136.915 ;
        RECT 2920.000 136.315 2955.000 136.915 ;
        RECT 3077.000 136.315 3112.000 136.915 ;
        RECT 3114.965 136.315 3188.035 136.915 ;
        RECT 3189.000 136.315 3224.000 136.915 ;
        RECT 3346.000 136.315 3381.000 136.915 ;
        RECT 3385.255 136.315 3588.000 136.915 ;
        RECT 0.000 131.065 198.120 136.315 ;
      LAYER met4 ;
        RECT 198.520 131.465 395.270 135.915 ;
      LAYER met4 ;
        RECT 395.670 131.065 467.330 136.315 ;
      LAYER met4 ;
        RECT 467.730 131.465 664.270 135.915 ;
      LAYER met4 ;
        RECT 664.670 131.065 736.330 136.315 ;
      LAYER met4 ;
        RECT 736.730 131.465 933.270 135.915 ;
      LAYER met4 ;
        RECT 933.670 131.065 1010.330 136.315 ;
      LAYER met4 ;
        RECT 1010.730 131.465 1207.270 135.915 ;
      LAYER met4 ;
        RECT 1207.670 131.065 1279.330 136.315 ;
      LAYER met4 ;
        RECT 1279.730 131.465 1476.270 135.915 ;
      LAYER met4 ;
        RECT 1476.670 131.065 1553.330 136.315 ;
      LAYER met4 ;
        RECT 1553.730 131.465 1750.270 135.915 ;
      LAYER met4 ;
        RECT 1750.670 131.065 1827.330 136.315 ;
      LAYER met4 ;
        RECT 1827.730 131.465 2024.270 135.915 ;
      LAYER met4 ;
        RECT 2024.670 131.065 2101.330 136.315 ;
      LAYER met4 ;
        RECT 2101.730 131.465 2298.270 135.915 ;
      LAYER met4 ;
        RECT 2298.670 131.065 2375.330 136.315 ;
      LAYER met4 ;
        RECT 2375.730 131.465 2572.270 135.915 ;
      LAYER met4 ;
        RECT 2572.670 131.065 2649.330 136.315 ;
      LAYER met4 ;
        RECT 2649.730 131.465 2846.270 135.915 ;
      LAYER met4 ;
        RECT 2846.670 131.065 2918.330 136.315 ;
      LAYER met4 ;
        RECT 2918.730 131.465 3115.270 135.915 ;
      LAYER met4 ;
        RECT 3115.670 131.065 3187.330 136.315 ;
      LAYER met4 ;
        RECT 3187.730 131.465 3385.270 135.915 ;
      LAYER met4 ;
        RECT 3385.670 131.065 3588.000 136.315 ;
        RECT 0.000 130.365 237.000 131.065 ;
        RECT 0.000 104.600 196.955 130.365 ;
        RECT 200.000 129.965 237.000 130.365 ;
        RECT 357.000 129.965 394.000 131.065 ;
        RECT 394.965 130.365 468.035 131.065 ;
      LAYER met4 ;
        RECT 197.355 105.000 201.000 129.965 ;
      LAYER met4 ;
        RECT 201.000 105.000 219.000 129.965 ;
      LAYER met4 ;
        RECT 219.000 105.000 221.000 129.965 ;
      LAYER met4 ;
        RECT 221.000 105.000 229.000 129.965 ;
      LAYER met4 ;
        RECT 229.000 105.000 231.000 129.965 ;
      LAYER met4 ;
        RECT 231.000 105.000 234.000 129.965 ;
      LAYER met4 ;
        RECT 234.000 105.000 358.000 129.965 ;
      LAYER met4 ;
        RECT 358.000 105.000 376.000 129.965 ;
      LAYER met4 ;
        RECT 376.000 105.000 378.000 129.965 ;
      LAYER met4 ;
        RECT 378.000 105.000 386.000 129.965 ;
      LAYER met4 ;
        RECT 386.000 105.000 388.000 129.965 ;
      LAYER met4 ;
        RECT 388.000 105.000 391.000 129.965 ;
      LAYER met4 ;
        RECT 391.000 105.000 395.270 129.965 ;
      LAYER met4 ;
        RECT 200.000 104.600 237.000 105.000 ;
        RECT 0.000 102.965 237.000 104.600 ;
        RECT 357.000 102.965 394.000 105.000 ;
        RECT 395.670 104.600 467.330 130.365 ;
        RECT 469.000 129.965 506.000 131.065 ;
        RECT 626.000 129.965 663.000 131.065 ;
        RECT 663.965 130.365 737.035 131.065 ;
      LAYER met4 ;
        RECT 467.730 105.000 470.000 129.965 ;
      LAYER met4 ;
        RECT 470.000 105.000 488.000 129.965 ;
      LAYER met4 ;
        RECT 488.000 105.000 490.000 129.965 ;
      LAYER met4 ;
        RECT 490.000 105.000 498.000 129.965 ;
      LAYER met4 ;
        RECT 498.000 105.000 500.000 129.965 ;
      LAYER met4 ;
        RECT 500.000 105.000 503.000 129.965 ;
      LAYER met4 ;
        RECT 503.000 105.000 627.000 129.965 ;
      LAYER met4 ;
        RECT 627.000 105.000 645.000 129.965 ;
      LAYER met4 ;
        RECT 645.000 105.000 647.000 129.965 ;
      LAYER met4 ;
        RECT 647.000 105.000 655.000 129.965 ;
      LAYER met4 ;
        RECT 655.000 105.000 657.000 129.965 ;
      LAYER met4 ;
        RECT 657.000 105.000 660.000 129.965 ;
      LAYER met4 ;
        RECT 660.000 105.000 664.270 129.965 ;
      LAYER met4 ;
        RECT 0.000 25.965 200.000 102.965 ;
        RECT 0.000 24.615 237.000 25.965 ;
        RECT 0.000 0.000 198.165 24.615 ;
        RECT 200.000 24.215 237.000 24.615 ;
        RECT 357.000 24.215 394.000 25.965 ;
        RECT 394.965 24.615 468.035 104.600 ;
        RECT 469.000 102.965 506.000 105.000 ;
        RECT 626.000 102.965 663.000 105.000 ;
        RECT 664.670 104.600 736.330 130.365 ;
        RECT 738.000 129.965 775.000 131.065 ;
        RECT 895.000 129.965 932.000 131.065 ;
        RECT 933.030 130.365 1011.035 131.065 ;
      LAYER met4 ;
        RECT 736.730 105.000 739.000 129.965 ;
      LAYER met4 ;
        RECT 739.000 105.000 757.000 129.965 ;
      LAYER met4 ;
        RECT 757.000 105.000 759.000 129.965 ;
      LAYER met4 ;
        RECT 759.000 105.000 767.000 129.965 ;
      LAYER met4 ;
        RECT 767.000 105.000 769.000 129.965 ;
      LAYER met4 ;
        RECT 769.000 105.000 772.000 129.965 ;
      LAYER met4 ;
        RECT 772.000 105.000 896.000 129.965 ;
      LAYER met4 ;
        RECT 896.000 105.000 914.000 129.965 ;
      LAYER met4 ;
        RECT 914.000 105.000 916.000 129.965 ;
      LAYER met4 ;
        RECT 916.000 105.000 924.000 129.965 ;
      LAYER met4 ;
        RECT 924.000 105.000 926.000 129.965 ;
      LAYER met4 ;
        RECT 926.000 105.000 929.000 129.965 ;
      LAYER met4 ;
        RECT 929.000 105.000 933.270 129.965 ;
        RECT 198.565 0.000 200.000 24.215 ;
      LAYER met4 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met4 ;
        RECT 394.000 0.000 395.270 24.215 ;
      LAYER met4 ;
        RECT 395.670 0.000 467.330 24.615 ;
        RECT 469.000 24.215 506.000 25.965 ;
        RECT 626.000 24.215 663.000 25.965 ;
        RECT 663.965 24.615 737.035 104.600 ;
        RECT 738.000 102.965 775.000 105.000 ;
        RECT 895.000 102.965 932.000 105.000 ;
        RECT 933.670 104.600 1010.330 130.365 ;
        RECT 1012.000 129.965 1049.000 131.065 ;
        RECT 1169.000 130.365 1318.000 131.065 ;
        RECT 1169.000 129.965 1206.000 130.365 ;
      LAYER met4 ;
        RECT 1010.730 105.000 1013.000 129.965 ;
      LAYER met4 ;
        RECT 1013.000 105.000 1031.000 129.965 ;
      LAYER met4 ;
        RECT 1031.000 105.000 1033.000 129.965 ;
      LAYER met4 ;
        RECT 1033.000 105.000 1041.000 129.965 ;
      LAYER met4 ;
        RECT 1041.000 105.000 1043.000 129.965 ;
      LAYER met4 ;
        RECT 1043.000 105.000 1046.000 129.965 ;
      LAYER met4 ;
        RECT 1046.000 105.000 1170.000 129.965 ;
      LAYER met4 ;
        RECT 1170.000 105.000 1188.000 129.965 ;
      LAYER met4 ;
        RECT 1188.000 105.000 1190.000 129.965 ;
      LAYER met4 ;
        RECT 1190.000 105.000 1198.000 129.965 ;
      LAYER met4 ;
        RECT 1198.000 105.000 1200.000 129.965 ;
      LAYER met4 ;
        RECT 1200.000 105.000 1203.000 129.965 ;
      LAYER met4 ;
        RECT 1203.000 105.000 1207.270 129.965 ;
        RECT 467.730 0.000 469.000 24.215 ;
      LAYER met4 ;
        RECT 469.000 0.000 663.000 24.215 ;
      LAYER met4 ;
        RECT 663.000 0.000 664.270 24.215 ;
      LAYER met4 ;
        RECT 664.670 0.000 736.330 24.615 ;
        RECT 738.000 24.215 775.000 25.965 ;
        RECT 895.000 24.215 932.000 25.965 ;
        RECT 933.030 24.615 1011.035 104.600 ;
        RECT 1012.000 102.965 1049.000 105.000 ;
        RECT 1169.000 104.600 1206.000 105.000 ;
        RECT 1207.670 104.600 1279.330 130.365 ;
        RECT 1281.000 129.965 1318.000 130.365 ;
        RECT 1438.000 129.965 1475.000 131.065 ;
        RECT 1476.030 130.365 1554.035 131.065 ;
      LAYER met4 ;
        RECT 1279.730 105.000 1282.000 129.965 ;
      LAYER met4 ;
        RECT 1282.000 105.000 1300.000 129.965 ;
      LAYER met4 ;
        RECT 1300.000 105.000 1302.000 129.965 ;
      LAYER met4 ;
        RECT 1302.000 105.000 1310.000 129.965 ;
      LAYER met4 ;
        RECT 1310.000 105.000 1312.000 129.965 ;
      LAYER met4 ;
        RECT 1312.000 105.000 1315.000 129.965 ;
      LAYER met4 ;
        RECT 1315.000 105.000 1439.000 129.965 ;
      LAYER met4 ;
        RECT 1439.000 105.000 1457.000 129.965 ;
      LAYER met4 ;
        RECT 1457.000 105.000 1459.000 129.965 ;
      LAYER met4 ;
        RECT 1459.000 105.000 1467.000 129.965 ;
      LAYER met4 ;
        RECT 1467.000 105.000 1469.000 129.965 ;
      LAYER met4 ;
        RECT 1469.000 105.000 1472.000 129.965 ;
      LAYER met4 ;
        RECT 1472.000 105.000 1476.270 129.965 ;
      LAYER met4 ;
        RECT 1281.000 104.600 1318.000 105.000 ;
        RECT 1169.000 102.965 1318.000 104.600 ;
        RECT 1438.000 102.965 1475.000 105.000 ;
        RECT 1476.670 104.600 1553.330 130.365 ;
        RECT 1555.000 129.965 1592.000 131.065 ;
        RECT 1712.000 129.965 1749.000 131.065 ;
        RECT 1750.030 130.365 1828.035 131.065 ;
      LAYER met4 ;
        RECT 1553.730 105.000 1556.000 129.965 ;
      LAYER met4 ;
        RECT 1556.000 105.000 1574.000 129.965 ;
      LAYER met4 ;
        RECT 1574.000 105.000 1576.000 129.965 ;
      LAYER met4 ;
        RECT 1576.000 105.000 1584.000 129.965 ;
      LAYER met4 ;
        RECT 1584.000 105.000 1586.000 129.965 ;
      LAYER met4 ;
        RECT 1586.000 105.000 1589.000 129.965 ;
      LAYER met4 ;
        RECT 1589.000 105.000 1713.000 129.965 ;
      LAYER met4 ;
        RECT 1713.000 105.000 1731.000 129.965 ;
      LAYER met4 ;
        RECT 1731.000 105.000 1733.000 129.965 ;
      LAYER met4 ;
        RECT 1733.000 105.000 1741.000 129.965 ;
      LAYER met4 ;
        RECT 1741.000 105.000 1743.000 129.965 ;
      LAYER met4 ;
        RECT 1743.000 105.000 1746.000 129.965 ;
      LAYER met4 ;
        RECT 1746.000 105.000 1750.270 129.965 ;
      LAYER met4 ;
        RECT 1206.000 25.965 1281.000 102.965 ;
      LAYER met4 ;
        RECT 736.730 0.000 738.000 24.215 ;
      LAYER met4 ;
        RECT 738.000 0.000 932.000 24.215 ;
      LAYER met4 ;
        RECT 932.000 0.000 933.270 24.215 ;
      LAYER met4 ;
        RECT 933.670 0.000 1010.330 24.615 ;
        RECT 1012.000 24.215 1049.000 25.965 ;
        RECT 1169.000 24.615 1318.000 25.965 ;
        RECT 1169.000 24.250 1206.000 24.615 ;
        RECT 1169.000 24.215 1206.215 24.250 ;
      LAYER met4 ;
        RECT 1010.730 0.000 1012.000 24.215 ;
      LAYER met4 ;
        RECT 1012.000 0.035 1204.530 24.215 ;
      LAYER met4 ;
        RECT 1204.530 0.035 1207.270 24.215 ;
      LAYER met4 ;
        RECT 1012.000 0.000 1206.000 0.035 ;
      LAYER met4 ;
        RECT 1206.000 0.000 1207.270 0.035 ;
      LAYER met4 ;
        RECT 1207.670 0.000 1279.330 24.615 ;
        RECT 1281.000 24.215 1318.000 24.615 ;
        RECT 1438.000 24.215 1475.000 25.965 ;
        RECT 1476.030 24.615 1554.035 104.600 ;
        RECT 1555.000 102.965 1592.000 105.000 ;
        RECT 1712.000 102.965 1749.000 105.000 ;
        RECT 1750.670 104.600 1827.330 130.365 ;
        RECT 1829.000 129.965 1866.000 131.065 ;
        RECT 1986.000 129.965 2023.000 131.065 ;
        RECT 2024.030 130.365 2102.035 131.065 ;
      LAYER met4 ;
        RECT 1827.730 105.000 1830.000 129.965 ;
      LAYER met4 ;
        RECT 1830.000 105.000 1848.000 129.965 ;
      LAYER met4 ;
        RECT 1848.000 105.000 1850.000 129.965 ;
      LAYER met4 ;
        RECT 1850.000 105.000 1858.000 129.965 ;
      LAYER met4 ;
        RECT 1858.000 105.000 1860.000 129.965 ;
      LAYER met4 ;
        RECT 1860.000 105.000 1863.000 129.965 ;
      LAYER met4 ;
        RECT 1863.000 105.000 1987.000 129.965 ;
      LAYER met4 ;
        RECT 1987.000 105.000 2005.000 129.965 ;
      LAYER met4 ;
        RECT 2005.000 105.000 2007.000 129.965 ;
      LAYER met4 ;
        RECT 2007.000 105.000 2015.000 129.965 ;
      LAYER met4 ;
        RECT 2015.000 105.000 2017.000 129.965 ;
      LAYER met4 ;
        RECT 2017.000 105.000 2020.000 129.965 ;
      LAYER met4 ;
        RECT 2020.000 105.000 2024.270 129.965 ;
        RECT 1279.730 0.000 1281.000 24.215 ;
      LAYER met4 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met4 ;
        RECT 1475.000 0.000 1476.270 24.215 ;
      LAYER met4 ;
        RECT 1476.670 0.000 1553.330 24.615 ;
        RECT 1555.000 24.215 1592.000 25.965 ;
        RECT 1712.000 24.215 1749.000 25.965 ;
        RECT 1750.030 24.615 1828.035 104.600 ;
        RECT 1829.000 102.965 1866.000 105.000 ;
        RECT 1986.000 102.965 2023.000 105.000 ;
        RECT 2024.670 104.600 2101.330 130.365 ;
        RECT 2103.000 129.965 2140.000 131.065 ;
        RECT 2260.000 129.965 2297.000 131.065 ;
        RECT 2298.030 130.365 2376.035 131.065 ;
      LAYER met4 ;
        RECT 2101.730 105.000 2104.000 129.965 ;
      LAYER met4 ;
        RECT 2104.000 105.000 2122.000 129.965 ;
      LAYER met4 ;
        RECT 2122.000 105.000 2124.000 129.965 ;
      LAYER met4 ;
        RECT 2124.000 105.000 2132.000 129.965 ;
      LAYER met4 ;
        RECT 2132.000 105.000 2134.000 129.965 ;
      LAYER met4 ;
        RECT 2134.000 105.000 2137.000 129.965 ;
      LAYER met4 ;
        RECT 2137.000 105.000 2261.000 129.965 ;
      LAYER met4 ;
        RECT 2261.000 105.000 2279.000 129.965 ;
      LAYER met4 ;
        RECT 2279.000 105.000 2281.000 129.965 ;
      LAYER met4 ;
        RECT 2281.000 105.000 2289.000 129.965 ;
      LAYER met4 ;
        RECT 2289.000 105.000 2291.000 129.965 ;
      LAYER met4 ;
        RECT 2291.000 105.000 2294.000 129.965 ;
      LAYER met4 ;
        RECT 2294.000 105.000 2298.270 129.965 ;
        RECT 1553.730 0.000 1555.000 24.215 ;
      LAYER met4 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met4 ;
        RECT 1749.000 0.000 1750.270 24.215 ;
      LAYER met4 ;
        RECT 1750.670 0.000 1827.330 24.615 ;
        RECT 1829.000 24.215 1866.000 25.965 ;
        RECT 1986.000 24.215 2023.000 25.965 ;
        RECT 2024.030 24.615 2102.035 104.600 ;
        RECT 2103.000 102.965 2140.000 105.000 ;
        RECT 2260.000 102.965 2297.000 105.000 ;
        RECT 2298.670 104.600 2375.330 130.365 ;
        RECT 2377.000 129.965 2414.000 131.065 ;
        RECT 2534.000 129.965 2571.000 131.065 ;
        RECT 2572.030 130.365 2650.035 131.065 ;
      LAYER met4 ;
        RECT 2375.730 105.000 2378.000 129.965 ;
      LAYER met4 ;
        RECT 2378.000 105.000 2396.000 129.965 ;
      LAYER met4 ;
        RECT 2396.000 105.000 2398.000 129.965 ;
      LAYER met4 ;
        RECT 2398.000 105.000 2406.000 129.965 ;
      LAYER met4 ;
        RECT 2406.000 105.000 2408.000 129.965 ;
      LAYER met4 ;
        RECT 2408.000 105.000 2411.000 129.965 ;
      LAYER met4 ;
        RECT 2411.000 105.000 2535.000 129.965 ;
      LAYER met4 ;
        RECT 2535.000 105.000 2553.000 129.965 ;
      LAYER met4 ;
        RECT 2553.000 105.000 2555.000 129.965 ;
      LAYER met4 ;
        RECT 2555.000 105.000 2563.000 129.965 ;
      LAYER met4 ;
        RECT 2563.000 105.000 2565.000 129.965 ;
      LAYER met4 ;
        RECT 2565.000 105.000 2568.000 129.965 ;
      LAYER met4 ;
        RECT 2568.000 105.000 2572.270 129.965 ;
        RECT 1827.730 0.000 1829.000 24.215 ;
      LAYER met4 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met4 ;
        RECT 2023.000 0.000 2024.270 24.215 ;
      LAYER met4 ;
        RECT 2024.670 0.000 2101.330 24.615 ;
        RECT 2103.000 24.215 2140.000 25.965 ;
        RECT 2260.000 24.215 2297.000 25.965 ;
        RECT 2298.030 24.615 2376.035 104.600 ;
        RECT 2377.000 102.965 2414.000 105.000 ;
        RECT 2534.000 102.965 2571.000 105.000 ;
        RECT 2572.670 104.600 2649.330 130.365 ;
        RECT 2651.000 129.965 2688.000 131.065 ;
        RECT 2808.000 129.965 2845.000 131.065 ;
        RECT 2845.965 130.365 2919.035 131.065 ;
      LAYER met4 ;
        RECT 2649.730 105.000 2652.000 129.965 ;
      LAYER met4 ;
        RECT 2652.000 105.000 2670.000 129.965 ;
      LAYER met4 ;
        RECT 2670.000 105.000 2672.000 129.965 ;
      LAYER met4 ;
        RECT 2672.000 105.000 2680.000 129.965 ;
      LAYER met4 ;
        RECT 2680.000 105.000 2682.000 129.965 ;
      LAYER met4 ;
        RECT 2682.000 105.000 2685.000 129.965 ;
      LAYER met4 ;
        RECT 2685.000 105.000 2809.000 129.965 ;
      LAYER met4 ;
        RECT 2809.000 105.000 2827.000 129.965 ;
      LAYER met4 ;
        RECT 2827.000 105.000 2829.000 129.965 ;
      LAYER met4 ;
        RECT 2829.000 105.000 2837.000 129.965 ;
      LAYER met4 ;
        RECT 2837.000 105.000 2839.000 129.965 ;
      LAYER met4 ;
        RECT 2839.000 105.000 2842.000 129.965 ;
      LAYER met4 ;
        RECT 2842.000 105.000 2846.270 129.965 ;
        RECT 2101.730 0.000 2103.000 24.215 ;
      LAYER met4 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met4 ;
        RECT 2297.000 0.000 2298.270 24.215 ;
      LAYER met4 ;
        RECT 2298.670 0.000 2375.330 24.615 ;
        RECT 2377.000 24.215 2414.000 25.965 ;
        RECT 2534.000 24.215 2571.000 25.965 ;
        RECT 2572.030 24.615 2650.035 104.600 ;
        RECT 2651.000 102.965 2688.000 105.000 ;
        RECT 2808.000 102.965 2845.000 105.000 ;
        RECT 2846.670 104.600 2918.330 130.365 ;
        RECT 2920.000 129.965 2957.000 131.065 ;
        RECT 3077.000 129.965 3114.000 131.065 ;
        RECT 3114.965 130.365 3188.035 131.065 ;
      LAYER met4 ;
        RECT 2918.730 105.000 2921.000 129.965 ;
      LAYER met4 ;
        RECT 2921.000 105.000 2939.000 129.965 ;
      LAYER met4 ;
        RECT 2939.000 105.000 2941.000 129.965 ;
      LAYER met4 ;
        RECT 2941.000 105.000 2949.000 129.965 ;
      LAYER met4 ;
        RECT 2949.000 105.000 2951.000 129.965 ;
      LAYER met4 ;
        RECT 2951.000 105.000 2954.000 129.965 ;
      LAYER met4 ;
        RECT 2954.000 105.000 3078.000 129.965 ;
      LAYER met4 ;
        RECT 3078.000 105.000 3096.000 129.965 ;
      LAYER met4 ;
        RECT 3096.000 105.000 3098.000 129.965 ;
      LAYER met4 ;
        RECT 3098.000 105.000 3106.000 129.965 ;
      LAYER met4 ;
        RECT 3106.000 105.000 3108.000 129.965 ;
      LAYER met4 ;
        RECT 3108.000 105.000 3111.000 129.965 ;
      LAYER met4 ;
        RECT 3111.000 105.000 3115.270 129.965 ;
        RECT 2375.730 0.000 2377.000 24.215 ;
      LAYER met4 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met4 ;
        RECT 2571.000 0.000 2572.270 24.215 ;
      LAYER met4 ;
        RECT 2572.670 0.000 2649.330 24.615 ;
        RECT 2651.000 24.215 2688.000 25.965 ;
        RECT 2808.000 24.215 2845.000 25.965 ;
        RECT 2845.965 24.615 2919.035 104.600 ;
        RECT 2920.000 102.965 2957.000 105.000 ;
        RECT 3077.000 102.965 3114.000 105.000 ;
        RECT 3115.670 104.600 3187.330 130.365 ;
        RECT 3189.000 129.965 3226.000 131.065 ;
        RECT 3346.000 129.965 3384.000 131.065 ;
        RECT 3385.255 130.365 3588.000 131.065 ;
      LAYER met4 ;
        RECT 3187.730 105.000 3190.000 129.965 ;
      LAYER met4 ;
        RECT 3190.000 105.000 3208.000 129.965 ;
      LAYER met4 ;
        RECT 3208.000 105.000 3210.000 129.965 ;
      LAYER met4 ;
        RECT 3210.000 105.000 3218.000 129.965 ;
      LAYER met4 ;
        RECT 3218.000 105.000 3220.000 129.965 ;
      LAYER met4 ;
        RECT 3220.000 105.000 3223.000 129.965 ;
      LAYER met4 ;
        RECT 3223.000 105.000 3347.000 129.965 ;
      LAYER met4 ;
        RECT 3347.000 105.000 3365.000 129.965 ;
      LAYER met4 ;
        RECT 3365.000 105.000 3367.000 129.965 ;
      LAYER met4 ;
        RECT 3367.000 105.000 3375.000 129.965 ;
      LAYER met4 ;
        RECT 3375.000 105.000 3377.000 129.965 ;
      LAYER met4 ;
        RECT 3377.000 105.000 3380.000 129.965 ;
      LAYER met4 ;
        RECT 3380.000 105.000 3385.855 129.965 ;
        RECT 2649.730 0.000 2651.000 24.215 ;
      LAYER met4 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met4 ;
        RECT 2845.000 0.000 2846.270 24.215 ;
      LAYER met4 ;
        RECT 2846.670 0.000 2918.330 24.615 ;
        RECT 2920.000 24.215 2957.000 25.965 ;
        RECT 3077.000 24.215 3114.000 25.965 ;
        RECT 3114.965 24.615 3188.035 104.600 ;
        RECT 3189.000 102.965 3226.000 105.000 ;
        RECT 3346.000 102.965 3384.000 105.000 ;
        RECT 3386.255 104.600 3588.000 130.365 ;
      LAYER met4 ;
        RECT 2918.730 0.000 2920.000 24.215 ;
      LAYER met4 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met4 ;
        RECT 3114.000 0.000 3115.270 24.215 ;
      LAYER met4 ;
        RECT 3115.670 0.000 3187.330 24.615 ;
        RECT 3189.000 24.215 3226.000 25.965 ;
        RECT 3346.000 24.215 3384.000 25.965 ;
        RECT 3385.255 24.615 3588.000 104.600 ;
      LAYER met4 ;
        RECT 3187.730 0.000 3189.000 24.215 ;
      LAYER met4 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met4 ;
        RECT 3384.000 0.000 3385.270 24.215 ;
      LAYER met4 ;
        RECT 3385.670 0.000 3588.000 24.615 ;
      LAYER met5 ;
        RECT 0.000 5084.585 204.000 5188.000 ;
      LAYER met5 ;
        RECT 204.000 5163.785 381.000 5188.000 ;
      LAYER met5 ;
        RECT 381.000 5156.610 461.000 5188.000 ;
      LAYER met5 ;
        RECT 461.000 5163.785 638.000 5188.000 ;
      LAYER met5 ;
        RECT 381.000 5090.960 390.600 5156.610 ;
        RECT 456.400 5090.960 461.000 5156.610 ;
        RECT 381.000 5084.585 461.000 5090.960 ;
        RECT 638.000 5156.610 718.000 5188.000 ;
      LAYER met5 ;
        RECT 718.000 5163.785 895.000 5188.000 ;
      LAYER met5 ;
        RECT 638.000 5090.960 647.600 5156.610 ;
        RECT 713.400 5090.960 718.000 5156.610 ;
        RECT 638.000 5084.585 718.000 5090.960 ;
        RECT 895.000 5156.610 975.000 5188.000 ;
      LAYER met5 ;
        RECT 975.000 5163.785 1152.000 5188.000 ;
      LAYER met5 ;
        RECT 895.000 5090.960 904.600 5156.610 ;
        RECT 970.400 5090.960 975.000 5156.610 ;
        RECT 895.000 5084.585 975.000 5090.960 ;
        RECT 1152.000 5156.610 1232.000 5188.000 ;
      LAYER met5 ;
        RECT 1232.000 5163.785 1410.000 5188.000 ;
      LAYER met5 ;
        RECT 1152.000 5090.960 1161.600 5156.610 ;
        RECT 1227.400 5090.960 1232.000 5156.610 ;
        RECT 1152.000 5084.585 1232.000 5090.960 ;
        RECT 1410.000 5156.610 1490.000 5188.000 ;
      LAYER met5 ;
        RECT 1490.000 5163.785 1667.000 5188.000 ;
      LAYER met5 ;
        RECT 1410.000 5090.960 1419.600 5156.610 ;
        RECT 1485.400 5090.960 1490.000 5156.610 ;
        RECT 1410.000 5084.585 1490.000 5090.960 ;
        RECT 1667.000 5155.545 1742.000 5188.000 ;
      LAYER met5 ;
        RECT 1742.000 5163.785 1919.000 5188.000 ;
      LAYER met5 ;
        RECT 1667.000 5091.520 1672.450 5155.545 ;
        RECT 1736.490 5091.520 1742.000 5155.545 ;
        RECT 1667.000 5084.585 1742.000 5091.520 ;
        RECT 1919.000 5156.610 1999.000 5188.000 ;
      LAYER met5 ;
        RECT 1999.000 5163.785 2364.000 5188.000 ;
      LAYER met5 ;
        RECT 1919.000 5090.960 1928.600 5156.610 ;
        RECT 1994.400 5090.960 1999.000 5156.610 ;
        RECT 1919.000 5084.585 1999.000 5090.960 ;
        RECT 2364.000 5156.610 2444.000 5188.000 ;
      LAYER met5 ;
        RECT 2444.000 5163.785 2621.000 5188.000 ;
      LAYER met5 ;
        RECT 2364.000 5090.960 2373.600 5156.610 ;
        RECT 2439.400 5090.960 2444.000 5156.610 ;
        RECT 2364.000 5084.585 2444.000 5090.960 ;
        RECT 2621.000 5156.610 2701.000 5188.000 ;
      LAYER met5 ;
        RECT 2701.000 5163.785 2878.000 5188.000 ;
      LAYER met5 ;
        RECT 2621.000 5090.960 2630.600 5156.610 ;
        RECT 2696.400 5090.960 2701.000 5156.610 ;
        RECT 2621.000 5084.585 2701.000 5090.960 ;
        RECT 2878.000 5155.545 2953.000 5188.000 ;
      LAYER met5 ;
        RECT 2953.000 5163.785 3130.000 5188.000 ;
      LAYER met5 ;
        RECT 2878.000 5091.520 2883.450 5155.545 ;
        RECT 2947.490 5091.520 2953.000 5155.545 ;
        RECT 2878.000 5084.585 2953.000 5091.520 ;
        RECT 3130.000 5156.610 3210.000 5188.000 ;
      LAYER met5 ;
        RECT 3210.000 5163.785 3388.000 5188.000 ;
      LAYER met5 ;
        RECT 3130.000 5090.960 3139.600 5156.610 ;
        RECT 3205.400 5090.960 3210.000 5156.610 ;
        RECT 3130.000 5084.585 3210.000 5090.960 ;
        RECT 3388.000 5084.585 3588.000 5188.000 ;
        RECT 0.000 5056.435 200.545 5084.585 ;
      LAYER met5 ;
        RECT 202.145 5058.035 205.000 5082.985 ;
      LAYER met5 ;
        RECT 206.600 5058.035 221.400 5082.985 ;
      LAYER met5 ;
        RECT 223.000 5058.035 225.000 5082.985 ;
      LAYER met5 ;
        RECT 226.600 5058.035 241.400 5082.985 ;
      LAYER met5 ;
        RECT 243.000 5058.035 245.000 5082.985 ;
      LAYER met5 ;
        RECT 246.600 5058.035 261.400 5082.985 ;
      LAYER met5 ;
        RECT 263.000 5058.035 265.000 5082.985 ;
      LAYER met5 ;
        RECT 266.600 5058.035 281.400 5082.985 ;
      LAYER met5 ;
        RECT 283.000 5058.035 285.000 5082.985 ;
      LAYER met5 ;
        RECT 286.600 5058.035 301.400 5082.985 ;
      LAYER met5 ;
        RECT 303.000 5058.035 305.000 5082.985 ;
      LAYER met5 ;
        RECT 306.600 5058.035 321.400 5082.985 ;
      LAYER met5 ;
        RECT 323.000 5058.035 325.000 5082.985 ;
      LAYER met5 ;
        RECT 326.600 5058.035 341.400 5082.985 ;
      LAYER met5 ;
        RECT 343.000 5058.035 345.000 5082.985 ;
      LAYER met5 ;
        RECT 346.600 5058.035 361.400 5082.985 ;
      LAYER met5 ;
        RECT 363.000 5058.035 365.000 5082.985 ;
      LAYER met5 ;
        RECT 366.600 5058.035 371.400 5082.985 ;
      LAYER met5 ;
        RECT 373.000 5058.035 375.000 5082.985 ;
        RECT 378.000 5058.035 382.270 5082.985 ;
      LAYER met5 ;
        RECT 0.000 5046.335 201.130 5056.435 ;
      LAYER met5 ;
        RECT 202.730 5052.185 382.270 5056.435 ;
        RECT 202.730 5046.335 382.270 5050.585 ;
      LAYER met5 ;
        RECT 0.000 5034.135 175.245 5046.335 ;
      LAYER met5 ;
        RECT 176.845 5035.735 382.270 5044.735 ;
      LAYER met5 ;
        RECT 0.000 5012.755 201.130 5034.135 ;
      LAYER met5 ;
        RECT 202.730 5029.685 382.270 5034.135 ;
        RECT 202.730 5024.840 382.270 5028.085 ;
        RECT 204.000 5024.835 381.000 5024.840 ;
        RECT 202.730 5019.985 382.270 5023.235 ;
        RECT 202.730 5013.935 382.270 5018.385 ;
      LAYER met5 ;
        RECT 0.000 4992.245 141.665 5012.755 ;
        RECT 0.000 4988.000 103.415 4992.245 ;
        RECT 131.565 4991.225 141.665 4992.245 ;
        RECT 131.565 4991.080 135.815 4991.225 ;
      LAYER met5 ;
        RECT 0.000 4851.000 24.215 4988.000 ;
        RECT 105.015 4985.000 129.965 4990.645 ;
        RECT 105.015 4980.000 129.965 4982.000 ;
      LAYER met5 ;
        RECT 105.015 4973.600 129.965 4978.400 ;
      LAYER met5 ;
        RECT 105.015 4970.000 129.965 4972.000 ;
      LAYER met5 ;
        RECT 105.015 4953.600 129.965 4968.400 ;
      LAYER met5 ;
        RECT 105.015 4950.000 129.965 4952.000 ;
      LAYER met5 ;
        RECT 105.015 4933.600 129.965 4948.400 ;
      LAYER met5 ;
        RECT 105.015 4930.000 129.965 4932.000 ;
      LAYER met5 ;
        RECT 105.015 4913.600 129.965 4928.400 ;
      LAYER met5 ;
        RECT 105.015 4910.000 129.965 4912.000 ;
      LAYER met5 ;
        RECT 105.015 4893.600 129.965 4908.400 ;
      LAYER met5 ;
        RECT 105.015 4890.000 129.965 4892.000 ;
      LAYER met5 ;
        RECT 105.015 4873.600 129.965 4888.400 ;
      LAYER met5 ;
        RECT 105.015 4870.000 129.965 4872.000 ;
      LAYER met5 ;
        RECT 105.015 4853.600 129.965 4868.400 ;
        RECT 0.000 4848.130 103.415 4851.000 ;
      LAYER met5 ;
        RECT 105.015 4849.730 129.965 4852.000 ;
        RECT 131.565 4849.730 135.815 4989.480 ;
        RECT 137.415 4849.730 141.665 4989.625 ;
        RECT 143.265 4849.730 152.265 5011.155 ;
      LAYER met5 ;
        RECT 153.865 5006.285 201.130 5012.755 ;
      LAYER met5 ;
        RECT 202.730 5007.885 382.270 5012.335 ;
      LAYER met5 ;
        RECT 383.870 5006.285 458.130 5084.585 ;
      LAYER met5 ;
        RECT 459.730 5058.035 462.000 5082.985 ;
      LAYER met5 ;
        RECT 463.600 5058.035 478.400 5082.985 ;
      LAYER met5 ;
        RECT 480.000 5058.035 482.000 5082.985 ;
      LAYER met5 ;
        RECT 483.600 5058.035 498.400 5082.985 ;
      LAYER met5 ;
        RECT 500.000 5058.035 502.000 5082.985 ;
      LAYER met5 ;
        RECT 503.600 5058.035 518.400 5082.985 ;
      LAYER met5 ;
        RECT 520.000 5058.035 522.000 5082.985 ;
      LAYER met5 ;
        RECT 523.600 5058.035 538.400 5082.985 ;
      LAYER met5 ;
        RECT 540.000 5058.035 542.000 5082.985 ;
      LAYER met5 ;
        RECT 543.600 5058.035 558.400 5082.985 ;
      LAYER met5 ;
        RECT 560.000 5058.035 562.000 5082.985 ;
      LAYER met5 ;
        RECT 563.600 5058.035 578.400 5082.985 ;
      LAYER met5 ;
        RECT 580.000 5058.035 582.000 5082.985 ;
      LAYER met5 ;
        RECT 583.600 5058.035 598.400 5082.985 ;
      LAYER met5 ;
        RECT 600.000 5058.035 602.000 5082.985 ;
      LAYER met5 ;
        RECT 603.600 5058.035 618.400 5082.985 ;
      LAYER met5 ;
        RECT 620.000 5058.035 622.000 5082.985 ;
      LAYER met5 ;
        RECT 623.600 5058.035 628.400 5082.985 ;
      LAYER met5 ;
        RECT 630.000 5058.035 632.000 5082.985 ;
        RECT 635.000 5058.035 639.270 5082.985 ;
        RECT 459.730 5052.185 639.270 5056.435 ;
        RECT 459.730 5046.335 639.270 5050.585 ;
        RECT 459.730 5035.735 639.270 5044.735 ;
        RECT 459.730 5029.685 639.270 5034.135 ;
        RECT 459.730 5024.840 639.270 5028.085 ;
        RECT 461.000 5024.835 638.000 5024.840 ;
        RECT 459.730 5019.985 639.270 5023.235 ;
        RECT 459.730 5013.935 639.270 5018.385 ;
        RECT 459.730 5007.885 639.270 5012.335 ;
      LAYER met5 ;
        RECT 640.870 5006.285 715.130 5084.585 ;
      LAYER met5 ;
        RECT 716.730 5058.035 719.000 5082.985 ;
      LAYER met5 ;
        RECT 720.600 5058.035 735.400 5082.985 ;
      LAYER met5 ;
        RECT 737.000 5058.035 739.000 5082.985 ;
      LAYER met5 ;
        RECT 740.600 5058.035 755.400 5082.985 ;
      LAYER met5 ;
        RECT 757.000 5058.035 759.000 5082.985 ;
      LAYER met5 ;
        RECT 760.600 5058.035 775.400 5082.985 ;
      LAYER met5 ;
        RECT 777.000 5058.035 779.000 5082.985 ;
      LAYER met5 ;
        RECT 780.600 5058.035 795.400 5082.985 ;
      LAYER met5 ;
        RECT 797.000 5058.035 799.000 5082.985 ;
      LAYER met5 ;
        RECT 800.600 5058.035 815.400 5082.985 ;
      LAYER met5 ;
        RECT 817.000 5058.035 819.000 5082.985 ;
      LAYER met5 ;
        RECT 820.600 5058.035 835.400 5082.985 ;
      LAYER met5 ;
        RECT 837.000 5058.035 839.000 5082.985 ;
      LAYER met5 ;
        RECT 840.600 5058.035 855.400 5082.985 ;
      LAYER met5 ;
        RECT 857.000 5058.035 859.000 5082.985 ;
      LAYER met5 ;
        RECT 860.600 5058.035 875.400 5082.985 ;
      LAYER met5 ;
        RECT 877.000 5058.035 879.000 5082.985 ;
      LAYER met5 ;
        RECT 880.600 5058.035 885.400 5082.985 ;
      LAYER met5 ;
        RECT 887.000 5058.035 889.000 5082.985 ;
        RECT 892.000 5058.035 896.270 5082.985 ;
        RECT 716.730 5052.185 896.270 5056.435 ;
        RECT 716.730 5046.335 896.270 5050.585 ;
        RECT 716.730 5035.735 896.270 5044.735 ;
        RECT 716.730 5029.685 896.270 5034.135 ;
        RECT 716.730 5024.840 896.270 5028.085 ;
        RECT 718.000 5024.835 895.000 5024.840 ;
        RECT 716.730 5019.985 896.270 5023.235 ;
        RECT 716.730 5013.935 896.270 5018.385 ;
        RECT 716.730 5007.885 896.270 5012.335 ;
      LAYER met5 ;
        RECT 897.870 5006.285 972.130 5084.585 ;
      LAYER met5 ;
        RECT 973.730 5058.035 976.000 5082.985 ;
      LAYER met5 ;
        RECT 977.600 5058.035 992.400 5082.985 ;
      LAYER met5 ;
        RECT 994.000 5058.035 996.000 5082.985 ;
      LAYER met5 ;
        RECT 997.600 5058.035 1012.400 5082.985 ;
      LAYER met5 ;
        RECT 1014.000 5058.035 1016.000 5082.985 ;
      LAYER met5 ;
        RECT 1017.600 5058.035 1032.400 5082.985 ;
      LAYER met5 ;
        RECT 1034.000 5058.035 1036.000 5082.985 ;
      LAYER met5 ;
        RECT 1037.600 5058.035 1052.400 5082.985 ;
      LAYER met5 ;
        RECT 1054.000 5058.035 1056.000 5082.985 ;
      LAYER met5 ;
        RECT 1057.600 5058.035 1072.400 5082.985 ;
      LAYER met5 ;
        RECT 1074.000 5058.035 1076.000 5082.985 ;
      LAYER met5 ;
        RECT 1077.600 5058.035 1092.400 5082.985 ;
      LAYER met5 ;
        RECT 1094.000 5058.035 1096.000 5082.985 ;
      LAYER met5 ;
        RECT 1097.600 5058.035 1112.400 5082.985 ;
      LAYER met5 ;
        RECT 1114.000 5058.035 1116.000 5082.985 ;
      LAYER met5 ;
        RECT 1117.600 5058.035 1132.400 5082.985 ;
      LAYER met5 ;
        RECT 1134.000 5058.035 1136.000 5082.985 ;
      LAYER met5 ;
        RECT 1137.600 5058.035 1142.400 5082.985 ;
      LAYER met5 ;
        RECT 1144.000 5058.035 1146.000 5082.985 ;
        RECT 1149.000 5058.035 1153.270 5082.985 ;
        RECT 973.730 5052.185 1153.270 5056.435 ;
        RECT 973.730 5046.335 1153.270 5050.585 ;
        RECT 973.730 5035.735 1153.270 5044.735 ;
        RECT 973.730 5029.685 1153.270 5034.135 ;
        RECT 973.730 5024.840 1153.270 5028.085 ;
        RECT 975.000 5024.835 1152.000 5024.840 ;
        RECT 973.730 5019.985 1153.270 5023.235 ;
        RECT 973.730 5013.935 1153.270 5018.385 ;
        RECT 973.730 5007.885 1153.270 5012.335 ;
      LAYER met5 ;
        RECT 1154.870 5006.285 1229.130 5084.585 ;
      LAYER met5 ;
        RECT 1230.730 5058.035 1233.000 5082.985 ;
      LAYER met5 ;
        RECT 1234.600 5058.035 1249.400 5082.985 ;
      LAYER met5 ;
        RECT 1251.000 5058.035 1253.000 5082.985 ;
      LAYER met5 ;
        RECT 1254.600 5058.035 1269.400 5082.985 ;
      LAYER met5 ;
        RECT 1271.000 5058.035 1273.000 5082.985 ;
      LAYER met5 ;
        RECT 1274.600 5058.035 1289.400 5082.985 ;
      LAYER met5 ;
        RECT 1291.000 5058.035 1293.000 5082.985 ;
      LAYER met5 ;
        RECT 1294.600 5058.035 1309.400 5082.985 ;
      LAYER met5 ;
        RECT 1311.000 5058.035 1313.000 5082.985 ;
      LAYER met5 ;
        RECT 1314.600 5058.035 1329.400 5082.985 ;
      LAYER met5 ;
        RECT 1331.000 5058.035 1333.000 5082.985 ;
      LAYER met5 ;
        RECT 1334.600 5058.035 1349.400 5082.985 ;
      LAYER met5 ;
        RECT 1351.000 5058.035 1353.000 5082.985 ;
      LAYER met5 ;
        RECT 1354.600 5058.035 1369.400 5082.985 ;
      LAYER met5 ;
        RECT 1371.000 5058.035 1373.000 5082.985 ;
      LAYER met5 ;
        RECT 1374.600 5058.035 1389.400 5082.985 ;
      LAYER met5 ;
        RECT 1391.000 5058.035 1393.000 5082.985 ;
      LAYER met5 ;
        RECT 1394.600 5058.035 1399.400 5082.985 ;
      LAYER met5 ;
        RECT 1401.000 5058.035 1403.000 5082.985 ;
        RECT 1406.000 5058.035 1411.270 5082.985 ;
        RECT 1230.730 5052.185 1411.270 5056.435 ;
        RECT 1230.730 5046.335 1411.270 5050.585 ;
        RECT 1230.730 5035.735 1411.270 5044.735 ;
        RECT 1230.730 5029.685 1411.270 5034.135 ;
        RECT 1230.730 5024.840 1411.270 5028.085 ;
        RECT 1232.000 5024.835 1410.000 5024.840 ;
        RECT 1230.730 5019.985 1411.270 5023.235 ;
        RECT 1230.730 5013.935 1411.270 5018.385 ;
        RECT 1230.730 5007.885 1411.270 5012.335 ;
      LAYER met5 ;
        RECT 1412.870 5006.285 1487.130 5084.585 ;
      LAYER met5 ;
        RECT 1488.730 5058.035 1491.000 5082.985 ;
      LAYER met5 ;
        RECT 1492.600 5058.035 1507.400 5082.985 ;
      LAYER met5 ;
        RECT 1509.000 5058.035 1511.000 5082.985 ;
      LAYER met5 ;
        RECT 1512.600 5058.035 1527.400 5082.985 ;
      LAYER met5 ;
        RECT 1529.000 5058.035 1531.000 5082.985 ;
      LAYER met5 ;
        RECT 1532.600 5058.035 1547.400 5082.985 ;
      LAYER met5 ;
        RECT 1549.000 5058.035 1551.000 5082.985 ;
      LAYER met5 ;
        RECT 1552.600 5058.035 1567.400 5082.985 ;
      LAYER met5 ;
        RECT 1569.000 5058.035 1571.000 5082.985 ;
      LAYER met5 ;
        RECT 1572.600 5058.035 1587.400 5082.985 ;
      LAYER met5 ;
        RECT 1589.000 5058.035 1591.000 5082.985 ;
      LAYER met5 ;
        RECT 1592.600 5058.035 1607.400 5082.985 ;
      LAYER met5 ;
        RECT 1609.000 5058.035 1611.000 5082.985 ;
      LAYER met5 ;
        RECT 1612.600 5058.035 1627.400 5082.985 ;
      LAYER met5 ;
        RECT 1629.000 5058.035 1631.000 5082.985 ;
      LAYER met5 ;
        RECT 1632.600 5058.035 1647.400 5082.985 ;
      LAYER met5 ;
        RECT 1649.000 5058.035 1651.000 5082.985 ;
      LAYER met5 ;
        RECT 1652.600 5058.035 1657.400 5082.985 ;
      LAYER met5 ;
        RECT 1659.000 5058.035 1661.000 5082.985 ;
        RECT 1664.000 5058.035 1668.270 5082.985 ;
        RECT 1488.730 5052.185 1668.270 5056.435 ;
        RECT 1488.730 5046.335 1668.270 5050.585 ;
        RECT 1488.730 5035.735 1668.270 5044.735 ;
        RECT 1488.730 5029.685 1668.270 5034.135 ;
        RECT 1488.730 5024.840 1668.270 5028.085 ;
      LAYER met5 ;
        RECT 1669.870 5024.840 1739.130 5084.585 ;
      LAYER met5 ;
        RECT 1740.730 5058.035 1743.000 5082.985 ;
      LAYER met5 ;
        RECT 1744.600 5058.035 1759.400 5082.985 ;
      LAYER met5 ;
        RECT 1761.000 5058.035 1763.000 5082.985 ;
      LAYER met5 ;
        RECT 1764.600 5058.035 1779.400 5082.985 ;
      LAYER met5 ;
        RECT 1781.000 5058.035 1783.000 5082.985 ;
      LAYER met5 ;
        RECT 1784.600 5058.035 1799.400 5082.985 ;
      LAYER met5 ;
        RECT 1801.000 5058.035 1803.000 5082.985 ;
      LAYER met5 ;
        RECT 1804.600 5058.035 1819.400 5082.985 ;
      LAYER met5 ;
        RECT 1821.000 5058.035 1823.000 5082.985 ;
      LAYER met5 ;
        RECT 1824.600 5058.035 1839.400 5082.985 ;
      LAYER met5 ;
        RECT 1841.000 5058.035 1843.000 5082.985 ;
      LAYER met5 ;
        RECT 1844.600 5058.035 1859.400 5082.985 ;
      LAYER met5 ;
        RECT 1861.000 5058.035 1863.000 5082.985 ;
      LAYER met5 ;
        RECT 1864.600 5058.035 1879.400 5082.985 ;
      LAYER met5 ;
        RECT 1881.000 5058.035 1883.000 5082.985 ;
      LAYER met5 ;
        RECT 1884.600 5058.035 1899.400 5082.985 ;
      LAYER met5 ;
        RECT 1901.000 5058.035 1903.000 5082.985 ;
      LAYER met5 ;
        RECT 1904.600 5058.035 1909.400 5082.985 ;
      LAYER met5 ;
        RECT 1911.000 5058.035 1913.000 5082.985 ;
        RECT 1916.000 5058.035 1920.270 5082.985 ;
        RECT 1740.730 5052.185 1920.270 5056.435 ;
        RECT 1740.730 5046.335 1920.270 5050.585 ;
        RECT 1740.730 5035.735 1920.270 5044.735 ;
        RECT 1740.730 5029.685 1920.270 5034.135 ;
        RECT 1740.730 5024.840 1920.270 5028.085 ;
        RECT 1490.000 5024.835 1667.000 5024.840 ;
      LAYER met5 ;
        RECT 1667.000 5024.835 1742.000 5024.840 ;
      LAYER met5 ;
        RECT 1742.000 5024.835 1919.000 5024.840 ;
        RECT 1488.730 5019.985 1668.270 5023.235 ;
        RECT 1488.730 5007.885 1668.270 5012.335 ;
      LAYER met5 ;
        RECT 1669.870 5006.285 1739.130 5024.835 ;
      LAYER met5 ;
        RECT 1740.730 5019.985 1920.270 5023.235 ;
        RECT 1740.730 5007.885 1920.270 5012.335 ;
      LAYER met5 ;
        RECT 1921.870 5006.285 1996.130 5084.585 ;
      LAYER met5 ;
        RECT 1997.730 5058.035 2000.000 5082.985 ;
      LAYER met5 ;
        RECT 2001.600 5058.035 2016.400 5082.985 ;
      LAYER met5 ;
        RECT 2018.000 5058.035 2020.000 5082.985 ;
      LAYER met5 ;
        RECT 2021.600 5058.035 2036.400 5082.985 ;
      LAYER met5 ;
        RECT 2038.000 5058.035 2040.000 5082.985 ;
      LAYER met5 ;
        RECT 2041.600 5058.035 2056.400 5082.985 ;
      LAYER met5 ;
        RECT 2058.000 5058.035 2060.000 5082.985 ;
      LAYER met5 ;
        RECT 2061.600 5058.035 2076.400 5082.985 ;
      LAYER met5 ;
        RECT 2078.000 5058.035 2080.000 5082.985 ;
      LAYER met5 ;
        RECT 2081.600 5058.035 2096.400 5082.985 ;
      LAYER met5 ;
        RECT 2098.000 5058.035 2100.000 5082.985 ;
      LAYER met5 ;
        RECT 2101.600 5058.035 2116.400 5082.985 ;
      LAYER met5 ;
        RECT 2118.000 5058.035 2120.000 5082.985 ;
      LAYER met5 ;
        RECT 2121.600 5058.035 2136.400 5082.985 ;
      LAYER met5 ;
        RECT 2138.000 5058.035 2140.000 5082.985 ;
      LAYER met5 ;
        RECT 2141.600 5058.035 2156.400 5082.985 ;
      LAYER met5 ;
        RECT 2158.000 5058.035 2160.000 5082.985 ;
      LAYER met5 ;
        RECT 2161.600 5058.035 2166.400 5082.985 ;
      LAYER met5 ;
        RECT 2168.000 5058.035 2170.000 5082.985 ;
        RECT 2173.000 5058.035 2187.000 5082.985 ;
      LAYER met5 ;
        RECT 2188.600 5058.035 2203.400 5082.985 ;
      LAYER met5 ;
        RECT 2205.000 5058.035 2207.000 5082.985 ;
      LAYER met5 ;
        RECT 2208.600 5058.035 2223.400 5082.985 ;
      LAYER met5 ;
        RECT 2225.000 5058.035 2227.000 5082.985 ;
      LAYER met5 ;
        RECT 2228.600 5058.035 2243.400 5082.985 ;
      LAYER met5 ;
        RECT 2245.000 5058.035 2247.000 5082.985 ;
      LAYER met5 ;
        RECT 2248.600 5058.035 2263.400 5082.985 ;
      LAYER met5 ;
        RECT 2265.000 5058.035 2267.000 5082.985 ;
      LAYER met5 ;
        RECT 2268.600 5058.035 2283.400 5082.985 ;
      LAYER met5 ;
        RECT 2285.000 5058.035 2287.000 5082.985 ;
      LAYER met5 ;
        RECT 2288.600 5058.035 2303.400 5082.985 ;
      LAYER met5 ;
        RECT 2305.000 5058.035 2307.000 5082.985 ;
      LAYER met5 ;
        RECT 2308.600 5058.035 2323.400 5082.985 ;
      LAYER met5 ;
        RECT 2325.000 5058.035 2327.000 5082.985 ;
      LAYER met5 ;
        RECT 2328.600 5058.035 2343.400 5082.985 ;
      LAYER met5 ;
        RECT 2345.000 5058.035 2347.000 5082.985 ;
      LAYER met5 ;
        RECT 2348.600 5058.035 2353.400 5082.985 ;
      LAYER met5 ;
        RECT 2355.000 5058.035 2357.000 5082.985 ;
        RECT 2360.000 5058.035 2365.270 5082.985 ;
        RECT 1997.730 5052.185 2365.270 5056.435 ;
        RECT 1997.730 5046.335 2365.270 5050.585 ;
        RECT 1997.730 5035.735 2176.000 5044.735 ;
        RECT 2181.000 5035.735 2365.270 5044.735 ;
        RECT 1997.730 5029.685 2181.000 5034.135 ;
        RECT 2186.000 5029.685 2365.270 5034.135 ;
        RECT 1997.730 5024.840 2176.000 5028.085 ;
        RECT 1999.000 5024.835 2176.000 5024.840 ;
        RECT 2181.000 5024.840 2365.270 5028.085 ;
        RECT 2181.000 5024.835 2364.000 5024.840 ;
        RECT 1997.730 5019.985 2365.270 5023.235 ;
        RECT 1997.730 5013.935 2365.270 5018.385 ;
        RECT 1997.730 5007.885 2365.270 5012.335 ;
      LAYER met5 ;
        RECT 2366.870 5006.285 2441.130 5084.585 ;
      LAYER met5 ;
        RECT 2442.730 5058.035 2445.000 5082.985 ;
      LAYER met5 ;
        RECT 2446.600 5058.035 2461.400 5082.985 ;
      LAYER met5 ;
        RECT 2463.000 5058.035 2465.000 5082.985 ;
      LAYER met5 ;
        RECT 2466.600 5058.035 2481.400 5082.985 ;
      LAYER met5 ;
        RECT 2483.000 5058.035 2485.000 5082.985 ;
      LAYER met5 ;
        RECT 2486.600 5058.035 2501.400 5082.985 ;
      LAYER met5 ;
        RECT 2503.000 5058.035 2505.000 5082.985 ;
      LAYER met5 ;
        RECT 2506.600 5058.035 2521.400 5082.985 ;
      LAYER met5 ;
        RECT 2523.000 5058.035 2525.000 5082.985 ;
      LAYER met5 ;
        RECT 2526.600 5058.035 2541.400 5082.985 ;
      LAYER met5 ;
        RECT 2543.000 5058.035 2545.000 5082.985 ;
      LAYER met5 ;
        RECT 2546.600 5058.035 2561.400 5082.985 ;
      LAYER met5 ;
        RECT 2563.000 5058.035 2565.000 5082.985 ;
      LAYER met5 ;
        RECT 2566.600 5058.035 2581.400 5082.985 ;
      LAYER met5 ;
        RECT 2583.000 5058.035 2585.000 5082.985 ;
      LAYER met5 ;
        RECT 2586.600 5058.035 2601.400 5082.985 ;
      LAYER met5 ;
        RECT 2603.000 5058.035 2605.000 5082.985 ;
      LAYER met5 ;
        RECT 2606.600 5058.035 2611.400 5082.985 ;
      LAYER met5 ;
        RECT 2613.000 5058.035 2615.000 5082.985 ;
        RECT 2618.000 5058.035 2622.270 5082.985 ;
        RECT 2442.730 5052.185 2622.270 5056.435 ;
        RECT 2442.730 5046.335 2622.270 5050.585 ;
        RECT 2442.730 5035.735 2622.270 5044.735 ;
        RECT 2442.730 5029.685 2622.270 5034.135 ;
        RECT 2442.730 5024.840 2622.270 5028.085 ;
        RECT 2444.000 5024.835 2621.000 5024.840 ;
        RECT 2442.730 5019.985 2622.270 5023.235 ;
        RECT 2442.730 5013.935 2622.270 5018.385 ;
        RECT 2442.730 5007.885 2622.270 5012.335 ;
      LAYER met5 ;
        RECT 2623.870 5006.285 2698.130 5084.585 ;
      LAYER met5 ;
        RECT 2699.730 5058.035 2702.000 5082.985 ;
      LAYER met5 ;
        RECT 2703.600 5058.035 2718.400 5082.985 ;
      LAYER met5 ;
        RECT 2720.000 5058.035 2722.000 5082.985 ;
      LAYER met5 ;
        RECT 2723.600 5058.035 2738.400 5082.985 ;
      LAYER met5 ;
        RECT 2740.000 5058.035 2742.000 5082.985 ;
      LAYER met5 ;
        RECT 2743.600 5058.035 2758.400 5082.985 ;
      LAYER met5 ;
        RECT 2760.000 5058.035 2762.000 5082.985 ;
      LAYER met5 ;
        RECT 2763.600 5058.035 2778.400 5082.985 ;
      LAYER met5 ;
        RECT 2780.000 5058.035 2782.000 5082.985 ;
      LAYER met5 ;
        RECT 2783.600 5058.035 2798.400 5082.985 ;
      LAYER met5 ;
        RECT 2800.000 5058.035 2802.000 5082.985 ;
      LAYER met5 ;
        RECT 2803.600 5058.035 2818.400 5082.985 ;
      LAYER met5 ;
        RECT 2820.000 5058.035 2822.000 5082.985 ;
      LAYER met5 ;
        RECT 2823.600 5058.035 2838.400 5082.985 ;
      LAYER met5 ;
        RECT 2840.000 5058.035 2842.000 5082.985 ;
      LAYER met5 ;
        RECT 2843.600 5058.035 2858.400 5082.985 ;
      LAYER met5 ;
        RECT 2860.000 5058.035 2862.000 5082.985 ;
      LAYER met5 ;
        RECT 2863.600 5058.035 2868.400 5082.985 ;
      LAYER met5 ;
        RECT 2870.000 5058.035 2872.000 5082.985 ;
        RECT 2875.000 5058.035 2879.270 5082.985 ;
        RECT 2699.730 5052.185 2879.270 5056.435 ;
        RECT 2699.730 5046.335 2879.270 5050.585 ;
        RECT 2699.730 5029.685 2879.270 5034.135 ;
      LAYER met5 ;
        RECT 2880.870 5024.840 2950.130 5084.585 ;
      LAYER met5 ;
        RECT 2951.730 5058.035 2954.000 5082.985 ;
      LAYER met5 ;
        RECT 2955.600 5058.035 2970.400 5082.985 ;
      LAYER met5 ;
        RECT 2972.000 5058.035 2974.000 5082.985 ;
      LAYER met5 ;
        RECT 2975.600 5058.035 2990.400 5082.985 ;
      LAYER met5 ;
        RECT 2992.000 5058.035 2994.000 5082.985 ;
      LAYER met5 ;
        RECT 2995.600 5058.035 3010.400 5082.985 ;
      LAYER met5 ;
        RECT 3012.000 5058.035 3014.000 5082.985 ;
      LAYER met5 ;
        RECT 3015.600 5058.035 3030.400 5082.985 ;
      LAYER met5 ;
        RECT 3032.000 5058.035 3034.000 5082.985 ;
      LAYER met5 ;
        RECT 3035.600 5058.035 3050.400 5082.985 ;
      LAYER met5 ;
        RECT 3052.000 5058.035 3054.000 5082.985 ;
      LAYER met5 ;
        RECT 3055.600 5058.035 3070.400 5082.985 ;
      LAYER met5 ;
        RECT 3072.000 5058.035 3074.000 5082.985 ;
      LAYER met5 ;
        RECT 3075.600 5058.035 3090.400 5082.985 ;
      LAYER met5 ;
        RECT 3092.000 5058.035 3094.000 5082.985 ;
      LAYER met5 ;
        RECT 3095.600 5058.035 3110.400 5082.985 ;
      LAYER met5 ;
        RECT 3112.000 5058.035 3114.000 5082.985 ;
      LAYER met5 ;
        RECT 3115.600 5058.035 3120.400 5082.985 ;
      LAYER met5 ;
        RECT 3122.000 5058.035 3124.000 5082.985 ;
        RECT 3127.000 5058.035 3131.270 5082.985 ;
        RECT 2951.730 5052.185 3131.270 5056.435 ;
        RECT 2951.730 5046.335 3131.270 5050.585 ;
        RECT 2951.730 5029.685 3131.270 5034.135 ;
      LAYER met5 ;
        RECT 2878.000 5024.835 2953.000 5024.840 ;
      LAYER met5 ;
        RECT 2699.730 5019.985 2879.270 5023.235 ;
        RECT 2699.730 5013.935 2879.270 5018.385 ;
        RECT 2699.730 5007.885 2879.270 5012.335 ;
      LAYER met5 ;
        RECT 2880.870 5006.285 2950.130 5024.835 ;
      LAYER met5 ;
        RECT 2951.730 5019.985 3131.270 5023.235 ;
        RECT 2951.730 5013.935 3131.270 5018.385 ;
        RECT 2951.730 5007.885 3131.270 5012.335 ;
      LAYER met5 ;
        RECT 3132.870 5006.285 3207.130 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5058.035 3211.000 5082.985 ;
      LAYER met5 ;
        RECT 3212.600 5058.035 3227.400 5082.985 ;
      LAYER met5 ;
        RECT 3229.000 5058.035 3231.000 5082.985 ;
      LAYER met5 ;
        RECT 3232.600 5058.035 3247.400 5082.985 ;
      LAYER met5 ;
        RECT 3249.000 5058.035 3251.000 5082.985 ;
      LAYER met5 ;
        RECT 3252.600 5058.035 3267.400 5082.985 ;
      LAYER met5 ;
        RECT 3269.000 5058.035 3271.000 5082.985 ;
      LAYER met5 ;
        RECT 3272.600 5058.035 3287.400 5082.985 ;
      LAYER met5 ;
        RECT 3289.000 5058.035 3291.000 5082.985 ;
      LAYER met5 ;
        RECT 3292.600 5058.035 3307.400 5082.985 ;
      LAYER met5 ;
        RECT 3309.000 5058.035 3311.000 5082.985 ;
      LAYER met5 ;
        RECT 3312.600 5058.035 3327.400 5082.985 ;
      LAYER met5 ;
        RECT 3329.000 5058.035 3331.000 5082.985 ;
      LAYER met5 ;
        RECT 3332.600 5058.035 3347.400 5082.985 ;
      LAYER met5 ;
        RECT 3349.000 5058.035 3351.000 5082.985 ;
      LAYER met5 ;
        RECT 3352.600 5058.035 3367.400 5082.985 ;
      LAYER met5 ;
        RECT 3369.000 5058.035 3371.000 5082.985 ;
      LAYER met5 ;
        RECT 3372.600 5058.035 3377.400 5082.985 ;
      LAYER met5 ;
        RECT 3379.000 5058.035 3381.000 5082.985 ;
        RECT 3384.000 5058.035 3390.645 5082.985 ;
      LAYER met5 ;
        RECT 3392.245 5056.435 3588.000 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5052.185 3389.480 5056.435 ;
      LAYER met5 ;
        RECT 3391.080 5052.185 3588.000 5056.435 ;
      LAYER met5 ;
        RECT 3208.730 5046.335 3389.625 5050.585 ;
      LAYER met5 ;
        RECT 3391.225 5046.335 3588.000 5052.185 ;
      LAYER met5 ;
        RECT 3208.730 5035.735 3411.155 5044.735 ;
      LAYER met5 ;
        RECT 3412.755 5034.135 3588.000 5046.335 ;
      LAYER met5 ;
        RECT 3208.730 5029.685 3389.475 5034.135 ;
      LAYER met5 ;
        RECT 3391.075 5028.085 3588.000 5034.135 ;
      LAYER met5 ;
        RECT 3208.730 5024.840 3389.335 5028.085 ;
        RECT 3210.000 5024.835 3389.335 5024.840 ;
      LAYER met5 ;
        RECT 3390.935 5024.835 3588.000 5028.085 ;
      LAYER met5 ;
        RECT 3208.730 5019.985 3389.385 5023.235 ;
      LAYER met5 ;
        RECT 3390.985 5019.985 3588.000 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5013.935 3389.600 5018.385 ;
      LAYER met5 ;
        RECT 3391.200 5012.755 3588.000 5019.985 ;
        RECT 3391.200 5012.335 3434.135 5012.755 ;
      LAYER met5 ;
        RECT 3208.730 5007.885 3389.525 5012.335 ;
      LAYER met5 ;
        RECT 3391.125 5006.285 3434.135 5012.335 ;
        RECT 153.865 5003.035 201.145 5006.285 ;
      LAYER met5 ;
        RECT 202.745 5003.035 381.965 5006.285 ;
      LAYER met5 ;
        RECT 383.565 5003.035 458.370 5006.285 ;
      LAYER met5 ;
        RECT 459.970 5003.035 638.965 5006.285 ;
      LAYER met5 ;
        RECT 640.565 5003.035 715.370 5006.285 ;
      LAYER met5 ;
        RECT 716.970 5003.035 895.965 5006.285 ;
      LAYER met5 ;
        RECT 897.565 5003.035 972.370 5006.285 ;
      LAYER met5 ;
        RECT 973.970 5003.035 1152.965 5006.285 ;
      LAYER met5 ;
        RECT 1154.565 5003.035 1229.370 5006.285 ;
      LAYER met5 ;
        RECT 1230.970 5003.035 1410.965 5006.285 ;
      LAYER met5 ;
        RECT 1412.565 5003.035 1487.370 5006.285 ;
      LAYER met5 ;
        RECT 1488.970 5003.035 1667.965 5006.285 ;
      LAYER met5 ;
        RECT 1669.565 5003.035 1739.435 5006.285 ;
      LAYER met5 ;
        RECT 1741.035 5003.035 1919.965 5006.285 ;
      LAYER met5 ;
        RECT 1921.565 5003.035 1996.370 5006.285 ;
      LAYER met5 ;
        RECT 1997.970 5003.035 2176.000 5006.285 ;
        RECT 2181.000 5003.035 2364.965 5006.285 ;
      LAYER met5 ;
        RECT 2366.565 5003.035 2441.370 5006.285 ;
      LAYER met5 ;
        RECT 2442.970 5003.035 2621.965 5006.285 ;
      LAYER met5 ;
        RECT 2623.565 5003.035 2698.370 5006.285 ;
      LAYER met5 ;
        RECT 2699.970 5003.035 2878.965 5006.285 ;
      LAYER met5 ;
        RECT 2880.565 5003.035 2950.435 5006.285 ;
      LAYER met5 ;
        RECT 2952.035 5003.035 3130.965 5006.285 ;
      LAYER met5 ;
        RECT 3132.565 5003.035 3207.370 5006.285 ;
      LAYER met5 ;
        RECT 3208.970 5003.035 3389.470 5006.285 ;
      LAYER met5 ;
        RECT 3391.070 5003.035 3434.135 5006.285 ;
        RECT 153.865 4993.385 201.130 5003.035 ;
      LAYER met5 ;
        RECT 202.730 4996.985 382.270 5001.435 ;
      LAYER met5 ;
        RECT 153.865 4991.200 184.965 4993.385 ;
        RECT 192.615 4991.950 201.130 4993.385 ;
        RECT 153.865 4991.075 168.015 4991.200 ;
        RECT 175.665 4991.125 184.965 4991.200 ;
        RECT 159.915 4990.985 168.015 4991.075 ;
        RECT 181.715 4991.070 184.965 4991.125 ;
        RECT 159.915 4990.935 163.165 4990.985 ;
      LAYER met5 ;
        RECT 153.865 4849.730 158.315 4989.475 ;
        RECT 159.915 4851.000 163.165 4989.335 ;
        RECT 159.915 4849.730 163.160 4851.000 ;
        RECT 164.765 4849.730 168.015 4989.385 ;
        RECT 169.615 4849.730 174.065 4989.600 ;
        RECT 175.665 4849.730 180.115 4989.525 ;
        RECT 181.715 4849.970 184.965 4989.470 ;
        RECT 186.565 4849.730 191.015 4991.785 ;
        RECT 192.615 4849.730 197.865 4990.350 ;
      LAYER met5 ;
        RECT 199.465 4990.135 201.130 4991.950 ;
      LAYER met5 ;
        RECT 202.730 4990.135 382.270 4995.385 ;
      LAYER met5 ;
        RECT 383.870 4990.135 458.130 5003.035 ;
      LAYER met5 ;
        RECT 459.730 4996.985 639.270 5001.435 ;
        RECT 459.730 4990.135 639.270 4995.385 ;
      LAYER met5 ;
        RECT 640.870 4990.135 715.130 5003.035 ;
      LAYER met5 ;
        RECT 716.730 4996.985 896.270 5001.435 ;
        RECT 716.730 4990.135 896.270 4995.385 ;
      LAYER met5 ;
        RECT 897.870 4990.135 972.130 5003.035 ;
      LAYER met5 ;
        RECT 973.730 4996.985 1153.270 5001.435 ;
        RECT 973.730 4990.135 1153.270 4995.385 ;
      LAYER met5 ;
        RECT 1154.870 4990.135 1229.130 5003.035 ;
      LAYER met5 ;
        RECT 1230.730 4996.985 1411.270 5001.435 ;
        RECT 1230.730 4990.135 1411.270 4995.385 ;
      LAYER met5 ;
        RECT 1412.870 4990.135 1487.130 5003.035 ;
      LAYER met5 ;
        RECT 1488.730 4996.985 1668.270 5001.435 ;
        RECT 1488.730 4990.135 1668.270 4995.385 ;
      LAYER met5 ;
        RECT 1669.870 4990.135 1739.130 5003.035 ;
      LAYER met5 ;
        RECT 1740.730 4996.985 1920.270 5001.435 ;
        RECT 1740.730 4990.135 1920.270 4995.385 ;
      LAYER met5 ;
        RECT 1921.870 4990.135 1996.130 5003.035 ;
      LAYER met5 ;
        RECT 1997.730 4996.985 2181.000 5001.435 ;
        RECT 2186.000 4996.985 2365.270 5001.435 ;
        RECT 1997.730 4990.135 2365.270 4995.385 ;
      LAYER met5 ;
        RECT 2366.870 4990.135 2441.130 5003.035 ;
      LAYER met5 ;
        RECT 2442.730 4996.985 2622.270 5001.435 ;
        RECT 2442.730 4990.135 2622.270 4995.385 ;
      LAYER met5 ;
        RECT 2623.870 4990.135 2698.130 5003.035 ;
      LAYER met5 ;
        RECT 2699.730 4996.985 2879.270 5001.435 ;
        RECT 2699.730 4990.135 2879.270 4995.385 ;
      LAYER met5 ;
        RECT 2880.870 4990.135 2950.130 5003.035 ;
      LAYER met5 ;
        RECT 2951.730 4996.985 3131.270 5001.435 ;
        RECT 2951.730 4990.135 3131.270 4995.385 ;
      LAYER met5 ;
        RECT 3132.870 4990.135 3207.130 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4996.985 3391.785 5001.435 ;
      LAYER met5 ;
        RECT 3393.385 4995.385 3434.135 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4990.135 3390.350 4995.385 ;
      LAYER met5 ;
        RECT 197.865 4989.600 201.130 4990.135 ;
        POLYGON 197.865 4989.600 199.465 4989.600 197.865 4988.000 ;
        RECT 199.465 4988.535 201.130 4989.600 ;
        POLYGON 3388.000 4990.135 3389.600 4990.135 3389.600 4988.535 ;
        RECT 3389.600 4988.535 3390.135 4990.135 ;
        RECT 3391.950 4988.535 3434.135 4995.385 ;
        RECT 199.465 4988.000 204.000 4988.535 ;
        RECT 3388.000 4986.870 3434.135 4988.535 ;
        RECT 3388.000 4984.000 3388.535 4986.870 ;
        RECT 3403.035 4986.855 3406.285 4986.870 ;
        RECT 181.715 4848.130 184.965 4848.370 ;
        RECT 0.000 4846.400 197.865 4848.130 ;
        RECT 0.000 4780.600 31.390 4846.400 ;
        RECT 97.040 4780.600 197.865 4846.400 ;
      LAYER met5 ;
        RECT 3390.135 4836.730 3395.385 4985.270 ;
        RECT 3396.985 4836.730 3401.435 4985.270 ;
        RECT 3403.035 4837.035 3406.285 4985.255 ;
        RECT 3407.885 4836.730 3412.335 4985.270 ;
        RECT 3413.935 4836.730 3418.385 4985.270 ;
        RECT 3419.985 4836.730 3423.235 4985.270 ;
        RECT 3424.840 4984.000 3428.085 4985.270 ;
        RECT 3424.835 4838.000 3428.085 4984.000 ;
        RECT 3424.840 4836.730 3428.085 4838.000 ;
        RECT 3429.685 4836.730 3434.135 4985.270 ;
        RECT 3435.735 4836.730 3444.735 5011.155 ;
      LAYER met5 ;
        RECT 3446.335 4987.455 3588.000 5012.755 ;
        RECT 3446.335 4986.870 3456.435 4987.455 ;
      LAYER met5 ;
        RECT 3446.335 4836.730 3450.585 4985.270 ;
        RECT 3452.185 4836.730 3456.435 4985.270 ;
        RECT 3458.035 4982.000 3482.985 4985.855 ;
      LAYER met5 ;
        RECT 3484.585 4984.000 3588.000 4987.455 ;
      LAYER met5 ;
        RECT 3458.035 4977.000 3482.985 4979.000 ;
      LAYER met5 ;
        RECT 3458.035 4960.600 3482.985 4975.400 ;
      LAYER met5 ;
        RECT 3458.035 4957.000 3482.985 4959.000 ;
      LAYER met5 ;
        RECT 3458.035 4940.600 3482.985 4955.400 ;
      LAYER met5 ;
        RECT 3458.035 4937.000 3482.985 4939.000 ;
      LAYER met5 ;
        RECT 3458.035 4920.600 3482.985 4935.400 ;
      LAYER met5 ;
        RECT 3458.035 4917.000 3482.985 4919.000 ;
      LAYER met5 ;
        RECT 3458.035 4900.600 3482.985 4915.400 ;
      LAYER met5 ;
        RECT 3458.035 4897.000 3482.985 4899.000 ;
      LAYER met5 ;
        RECT 3458.035 4880.600 3482.985 4895.400 ;
      LAYER met5 ;
        RECT 3458.035 4877.000 3482.985 4879.000 ;
      LAYER met5 ;
        RECT 3458.035 4860.600 3482.985 4875.400 ;
      LAYER met5 ;
        RECT 3458.035 4857.000 3482.985 4859.000 ;
      LAYER met5 ;
        RECT 3458.035 4840.600 3482.985 4855.400 ;
      LAYER met5 ;
        RECT 3458.035 4836.730 3482.985 4839.000 ;
        RECT 3563.785 4838.000 3588.000 4984.000 ;
      LAYER met5 ;
        RECT 3403.035 4835.130 3406.285 4835.435 ;
        RECT 3484.585 4835.130 3588.000 4838.000 ;
        RECT 0.000 4773.870 197.865 4780.600 ;
        RECT 3390.135 4828.400 3588.000 4835.130 ;
        RECT 0.000 4771.000 103.415 4773.870 ;
        RECT 181.715 4773.565 184.965 4773.870 ;
      LAYER met5 ;
        RECT 0.000 4635.000 24.215 4771.000 ;
        RECT 105.015 4769.000 129.965 4772.270 ;
        RECT 105.015 4764.000 129.965 4766.000 ;
      LAYER met5 ;
        RECT 105.015 4757.600 129.965 4762.400 ;
      LAYER met5 ;
        RECT 105.015 4754.000 129.965 4756.000 ;
      LAYER met5 ;
        RECT 105.015 4737.600 129.965 4752.400 ;
      LAYER met5 ;
        RECT 105.015 4734.000 129.965 4736.000 ;
      LAYER met5 ;
        RECT 105.015 4717.600 129.965 4732.400 ;
      LAYER met5 ;
        RECT 105.015 4714.000 129.965 4716.000 ;
      LAYER met5 ;
        RECT 105.015 4697.600 129.965 4712.400 ;
      LAYER met5 ;
        RECT 105.015 4694.000 129.965 4696.000 ;
      LAYER met5 ;
        RECT 105.015 4677.600 129.965 4692.400 ;
      LAYER met5 ;
        RECT 105.015 4674.000 129.965 4676.000 ;
      LAYER met5 ;
        RECT 105.015 4657.600 129.965 4672.400 ;
      LAYER met5 ;
        RECT 105.015 4654.000 129.965 4656.000 ;
      LAYER met5 ;
        RECT 105.015 4637.600 129.965 4652.400 ;
        RECT 0.000 4632.130 103.415 4635.000 ;
      LAYER met5 ;
        RECT 105.015 4633.730 129.965 4636.000 ;
        RECT 131.565 4633.730 135.815 4772.270 ;
        RECT 137.415 4633.730 141.665 4772.270 ;
        RECT 143.265 4633.730 152.265 4772.270 ;
        RECT 153.865 4633.730 158.315 4772.270 ;
        RECT 159.915 4771.000 163.160 4772.270 ;
        RECT 159.915 4635.000 163.165 4771.000 ;
        RECT 159.915 4633.730 163.160 4635.000 ;
      LAYER met5 ;
        RECT 163.160 4632.130 163.165 4635.000 ;
      LAYER met5 ;
        RECT 164.765 4633.730 168.015 4772.270 ;
        RECT 169.615 4633.730 174.065 4772.270 ;
        RECT 175.665 4633.730 180.115 4772.270 ;
        RECT 181.715 4634.035 184.965 4771.965 ;
        RECT 192.615 4633.730 197.865 4772.270 ;
      LAYER met5 ;
        RECT 3390.135 4762.600 3490.960 4828.400 ;
        RECT 3556.610 4762.600 3588.000 4828.400 ;
        RECT 3390.135 4760.870 3588.000 4762.600 ;
        RECT 3403.035 4760.630 3406.285 4760.870 ;
        RECT 181.715 4632.130 184.965 4632.435 ;
        RECT 0.000 4626.270 197.865 4632.130 ;
        RECT 0.000 4568.670 29.235 4626.270 ;
        RECT 99.700 4568.670 197.865 4626.270 ;
      LAYER met5 ;
        RECT 3390.135 4611.730 3395.385 4759.270 ;
        RECT 3403.035 4612.035 3406.285 4759.030 ;
        RECT 3407.885 4611.730 3412.335 4759.270 ;
        RECT 3413.935 4611.730 3418.385 4759.270 ;
        RECT 3419.985 4611.730 3423.235 4759.270 ;
        RECT 3424.840 4758.000 3428.085 4759.270 ;
        RECT 3424.835 4613.000 3428.085 4758.000 ;
      LAYER met5 ;
        RECT 3403.035 4610.130 3406.285 4610.435 ;
        RECT 3424.835 4610.130 3424.840 4613.000 ;
      LAYER met5 ;
        RECT 3424.840 4611.730 3428.085 4613.000 ;
        RECT 3429.685 4611.730 3434.135 4759.270 ;
        RECT 3435.735 4611.730 3444.735 4759.270 ;
        RECT 3446.335 4611.730 3450.585 4759.270 ;
        RECT 3452.185 4611.730 3456.435 4759.270 ;
        RECT 3458.035 4757.000 3482.985 4759.270 ;
      LAYER met5 ;
        RECT 3484.585 4758.000 3588.000 4760.870 ;
      LAYER met5 ;
        RECT 3458.035 4752.000 3482.985 4754.000 ;
      LAYER met5 ;
        RECT 3458.035 4735.600 3482.985 4750.400 ;
      LAYER met5 ;
        RECT 3458.035 4732.000 3482.985 4734.000 ;
      LAYER met5 ;
        RECT 3458.035 4715.600 3482.985 4730.400 ;
      LAYER met5 ;
        RECT 3458.035 4712.000 3482.985 4714.000 ;
      LAYER met5 ;
        RECT 3458.035 4695.600 3482.985 4710.400 ;
      LAYER met5 ;
        RECT 3458.035 4692.000 3482.985 4694.000 ;
      LAYER met5 ;
        RECT 3458.035 4675.600 3482.985 4690.400 ;
      LAYER met5 ;
        RECT 3458.035 4672.000 3482.985 4674.000 ;
      LAYER met5 ;
        RECT 3458.035 4655.600 3482.985 4670.400 ;
      LAYER met5 ;
        RECT 3458.035 4652.000 3482.985 4654.000 ;
      LAYER met5 ;
        RECT 3458.035 4635.600 3482.985 4650.400 ;
      LAYER met5 ;
        RECT 3458.035 4632.000 3482.985 4634.000 ;
      LAYER met5 ;
        RECT 3458.035 4615.600 3482.985 4630.400 ;
      LAYER met5 ;
        RECT 3458.035 4611.730 3482.985 4614.000 ;
        RECT 3563.785 4613.000 3588.000 4758.000 ;
      LAYER met5 ;
        RECT 3484.585 4610.130 3588.000 4613.000 ;
        RECT 0.000 4562.870 197.865 4568.670 ;
        RECT 3390.135 4604.330 3588.000 4610.130 ;
        RECT 0.000 4560.000 103.415 4562.870 ;
      LAYER met5 ;
        RECT 0.000 4424.000 24.215 4560.000 ;
        RECT 105.015 4558.000 129.965 4561.270 ;
        RECT 105.015 4553.000 129.965 4555.000 ;
      LAYER met5 ;
        RECT 105.015 4546.600 129.965 4551.400 ;
      LAYER met5 ;
        RECT 105.015 4543.000 129.965 4545.000 ;
      LAYER met5 ;
        RECT 105.015 4526.600 129.965 4541.400 ;
      LAYER met5 ;
        RECT 105.015 4523.000 129.965 4525.000 ;
      LAYER met5 ;
        RECT 105.015 4506.600 129.965 4521.400 ;
      LAYER met5 ;
        RECT 105.015 4503.000 129.965 4505.000 ;
      LAYER met5 ;
        RECT 105.015 4486.600 129.965 4501.400 ;
      LAYER met5 ;
        RECT 105.015 4483.000 129.965 4485.000 ;
      LAYER met5 ;
        RECT 105.015 4466.600 129.965 4481.400 ;
      LAYER met5 ;
        RECT 105.015 4463.000 129.965 4465.000 ;
      LAYER met5 ;
        RECT 105.015 4446.600 129.965 4461.400 ;
      LAYER met5 ;
        RECT 105.015 4443.000 129.965 4445.000 ;
      LAYER met5 ;
        RECT 105.015 4426.600 129.965 4441.400 ;
        RECT 0.000 4421.130 103.415 4424.000 ;
      LAYER met5 ;
        RECT 105.015 4422.730 129.965 4425.000 ;
        RECT 131.565 4422.730 135.815 4561.270 ;
        RECT 137.415 4422.730 141.665 4561.270 ;
        RECT 143.265 4422.730 152.265 4561.270 ;
        RECT 153.865 4422.730 158.315 4561.270 ;
        RECT 159.915 4560.000 163.160 4561.270 ;
      LAYER met5 ;
        RECT 163.160 4560.000 163.165 4562.870 ;
        RECT 181.715 4562.565 184.965 4562.870 ;
      LAYER met5 ;
        RECT 159.915 4424.000 163.165 4560.000 ;
        RECT 159.915 4422.730 163.160 4424.000 ;
      LAYER met5 ;
        RECT 163.160 4421.130 163.165 4424.000 ;
      LAYER met5 ;
        RECT 164.765 4422.730 168.015 4561.270 ;
        RECT 169.615 4422.730 174.065 4561.270 ;
        RECT 175.665 4422.730 180.115 4561.270 ;
        RECT 181.715 4423.035 184.965 4560.965 ;
        RECT 192.615 4422.730 197.865 4561.270 ;
      LAYER met5 ;
        RECT 3390.135 4546.730 3488.300 4604.330 ;
        RECT 3558.765 4546.730 3588.000 4604.330 ;
        RECT 3390.135 4540.870 3588.000 4546.730 ;
        RECT 3403.035 4540.565 3406.285 4540.870 ;
        RECT 181.715 4421.130 184.965 4421.435 ;
        RECT 0.000 4418.490 197.865 4421.130 ;
        RECT 0.000 4354.450 32.455 4418.490 ;
      LAYER met5 ;
        RECT 34.055 4356.050 94.880 4416.890 ;
      LAYER met5 ;
        RECT 96.480 4354.450 197.865 4418.490 ;
      LAYER met5 ;
        RECT 3390.135 4390.730 3395.385 4539.270 ;
        RECT 3403.035 4391.035 3406.285 4538.965 ;
        RECT 3407.885 4390.730 3412.335 4539.270 ;
        RECT 3413.935 4390.730 3418.385 4539.270 ;
        RECT 3419.985 4390.730 3423.235 4539.270 ;
      LAYER met5 ;
        RECT 3424.835 4538.000 3424.840 4540.870 ;
      LAYER met5 ;
        RECT 3424.840 4538.000 3428.085 4539.270 ;
        RECT 3424.835 4392.000 3428.085 4538.000 ;
        RECT 3424.840 4390.730 3428.085 4392.000 ;
        RECT 3429.685 4390.730 3434.135 4539.270 ;
        RECT 3435.735 4390.730 3444.735 4539.270 ;
        RECT 3446.335 4390.730 3450.585 4539.270 ;
        RECT 3452.185 4390.730 3456.435 4539.270 ;
        RECT 3458.035 4536.000 3482.985 4539.270 ;
      LAYER met5 ;
        RECT 3484.585 4538.000 3588.000 4540.870 ;
      LAYER met5 ;
        RECT 3458.035 4531.000 3482.985 4533.000 ;
      LAYER met5 ;
        RECT 3458.035 4514.600 3482.985 4529.400 ;
      LAYER met5 ;
        RECT 3458.035 4511.000 3482.985 4513.000 ;
      LAYER met5 ;
        RECT 3458.035 4494.600 3482.985 4509.400 ;
      LAYER met5 ;
        RECT 3458.035 4491.000 3482.985 4493.000 ;
      LAYER met5 ;
        RECT 3458.035 4474.600 3482.985 4489.400 ;
      LAYER met5 ;
        RECT 3458.035 4471.000 3482.985 4473.000 ;
      LAYER met5 ;
        RECT 3458.035 4454.600 3482.985 4469.400 ;
      LAYER met5 ;
        RECT 3458.035 4451.000 3482.985 4453.000 ;
      LAYER met5 ;
        RECT 3458.035 4434.600 3482.985 4449.400 ;
      LAYER met5 ;
        RECT 3458.035 4431.000 3482.985 4433.000 ;
      LAYER met5 ;
        RECT 3458.035 4414.600 3482.985 4429.400 ;
      LAYER met5 ;
        RECT 3458.035 4411.000 3482.985 4413.000 ;
      LAYER met5 ;
        RECT 3458.035 4394.600 3482.985 4409.400 ;
      LAYER met5 ;
        RECT 3458.035 4390.730 3482.985 4393.000 ;
        RECT 3563.785 4392.000 3588.000 4538.000 ;
      LAYER met5 ;
        RECT 3403.035 4389.130 3406.285 4389.435 ;
        RECT 3484.585 4389.130 3588.000 4392.000 ;
        RECT 0.000 4351.870 197.865 4354.450 ;
        RECT 3390.135 4382.400 3588.000 4389.130 ;
        RECT 0.000 4349.000 103.415 4351.870 ;
      LAYER met5 ;
        RECT 0.000 4213.000 24.215 4349.000 ;
        RECT 105.015 4347.000 129.965 4350.270 ;
        RECT 105.015 4342.000 129.965 4344.000 ;
      LAYER met5 ;
        RECT 105.015 4335.600 129.965 4340.400 ;
      LAYER met5 ;
        RECT 105.015 4332.000 129.965 4334.000 ;
      LAYER met5 ;
        RECT 105.015 4315.600 129.965 4330.400 ;
      LAYER met5 ;
        RECT 105.015 4312.000 129.965 4314.000 ;
      LAYER met5 ;
        RECT 105.015 4295.600 129.965 4310.400 ;
      LAYER met5 ;
        RECT 105.015 4292.000 129.965 4294.000 ;
      LAYER met5 ;
        RECT 105.015 4275.600 129.965 4290.400 ;
      LAYER met5 ;
        RECT 105.015 4272.000 129.965 4274.000 ;
      LAYER met5 ;
        RECT 105.015 4255.600 129.965 4270.400 ;
      LAYER met5 ;
        RECT 105.015 4252.000 129.965 4254.000 ;
      LAYER met5 ;
        RECT 105.015 4235.600 129.965 4250.400 ;
      LAYER met5 ;
        RECT 105.015 4232.000 129.965 4234.000 ;
      LAYER met5 ;
        RECT 105.015 4215.600 129.965 4230.400 ;
        RECT 0.000 4210.130 103.415 4213.000 ;
      LAYER met5 ;
        RECT 105.015 4211.730 129.965 4214.000 ;
        RECT 131.565 4211.730 135.815 4350.270 ;
        RECT 137.415 4211.730 141.665 4350.270 ;
        RECT 153.865 4211.730 158.315 4350.270 ;
      LAYER met5 ;
        RECT 163.160 4349.000 163.165 4351.870 ;
        RECT 181.715 4351.565 184.965 4351.870 ;
        RECT 163.160 4210.130 163.165 4213.000 ;
      LAYER met5 ;
        RECT 164.765 4211.730 168.015 4350.270 ;
        RECT 169.615 4211.730 174.065 4350.270 ;
        RECT 175.665 4211.730 180.115 4350.270 ;
        RECT 181.715 4212.035 184.965 4349.965 ;
        RECT 186.565 4211.730 191.015 4350.270 ;
        RECT 192.615 4211.730 197.865 4350.270 ;
      LAYER met5 ;
        RECT 3390.135 4316.600 3490.960 4382.400 ;
        RECT 3556.610 4316.600 3588.000 4382.400 ;
        RECT 3390.135 4314.870 3588.000 4316.600 ;
        RECT 3403.035 4314.630 3406.285 4314.870 ;
        RECT 181.715 4210.130 184.965 4210.435 ;
        RECT 0.000 4207.490 197.865 4210.130 ;
        RECT 0.000 4143.450 32.455 4207.490 ;
        RECT 96.480 4143.450 197.865 4207.490 ;
      LAYER met5 ;
        RECT 3390.135 4165.730 3395.385 4313.270 ;
        RECT 3396.985 4165.730 3401.435 4313.270 ;
        RECT 3407.885 4165.730 3412.335 4313.270 ;
        RECT 3413.935 4165.730 3418.385 4313.270 ;
        RECT 3419.985 4165.730 3423.235 4313.270 ;
        RECT 3424.840 4312.000 3428.085 4313.270 ;
        RECT 3424.835 4167.000 3428.085 4312.000 ;
      LAYER met5 ;
        RECT 3403.035 4164.130 3406.285 4164.435 ;
        RECT 3424.835 4164.130 3424.840 4167.000 ;
      LAYER met5 ;
        RECT 3424.840 4165.730 3428.085 4167.000 ;
        RECT 3429.685 4165.730 3434.135 4313.270 ;
        RECT 3435.735 4165.730 3444.735 4313.270 ;
        RECT 3446.335 4165.730 3450.585 4313.270 ;
        RECT 3452.185 4165.730 3456.435 4313.270 ;
        RECT 3458.035 4311.000 3482.985 4313.270 ;
      LAYER met5 ;
        RECT 3484.585 4312.000 3588.000 4314.870 ;
      LAYER met5 ;
        RECT 3458.035 4306.000 3482.985 4308.000 ;
      LAYER met5 ;
        RECT 3458.035 4289.600 3482.985 4304.400 ;
      LAYER met5 ;
        RECT 3458.035 4286.000 3482.985 4288.000 ;
      LAYER met5 ;
        RECT 3458.035 4269.600 3482.985 4284.400 ;
      LAYER met5 ;
        RECT 3458.035 4266.000 3482.985 4268.000 ;
      LAYER met5 ;
        RECT 3458.035 4249.600 3482.985 4264.400 ;
      LAYER met5 ;
        RECT 3458.035 4246.000 3482.985 4248.000 ;
      LAYER met5 ;
        RECT 3458.035 4229.600 3482.985 4244.400 ;
      LAYER met5 ;
        RECT 3458.035 4226.000 3482.985 4228.000 ;
      LAYER met5 ;
        RECT 3458.035 4209.600 3482.985 4224.400 ;
      LAYER met5 ;
        RECT 3458.035 4206.000 3482.985 4208.000 ;
      LAYER met5 ;
        RECT 3458.035 4189.600 3482.985 4204.400 ;
      LAYER met5 ;
        RECT 3458.035 4186.000 3482.985 4188.000 ;
      LAYER met5 ;
        RECT 3458.035 4169.600 3482.985 4184.400 ;
      LAYER met5 ;
        RECT 3458.035 4165.730 3482.985 4168.000 ;
        RECT 3563.785 4167.000 3588.000 4312.000 ;
      LAYER met5 ;
        RECT 3484.585 4164.130 3588.000 4167.000 ;
        RECT 0.000 4140.870 197.865 4143.450 ;
        RECT 3390.135 4161.550 3588.000 4164.130 ;
        RECT 0.000 4138.000 103.415 4140.870 ;
      LAYER met5 ;
        RECT 0.000 4002.000 24.215 4138.000 ;
        RECT 105.015 4136.000 129.965 4139.270 ;
        RECT 105.015 4131.000 129.965 4133.000 ;
      LAYER met5 ;
        RECT 105.015 4124.600 129.965 4129.400 ;
      LAYER met5 ;
        RECT 105.015 4121.000 129.965 4123.000 ;
      LAYER met5 ;
        RECT 105.015 4104.600 129.965 4119.400 ;
      LAYER met5 ;
        RECT 105.015 4101.000 129.965 4103.000 ;
      LAYER met5 ;
        RECT 105.015 4084.600 129.965 4099.400 ;
      LAYER met5 ;
        RECT 105.015 4081.000 129.965 4083.000 ;
      LAYER met5 ;
        RECT 105.015 4064.600 129.965 4079.400 ;
      LAYER met5 ;
        RECT 105.015 4061.000 129.965 4063.000 ;
      LAYER met5 ;
        RECT 105.015 4044.600 129.965 4059.400 ;
      LAYER met5 ;
        RECT 105.015 4041.000 129.965 4043.000 ;
      LAYER met5 ;
        RECT 105.015 4024.600 129.965 4039.400 ;
      LAYER met5 ;
        RECT 105.015 4021.000 129.965 4023.000 ;
      LAYER met5 ;
        RECT 105.015 4004.600 129.965 4019.400 ;
        RECT 0.000 3999.130 103.415 4002.000 ;
      LAYER met5 ;
        RECT 105.015 4000.730 129.965 4003.000 ;
        RECT 131.565 4000.730 135.815 4139.270 ;
        RECT 137.415 4000.730 141.665 4139.270 ;
        RECT 153.865 4000.730 158.315 4139.270 ;
      LAYER met5 ;
        RECT 163.160 4138.000 163.165 4140.870 ;
        RECT 181.715 4140.565 184.965 4140.870 ;
      LAYER met5 ;
        RECT 164.765 4000.730 168.015 4139.270 ;
        RECT 169.615 4000.730 174.065 4139.270 ;
        RECT 175.665 4000.730 180.115 4139.270 ;
        RECT 181.715 4000.970 184.965 4138.965 ;
        RECT 186.565 4000.730 191.015 4139.270 ;
        RECT 192.615 4000.730 197.865 4139.270 ;
      LAYER met5 ;
        RECT 3390.135 4097.510 3491.520 4161.550 ;
        RECT 3555.545 4097.510 3588.000 4161.550 ;
        RECT 3390.135 4094.870 3588.000 4097.510 ;
        RECT 3403.035 4094.565 3406.285 4094.870 ;
        RECT 181.715 3999.130 184.965 3999.370 ;
        RECT 0.000 3997.400 197.865 3999.130 ;
        RECT 0.000 3931.600 31.390 3997.400 ;
        RECT 97.040 3931.600 197.865 3997.400 ;
      LAYER met5 ;
        RECT 3390.135 3944.730 3395.385 4093.270 ;
        RECT 3396.985 3944.730 3401.435 4093.270 ;
        RECT 3407.885 3944.730 3412.335 4093.270 ;
        RECT 3413.935 3944.730 3418.385 4093.270 ;
        RECT 3419.985 3944.730 3423.235 4093.270 ;
      LAYER met5 ;
        RECT 3424.835 4092.000 3424.840 4094.870 ;
      LAYER met5 ;
        RECT 3424.840 4092.000 3428.085 4093.270 ;
        RECT 3424.835 3946.000 3428.085 4092.000 ;
        RECT 3424.840 3944.730 3428.085 3946.000 ;
        RECT 3429.685 3944.730 3434.135 4093.270 ;
        RECT 3435.735 3944.730 3444.735 4093.270 ;
        RECT 3446.335 3944.730 3450.585 4093.270 ;
        RECT 3452.185 3944.730 3456.435 4093.270 ;
        RECT 3458.035 4090.000 3482.985 4093.270 ;
      LAYER met5 ;
        RECT 3484.585 4092.000 3588.000 4094.870 ;
      LAYER met5 ;
        RECT 3458.035 4085.000 3482.985 4087.000 ;
      LAYER met5 ;
        RECT 3458.035 4068.600 3482.985 4083.400 ;
      LAYER met5 ;
        RECT 3458.035 4065.000 3482.985 4067.000 ;
      LAYER met5 ;
        RECT 3458.035 4048.600 3482.985 4063.400 ;
      LAYER met5 ;
        RECT 3458.035 4045.000 3482.985 4047.000 ;
      LAYER met5 ;
        RECT 3458.035 4028.600 3482.985 4043.400 ;
      LAYER met5 ;
        RECT 3458.035 4025.000 3482.985 4027.000 ;
      LAYER met5 ;
        RECT 3458.035 4008.600 3482.985 4023.400 ;
      LAYER met5 ;
        RECT 3458.035 4005.000 3482.985 4007.000 ;
      LAYER met5 ;
        RECT 3458.035 3988.600 3482.985 4003.400 ;
      LAYER met5 ;
        RECT 3458.035 3985.000 3482.985 3987.000 ;
      LAYER met5 ;
        RECT 3458.035 3968.600 3482.985 3983.400 ;
      LAYER met5 ;
        RECT 3458.035 3965.000 3482.985 3967.000 ;
      LAYER met5 ;
        RECT 3458.035 3948.600 3482.985 3963.400 ;
      LAYER met5 ;
        RECT 3458.035 3944.730 3482.985 3947.000 ;
        RECT 3563.785 3946.000 3588.000 4092.000 ;
      LAYER met5 ;
        RECT 3403.035 3943.130 3406.285 3943.435 ;
        RECT 3484.585 3943.130 3588.000 3946.000 ;
        RECT 0.000 3924.870 197.865 3931.600 ;
        RECT 3390.135 3936.400 3588.000 3943.130 ;
        RECT 0.000 3922.000 103.415 3924.870 ;
        RECT 181.715 3924.565 184.965 3924.870 ;
      LAYER met5 ;
        RECT 0.000 3786.000 24.215 3922.000 ;
        RECT 105.015 3920.000 129.965 3923.270 ;
        RECT 105.015 3915.000 129.965 3917.000 ;
      LAYER met5 ;
        RECT 105.015 3908.600 129.965 3913.400 ;
      LAYER met5 ;
        RECT 105.015 3905.000 129.965 3907.000 ;
      LAYER met5 ;
        RECT 105.015 3888.600 129.965 3903.400 ;
      LAYER met5 ;
        RECT 105.015 3885.000 129.965 3887.000 ;
      LAYER met5 ;
        RECT 105.015 3868.600 129.965 3883.400 ;
      LAYER met5 ;
        RECT 105.015 3865.000 129.965 3867.000 ;
      LAYER met5 ;
        RECT 105.015 3848.600 129.965 3863.400 ;
      LAYER met5 ;
        RECT 105.015 3845.000 129.965 3847.000 ;
      LAYER met5 ;
        RECT 105.015 3828.600 129.965 3843.400 ;
      LAYER met5 ;
        RECT 105.015 3825.000 129.965 3827.000 ;
      LAYER met5 ;
        RECT 105.015 3808.600 129.965 3823.400 ;
      LAYER met5 ;
        RECT 105.015 3805.000 129.965 3807.000 ;
      LAYER met5 ;
        RECT 105.015 3788.600 129.965 3803.400 ;
        RECT 0.000 3783.130 103.415 3786.000 ;
      LAYER met5 ;
        RECT 105.015 3784.730 129.965 3787.000 ;
        RECT 131.565 3784.730 135.815 3923.270 ;
        RECT 137.415 3784.730 141.665 3923.270 ;
        RECT 143.265 3784.730 152.265 3923.270 ;
        RECT 153.865 3784.730 158.315 3923.270 ;
        RECT 159.915 3922.000 163.160 3923.270 ;
        RECT 159.915 3786.000 163.165 3922.000 ;
        RECT 159.915 3784.730 163.160 3786.000 ;
        RECT 164.765 3784.730 168.015 3923.270 ;
        RECT 169.615 3784.730 174.065 3923.270 ;
        RECT 175.665 3784.730 180.115 3923.270 ;
        RECT 181.715 3784.970 184.965 3922.965 ;
        RECT 186.565 3784.730 191.015 3923.270 ;
        RECT 192.615 3784.730 197.865 3923.270 ;
      LAYER met5 ;
        RECT 3390.135 3870.600 3490.960 3936.400 ;
        RECT 3556.610 3870.600 3588.000 3936.400 ;
        RECT 3390.135 3868.870 3588.000 3870.600 ;
        RECT 3403.035 3868.630 3406.285 3868.870 ;
        RECT 181.715 3783.130 184.965 3783.370 ;
        RECT 0.000 3781.400 197.865 3783.130 ;
        RECT 0.000 3715.600 31.390 3781.400 ;
        RECT 97.040 3715.600 197.865 3781.400 ;
      LAYER met5 ;
        RECT 3390.135 3719.730 3395.385 3867.270 ;
        RECT 3396.985 3719.730 3401.435 3867.270 ;
        RECT 3403.035 3720.035 3406.285 3867.030 ;
        RECT 3407.885 3719.730 3412.335 3867.270 ;
        RECT 3413.935 3719.730 3418.385 3867.270 ;
        RECT 3419.985 3719.730 3423.235 3867.270 ;
        RECT 3424.840 3866.000 3428.085 3867.270 ;
        RECT 3424.835 3721.000 3428.085 3866.000 ;
        RECT 3424.840 3719.730 3428.085 3721.000 ;
        RECT 3429.685 3719.730 3434.135 3867.270 ;
        RECT 3435.735 3719.730 3444.735 3867.270 ;
        RECT 3446.335 3719.730 3450.585 3867.270 ;
        RECT 3452.185 3719.730 3456.435 3867.270 ;
        RECT 3458.035 3865.000 3482.985 3867.270 ;
      LAYER met5 ;
        RECT 3484.585 3866.000 3588.000 3868.870 ;
      LAYER met5 ;
        RECT 3458.035 3860.000 3482.985 3862.000 ;
      LAYER met5 ;
        RECT 3458.035 3843.600 3482.985 3858.400 ;
      LAYER met5 ;
        RECT 3458.035 3840.000 3482.985 3842.000 ;
      LAYER met5 ;
        RECT 3458.035 3823.600 3482.985 3838.400 ;
      LAYER met5 ;
        RECT 3458.035 3820.000 3482.985 3822.000 ;
      LAYER met5 ;
        RECT 3458.035 3803.600 3482.985 3818.400 ;
      LAYER met5 ;
        RECT 3458.035 3800.000 3482.985 3802.000 ;
      LAYER met5 ;
        RECT 3458.035 3783.600 3482.985 3798.400 ;
      LAYER met5 ;
        RECT 3458.035 3780.000 3482.985 3782.000 ;
      LAYER met5 ;
        RECT 3458.035 3763.600 3482.985 3778.400 ;
      LAYER met5 ;
        RECT 3458.035 3760.000 3482.985 3762.000 ;
      LAYER met5 ;
        RECT 3458.035 3743.600 3482.985 3758.400 ;
      LAYER met5 ;
        RECT 3458.035 3740.000 3482.985 3742.000 ;
      LAYER met5 ;
        RECT 3458.035 3723.600 3482.985 3738.400 ;
      LAYER met5 ;
        RECT 3458.035 3719.730 3482.985 3722.000 ;
        RECT 3563.785 3721.000 3588.000 3866.000 ;
      LAYER met5 ;
        RECT 3403.035 3718.130 3406.285 3718.435 ;
        RECT 3484.585 3718.130 3588.000 3721.000 ;
        RECT 0.000 3708.870 197.865 3715.600 ;
        RECT 3390.135 3711.400 3588.000 3718.130 ;
        RECT 0.000 3706.000 103.415 3708.870 ;
        RECT 181.715 3708.565 184.965 3708.870 ;
      LAYER met5 ;
        RECT 0.000 3570.000 24.215 3706.000 ;
        RECT 105.015 3704.000 129.965 3707.270 ;
        RECT 105.015 3699.000 129.965 3701.000 ;
      LAYER met5 ;
        RECT 105.015 3692.600 129.965 3697.400 ;
      LAYER met5 ;
        RECT 105.015 3689.000 129.965 3691.000 ;
      LAYER met5 ;
        RECT 105.015 3672.600 129.965 3687.400 ;
      LAYER met5 ;
        RECT 105.015 3669.000 129.965 3671.000 ;
      LAYER met5 ;
        RECT 105.015 3652.600 129.965 3667.400 ;
      LAYER met5 ;
        RECT 105.015 3649.000 129.965 3651.000 ;
      LAYER met5 ;
        RECT 105.015 3632.600 129.965 3647.400 ;
      LAYER met5 ;
        RECT 105.015 3629.000 129.965 3631.000 ;
      LAYER met5 ;
        RECT 105.015 3612.600 129.965 3627.400 ;
      LAYER met5 ;
        RECT 105.015 3609.000 129.965 3611.000 ;
      LAYER met5 ;
        RECT 105.015 3592.600 129.965 3607.400 ;
      LAYER met5 ;
        RECT 105.015 3589.000 129.965 3591.000 ;
      LAYER met5 ;
        RECT 105.015 3572.600 129.965 3587.400 ;
        RECT 0.000 3567.130 103.415 3570.000 ;
      LAYER met5 ;
        RECT 105.015 3568.730 129.965 3571.000 ;
        RECT 131.565 3568.730 135.815 3707.270 ;
        RECT 137.415 3568.730 141.665 3707.270 ;
        RECT 143.265 3568.730 152.265 3707.270 ;
        RECT 153.865 3568.730 158.315 3707.270 ;
        RECT 159.915 3706.000 163.160 3707.270 ;
        RECT 159.915 3570.000 163.165 3706.000 ;
        RECT 159.915 3568.730 163.160 3570.000 ;
        RECT 164.765 3568.730 168.015 3707.270 ;
        RECT 169.615 3568.730 174.065 3707.270 ;
        RECT 175.665 3568.730 180.115 3707.270 ;
        RECT 181.715 3568.970 184.965 3706.965 ;
        RECT 186.565 3568.730 191.015 3707.270 ;
        RECT 192.615 3568.730 197.865 3707.270 ;
      LAYER met5 ;
        RECT 3390.135 3645.600 3490.960 3711.400 ;
        RECT 3556.610 3645.600 3588.000 3711.400 ;
        RECT 3390.135 3643.870 3588.000 3645.600 ;
        RECT 3403.035 3643.630 3406.285 3643.870 ;
        RECT 181.715 3567.130 184.965 3567.370 ;
        RECT 0.000 3565.400 197.865 3567.130 ;
        RECT 0.000 3499.600 31.390 3565.400 ;
        RECT 97.040 3499.600 197.865 3565.400 ;
        RECT 0.000 3492.870 197.865 3499.600 ;
      LAYER met5 ;
        RECT 3390.135 3494.730 3395.385 3642.270 ;
        RECT 3396.985 3494.730 3401.435 3642.270 ;
        RECT 3403.035 3495.035 3406.285 3642.030 ;
        RECT 3407.885 3494.730 3412.335 3642.270 ;
        RECT 3413.935 3494.730 3418.385 3642.270 ;
        RECT 3419.985 3494.730 3423.235 3642.270 ;
        RECT 3424.840 3641.000 3428.085 3642.270 ;
        RECT 3424.835 3496.000 3428.085 3641.000 ;
        RECT 3424.840 3494.730 3428.085 3496.000 ;
        RECT 3429.685 3494.730 3434.135 3642.270 ;
        RECT 3435.735 3494.730 3444.735 3642.270 ;
        RECT 3446.335 3494.730 3450.585 3642.270 ;
        RECT 3452.185 3494.730 3456.435 3642.270 ;
        RECT 3458.035 3640.000 3482.985 3642.270 ;
      LAYER met5 ;
        RECT 3484.585 3641.000 3588.000 3643.870 ;
      LAYER met5 ;
        RECT 3458.035 3635.000 3482.985 3637.000 ;
      LAYER met5 ;
        RECT 3458.035 3618.600 3482.985 3633.400 ;
      LAYER met5 ;
        RECT 3458.035 3615.000 3482.985 3617.000 ;
      LAYER met5 ;
        RECT 3458.035 3598.600 3482.985 3613.400 ;
      LAYER met5 ;
        RECT 3458.035 3595.000 3482.985 3597.000 ;
      LAYER met5 ;
        RECT 3458.035 3578.600 3482.985 3593.400 ;
      LAYER met5 ;
        RECT 3458.035 3575.000 3482.985 3577.000 ;
      LAYER met5 ;
        RECT 3458.035 3558.600 3482.985 3573.400 ;
      LAYER met5 ;
        RECT 3458.035 3555.000 3482.985 3557.000 ;
      LAYER met5 ;
        RECT 3458.035 3538.600 3482.985 3553.400 ;
      LAYER met5 ;
        RECT 3458.035 3535.000 3482.985 3537.000 ;
      LAYER met5 ;
        RECT 3458.035 3518.600 3482.985 3533.400 ;
      LAYER met5 ;
        RECT 3458.035 3515.000 3482.985 3517.000 ;
      LAYER met5 ;
        RECT 3458.035 3498.600 3482.985 3513.400 ;
      LAYER met5 ;
        RECT 3458.035 3494.730 3482.985 3497.000 ;
        RECT 3563.785 3496.000 3588.000 3641.000 ;
      LAYER met5 ;
        RECT 3403.035 3493.130 3406.285 3493.435 ;
        RECT 3484.585 3493.130 3588.000 3496.000 ;
        RECT 0.000 3490.000 103.415 3492.870 ;
        RECT 181.715 3492.565 184.965 3492.870 ;
      LAYER met5 ;
        RECT 0.000 3354.000 24.215 3490.000 ;
        RECT 105.015 3488.000 129.965 3491.270 ;
        RECT 105.015 3483.000 129.965 3485.000 ;
      LAYER met5 ;
        RECT 105.015 3476.600 129.965 3481.400 ;
      LAYER met5 ;
        RECT 105.015 3473.000 129.965 3475.000 ;
      LAYER met5 ;
        RECT 105.015 3456.600 129.965 3471.400 ;
      LAYER met5 ;
        RECT 105.015 3453.000 129.965 3455.000 ;
      LAYER met5 ;
        RECT 105.015 3436.600 129.965 3451.400 ;
      LAYER met5 ;
        RECT 105.015 3433.000 129.965 3435.000 ;
      LAYER met5 ;
        RECT 105.015 3416.600 129.965 3431.400 ;
      LAYER met5 ;
        RECT 105.015 3413.000 129.965 3415.000 ;
      LAYER met5 ;
        RECT 105.015 3396.600 129.965 3411.400 ;
      LAYER met5 ;
        RECT 105.015 3393.000 129.965 3395.000 ;
      LAYER met5 ;
        RECT 105.015 3376.600 129.965 3391.400 ;
      LAYER met5 ;
        RECT 105.015 3373.000 129.965 3375.000 ;
      LAYER met5 ;
        RECT 105.015 3356.600 129.965 3371.400 ;
        RECT 0.000 3351.130 103.415 3354.000 ;
      LAYER met5 ;
        RECT 105.015 3352.730 129.965 3355.000 ;
        RECT 131.565 3352.730 135.815 3491.270 ;
        RECT 137.415 3352.730 141.665 3491.270 ;
        RECT 143.265 3352.730 152.265 3491.270 ;
        RECT 153.865 3352.730 158.315 3491.270 ;
        RECT 159.915 3490.000 163.160 3491.270 ;
        RECT 159.915 3354.000 163.165 3490.000 ;
        RECT 159.915 3352.730 163.160 3354.000 ;
        RECT 164.765 3352.730 168.015 3491.270 ;
        RECT 169.615 3352.730 174.065 3491.270 ;
        RECT 175.665 3352.730 180.115 3491.270 ;
        RECT 181.715 3352.970 184.965 3490.965 ;
        RECT 186.565 3352.730 191.015 3491.270 ;
        RECT 192.615 3352.730 197.865 3491.270 ;
      LAYER met5 ;
        RECT 3390.135 3486.400 3588.000 3493.130 ;
        RECT 3390.135 3420.600 3490.960 3486.400 ;
        RECT 3556.610 3420.600 3588.000 3486.400 ;
        RECT 3390.135 3418.870 3588.000 3420.600 ;
        RECT 3403.035 3418.630 3406.285 3418.870 ;
        RECT 181.715 3351.130 184.965 3351.370 ;
        RECT 0.000 3349.400 197.865 3351.130 ;
        RECT 0.000 3283.600 31.390 3349.400 ;
        RECT 97.040 3283.600 197.865 3349.400 ;
        RECT 0.000 3276.870 197.865 3283.600 ;
        RECT 0.000 3274.000 103.415 3276.870 ;
        RECT 181.715 3276.565 184.965 3276.870 ;
      LAYER met5 ;
        RECT 0.000 3138.000 24.215 3274.000 ;
        RECT 105.015 3272.000 129.965 3275.270 ;
        RECT 105.015 3267.000 129.965 3269.000 ;
      LAYER met5 ;
        RECT 105.015 3260.600 129.965 3265.400 ;
      LAYER met5 ;
        RECT 105.015 3257.000 129.965 3259.000 ;
      LAYER met5 ;
        RECT 105.015 3240.600 129.965 3255.400 ;
      LAYER met5 ;
        RECT 105.015 3237.000 129.965 3239.000 ;
      LAYER met5 ;
        RECT 105.015 3220.600 129.965 3235.400 ;
      LAYER met5 ;
        RECT 105.015 3217.000 129.965 3219.000 ;
      LAYER met5 ;
        RECT 105.015 3200.600 129.965 3215.400 ;
      LAYER met5 ;
        RECT 105.015 3197.000 129.965 3199.000 ;
      LAYER met5 ;
        RECT 105.015 3180.600 129.965 3195.400 ;
      LAYER met5 ;
        RECT 105.015 3177.000 129.965 3179.000 ;
      LAYER met5 ;
        RECT 105.015 3160.600 129.965 3175.400 ;
      LAYER met5 ;
        RECT 105.015 3157.000 129.965 3159.000 ;
      LAYER met5 ;
        RECT 105.015 3140.600 129.965 3155.400 ;
        RECT 0.000 3135.130 103.415 3138.000 ;
      LAYER met5 ;
        RECT 105.015 3136.730 129.965 3139.000 ;
        RECT 131.565 3136.730 135.815 3275.270 ;
        RECT 137.415 3136.730 141.665 3275.270 ;
        RECT 143.265 3136.730 152.265 3275.270 ;
        RECT 153.865 3136.730 158.315 3275.270 ;
        RECT 159.915 3274.000 163.160 3275.270 ;
        RECT 159.915 3138.000 163.165 3274.000 ;
        RECT 159.915 3136.730 163.160 3138.000 ;
        RECT 164.765 3136.730 168.015 3275.270 ;
        RECT 169.615 3136.730 174.065 3275.270 ;
        RECT 175.665 3136.730 180.115 3275.270 ;
        RECT 181.715 3136.970 184.965 3274.965 ;
        RECT 186.565 3136.730 191.015 3275.270 ;
        RECT 192.615 3136.730 197.865 3275.270 ;
        RECT 3390.135 3268.730 3395.385 3417.270 ;
        RECT 3396.985 3268.730 3401.435 3417.270 ;
        RECT 3403.035 3269.035 3406.285 3417.030 ;
        RECT 3407.885 3268.730 3412.335 3417.270 ;
        RECT 3413.935 3268.730 3418.385 3417.270 ;
        RECT 3419.985 3268.730 3423.235 3417.270 ;
        RECT 3424.840 3416.000 3428.085 3417.270 ;
        RECT 3424.835 3270.000 3428.085 3416.000 ;
        RECT 3424.840 3268.730 3428.085 3270.000 ;
        RECT 3429.685 3268.730 3434.135 3417.270 ;
        RECT 3435.735 3268.730 3444.735 3417.270 ;
        RECT 3446.335 3268.730 3450.585 3417.270 ;
        RECT 3452.185 3268.730 3456.435 3417.270 ;
        RECT 3458.035 3414.000 3482.985 3417.270 ;
      LAYER met5 ;
        RECT 3484.585 3416.000 3588.000 3418.870 ;
      LAYER met5 ;
        RECT 3458.035 3409.000 3482.985 3411.000 ;
      LAYER met5 ;
        RECT 3458.035 3392.600 3482.985 3407.400 ;
      LAYER met5 ;
        RECT 3458.035 3389.000 3482.985 3391.000 ;
      LAYER met5 ;
        RECT 3458.035 3372.600 3482.985 3387.400 ;
      LAYER met5 ;
        RECT 3458.035 3369.000 3482.985 3371.000 ;
      LAYER met5 ;
        RECT 3458.035 3352.600 3482.985 3367.400 ;
      LAYER met5 ;
        RECT 3458.035 3349.000 3482.985 3351.000 ;
      LAYER met5 ;
        RECT 3458.035 3332.600 3482.985 3347.400 ;
      LAYER met5 ;
        RECT 3458.035 3329.000 3482.985 3331.000 ;
      LAYER met5 ;
        RECT 3458.035 3312.600 3482.985 3327.400 ;
      LAYER met5 ;
        RECT 3458.035 3309.000 3482.985 3311.000 ;
      LAYER met5 ;
        RECT 3458.035 3292.600 3482.985 3307.400 ;
      LAYER met5 ;
        RECT 3458.035 3289.000 3482.985 3291.000 ;
      LAYER met5 ;
        RECT 3458.035 3272.600 3482.985 3287.400 ;
      LAYER met5 ;
        RECT 3458.035 3268.730 3482.985 3271.000 ;
        RECT 3563.785 3270.000 3588.000 3416.000 ;
      LAYER met5 ;
        RECT 3403.035 3267.130 3406.285 3267.435 ;
        RECT 3484.585 3267.130 3588.000 3270.000 ;
        RECT 3390.135 3260.400 3588.000 3267.130 ;
        RECT 3390.135 3194.600 3490.960 3260.400 ;
        RECT 3556.610 3194.600 3588.000 3260.400 ;
        RECT 3390.135 3192.870 3588.000 3194.600 ;
        RECT 3403.035 3192.630 3406.285 3192.870 ;
        RECT 181.715 3135.130 184.965 3135.370 ;
        RECT 0.000 3133.400 197.865 3135.130 ;
        RECT 0.000 3067.600 31.390 3133.400 ;
        RECT 97.040 3067.600 197.865 3133.400 ;
        RECT 0.000 3060.870 197.865 3067.600 ;
        RECT 0.000 3058.000 103.415 3060.870 ;
        RECT 181.715 3060.565 184.965 3060.870 ;
      LAYER met5 ;
        RECT 0.000 2922.000 24.215 3058.000 ;
        RECT 105.015 3056.000 129.965 3059.270 ;
        RECT 105.015 3051.000 129.965 3053.000 ;
      LAYER met5 ;
        RECT 105.015 3044.600 129.965 3049.400 ;
      LAYER met5 ;
        RECT 105.015 3041.000 129.965 3043.000 ;
      LAYER met5 ;
        RECT 105.015 3024.600 129.965 3039.400 ;
      LAYER met5 ;
        RECT 105.015 3021.000 129.965 3023.000 ;
      LAYER met5 ;
        RECT 105.015 3004.600 129.965 3019.400 ;
      LAYER met5 ;
        RECT 105.015 3001.000 129.965 3003.000 ;
      LAYER met5 ;
        RECT 105.015 2984.600 129.965 2999.400 ;
      LAYER met5 ;
        RECT 105.015 2981.000 129.965 2983.000 ;
      LAYER met5 ;
        RECT 105.015 2964.600 129.965 2979.400 ;
      LAYER met5 ;
        RECT 105.015 2961.000 129.965 2963.000 ;
      LAYER met5 ;
        RECT 105.015 2944.600 129.965 2959.400 ;
      LAYER met5 ;
        RECT 105.015 2941.000 129.965 2943.000 ;
      LAYER met5 ;
        RECT 105.015 2924.600 129.965 2939.400 ;
        RECT 0.000 2919.130 103.415 2922.000 ;
      LAYER met5 ;
        RECT 105.015 2920.730 129.965 2923.000 ;
        RECT 131.565 2920.730 135.815 3059.270 ;
        RECT 137.415 2920.730 141.665 3059.270 ;
        RECT 143.265 2920.730 152.265 3059.270 ;
        RECT 153.865 2920.730 158.315 3059.270 ;
        RECT 159.915 3058.000 163.160 3059.270 ;
        RECT 159.915 2922.000 163.165 3058.000 ;
        RECT 159.915 2920.730 163.160 2922.000 ;
        RECT 164.765 2920.730 168.015 3059.270 ;
        RECT 169.615 2920.730 174.065 3059.270 ;
        RECT 175.665 2920.730 180.115 3059.270 ;
        RECT 181.715 2920.970 184.965 3058.965 ;
        RECT 186.565 2920.730 191.015 3059.270 ;
        RECT 192.615 2920.730 197.865 3059.270 ;
        RECT 3390.135 3043.730 3395.385 3191.270 ;
        RECT 3396.985 3043.730 3401.435 3191.270 ;
        RECT 3403.035 3044.035 3406.285 3191.030 ;
        RECT 3407.885 3043.730 3412.335 3191.270 ;
        RECT 3413.935 3043.730 3418.385 3191.270 ;
        RECT 3419.985 3043.730 3423.235 3191.270 ;
        RECT 3424.840 3190.000 3428.085 3191.270 ;
        RECT 3424.835 3045.000 3428.085 3190.000 ;
        RECT 3424.840 3043.730 3428.085 3045.000 ;
        RECT 3429.685 3043.730 3434.135 3191.270 ;
        RECT 3435.735 3043.730 3444.735 3191.270 ;
        RECT 3446.335 3043.730 3450.585 3191.270 ;
        RECT 3452.185 3043.730 3456.435 3191.270 ;
        RECT 3458.035 3189.000 3482.985 3191.270 ;
      LAYER met5 ;
        RECT 3484.585 3190.000 3588.000 3192.870 ;
      LAYER met5 ;
        RECT 3458.035 3184.000 3482.985 3186.000 ;
      LAYER met5 ;
        RECT 3458.035 3167.600 3482.985 3182.400 ;
      LAYER met5 ;
        RECT 3458.035 3164.000 3482.985 3166.000 ;
      LAYER met5 ;
        RECT 3458.035 3147.600 3482.985 3162.400 ;
      LAYER met5 ;
        RECT 3458.035 3144.000 3482.985 3146.000 ;
      LAYER met5 ;
        RECT 3458.035 3127.600 3482.985 3142.400 ;
      LAYER met5 ;
        RECT 3458.035 3124.000 3482.985 3126.000 ;
      LAYER met5 ;
        RECT 3458.035 3107.600 3482.985 3122.400 ;
      LAYER met5 ;
        RECT 3458.035 3104.000 3482.985 3106.000 ;
      LAYER met5 ;
        RECT 3458.035 3087.600 3482.985 3102.400 ;
      LAYER met5 ;
        RECT 3458.035 3084.000 3482.985 3086.000 ;
      LAYER met5 ;
        RECT 3458.035 3067.600 3482.985 3082.400 ;
      LAYER met5 ;
        RECT 3458.035 3064.000 3482.985 3066.000 ;
      LAYER met5 ;
        RECT 3458.035 3047.600 3482.985 3062.400 ;
      LAYER met5 ;
        RECT 3458.035 3043.730 3482.985 3046.000 ;
        RECT 3563.785 3045.000 3588.000 3190.000 ;
      LAYER met5 ;
        RECT 3403.035 3042.130 3406.285 3042.435 ;
        RECT 3484.585 3042.130 3588.000 3045.000 ;
        RECT 3390.135 3035.400 3588.000 3042.130 ;
        RECT 3390.135 2969.600 3490.960 3035.400 ;
        RECT 3556.610 2969.600 3588.000 3035.400 ;
        RECT 3390.135 2967.870 3588.000 2969.600 ;
        RECT 3403.035 2967.630 3406.285 2967.870 ;
        RECT 181.715 2919.130 184.965 2919.370 ;
        RECT 0.000 2917.400 197.865 2919.130 ;
        RECT 0.000 2851.600 31.390 2917.400 ;
        RECT 97.040 2851.600 197.865 2917.400 ;
        RECT 0.000 2844.870 197.865 2851.600 ;
        RECT 0.000 2842.000 103.415 2844.870 ;
        RECT 181.715 2844.565 184.965 2844.870 ;
      LAYER met5 ;
        RECT 0.000 2706.000 24.215 2842.000 ;
        RECT 105.015 2840.000 129.965 2843.270 ;
        RECT 105.015 2835.000 129.965 2837.000 ;
      LAYER met5 ;
        RECT 105.015 2828.600 129.965 2833.400 ;
      LAYER met5 ;
        RECT 105.015 2825.000 129.965 2827.000 ;
      LAYER met5 ;
        RECT 105.015 2808.600 129.965 2823.400 ;
      LAYER met5 ;
        RECT 105.015 2805.000 129.965 2807.000 ;
      LAYER met5 ;
        RECT 105.015 2788.600 129.965 2803.400 ;
      LAYER met5 ;
        RECT 105.015 2785.000 129.965 2787.000 ;
      LAYER met5 ;
        RECT 105.015 2768.600 129.965 2783.400 ;
      LAYER met5 ;
        RECT 105.015 2765.000 129.965 2767.000 ;
      LAYER met5 ;
        RECT 105.015 2748.600 129.965 2763.400 ;
      LAYER met5 ;
        RECT 105.015 2745.000 129.965 2747.000 ;
      LAYER met5 ;
        RECT 105.015 2728.600 129.965 2743.400 ;
      LAYER met5 ;
        RECT 105.015 2725.000 129.965 2727.000 ;
      LAYER met5 ;
        RECT 105.015 2708.600 129.965 2723.400 ;
        RECT 0.000 2703.130 103.415 2706.000 ;
      LAYER met5 ;
        RECT 105.015 2704.730 129.965 2707.000 ;
        RECT 131.565 2704.730 135.815 2843.270 ;
        RECT 137.415 2704.730 141.665 2843.270 ;
        RECT 143.265 2704.730 152.265 2843.270 ;
        RECT 153.865 2704.730 158.315 2843.270 ;
        RECT 159.915 2842.000 163.160 2843.270 ;
        RECT 159.915 2706.000 163.165 2842.000 ;
        RECT 159.915 2704.730 163.160 2706.000 ;
        RECT 164.765 2704.730 168.015 2843.270 ;
        RECT 169.615 2704.730 174.065 2843.270 ;
        RECT 175.665 2704.730 180.115 2843.270 ;
        RECT 181.715 2704.970 184.965 2842.965 ;
        RECT 186.565 2704.730 191.015 2843.270 ;
        RECT 192.615 2704.730 197.865 2843.270 ;
        RECT 3390.135 2817.730 3395.385 2966.270 ;
        RECT 3396.985 2817.730 3401.435 2966.270 ;
        RECT 3403.035 2818.035 3406.285 2966.030 ;
        RECT 3407.885 2817.730 3412.335 2966.270 ;
        RECT 3413.935 2817.730 3418.385 2966.270 ;
        RECT 3419.985 2817.730 3423.235 2966.270 ;
        RECT 3424.840 2965.000 3428.085 2966.270 ;
        RECT 3424.835 2819.000 3428.085 2965.000 ;
        RECT 3424.840 2817.730 3428.085 2819.000 ;
        RECT 3429.685 2817.730 3434.135 2966.270 ;
        RECT 3435.735 2817.730 3444.735 2966.270 ;
        RECT 3446.335 2817.730 3450.585 2966.270 ;
        RECT 3452.185 2817.730 3456.435 2966.270 ;
        RECT 3458.035 2963.000 3482.985 2966.270 ;
      LAYER met5 ;
        RECT 3484.585 2965.000 3588.000 2967.870 ;
      LAYER met5 ;
        RECT 3458.035 2958.000 3482.985 2960.000 ;
      LAYER met5 ;
        RECT 3458.035 2941.600 3482.985 2956.400 ;
      LAYER met5 ;
        RECT 3458.035 2938.000 3482.985 2940.000 ;
      LAYER met5 ;
        RECT 3458.035 2921.600 3482.985 2936.400 ;
      LAYER met5 ;
        RECT 3458.035 2918.000 3482.985 2920.000 ;
      LAYER met5 ;
        RECT 3458.035 2901.600 3482.985 2916.400 ;
      LAYER met5 ;
        RECT 3458.035 2898.000 3482.985 2900.000 ;
      LAYER met5 ;
        RECT 3458.035 2881.600 3482.985 2896.400 ;
      LAYER met5 ;
        RECT 3458.035 2878.000 3482.985 2880.000 ;
      LAYER met5 ;
        RECT 3458.035 2861.600 3482.985 2876.400 ;
      LAYER met5 ;
        RECT 3458.035 2858.000 3482.985 2860.000 ;
      LAYER met5 ;
        RECT 3458.035 2841.600 3482.985 2856.400 ;
      LAYER met5 ;
        RECT 3458.035 2838.000 3482.985 2840.000 ;
      LAYER met5 ;
        RECT 3458.035 2821.600 3482.985 2836.400 ;
      LAYER met5 ;
        RECT 3458.035 2817.730 3482.985 2820.000 ;
        RECT 3563.785 2819.000 3588.000 2965.000 ;
      LAYER met5 ;
        RECT 3403.035 2816.130 3406.285 2816.435 ;
        RECT 3484.585 2816.130 3588.000 2819.000 ;
        RECT 3390.135 2809.400 3588.000 2816.130 ;
        RECT 3390.135 2743.600 3490.960 2809.400 ;
        RECT 3556.610 2743.600 3588.000 2809.400 ;
        RECT 3390.135 2741.870 3588.000 2743.600 ;
        RECT 3403.035 2741.630 3406.285 2741.870 ;
        RECT 181.715 2703.130 184.965 2703.370 ;
        RECT 0.000 2701.400 197.865 2703.130 ;
        RECT 0.000 2635.600 31.390 2701.400 ;
        RECT 97.040 2635.600 197.865 2701.400 ;
        RECT 0.000 2628.870 197.865 2635.600 ;
        RECT 0.000 2626.000 103.415 2628.870 ;
        RECT 181.715 2628.565 184.965 2628.870 ;
      LAYER met5 ;
        RECT 0.000 2490.000 24.215 2626.000 ;
        RECT 105.015 2624.000 129.965 2627.270 ;
        RECT 105.015 2619.000 129.965 2621.000 ;
      LAYER met5 ;
        RECT 105.015 2612.600 129.965 2617.400 ;
      LAYER met5 ;
        RECT 105.015 2609.000 129.965 2611.000 ;
      LAYER met5 ;
        RECT 105.015 2592.600 129.965 2607.400 ;
      LAYER met5 ;
        RECT 105.015 2589.000 129.965 2591.000 ;
      LAYER met5 ;
        RECT 105.015 2572.600 129.965 2587.400 ;
      LAYER met5 ;
        RECT 105.015 2569.000 129.965 2571.000 ;
      LAYER met5 ;
        RECT 105.015 2552.600 129.965 2567.400 ;
      LAYER met5 ;
        RECT 105.015 2549.000 129.965 2551.000 ;
      LAYER met5 ;
        RECT 105.015 2532.600 129.965 2547.400 ;
      LAYER met5 ;
        RECT 105.015 2529.000 129.965 2531.000 ;
      LAYER met5 ;
        RECT 105.015 2512.600 129.965 2527.400 ;
      LAYER met5 ;
        RECT 105.015 2509.000 129.965 2511.000 ;
      LAYER met5 ;
        RECT 105.015 2492.600 129.965 2507.400 ;
        RECT 0.000 2487.130 103.415 2490.000 ;
      LAYER met5 ;
        RECT 105.015 2488.730 129.965 2491.000 ;
        RECT 131.565 2488.730 135.815 2627.270 ;
        RECT 137.415 2488.730 141.665 2627.270 ;
        RECT 143.265 2488.730 152.265 2627.270 ;
        RECT 153.865 2488.730 158.315 2627.270 ;
        RECT 159.915 2626.000 163.160 2627.270 ;
        RECT 159.915 2490.000 163.165 2626.000 ;
        RECT 159.915 2488.730 163.160 2490.000 ;
      LAYER met5 ;
        RECT 163.160 2487.130 163.165 2490.000 ;
      LAYER met5 ;
        RECT 164.765 2488.730 168.015 2627.270 ;
        RECT 169.615 2488.730 174.065 2627.270 ;
        RECT 175.665 2488.730 180.115 2627.270 ;
        RECT 186.565 2488.730 191.015 2627.270 ;
        RECT 192.615 2488.730 197.865 2627.270 ;
        RECT 3390.135 2592.730 3395.385 2740.270 ;
        RECT 3396.985 2592.730 3401.435 2740.270 ;
        RECT 3403.035 2593.035 3406.285 2740.030 ;
        RECT 3407.885 2592.730 3412.335 2740.270 ;
        RECT 3413.935 2592.730 3418.385 2740.270 ;
        RECT 3419.985 2592.730 3423.235 2740.270 ;
        RECT 3424.840 2739.000 3428.085 2740.270 ;
        RECT 3424.835 2594.000 3428.085 2739.000 ;
      LAYER met5 ;
        RECT 3403.035 2591.130 3406.285 2591.435 ;
        RECT 3424.835 2591.130 3424.840 2594.000 ;
      LAYER met5 ;
        RECT 3424.840 2592.730 3428.085 2594.000 ;
        RECT 3429.685 2592.730 3434.135 2740.270 ;
        RECT 3435.735 2592.730 3444.735 2740.270 ;
        RECT 3446.335 2592.730 3450.585 2740.270 ;
        RECT 3452.185 2592.730 3456.435 2740.270 ;
        RECT 3458.035 2738.000 3482.985 2740.270 ;
      LAYER met5 ;
        RECT 3484.585 2739.000 3588.000 2741.870 ;
      LAYER met5 ;
        RECT 3458.035 2733.000 3482.985 2735.000 ;
      LAYER met5 ;
        RECT 3458.035 2716.600 3482.985 2731.400 ;
      LAYER met5 ;
        RECT 3458.035 2713.000 3482.985 2715.000 ;
      LAYER met5 ;
        RECT 3458.035 2696.600 3482.985 2711.400 ;
      LAYER met5 ;
        RECT 3458.035 2693.000 3482.985 2695.000 ;
      LAYER met5 ;
        RECT 3458.035 2676.600 3482.985 2691.400 ;
      LAYER met5 ;
        RECT 3458.035 2673.000 3482.985 2675.000 ;
      LAYER met5 ;
        RECT 3458.035 2656.600 3482.985 2671.400 ;
      LAYER met5 ;
        RECT 3458.035 2653.000 3482.985 2655.000 ;
      LAYER met5 ;
        RECT 3458.035 2636.600 3482.985 2651.400 ;
      LAYER met5 ;
        RECT 3458.035 2633.000 3482.985 2635.000 ;
      LAYER met5 ;
        RECT 3458.035 2616.600 3482.985 2631.400 ;
      LAYER met5 ;
        RECT 3458.035 2613.000 3482.985 2615.000 ;
      LAYER met5 ;
        RECT 3458.035 2596.600 3482.985 2611.400 ;
      LAYER met5 ;
        RECT 3458.035 2592.730 3482.985 2595.000 ;
        RECT 3563.785 2594.000 3588.000 2739.000 ;
      LAYER met5 ;
        RECT 3484.585 2591.130 3588.000 2594.000 ;
        RECT 3390.135 2588.550 3588.000 2591.130 ;
        RECT 3390.135 2524.510 3491.520 2588.550 ;
      LAYER met5 ;
        RECT 3493.120 2526.110 3553.945 2586.950 ;
      LAYER met5 ;
        RECT 3555.545 2524.510 3588.000 2588.550 ;
        RECT 3390.135 2521.870 3588.000 2524.510 ;
        RECT 3403.035 2521.565 3406.285 2521.870 ;
        RECT 181.715 2487.130 184.965 2487.435 ;
        RECT 0.000 2484.490 197.865 2487.130 ;
        RECT 0.000 2420.450 32.455 2484.490 ;
        RECT 96.480 2420.450 197.865 2484.490 ;
        RECT 0.000 2417.870 197.865 2420.450 ;
        RECT 0.000 2415.000 103.415 2417.870 ;
      LAYER met5 ;
        RECT 0.000 2279.000 24.215 2415.000 ;
        RECT 105.015 2413.000 129.965 2416.270 ;
        RECT 105.015 2408.000 129.965 2410.000 ;
      LAYER met5 ;
        RECT 105.015 2401.600 129.965 2406.400 ;
      LAYER met5 ;
        RECT 105.015 2398.000 129.965 2400.000 ;
      LAYER met5 ;
        RECT 105.015 2381.600 129.965 2396.400 ;
      LAYER met5 ;
        RECT 105.015 2378.000 129.965 2380.000 ;
      LAYER met5 ;
        RECT 105.015 2361.600 129.965 2376.400 ;
      LAYER met5 ;
        RECT 105.015 2358.000 129.965 2360.000 ;
      LAYER met5 ;
        RECT 105.015 2341.600 129.965 2356.400 ;
      LAYER met5 ;
        RECT 105.015 2338.000 129.965 2340.000 ;
      LAYER met5 ;
        RECT 105.015 2321.600 129.965 2336.400 ;
      LAYER met5 ;
        RECT 105.015 2318.000 129.965 2320.000 ;
      LAYER met5 ;
        RECT 105.015 2301.600 129.965 2316.400 ;
      LAYER met5 ;
        RECT 105.015 2298.000 129.965 2300.000 ;
      LAYER met5 ;
        RECT 105.015 2281.600 129.965 2296.400 ;
        RECT 0.000 2276.130 103.415 2279.000 ;
      LAYER met5 ;
        RECT 105.015 2277.730 129.965 2280.000 ;
        RECT 131.565 2277.730 135.815 2416.270 ;
        RECT 137.415 2277.730 141.665 2416.270 ;
        RECT 143.265 2277.730 152.265 2416.270 ;
        RECT 159.915 2415.000 163.160 2416.270 ;
      LAYER met5 ;
        RECT 163.160 2415.000 163.165 2417.870 ;
        RECT 181.715 2417.565 184.965 2417.870 ;
      LAYER met5 ;
        RECT 159.915 2279.000 163.165 2415.000 ;
        RECT 159.915 2277.730 163.160 2279.000 ;
      LAYER met5 ;
        RECT 163.160 2276.130 163.165 2279.000 ;
      LAYER met5 ;
        RECT 164.765 2277.730 168.015 2416.270 ;
        RECT 169.615 2277.730 174.065 2416.270 ;
        RECT 175.665 2277.730 180.115 2416.270 ;
        RECT 186.565 2277.730 191.015 2416.270 ;
        RECT 192.615 2277.730 197.865 2416.270 ;
        RECT 3390.135 2372.730 3395.385 2520.270 ;
        RECT 3396.985 2372.730 3401.435 2520.270 ;
        RECT 3403.035 2373.035 3406.285 2519.965 ;
        RECT 3407.885 2372.730 3412.335 2520.270 ;
        RECT 3413.935 2372.730 3418.385 2520.270 ;
        RECT 3419.985 2372.730 3423.235 2520.270 ;
      LAYER met5 ;
        RECT 3424.835 2519.000 3424.840 2521.870 ;
      LAYER met5 ;
        RECT 3424.840 2519.000 3428.085 2520.270 ;
        RECT 3424.835 2374.000 3428.085 2519.000 ;
      LAYER met5 ;
        RECT 3403.035 2371.130 3406.285 2371.435 ;
        RECT 3424.835 2371.130 3424.840 2374.000 ;
      LAYER met5 ;
        RECT 3424.840 2372.730 3428.085 2374.000 ;
        RECT 3435.735 2372.730 3444.735 2520.270 ;
        RECT 3446.335 2372.730 3450.585 2520.270 ;
        RECT 3452.185 2372.730 3456.435 2520.270 ;
        RECT 3458.035 2518.000 3482.985 2520.270 ;
      LAYER met5 ;
        RECT 3484.585 2519.000 3588.000 2521.870 ;
      LAYER met5 ;
        RECT 3458.035 2513.000 3482.985 2515.000 ;
      LAYER met5 ;
        RECT 3458.035 2496.600 3482.985 2511.400 ;
      LAYER met5 ;
        RECT 3458.035 2493.000 3482.985 2495.000 ;
      LAYER met5 ;
        RECT 3458.035 2476.600 3482.985 2491.400 ;
      LAYER met5 ;
        RECT 3458.035 2473.000 3482.985 2475.000 ;
      LAYER met5 ;
        RECT 3458.035 2456.600 3482.985 2471.400 ;
      LAYER met5 ;
        RECT 3458.035 2453.000 3482.985 2455.000 ;
      LAYER met5 ;
        RECT 3458.035 2436.600 3482.985 2451.400 ;
      LAYER met5 ;
        RECT 3458.035 2433.000 3482.985 2435.000 ;
      LAYER met5 ;
        RECT 3458.035 2416.600 3482.985 2431.400 ;
      LAYER met5 ;
        RECT 3458.035 2413.000 3482.985 2415.000 ;
      LAYER met5 ;
        RECT 3458.035 2396.600 3482.985 2411.400 ;
      LAYER met5 ;
        RECT 3458.035 2393.000 3482.985 2395.000 ;
      LAYER met5 ;
        RECT 3458.035 2376.600 3482.985 2391.400 ;
      LAYER met5 ;
        RECT 3458.035 2372.730 3482.985 2375.000 ;
        RECT 3563.785 2374.000 3588.000 2519.000 ;
      LAYER met5 ;
        RECT 3484.585 2371.130 3588.000 2374.000 ;
        RECT 3390.135 2365.330 3588.000 2371.130 ;
        RECT 3390.135 2307.730 3488.300 2365.330 ;
        RECT 3558.765 2307.730 3588.000 2365.330 ;
        RECT 3390.135 2301.870 3588.000 2307.730 ;
        RECT 3403.035 2301.565 3406.285 2301.870 ;
        RECT 181.715 2276.130 184.965 2276.435 ;
        RECT 0.000 2270.270 197.865 2276.130 ;
        RECT 0.000 2212.670 29.235 2270.270 ;
        RECT 99.700 2212.670 197.865 2270.270 ;
        RECT 0.000 2206.870 197.865 2212.670 ;
        RECT 0.000 2204.000 103.415 2206.870 ;
      LAYER met5 ;
        RECT 0.000 2068.000 24.215 2204.000 ;
        RECT 105.015 2202.000 129.965 2205.270 ;
        RECT 105.015 2197.000 129.965 2199.000 ;
      LAYER met5 ;
        RECT 105.015 2190.600 129.965 2195.400 ;
      LAYER met5 ;
        RECT 105.015 2187.000 129.965 2189.000 ;
      LAYER met5 ;
        RECT 105.015 2170.600 129.965 2185.400 ;
      LAYER met5 ;
        RECT 105.015 2167.000 129.965 2169.000 ;
      LAYER met5 ;
        RECT 105.015 2150.600 129.965 2165.400 ;
      LAYER met5 ;
        RECT 105.015 2147.000 129.965 2149.000 ;
      LAYER met5 ;
        RECT 105.015 2130.600 129.965 2145.400 ;
      LAYER met5 ;
        RECT 105.015 2127.000 129.965 2129.000 ;
      LAYER met5 ;
        RECT 105.015 2110.600 129.965 2125.400 ;
      LAYER met5 ;
        RECT 105.015 2107.000 129.965 2109.000 ;
      LAYER met5 ;
        RECT 105.015 2090.600 129.965 2105.400 ;
      LAYER met5 ;
        RECT 105.015 2087.000 129.965 2089.000 ;
      LAYER met5 ;
        RECT 105.015 2070.600 129.965 2085.400 ;
        RECT 0.000 2065.130 103.415 2068.000 ;
      LAYER met5 ;
        RECT 105.015 2066.730 129.965 2069.000 ;
        RECT 131.565 2066.730 135.815 2205.270 ;
        RECT 137.415 2066.730 141.665 2205.270 ;
        RECT 143.265 2066.730 152.265 2205.270 ;
        RECT 159.915 2204.000 163.160 2205.270 ;
      LAYER met5 ;
        RECT 163.160 2204.000 163.165 2206.870 ;
        RECT 181.715 2206.565 184.965 2206.870 ;
      LAYER met5 ;
        RECT 159.915 2068.000 163.165 2204.000 ;
        RECT 159.915 2066.730 163.160 2068.000 ;
        RECT 164.765 2066.730 168.015 2205.270 ;
        RECT 169.615 2066.730 174.065 2205.270 ;
        RECT 175.665 2066.730 180.115 2205.270 ;
        RECT 181.715 2066.970 184.965 2204.965 ;
        RECT 186.565 2066.730 191.015 2205.270 ;
        RECT 192.615 2066.730 197.865 2205.270 ;
        RECT 3390.135 2151.730 3395.385 2300.270 ;
        RECT 3396.985 2151.730 3401.435 2300.270 ;
        RECT 3403.035 2152.035 3406.285 2299.965 ;
        RECT 3407.885 2151.730 3412.335 2300.270 ;
        RECT 3413.935 2151.730 3418.385 2300.270 ;
        RECT 3419.985 2151.730 3423.235 2300.270 ;
      LAYER met5 ;
        RECT 3424.835 2299.000 3424.840 2301.870 ;
      LAYER met5 ;
        RECT 3424.840 2299.000 3428.085 2300.270 ;
        RECT 3424.835 2153.000 3428.085 2299.000 ;
      LAYER met5 ;
        RECT 3403.035 2150.130 3406.285 2150.435 ;
        RECT 3424.835 2150.130 3424.840 2153.000 ;
      LAYER met5 ;
        RECT 3424.840 2151.730 3428.085 2153.000 ;
        RECT 3435.735 2151.730 3444.735 2300.270 ;
        RECT 3446.335 2151.730 3450.585 2300.270 ;
        RECT 3452.185 2151.730 3456.435 2300.270 ;
        RECT 3458.035 2297.000 3482.985 2300.270 ;
      LAYER met5 ;
        RECT 3484.585 2299.000 3588.000 2301.870 ;
      LAYER met5 ;
        RECT 3458.035 2292.000 3482.985 2294.000 ;
      LAYER met5 ;
        RECT 3458.035 2275.600 3482.985 2290.400 ;
      LAYER met5 ;
        RECT 3458.035 2272.000 3482.985 2274.000 ;
      LAYER met5 ;
        RECT 3458.035 2255.600 3482.985 2270.400 ;
      LAYER met5 ;
        RECT 3458.035 2252.000 3482.985 2254.000 ;
      LAYER met5 ;
        RECT 3458.035 2235.600 3482.985 2250.400 ;
      LAYER met5 ;
        RECT 3458.035 2232.000 3482.985 2234.000 ;
      LAYER met5 ;
        RECT 3458.035 2215.600 3482.985 2230.400 ;
      LAYER met5 ;
        RECT 3458.035 2212.000 3482.985 2214.000 ;
      LAYER met5 ;
        RECT 3458.035 2195.600 3482.985 2210.400 ;
      LAYER met5 ;
        RECT 3458.035 2192.000 3482.985 2194.000 ;
      LAYER met5 ;
        RECT 3458.035 2175.600 3482.985 2190.400 ;
      LAYER met5 ;
        RECT 3458.035 2172.000 3482.985 2174.000 ;
      LAYER met5 ;
        RECT 3458.035 2155.600 3482.985 2170.400 ;
      LAYER met5 ;
        RECT 3458.035 2151.730 3482.985 2154.000 ;
        RECT 3563.785 2153.000 3588.000 2299.000 ;
      LAYER met5 ;
        RECT 3484.585 2150.130 3588.000 2153.000 ;
        RECT 3390.135 2147.550 3588.000 2150.130 ;
        RECT 3390.135 2083.510 3491.520 2147.550 ;
      LAYER met5 ;
        RECT 3493.120 2085.110 3553.945 2145.950 ;
      LAYER met5 ;
        RECT 3555.545 2083.510 3588.000 2147.550 ;
        RECT 3390.135 2080.870 3588.000 2083.510 ;
        RECT 3403.035 2080.565 3406.285 2080.870 ;
        RECT 181.715 2065.130 184.965 2065.370 ;
        RECT 0.000 2063.400 197.865 2065.130 ;
        RECT 0.000 1997.600 31.390 2063.400 ;
        RECT 97.040 1997.600 197.865 2063.400 ;
        RECT 0.000 1990.870 197.865 1997.600 ;
        RECT 0.000 1988.000 103.415 1990.870 ;
        RECT 181.715 1990.565 184.965 1990.870 ;
      LAYER met5 ;
        RECT 0.000 1852.000 24.215 1988.000 ;
        RECT 105.015 1986.000 129.965 1989.270 ;
        RECT 105.015 1981.000 129.965 1983.000 ;
      LAYER met5 ;
        RECT 105.015 1974.600 129.965 1979.400 ;
      LAYER met5 ;
        RECT 105.015 1971.000 129.965 1973.000 ;
      LAYER met5 ;
        RECT 105.015 1954.600 129.965 1969.400 ;
      LAYER met5 ;
        RECT 105.015 1951.000 129.965 1953.000 ;
      LAYER met5 ;
        RECT 105.015 1934.600 129.965 1949.400 ;
      LAYER met5 ;
        RECT 105.015 1931.000 129.965 1933.000 ;
      LAYER met5 ;
        RECT 105.015 1914.600 129.965 1929.400 ;
      LAYER met5 ;
        RECT 105.015 1911.000 129.965 1913.000 ;
      LAYER met5 ;
        RECT 105.015 1894.600 129.965 1909.400 ;
      LAYER met5 ;
        RECT 105.015 1891.000 129.965 1893.000 ;
      LAYER met5 ;
        RECT 105.015 1874.600 129.965 1889.400 ;
      LAYER met5 ;
        RECT 105.015 1871.000 129.965 1873.000 ;
      LAYER met5 ;
        RECT 105.015 1854.600 129.965 1869.400 ;
        RECT 0.000 1849.130 103.415 1852.000 ;
      LAYER met5 ;
        RECT 105.015 1850.730 129.965 1853.000 ;
        RECT 131.565 1850.730 135.815 1989.270 ;
        RECT 137.415 1850.730 141.665 1989.270 ;
        RECT 143.265 1850.730 152.265 1989.270 ;
        RECT 153.865 1850.730 158.315 1989.270 ;
        RECT 159.915 1988.000 163.160 1989.270 ;
        RECT 159.915 1852.000 163.165 1988.000 ;
        RECT 159.915 1850.730 163.160 1852.000 ;
        RECT 164.765 1850.730 168.015 1989.270 ;
        RECT 169.615 1850.730 174.065 1989.270 ;
        RECT 175.665 1850.730 180.115 1989.270 ;
        RECT 181.715 1850.970 184.965 1988.965 ;
        RECT 186.565 1850.730 191.015 1989.270 ;
        RECT 192.615 1850.730 197.865 1989.270 ;
        RECT 3390.135 1931.730 3395.385 2079.270 ;
        RECT 3396.985 1931.730 3401.435 2079.270 ;
        RECT 3403.035 1932.035 3406.285 2078.965 ;
        RECT 3407.885 1931.730 3412.335 2079.270 ;
        RECT 3413.935 1931.730 3418.385 2079.270 ;
        RECT 3419.985 1931.730 3423.235 2079.270 ;
      LAYER met5 ;
        RECT 3424.835 2078.000 3424.840 2080.870 ;
      LAYER met5 ;
        RECT 3424.840 2078.000 3428.085 2079.270 ;
        RECT 3424.835 1933.000 3428.085 2078.000 ;
        RECT 3424.840 1931.730 3428.085 1933.000 ;
        RECT 3429.685 1931.730 3434.135 2079.270 ;
        RECT 3435.735 1931.730 3444.735 2079.270 ;
        RECT 3446.335 1931.730 3450.585 2079.270 ;
        RECT 3452.185 1931.730 3456.435 2079.270 ;
        RECT 3458.035 2077.000 3482.985 2079.270 ;
      LAYER met5 ;
        RECT 3484.585 2078.000 3588.000 2080.870 ;
      LAYER met5 ;
        RECT 3458.035 2072.000 3482.985 2074.000 ;
      LAYER met5 ;
        RECT 3458.035 2055.600 3482.985 2070.400 ;
      LAYER met5 ;
        RECT 3458.035 2052.000 3482.985 2054.000 ;
      LAYER met5 ;
        RECT 3458.035 2035.600 3482.985 2050.400 ;
      LAYER met5 ;
        RECT 3458.035 2032.000 3482.985 2034.000 ;
      LAYER met5 ;
        RECT 3458.035 2015.600 3482.985 2030.400 ;
      LAYER met5 ;
        RECT 3458.035 2012.000 3482.985 2014.000 ;
      LAYER met5 ;
        RECT 3458.035 1995.600 3482.985 2010.400 ;
      LAYER met5 ;
        RECT 3458.035 1992.000 3482.985 1994.000 ;
      LAYER met5 ;
        RECT 3458.035 1975.600 3482.985 1990.400 ;
      LAYER met5 ;
        RECT 3458.035 1972.000 3482.985 1974.000 ;
      LAYER met5 ;
        RECT 3458.035 1955.600 3482.985 1970.400 ;
      LAYER met5 ;
        RECT 3458.035 1952.000 3482.985 1954.000 ;
      LAYER met5 ;
        RECT 3458.035 1935.600 3482.985 1950.400 ;
      LAYER met5 ;
        RECT 3458.035 1931.730 3482.985 1934.000 ;
        RECT 3563.785 1933.000 3588.000 2078.000 ;
      LAYER met5 ;
        RECT 3403.035 1930.130 3406.285 1930.435 ;
        RECT 3484.585 1930.130 3588.000 1933.000 ;
        RECT 3390.135 1923.400 3588.000 1930.130 ;
        RECT 3390.135 1857.600 3490.960 1923.400 ;
        RECT 3556.610 1857.600 3588.000 1923.400 ;
        RECT 3390.135 1855.870 3588.000 1857.600 ;
        RECT 3403.035 1855.630 3406.285 1855.870 ;
        RECT 181.715 1849.130 184.965 1849.370 ;
        RECT 0.000 1847.400 197.865 1849.130 ;
        RECT 0.000 1781.600 31.390 1847.400 ;
        RECT 97.040 1781.600 197.865 1847.400 ;
        RECT 0.000 1774.870 197.865 1781.600 ;
        RECT 0.000 1772.000 103.415 1774.870 ;
        RECT 181.715 1774.565 184.965 1774.870 ;
      LAYER met5 ;
        RECT 0.000 1636.000 24.215 1772.000 ;
        RECT 105.015 1770.000 129.965 1773.270 ;
        RECT 105.015 1765.000 129.965 1767.000 ;
      LAYER met5 ;
        RECT 105.015 1758.600 129.965 1763.400 ;
      LAYER met5 ;
        RECT 105.015 1755.000 129.965 1757.000 ;
      LAYER met5 ;
        RECT 105.015 1738.600 129.965 1753.400 ;
      LAYER met5 ;
        RECT 105.015 1735.000 129.965 1737.000 ;
      LAYER met5 ;
        RECT 105.015 1718.600 129.965 1733.400 ;
      LAYER met5 ;
        RECT 105.015 1715.000 129.965 1717.000 ;
      LAYER met5 ;
        RECT 105.015 1698.600 129.965 1713.400 ;
      LAYER met5 ;
        RECT 105.015 1695.000 129.965 1697.000 ;
      LAYER met5 ;
        RECT 105.015 1678.600 129.965 1693.400 ;
      LAYER met5 ;
        RECT 105.015 1675.000 129.965 1677.000 ;
      LAYER met5 ;
        RECT 105.015 1658.600 129.965 1673.400 ;
      LAYER met5 ;
        RECT 105.015 1655.000 129.965 1657.000 ;
      LAYER met5 ;
        RECT 105.015 1638.600 129.965 1653.400 ;
        RECT 0.000 1633.130 103.415 1636.000 ;
      LAYER met5 ;
        RECT 105.015 1634.730 129.965 1637.000 ;
        RECT 131.565 1634.730 135.815 1773.270 ;
        RECT 137.415 1634.730 141.665 1773.270 ;
        RECT 143.265 1634.730 152.265 1773.270 ;
        RECT 153.865 1634.730 158.315 1773.270 ;
        RECT 159.915 1772.000 163.160 1773.270 ;
        RECT 159.915 1636.000 163.165 1772.000 ;
        RECT 159.915 1634.730 163.160 1636.000 ;
        RECT 164.765 1634.730 168.015 1773.270 ;
        RECT 169.615 1634.730 174.065 1773.270 ;
        RECT 175.665 1634.730 180.115 1773.270 ;
        RECT 181.715 1634.970 184.965 1772.965 ;
        RECT 186.565 1634.730 191.015 1773.270 ;
        RECT 192.615 1634.730 197.865 1773.270 ;
        RECT 3390.135 1705.730 3395.385 1854.270 ;
        RECT 3396.985 1705.730 3401.435 1854.270 ;
        RECT 3403.035 1706.035 3406.285 1854.030 ;
        RECT 3407.885 1705.730 3412.335 1854.270 ;
        RECT 3413.935 1705.730 3418.385 1854.270 ;
        RECT 3419.985 1705.730 3423.235 1854.270 ;
        RECT 3424.840 1853.000 3428.085 1854.270 ;
        RECT 3424.835 1707.000 3428.085 1853.000 ;
        RECT 3424.840 1705.730 3428.085 1707.000 ;
        RECT 3429.685 1705.730 3434.135 1854.270 ;
        RECT 3435.735 1705.730 3444.735 1854.270 ;
        RECT 3446.335 1705.730 3450.585 1854.270 ;
        RECT 3452.185 1705.730 3456.435 1854.270 ;
        RECT 3458.035 1851.000 3482.985 1854.270 ;
      LAYER met5 ;
        RECT 3484.585 1853.000 3588.000 1855.870 ;
      LAYER met5 ;
        RECT 3458.035 1846.000 3482.985 1848.000 ;
      LAYER met5 ;
        RECT 3458.035 1829.600 3482.985 1844.400 ;
      LAYER met5 ;
        RECT 3458.035 1826.000 3482.985 1828.000 ;
      LAYER met5 ;
        RECT 3458.035 1809.600 3482.985 1824.400 ;
      LAYER met5 ;
        RECT 3458.035 1806.000 3482.985 1808.000 ;
      LAYER met5 ;
        RECT 3458.035 1789.600 3482.985 1804.400 ;
      LAYER met5 ;
        RECT 3458.035 1786.000 3482.985 1788.000 ;
      LAYER met5 ;
        RECT 3458.035 1769.600 3482.985 1784.400 ;
      LAYER met5 ;
        RECT 3458.035 1766.000 3482.985 1768.000 ;
      LAYER met5 ;
        RECT 3458.035 1749.600 3482.985 1764.400 ;
      LAYER met5 ;
        RECT 3458.035 1746.000 3482.985 1748.000 ;
      LAYER met5 ;
        RECT 3458.035 1729.600 3482.985 1744.400 ;
      LAYER met5 ;
        RECT 3458.035 1726.000 3482.985 1728.000 ;
      LAYER met5 ;
        RECT 3458.035 1709.600 3482.985 1724.400 ;
      LAYER met5 ;
        RECT 3458.035 1705.730 3482.985 1708.000 ;
        RECT 3563.785 1707.000 3588.000 1853.000 ;
      LAYER met5 ;
        RECT 3403.035 1704.130 3406.285 1704.435 ;
        RECT 3484.585 1704.130 3588.000 1707.000 ;
        RECT 3390.135 1697.400 3588.000 1704.130 ;
        RECT 181.715 1633.130 184.965 1633.370 ;
        RECT 0.000 1631.400 197.865 1633.130 ;
        RECT 0.000 1565.600 31.390 1631.400 ;
        RECT 97.040 1565.600 197.865 1631.400 ;
        RECT 3390.135 1631.600 3490.960 1697.400 ;
        RECT 3556.610 1631.600 3588.000 1697.400 ;
        RECT 3390.135 1629.870 3588.000 1631.600 ;
        RECT 3403.035 1629.630 3406.285 1629.870 ;
        RECT 0.000 1558.870 197.865 1565.600 ;
        RECT 0.000 1556.000 103.415 1558.870 ;
        RECT 181.715 1558.565 184.965 1558.870 ;
      LAYER met5 ;
        RECT 0.000 1420.000 24.215 1556.000 ;
        RECT 105.015 1554.000 129.965 1557.270 ;
        RECT 105.015 1549.000 129.965 1551.000 ;
      LAYER met5 ;
        RECT 105.015 1542.600 129.965 1547.400 ;
      LAYER met5 ;
        RECT 105.015 1539.000 129.965 1541.000 ;
      LAYER met5 ;
        RECT 105.015 1522.600 129.965 1537.400 ;
      LAYER met5 ;
        RECT 105.015 1519.000 129.965 1521.000 ;
      LAYER met5 ;
        RECT 105.015 1502.600 129.965 1517.400 ;
      LAYER met5 ;
        RECT 105.015 1499.000 129.965 1501.000 ;
      LAYER met5 ;
        RECT 105.015 1482.600 129.965 1497.400 ;
      LAYER met5 ;
        RECT 105.015 1479.000 129.965 1481.000 ;
      LAYER met5 ;
        RECT 105.015 1462.600 129.965 1477.400 ;
      LAYER met5 ;
        RECT 105.015 1459.000 129.965 1461.000 ;
      LAYER met5 ;
        RECT 105.015 1442.600 129.965 1457.400 ;
      LAYER met5 ;
        RECT 105.015 1439.000 129.965 1441.000 ;
      LAYER met5 ;
        RECT 105.015 1422.600 129.965 1437.400 ;
        RECT 0.000 1417.130 103.415 1420.000 ;
      LAYER met5 ;
        RECT 105.015 1418.730 129.965 1421.000 ;
        RECT 131.565 1418.730 135.815 1557.270 ;
        RECT 137.415 1418.730 141.665 1557.270 ;
        RECT 143.265 1418.730 152.265 1557.270 ;
        RECT 153.865 1418.730 158.315 1557.270 ;
        RECT 159.915 1556.000 163.160 1557.270 ;
        RECT 159.915 1420.000 163.165 1556.000 ;
        RECT 159.915 1418.730 163.160 1420.000 ;
        RECT 164.765 1418.730 168.015 1557.270 ;
        RECT 169.615 1418.730 174.065 1557.270 ;
        RECT 175.665 1418.730 180.115 1557.270 ;
        RECT 181.715 1418.970 184.965 1556.965 ;
        RECT 186.565 1418.730 191.015 1557.270 ;
        RECT 192.615 1418.730 197.865 1557.270 ;
        RECT 3390.135 1480.730 3395.385 1628.270 ;
        RECT 3396.985 1480.730 3401.435 1628.270 ;
        RECT 3403.035 1481.035 3406.285 1628.030 ;
        RECT 3407.885 1480.730 3412.335 1628.270 ;
        RECT 3413.935 1480.730 3418.385 1628.270 ;
        RECT 3419.985 1480.730 3423.235 1628.270 ;
        RECT 3424.840 1627.000 3428.085 1628.270 ;
        RECT 3424.835 1482.000 3428.085 1627.000 ;
        RECT 3424.840 1480.730 3428.085 1482.000 ;
        RECT 3429.685 1480.730 3434.135 1628.270 ;
        RECT 3435.735 1480.730 3444.735 1628.270 ;
        RECT 3446.335 1480.730 3450.585 1628.270 ;
        RECT 3452.185 1480.730 3456.435 1628.270 ;
        RECT 3458.035 1626.000 3482.985 1628.270 ;
      LAYER met5 ;
        RECT 3484.585 1627.000 3588.000 1629.870 ;
      LAYER met5 ;
        RECT 3458.035 1621.000 3482.985 1623.000 ;
      LAYER met5 ;
        RECT 3458.035 1604.600 3482.985 1619.400 ;
      LAYER met5 ;
        RECT 3458.035 1601.000 3482.985 1603.000 ;
      LAYER met5 ;
        RECT 3458.035 1584.600 3482.985 1599.400 ;
      LAYER met5 ;
        RECT 3458.035 1581.000 3482.985 1583.000 ;
      LAYER met5 ;
        RECT 3458.035 1564.600 3482.985 1579.400 ;
      LAYER met5 ;
        RECT 3458.035 1561.000 3482.985 1563.000 ;
      LAYER met5 ;
        RECT 3458.035 1544.600 3482.985 1559.400 ;
      LAYER met5 ;
        RECT 3458.035 1541.000 3482.985 1543.000 ;
      LAYER met5 ;
        RECT 3458.035 1524.600 3482.985 1539.400 ;
      LAYER met5 ;
        RECT 3458.035 1521.000 3482.985 1523.000 ;
      LAYER met5 ;
        RECT 3458.035 1504.600 3482.985 1519.400 ;
      LAYER met5 ;
        RECT 3458.035 1501.000 3482.985 1503.000 ;
      LAYER met5 ;
        RECT 3458.035 1484.600 3482.985 1499.400 ;
      LAYER met5 ;
        RECT 3458.035 1480.730 3482.985 1483.000 ;
        RECT 3563.785 1482.000 3588.000 1627.000 ;
      LAYER met5 ;
        RECT 3403.035 1479.130 3406.285 1479.435 ;
        RECT 3484.585 1479.130 3588.000 1482.000 ;
        RECT 3390.135 1472.400 3588.000 1479.130 ;
        RECT 181.715 1417.130 184.965 1417.370 ;
        RECT 0.000 1415.400 197.865 1417.130 ;
        RECT 0.000 1349.600 31.390 1415.400 ;
        RECT 97.040 1349.600 197.865 1415.400 ;
        RECT 3390.135 1406.600 3490.960 1472.400 ;
        RECT 3556.610 1406.600 3588.000 1472.400 ;
        RECT 3390.135 1404.870 3588.000 1406.600 ;
        RECT 3403.035 1404.630 3406.285 1404.870 ;
        RECT 0.000 1342.870 197.865 1349.600 ;
        RECT 0.000 1340.000 103.415 1342.870 ;
        RECT 181.715 1342.565 184.965 1342.870 ;
      LAYER met5 ;
        RECT 0.000 1204.000 24.215 1340.000 ;
        RECT 105.015 1338.000 129.965 1341.270 ;
        RECT 105.015 1333.000 129.965 1335.000 ;
      LAYER met5 ;
        RECT 105.015 1326.600 129.965 1331.400 ;
      LAYER met5 ;
        RECT 105.015 1323.000 129.965 1325.000 ;
      LAYER met5 ;
        RECT 105.015 1306.600 129.965 1321.400 ;
      LAYER met5 ;
        RECT 105.015 1303.000 129.965 1305.000 ;
      LAYER met5 ;
        RECT 105.015 1286.600 129.965 1301.400 ;
      LAYER met5 ;
        RECT 105.015 1283.000 129.965 1285.000 ;
      LAYER met5 ;
        RECT 105.015 1266.600 129.965 1281.400 ;
      LAYER met5 ;
        RECT 105.015 1263.000 129.965 1265.000 ;
      LAYER met5 ;
        RECT 105.015 1246.600 129.965 1261.400 ;
      LAYER met5 ;
        RECT 105.015 1243.000 129.965 1245.000 ;
      LAYER met5 ;
        RECT 105.015 1226.600 129.965 1241.400 ;
      LAYER met5 ;
        RECT 105.015 1223.000 129.965 1225.000 ;
      LAYER met5 ;
        RECT 105.015 1206.600 129.965 1221.400 ;
        RECT 0.000 1201.130 103.415 1204.000 ;
      LAYER met5 ;
        RECT 105.015 1202.730 129.965 1205.000 ;
        RECT 131.565 1202.730 135.815 1341.270 ;
        RECT 137.415 1202.730 141.665 1341.270 ;
        RECT 143.265 1202.730 152.265 1341.270 ;
        RECT 153.865 1202.730 158.315 1341.270 ;
        RECT 159.915 1340.000 163.160 1341.270 ;
        RECT 159.915 1204.000 163.165 1340.000 ;
        RECT 159.915 1202.730 163.160 1204.000 ;
        RECT 164.765 1202.730 168.015 1341.270 ;
        RECT 169.615 1202.730 174.065 1341.270 ;
        RECT 175.665 1202.730 180.115 1341.270 ;
        RECT 181.715 1202.970 184.965 1340.965 ;
        RECT 186.565 1202.730 191.015 1341.270 ;
        RECT 192.615 1202.730 197.865 1341.270 ;
        RECT 3390.135 1255.730 3395.385 1403.270 ;
        RECT 3396.985 1255.730 3401.435 1403.270 ;
        RECT 3403.035 1256.035 3406.285 1403.030 ;
        RECT 3407.885 1255.730 3412.335 1403.270 ;
        RECT 3413.935 1255.730 3418.385 1403.270 ;
        RECT 3419.985 1255.730 3423.235 1403.270 ;
        RECT 3424.840 1402.000 3428.085 1403.270 ;
        RECT 3424.835 1257.000 3428.085 1402.000 ;
        RECT 3424.840 1255.730 3428.085 1257.000 ;
        RECT 3429.685 1255.730 3434.135 1403.270 ;
        RECT 3435.735 1255.730 3444.735 1403.270 ;
        RECT 3446.335 1255.730 3450.585 1403.270 ;
        RECT 3452.185 1255.730 3456.435 1403.270 ;
        RECT 3458.035 1401.000 3482.985 1403.270 ;
      LAYER met5 ;
        RECT 3484.585 1402.000 3588.000 1404.870 ;
      LAYER met5 ;
        RECT 3458.035 1396.000 3482.985 1398.000 ;
      LAYER met5 ;
        RECT 3458.035 1379.600 3482.985 1394.400 ;
      LAYER met5 ;
        RECT 3458.035 1376.000 3482.985 1378.000 ;
      LAYER met5 ;
        RECT 3458.035 1359.600 3482.985 1374.400 ;
      LAYER met5 ;
        RECT 3458.035 1356.000 3482.985 1358.000 ;
      LAYER met5 ;
        RECT 3458.035 1339.600 3482.985 1354.400 ;
      LAYER met5 ;
        RECT 3458.035 1336.000 3482.985 1338.000 ;
      LAYER met5 ;
        RECT 3458.035 1319.600 3482.985 1334.400 ;
      LAYER met5 ;
        RECT 3458.035 1316.000 3482.985 1318.000 ;
      LAYER met5 ;
        RECT 3458.035 1299.600 3482.985 1314.400 ;
      LAYER met5 ;
        RECT 3458.035 1296.000 3482.985 1298.000 ;
      LAYER met5 ;
        RECT 3458.035 1279.600 3482.985 1294.400 ;
      LAYER met5 ;
        RECT 3458.035 1276.000 3482.985 1278.000 ;
      LAYER met5 ;
        RECT 3458.035 1259.600 3482.985 1274.400 ;
      LAYER met5 ;
        RECT 3458.035 1255.730 3482.985 1258.000 ;
        RECT 3563.785 1257.000 3588.000 1402.000 ;
      LAYER met5 ;
        RECT 3403.035 1254.130 3406.285 1254.435 ;
        RECT 3484.585 1254.130 3588.000 1257.000 ;
        RECT 3390.135 1247.400 3588.000 1254.130 ;
        RECT 181.715 1201.130 184.965 1201.370 ;
        RECT 0.000 1199.400 197.865 1201.130 ;
        RECT 0.000 1133.600 31.390 1199.400 ;
        RECT 97.040 1133.600 197.865 1199.400 ;
        RECT 3390.135 1181.600 3490.960 1247.400 ;
        RECT 3556.610 1181.600 3588.000 1247.400 ;
        RECT 3390.135 1179.870 3588.000 1181.600 ;
        RECT 3403.035 1179.630 3406.285 1179.870 ;
        RECT 0.000 1126.870 197.865 1133.600 ;
        RECT 0.000 1124.000 103.415 1126.870 ;
        RECT 181.715 1126.565 184.965 1126.870 ;
      LAYER met5 ;
        RECT 0.000 988.000 24.215 1124.000 ;
        RECT 105.015 1122.000 129.965 1125.270 ;
        RECT 105.015 1117.000 129.965 1119.000 ;
      LAYER met5 ;
        RECT 105.015 1110.600 129.965 1115.400 ;
      LAYER met5 ;
        RECT 105.015 1107.000 129.965 1109.000 ;
      LAYER met5 ;
        RECT 105.015 1090.600 129.965 1105.400 ;
      LAYER met5 ;
        RECT 105.015 1087.000 129.965 1089.000 ;
      LAYER met5 ;
        RECT 105.015 1070.600 129.965 1085.400 ;
      LAYER met5 ;
        RECT 105.015 1067.000 129.965 1069.000 ;
      LAYER met5 ;
        RECT 105.015 1050.600 129.965 1065.400 ;
      LAYER met5 ;
        RECT 105.015 1047.000 129.965 1049.000 ;
      LAYER met5 ;
        RECT 105.015 1030.600 129.965 1045.400 ;
      LAYER met5 ;
        RECT 105.015 1027.000 129.965 1029.000 ;
      LAYER met5 ;
        RECT 105.015 1010.600 129.965 1025.400 ;
      LAYER met5 ;
        RECT 105.015 1007.000 129.965 1009.000 ;
      LAYER met5 ;
        RECT 105.015 990.600 129.965 1005.400 ;
        RECT 0.000 985.130 103.415 988.000 ;
      LAYER met5 ;
        RECT 105.015 986.730 129.965 989.000 ;
        RECT 131.565 986.730 135.815 1125.270 ;
        RECT 137.415 986.730 141.665 1125.270 ;
        RECT 143.265 986.730 152.265 1125.270 ;
        RECT 153.865 986.730 158.315 1125.270 ;
        RECT 159.915 1124.000 163.160 1125.270 ;
        RECT 159.915 988.000 163.165 1124.000 ;
        RECT 159.915 986.730 163.160 988.000 ;
        RECT 164.765 986.730 168.015 1125.270 ;
        RECT 169.615 986.730 174.065 1125.270 ;
        RECT 175.665 986.730 180.115 1125.270 ;
        RECT 181.715 986.970 184.965 1124.965 ;
        RECT 186.565 986.730 191.015 1125.270 ;
        RECT 192.615 986.730 197.865 1125.270 ;
        RECT 3390.135 1029.730 3395.385 1178.270 ;
        RECT 3396.985 1029.730 3401.435 1178.270 ;
        RECT 3403.035 1030.035 3406.285 1178.030 ;
        RECT 3407.885 1029.730 3412.335 1178.270 ;
        RECT 3413.935 1029.730 3418.385 1178.270 ;
        RECT 3419.985 1029.730 3423.235 1178.270 ;
        RECT 3424.840 1177.000 3428.085 1178.270 ;
        RECT 3424.835 1031.000 3428.085 1177.000 ;
        RECT 3424.840 1029.730 3428.085 1031.000 ;
        RECT 3429.685 1029.730 3434.135 1178.270 ;
        RECT 3435.735 1029.730 3444.735 1178.270 ;
        RECT 3446.335 1029.730 3450.585 1178.270 ;
        RECT 3452.185 1029.730 3456.435 1178.270 ;
        RECT 3458.035 1175.000 3482.985 1178.270 ;
      LAYER met5 ;
        RECT 3484.585 1177.000 3588.000 1179.870 ;
      LAYER met5 ;
        RECT 3458.035 1170.000 3482.985 1172.000 ;
      LAYER met5 ;
        RECT 3458.035 1153.600 3482.985 1168.400 ;
      LAYER met5 ;
        RECT 3458.035 1150.000 3482.985 1152.000 ;
      LAYER met5 ;
        RECT 3458.035 1133.600 3482.985 1148.400 ;
      LAYER met5 ;
        RECT 3458.035 1130.000 3482.985 1132.000 ;
      LAYER met5 ;
        RECT 3458.035 1113.600 3482.985 1128.400 ;
      LAYER met5 ;
        RECT 3458.035 1110.000 3482.985 1112.000 ;
      LAYER met5 ;
        RECT 3458.035 1093.600 3482.985 1108.400 ;
      LAYER met5 ;
        RECT 3458.035 1090.000 3482.985 1092.000 ;
      LAYER met5 ;
        RECT 3458.035 1073.600 3482.985 1088.400 ;
      LAYER met5 ;
        RECT 3458.035 1070.000 3482.985 1072.000 ;
      LAYER met5 ;
        RECT 3458.035 1053.600 3482.985 1068.400 ;
      LAYER met5 ;
        RECT 3458.035 1050.000 3482.985 1052.000 ;
      LAYER met5 ;
        RECT 3458.035 1033.600 3482.985 1048.400 ;
      LAYER met5 ;
        RECT 3458.035 1029.730 3482.985 1032.000 ;
        RECT 3563.785 1031.000 3588.000 1177.000 ;
      LAYER met5 ;
        RECT 3403.035 1028.130 3406.285 1028.435 ;
        RECT 3484.585 1028.130 3588.000 1031.000 ;
        RECT 3390.135 1021.400 3588.000 1028.130 ;
        RECT 181.715 985.130 184.965 985.370 ;
        RECT 0.000 983.400 197.865 985.130 ;
        RECT 0.000 917.600 31.390 983.400 ;
        RECT 97.040 917.600 197.865 983.400 ;
        RECT 3390.135 955.600 3490.960 1021.400 ;
        RECT 3556.610 955.600 3588.000 1021.400 ;
        RECT 3390.135 953.870 3588.000 955.600 ;
        RECT 3403.035 953.630 3406.285 953.870 ;
        RECT 0.000 910.870 197.865 917.600 ;
        RECT 0.000 908.000 103.415 910.870 ;
        RECT 181.715 910.565 184.965 910.870 ;
      LAYER met5 ;
        RECT 0.000 626.000 24.215 908.000 ;
        RECT 105.015 906.000 129.965 909.270 ;
        RECT 105.015 901.000 129.965 903.000 ;
      LAYER met5 ;
        RECT 105.015 894.600 129.965 899.400 ;
      LAYER met5 ;
        RECT 105.015 891.000 129.965 893.000 ;
      LAYER met5 ;
        RECT 105.015 874.600 129.965 889.400 ;
      LAYER met5 ;
        RECT 105.015 871.000 129.965 873.000 ;
      LAYER met5 ;
        RECT 105.015 854.600 129.965 869.400 ;
      LAYER met5 ;
        RECT 105.015 851.000 129.965 853.000 ;
      LAYER met5 ;
        RECT 105.015 834.600 129.965 849.400 ;
      LAYER met5 ;
        RECT 105.015 831.000 129.965 833.000 ;
      LAYER met5 ;
        RECT 105.015 814.600 129.965 829.400 ;
      LAYER met5 ;
        RECT 105.015 811.000 129.965 813.000 ;
      LAYER met5 ;
        RECT 105.015 794.600 129.965 809.400 ;
      LAYER met5 ;
        RECT 105.015 791.000 129.965 793.000 ;
      LAYER met5 ;
        RECT 105.015 774.600 129.965 789.400 ;
      LAYER met5 ;
        RECT 105.015 760.000 129.965 773.000 ;
        RECT 105.015 755.000 129.965 757.000 ;
      LAYER met5 ;
        RECT 105.015 748.600 129.965 753.400 ;
      LAYER met5 ;
        RECT 105.015 745.000 129.965 747.000 ;
      LAYER met5 ;
        RECT 105.015 728.600 129.965 743.400 ;
      LAYER met5 ;
        RECT 105.015 725.000 129.965 727.000 ;
      LAYER met5 ;
        RECT 105.015 708.600 129.965 723.400 ;
      LAYER met5 ;
        RECT 105.015 705.000 129.965 707.000 ;
      LAYER met5 ;
        RECT 105.015 688.600 129.965 703.400 ;
      LAYER met5 ;
        RECT 105.015 685.000 129.965 687.000 ;
      LAYER met5 ;
        RECT 105.015 668.600 129.965 683.400 ;
      LAYER met5 ;
        RECT 105.015 665.000 129.965 667.000 ;
      LAYER met5 ;
        RECT 105.015 648.600 129.965 663.400 ;
      LAYER met5 ;
        RECT 105.015 645.000 129.965 647.000 ;
      LAYER met5 ;
        RECT 105.015 628.600 129.965 643.400 ;
        RECT 0.000 623.130 103.415 626.000 ;
      LAYER met5 ;
        RECT 131.565 624.730 135.815 909.270 ;
        RECT 137.415 624.730 141.665 909.270 ;
        RECT 143.265 767.000 152.265 909.270 ;
        RECT 153.865 772.000 158.315 909.270 ;
        RECT 159.915 908.000 163.160 909.270 ;
        RECT 159.915 767.000 163.165 908.000 ;
        RECT 143.265 624.730 152.265 762.000 ;
        RECT 153.865 624.730 158.315 767.000 ;
        RECT 159.915 626.000 163.165 762.000 ;
        RECT 159.915 624.730 163.160 626.000 ;
      LAYER met5 ;
        RECT 163.160 623.130 163.165 626.000 ;
      LAYER met5 ;
        RECT 164.765 624.730 168.015 909.270 ;
        RECT 169.615 624.730 174.065 909.270 ;
        RECT 181.715 767.000 184.965 908.965 ;
        RECT 186.565 772.000 191.015 909.270 ;
        RECT 181.715 625.035 184.965 762.000 ;
        RECT 186.565 624.730 191.015 767.000 ;
        RECT 192.615 624.730 197.865 909.270 ;
        RECT 3390.135 804.730 3395.385 952.270 ;
        RECT 3396.985 804.730 3401.435 952.270 ;
        RECT 3403.035 805.035 3406.285 952.030 ;
        RECT 3407.885 804.730 3412.335 952.270 ;
        RECT 3413.935 804.730 3418.385 952.270 ;
        RECT 3419.985 804.730 3423.235 952.270 ;
        RECT 3424.840 951.000 3428.085 952.270 ;
        RECT 3424.835 806.000 3428.085 951.000 ;
        RECT 3424.840 804.730 3428.085 806.000 ;
        RECT 3429.685 804.730 3434.135 952.270 ;
        RECT 3435.735 804.730 3444.735 952.270 ;
        RECT 3446.335 804.730 3450.585 952.270 ;
        RECT 3452.185 804.730 3456.435 952.270 ;
        RECT 3458.035 950.000 3482.985 952.270 ;
      LAYER met5 ;
        RECT 3484.585 951.000 3588.000 953.870 ;
      LAYER met5 ;
        RECT 3458.035 945.000 3482.985 947.000 ;
      LAYER met5 ;
        RECT 3458.035 928.600 3482.985 943.400 ;
      LAYER met5 ;
        RECT 3458.035 925.000 3482.985 927.000 ;
      LAYER met5 ;
        RECT 3458.035 908.600 3482.985 923.400 ;
      LAYER met5 ;
        RECT 3458.035 905.000 3482.985 907.000 ;
      LAYER met5 ;
        RECT 3458.035 888.600 3482.985 903.400 ;
      LAYER met5 ;
        RECT 3458.035 885.000 3482.985 887.000 ;
      LAYER met5 ;
        RECT 3458.035 868.600 3482.985 883.400 ;
      LAYER met5 ;
        RECT 3458.035 865.000 3482.985 867.000 ;
      LAYER met5 ;
        RECT 3458.035 848.600 3482.985 863.400 ;
      LAYER met5 ;
        RECT 3458.035 845.000 3482.985 847.000 ;
      LAYER met5 ;
        RECT 3458.035 828.600 3482.985 843.400 ;
      LAYER met5 ;
        RECT 3458.035 825.000 3482.985 827.000 ;
      LAYER met5 ;
        RECT 3458.035 808.600 3482.985 823.400 ;
      LAYER met5 ;
        RECT 3458.035 804.730 3482.985 807.000 ;
        RECT 3563.785 806.000 3588.000 951.000 ;
      LAYER met5 ;
        RECT 3403.035 803.130 3406.285 803.435 ;
        RECT 3484.585 803.130 3588.000 806.000 ;
        RECT 3390.135 796.400 3588.000 803.130 ;
        RECT 3390.135 730.600 3490.960 796.400 ;
        RECT 3556.610 730.600 3588.000 796.400 ;
        RECT 3390.135 728.870 3588.000 730.600 ;
        RECT 3403.035 728.630 3406.285 728.870 ;
        RECT 181.715 623.130 184.965 623.435 ;
        RECT 0.000 620.490 197.865 623.130 ;
        RECT 0.000 556.450 32.455 620.490 ;
        RECT 96.480 556.450 197.865 620.490 ;
      LAYER met5 ;
        RECT 3390.135 578.730 3395.385 727.270 ;
        RECT 3396.985 578.730 3401.435 727.270 ;
        RECT 3403.035 579.035 3406.285 727.030 ;
        RECT 3407.885 578.730 3412.335 727.270 ;
        RECT 3413.935 578.730 3418.385 727.270 ;
        RECT 3419.985 578.730 3423.235 727.270 ;
        RECT 3424.840 726.000 3428.085 727.270 ;
        RECT 3424.835 580.000 3428.085 726.000 ;
        RECT 3424.840 578.730 3428.085 580.000 ;
        RECT 3429.685 578.730 3434.135 727.270 ;
        RECT 3435.735 578.730 3444.735 727.270 ;
        RECT 3446.335 578.730 3450.585 727.270 ;
        RECT 3452.185 578.730 3456.435 727.270 ;
        RECT 3458.035 724.000 3482.985 727.270 ;
      LAYER met5 ;
        RECT 3484.585 726.000 3588.000 728.870 ;
      LAYER met5 ;
        RECT 3458.035 719.000 3482.985 721.000 ;
      LAYER met5 ;
        RECT 3458.035 702.600 3482.985 717.400 ;
      LAYER met5 ;
        RECT 3458.035 699.000 3482.985 701.000 ;
      LAYER met5 ;
        RECT 3458.035 682.600 3482.985 697.400 ;
      LAYER met5 ;
        RECT 3458.035 679.000 3482.985 681.000 ;
      LAYER met5 ;
        RECT 3458.035 662.600 3482.985 677.400 ;
      LAYER met5 ;
        RECT 3458.035 659.000 3482.985 661.000 ;
      LAYER met5 ;
        RECT 3458.035 642.600 3482.985 657.400 ;
      LAYER met5 ;
        RECT 3458.035 639.000 3482.985 641.000 ;
      LAYER met5 ;
        RECT 3458.035 622.600 3482.985 637.400 ;
      LAYER met5 ;
        RECT 3458.035 619.000 3482.985 621.000 ;
      LAYER met5 ;
        RECT 3458.035 602.600 3482.985 617.400 ;
      LAYER met5 ;
        RECT 3458.035 599.000 3482.985 601.000 ;
      LAYER met5 ;
        RECT 3458.035 582.600 3482.985 597.400 ;
      LAYER met5 ;
        RECT 3458.035 578.730 3482.985 581.000 ;
        RECT 3563.785 580.000 3588.000 726.000 ;
      LAYER met5 ;
        RECT 3403.035 577.130 3406.285 577.435 ;
        RECT 3484.585 577.130 3588.000 580.000 ;
        RECT 0.000 553.870 197.865 556.450 ;
        RECT 3390.135 570.400 3588.000 577.130 ;
        RECT 0.000 551.000 103.415 553.870 ;
      LAYER met5 ;
        RECT 0.000 415.000 24.215 551.000 ;
        RECT 105.015 544.000 129.965 546.000 ;
      LAYER met5 ;
        RECT 105.015 537.600 129.965 542.400 ;
      LAYER met5 ;
        RECT 105.015 534.000 129.965 536.000 ;
      LAYER met5 ;
        RECT 105.015 517.600 129.965 532.400 ;
      LAYER met5 ;
        RECT 105.015 514.000 129.965 516.000 ;
      LAYER met5 ;
        RECT 105.015 497.600 129.965 512.400 ;
      LAYER met5 ;
        RECT 105.015 494.000 129.965 496.000 ;
      LAYER met5 ;
        RECT 105.015 477.600 129.965 492.400 ;
      LAYER met5 ;
        RECT 105.015 474.000 129.965 476.000 ;
      LAYER met5 ;
        RECT 105.015 457.600 129.965 472.400 ;
      LAYER met5 ;
        RECT 105.015 454.000 129.965 456.000 ;
      LAYER met5 ;
        RECT 105.015 437.600 129.965 452.400 ;
      LAYER met5 ;
        RECT 105.015 434.000 129.965 436.000 ;
      LAYER met5 ;
        RECT 105.015 417.600 129.965 432.400 ;
        RECT 0.000 412.130 103.415 415.000 ;
      LAYER met5 ;
        RECT 105.015 413.730 129.965 416.000 ;
        RECT 131.565 413.730 135.815 552.270 ;
        RECT 137.415 413.730 141.665 552.270 ;
        RECT 143.265 413.730 152.265 552.270 ;
        RECT 153.865 413.730 158.315 552.270 ;
        RECT 159.915 551.000 163.160 552.270 ;
      LAYER met5 ;
        RECT 163.160 551.000 163.165 553.870 ;
        RECT 181.715 553.565 184.965 553.870 ;
      LAYER met5 ;
        RECT 159.915 415.000 163.165 551.000 ;
        RECT 159.915 413.730 163.160 415.000 ;
        RECT 164.765 413.730 168.015 552.270 ;
        RECT 169.615 413.730 174.065 552.270 ;
        RECT 181.715 414.035 184.965 551.965 ;
        RECT 192.615 413.730 197.865 552.270 ;
      LAYER met5 ;
        RECT 3390.135 504.600 3490.960 570.400 ;
        RECT 3556.610 504.600 3588.000 570.400 ;
        RECT 3390.135 502.870 3588.000 504.600 ;
        RECT 3403.035 502.630 3406.285 502.870 ;
        RECT 181.715 412.130 184.965 412.435 ;
        RECT 0.000 406.270 197.865 412.130 ;
        RECT 0.000 348.670 29.235 406.270 ;
        RECT 99.700 348.670 197.865 406.270 ;
        RECT 0.000 342.870 197.865 348.670 ;
        RECT 0.000 340.000 103.415 342.870 ;
        RECT 181.715 342.565 184.965 342.870 ;
      LAYER met5 ;
        RECT 0.000 204.000 24.215 340.000 ;
        RECT 105.015 338.000 129.965 341.270 ;
        RECT 105.015 333.000 129.965 335.000 ;
      LAYER met5 ;
        RECT 105.015 326.600 129.965 331.400 ;
      LAYER met5 ;
        RECT 105.015 323.000 129.965 325.000 ;
      LAYER met5 ;
        RECT 105.015 306.600 129.965 321.400 ;
      LAYER met5 ;
        RECT 105.015 303.000 129.965 305.000 ;
      LAYER met5 ;
        RECT 105.015 286.600 129.965 301.400 ;
      LAYER met5 ;
        RECT 105.015 283.000 129.965 285.000 ;
      LAYER met5 ;
        RECT 105.015 266.600 129.965 281.400 ;
      LAYER met5 ;
        RECT 105.015 263.000 129.965 265.000 ;
      LAYER met5 ;
        RECT 105.015 246.600 129.965 261.400 ;
      LAYER met5 ;
        RECT 105.015 243.000 129.965 245.000 ;
      LAYER met5 ;
        RECT 105.015 226.600 129.965 241.400 ;
      LAYER met5 ;
        RECT 105.015 223.000 129.965 225.000 ;
      LAYER met5 ;
        RECT 105.015 206.600 129.965 221.400 ;
        RECT 0.000 200.545 103.415 204.000 ;
      LAYER met5 ;
        RECT 105.015 202.145 129.965 205.000 ;
        RECT 131.565 202.730 135.815 341.270 ;
        RECT 137.415 202.730 141.665 341.270 ;
      LAYER met5 ;
        RECT 131.565 200.545 141.665 201.130 ;
        RECT 0.000 175.245 141.665 200.545 ;
      LAYER met5 ;
        RECT 143.265 176.845 152.265 341.270 ;
        RECT 153.865 202.730 158.315 341.270 ;
        RECT 159.915 340.000 163.160 341.270 ;
        RECT 159.915 204.000 163.165 340.000 ;
        RECT 159.915 202.730 163.160 204.000 ;
        RECT 164.765 202.730 168.015 341.270 ;
        RECT 169.615 202.730 174.065 341.270 ;
        RECT 175.665 202.730 180.115 341.270 ;
        RECT 181.715 202.745 184.965 340.965 ;
        RECT 192.615 202.730 197.865 341.270 ;
      LAYER met5 ;
        RECT 181.715 201.130 184.965 201.145 ;
        RECT 199.465 201.130 200.000 204.000 ;
        RECT 153.865 199.465 200.000 201.130 ;
        RECT 3384.000 199.465 3388.535 200.000 ;
        RECT 153.865 192.615 196.050 199.465 ;
        RECT 197.865 197.865 198.400 199.465 ;
        POLYGON 198.400 199.465 200.000 197.865 198.400 197.865 ;
        RECT 3386.870 198.400 3388.535 199.465 ;
        POLYGON 3390.135 200.000 3390.135 198.400 3388.535 198.400 ;
        RECT 3386.870 197.865 3390.135 198.400 ;
      LAYER met5 ;
        RECT 197.650 192.615 395.270 197.865 ;
      LAYER met5 ;
        RECT 153.865 184.965 194.615 192.615 ;
      LAYER met5 ;
        RECT 237.000 191.015 357.000 192.615 ;
        RECT 196.215 186.565 395.270 191.015 ;
      LAYER met5 ;
        RECT 396.870 184.965 466.130 197.865 ;
      LAYER met5 ;
        RECT 467.730 192.615 664.270 197.865 ;
        RECT 506.000 191.015 626.000 192.615 ;
        RECT 467.730 186.565 664.270 191.015 ;
      LAYER met5 ;
        RECT 665.870 184.965 735.130 197.865 ;
      LAYER met5 ;
        RECT 736.730 192.615 933.270 197.865 ;
        RECT 775.000 191.015 895.000 192.615 ;
        RECT 736.730 186.565 933.270 191.015 ;
      LAYER met5 ;
        RECT 934.870 184.965 1009.130 197.865 ;
      LAYER met5 ;
        RECT 1010.730 192.615 1207.270 197.865 ;
        RECT 1049.000 191.015 1169.000 192.615 ;
        RECT 1010.730 186.565 1207.270 191.015 ;
      LAYER met5 ;
        RECT 1208.870 184.965 1278.130 197.865 ;
      LAYER met5 ;
        RECT 1279.730 192.615 1476.270 197.865 ;
        RECT 1318.000 191.015 1438.000 192.615 ;
        RECT 1279.730 186.565 1476.270 191.015 ;
      LAYER met5 ;
        RECT 1477.870 184.965 1552.130 197.865 ;
      LAYER met5 ;
        RECT 1553.730 192.615 1750.270 197.865 ;
        RECT 1592.000 191.015 1712.000 192.615 ;
        RECT 1553.730 186.565 1750.270 191.015 ;
      LAYER met5 ;
        RECT 1751.870 184.965 1826.130 197.865 ;
      LAYER met5 ;
        RECT 1827.730 192.615 2024.270 197.865 ;
        RECT 1866.000 191.015 1986.000 192.615 ;
        RECT 1827.730 186.565 2024.270 191.015 ;
      LAYER met5 ;
        RECT 2025.870 184.965 2100.130 197.865 ;
      LAYER met5 ;
        RECT 2101.730 192.615 2298.270 197.865 ;
        RECT 2140.000 191.015 2260.000 192.615 ;
        RECT 2101.730 186.565 2298.270 191.015 ;
      LAYER met5 ;
        RECT 2299.870 184.965 2374.130 197.865 ;
      LAYER met5 ;
        RECT 2375.730 192.615 2572.270 197.865 ;
        RECT 2414.000 191.015 2534.000 192.615 ;
        RECT 2375.730 186.565 2572.270 191.015 ;
      LAYER met5 ;
        RECT 2573.870 184.965 2648.130 197.865 ;
      LAYER met5 ;
        RECT 2649.730 192.615 2846.270 197.865 ;
        RECT 2688.000 191.015 2808.000 192.615 ;
        RECT 2649.730 186.565 2846.270 191.015 ;
      LAYER met5 ;
        RECT 2847.870 184.965 2917.130 197.865 ;
      LAYER met5 ;
        RECT 2918.730 192.615 3115.270 197.865 ;
        RECT 2957.000 191.015 3077.000 192.615 ;
        RECT 2918.730 186.565 3115.270 191.015 ;
      LAYER met5 ;
        RECT 3116.870 184.965 3186.130 197.865 ;
      LAYER met5 ;
        RECT 3187.730 192.615 3385.270 197.865 ;
      LAYER met5 ;
        RECT 3386.870 196.050 3388.535 197.865 ;
      LAYER met5 ;
        RECT 3390.135 197.650 3395.385 501.270 ;
        RECT 3396.985 355.000 3401.435 501.270 ;
        RECT 3403.035 350.000 3406.285 501.030 ;
        RECT 3396.985 196.215 3401.435 350.000 ;
        RECT 3403.035 198.530 3406.285 345.000 ;
        RECT 3407.885 198.475 3412.335 501.270 ;
        RECT 3413.935 198.400 3418.385 501.270 ;
        RECT 3419.985 198.615 3423.235 501.270 ;
        RECT 3424.840 500.000 3428.085 501.270 ;
        RECT 3424.835 350.000 3428.085 500.000 ;
        RECT 3429.685 355.000 3434.135 501.270 ;
        RECT 3435.735 350.000 3444.735 501.270 ;
        RECT 3424.835 198.665 3428.085 345.000 ;
        RECT 3429.685 198.525 3434.135 350.000 ;
      LAYER met5 ;
        RECT 3424.835 197.015 3428.085 197.065 ;
        RECT 3403.035 196.875 3406.285 196.930 ;
        RECT 3419.985 196.925 3428.085 197.015 ;
        RECT 3403.035 196.800 3412.335 196.875 ;
        RECT 3419.985 196.800 3434.135 196.925 ;
        RECT 3386.870 194.615 3395.385 196.050 ;
        RECT 3403.035 194.615 3434.135 196.800 ;
      LAYER met5 ;
        RECT 3226.000 191.015 3346.000 192.615 ;
        RECT 3187.730 186.565 3385.270 191.015 ;
      LAYER met5 ;
        RECT 3386.870 184.965 3434.135 194.615 ;
        RECT 153.865 181.715 196.930 184.965 ;
      LAYER met5 ;
        RECT 198.530 181.715 394.965 184.965 ;
      LAYER met5 ;
        RECT 396.565 181.715 466.435 184.965 ;
      LAYER met5 ;
        RECT 468.035 181.715 663.965 184.965 ;
      LAYER met5 ;
        RECT 665.565 181.715 735.435 184.965 ;
      LAYER met5 ;
        RECT 737.035 181.715 933.030 184.965 ;
      LAYER met5 ;
        RECT 934.630 181.715 1009.435 184.965 ;
      LAYER met5 ;
        RECT 1011.035 181.715 1206.965 184.965 ;
      LAYER met5 ;
        RECT 1208.565 181.715 1278.435 184.965 ;
      LAYER met5 ;
        RECT 1280.035 181.715 1476.030 184.965 ;
      LAYER met5 ;
        RECT 1477.630 181.715 1552.435 184.965 ;
      LAYER met5 ;
        RECT 1554.035 181.715 1750.030 184.965 ;
      LAYER met5 ;
        RECT 1751.630 181.715 1826.435 184.965 ;
      LAYER met5 ;
        RECT 1828.035 181.715 2024.030 184.965 ;
      LAYER met5 ;
        RECT 2025.630 181.715 2100.435 184.965 ;
      LAYER met5 ;
        RECT 2102.035 181.715 2298.030 184.965 ;
      LAYER met5 ;
        RECT 2299.630 181.715 2374.435 184.965 ;
      LAYER met5 ;
        RECT 2376.035 181.715 2572.030 184.965 ;
      LAYER met5 ;
        RECT 2573.630 181.715 2648.435 184.965 ;
      LAYER met5 ;
        RECT 2650.035 181.715 2845.965 184.965 ;
      LAYER met5 ;
        RECT 2847.565 181.715 2917.435 184.965 ;
        RECT 3116.565 181.715 3186.435 184.965 ;
        RECT 3386.855 181.715 3434.135 184.965 ;
        RECT 153.865 175.665 196.875 181.715 ;
      LAYER met5 ;
        RECT 198.475 175.665 395.270 180.115 ;
      LAYER met5 ;
        RECT 153.865 175.245 196.800 175.665 ;
        RECT 0.000 168.015 196.800 175.245 ;
      LAYER met5 ;
        RECT 198.400 169.615 395.270 174.065 ;
      LAYER met5 ;
        RECT 0.000 163.165 197.015 168.015 ;
      LAYER met5 ;
        RECT 198.615 164.765 395.270 168.015 ;
      LAYER met5 ;
        RECT 396.870 163.165 466.130 181.715 ;
      LAYER met5 ;
        RECT 467.730 175.665 664.270 180.115 ;
        RECT 467.730 169.615 664.270 174.065 ;
        RECT 467.730 164.765 664.270 168.015 ;
      LAYER met5 ;
        RECT 0.000 159.915 197.065 163.165 ;
        RECT 394.000 163.160 469.000 163.165 ;
        RECT 0.000 153.865 196.925 159.915 ;
      LAYER met5 ;
        RECT 198.525 153.865 395.270 158.315 ;
      LAYER met5 ;
        RECT 0.000 141.665 175.245 153.865 ;
        RECT 0.000 135.815 196.775 141.665 ;
      LAYER met5 ;
        RECT 198.375 137.415 395.270 141.665 ;
      LAYER met5 ;
        RECT 0.000 131.565 196.920 135.815 ;
      LAYER met5 ;
        RECT 198.520 131.565 395.270 135.815 ;
      LAYER met5 ;
        RECT 0.000 103.415 195.755 131.565 ;
      LAYER met5 ;
        RECT 197.355 105.015 201.000 129.965 ;
      LAYER met5 ;
        RECT 202.600 105.015 217.400 129.965 ;
      LAYER met5 ;
        RECT 219.000 105.015 221.000 129.965 ;
      LAYER met5 ;
        RECT 222.600 105.015 227.400 129.965 ;
      LAYER met5 ;
        RECT 229.000 105.015 231.000 129.965 ;
        RECT 234.000 105.015 358.000 129.965 ;
      LAYER met5 ;
        RECT 359.600 105.015 374.400 129.965 ;
      LAYER met5 ;
        RECT 376.000 105.015 378.000 129.965 ;
      LAYER met5 ;
        RECT 379.600 105.015 384.400 129.965 ;
      LAYER met5 ;
        RECT 386.000 105.015 388.000 129.965 ;
        RECT 391.000 105.015 395.270 129.965 ;
      LAYER met5 ;
        RECT 396.870 103.415 466.130 163.160 ;
      LAYER met5 ;
        RECT 467.730 153.865 664.270 158.315 ;
        RECT 467.730 137.415 664.270 141.665 ;
        RECT 467.730 131.565 664.270 135.815 ;
        RECT 467.730 105.015 470.000 129.965 ;
      LAYER met5 ;
        RECT 471.600 105.015 486.400 129.965 ;
      LAYER met5 ;
        RECT 488.000 105.015 490.000 129.965 ;
      LAYER met5 ;
        RECT 491.600 105.015 496.400 129.965 ;
      LAYER met5 ;
        RECT 498.000 105.015 500.000 129.965 ;
        RECT 503.000 105.015 627.000 129.965 ;
      LAYER met5 ;
        RECT 628.600 105.015 643.400 129.965 ;
      LAYER met5 ;
        RECT 645.000 105.015 647.000 129.965 ;
      LAYER met5 ;
        RECT 648.600 105.015 653.400 129.965 ;
      LAYER met5 ;
        RECT 655.000 105.015 657.000 129.965 ;
        RECT 660.000 105.015 664.270 129.965 ;
      LAYER met5 ;
        RECT 665.870 103.415 735.130 181.715 ;
      LAYER met5 ;
        RECT 736.730 175.665 933.270 180.115 ;
        RECT 736.730 169.615 933.270 174.065 ;
        RECT 736.730 164.765 933.270 168.015 ;
        RECT 738.000 163.160 932.000 163.165 ;
        RECT 736.730 159.915 933.270 163.160 ;
        RECT 736.730 153.865 933.270 158.315 ;
        RECT 736.730 143.265 933.270 152.265 ;
        RECT 736.730 137.415 933.270 141.665 ;
        RECT 736.730 131.565 933.270 135.815 ;
        RECT 736.730 105.015 739.000 129.965 ;
      LAYER met5 ;
        RECT 740.600 105.015 755.400 129.965 ;
      LAYER met5 ;
        RECT 757.000 105.015 759.000 129.965 ;
      LAYER met5 ;
        RECT 760.600 105.015 765.400 129.965 ;
      LAYER met5 ;
        RECT 767.000 105.015 769.000 129.965 ;
        RECT 772.000 105.015 896.000 129.965 ;
      LAYER met5 ;
        RECT 897.600 105.015 912.400 129.965 ;
      LAYER met5 ;
        RECT 914.000 105.015 916.000 129.965 ;
      LAYER met5 ;
        RECT 917.600 105.015 922.400 129.965 ;
      LAYER met5 ;
        RECT 924.000 105.015 926.000 129.965 ;
        RECT 929.000 105.015 933.270 129.965 ;
      LAYER met5 ;
        RECT 934.870 103.415 1009.130 181.715 ;
      LAYER met5 ;
        RECT 1010.730 175.665 1207.270 180.115 ;
        RECT 1010.730 169.615 1207.270 174.065 ;
        RECT 1010.730 164.765 1207.270 168.015 ;
        RECT 1012.000 163.160 1206.000 163.165 ;
        RECT 1010.730 159.915 1207.270 163.160 ;
        RECT 1010.730 143.265 1207.270 152.265 ;
        RECT 1010.730 137.415 1207.270 141.665 ;
        RECT 1010.730 131.565 1207.270 135.815 ;
        RECT 1010.730 105.015 1013.000 129.965 ;
      LAYER met5 ;
        RECT 1014.600 105.015 1029.400 129.965 ;
      LAYER met5 ;
        RECT 1031.000 105.015 1033.000 129.965 ;
      LAYER met5 ;
        RECT 1034.600 105.015 1039.400 129.965 ;
      LAYER met5 ;
        RECT 1041.000 105.015 1043.000 129.965 ;
        RECT 1046.000 105.015 1170.000 129.965 ;
      LAYER met5 ;
        RECT 1171.600 105.015 1186.400 129.965 ;
      LAYER met5 ;
        RECT 1188.000 105.015 1190.000 129.965 ;
      LAYER met5 ;
        RECT 1191.600 105.015 1196.400 129.965 ;
      LAYER met5 ;
        RECT 1198.000 105.015 1200.000 129.965 ;
        RECT 1203.000 105.015 1207.270 129.965 ;
      LAYER met5 ;
        RECT 1208.870 103.415 1278.130 181.715 ;
      LAYER met5 ;
        RECT 1279.730 175.665 1476.270 180.115 ;
        RECT 1279.730 169.615 1476.270 174.065 ;
        RECT 1279.730 164.765 1476.270 168.015 ;
        RECT 1281.000 163.160 1475.000 163.165 ;
        RECT 1279.730 159.915 1476.270 163.160 ;
        RECT 1279.730 143.265 1476.270 152.265 ;
        RECT 1279.730 137.415 1476.270 141.665 ;
        RECT 1279.730 131.565 1476.270 135.815 ;
        RECT 1279.730 105.015 1282.000 129.965 ;
      LAYER met5 ;
        RECT 1283.600 105.015 1298.400 129.965 ;
      LAYER met5 ;
        RECT 1300.000 105.015 1302.000 129.965 ;
      LAYER met5 ;
        RECT 1303.600 105.015 1308.400 129.965 ;
      LAYER met5 ;
        RECT 1310.000 105.015 1312.000 129.965 ;
        RECT 1315.000 105.015 1439.000 129.965 ;
      LAYER met5 ;
        RECT 1440.600 105.015 1455.400 129.965 ;
      LAYER met5 ;
        RECT 1457.000 105.015 1459.000 129.965 ;
      LAYER met5 ;
        RECT 1460.600 105.015 1465.400 129.965 ;
      LAYER met5 ;
        RECT 1467.000 105.015 1469.000 129.965 ;
        RECT 1472.000 105.015 1476.270 129.965 ;
      LAYER met5 ;
        RECT 1477.870 103.415 1552.130 181.715 ;
      LAYER met5 ;
        RECT 1553.730 175.665 1750.270 180.115 ;
        RECT 1553.730 169.615 1750.270 174.065 ;
        RECT 1553.730 164.765 1750.270 168.015 ;
        RECT 1555.000 163.160 1749.000 163.165 ;
        RECT 1553.730 159.915 1750.270 163.160 ;
        RECT 1553.730 153.865 1750.270 158.315 ;
        RECT 1553.730 143.265 1750.270 152.265 ;
        RECT 1553.730 137.415 1750.270 141.665 ;
        RECT 1553.730 131.565 1750.270 135.815 ;
        RECT 1553.730 105.015 1556.000 129.965 ;
      LAYER met5 ;
        RECT 1557.600 105.015 1572.400 129.965 ;
      LAYER met5 ;
        RECT 1574.000 105.015 1576.000 129.965 ;
      LAYER met5 ;
        RECT 1577.600 105.015 1582.400 129.965 ;
      LAYER met5 ;
        RECT 1584.000 105.015 1586.000 129.965 ;
        RECT 1589.000 105.015 1713.000 129.965 ;
      LAYER met5 ;
        RECT 1714.600 105.015 1729.400 129.965 ;
      LAYER met5 ;
        RECT 1731.000 105.015 1733.000 129.965 ;
      LAYER met5 ;
        RECT 1734.600 105.015 1739.400 129.965 ;
      LAYER met5 ;
        RECT 1741.000 105.015 1743.000 129.965 ;
        RECT 1746.000 105.015 1750.270 129.965 ;
      LAYER met5 ;
        RECT 1751.870 103.415 1826.130 181.715 ;
      LAYER met5 ;
        RECT 1827.730 175.665 2024.270 180.115 ;
        RECT 1827.730 169.615 2024.270 174.065 ;
        RECT 1827.730 164.765 2024.270 168.015 ;
        RECT 1829.000 163.160 2023.000 163.165 ;
        RECT 1827.730 159.915 2024.270 163.160 ;
        RECT 1827.730 153.865 2024.270 158.315 ;
        RECT 1827.730 143.265 2024.270 152.265 ;
        RECT 1827.730 137.415 2024.270 141.665 ;
        RECT 1827.730 131.565 2024.270 135.815 ;
        RECT 1827.730 105.015 1830.000 129.965 ;
      LAYER met5 ;
        RECT 1831.600 105.015 1846.400 129.965 ;
      LAYER met5 ;
        RECT 1848.000 105.015 1850.000 129.965 ;
      LAYER met5 ;
        RECT 1851.600 105.015 1856.400 129.965 ;
      LAYER met5 ;
        RECT 1858.000 105.015 1860.000 129.965 ;
        RECT 1863.000 105.015 1987.000 129.965 ;
      LAYER met5 ;
        RECT 1988.600 105.015 2003.400 129.965 ;
      LAYER met5 ;
        RECT 2005.000 105.015 2007.000 129.965 ;
      LAYER met5 ;
        RECT 2008.600 105.015 2013.400 129.965 ;
      LAYER met5 ;
        RECT 2015.000 105.015 2017.000 129.965 ;
        RECT 2020.000 105.015 2024.270 129.965 ;
      LAYER met5 ;
        RECT 2025.870 103.415 2100.130 181.715 ;
      LAYER met5 ;
        RECT 2101.730 175.665 2298.270 180.115 ;
        RECT 2101.730 169.615 2298.270 174.065 ;
        RECT 2101.730 164.765 2298.270 168.015 ;
        RECT 2103.000 163.160 2297.000 163.165 ;
        RECT 2101.730 159.915 2298.270 163.160 ;
        RECT 2101.730 153.865 2298.270 158.315 ;
        RECT 2101.730 143.265 2298.270 152.265 ;
        RECT 2101.730 137.415 2298.270 141.665 ;
        RECT 2101.730 131.565 2298.270 135.815 ;
        RECT 2101.730 105.015 2104.000 129.965 ;
      LAYER met5 ;
        RECT 2105.600 105.015 2120.400 129.965 ;
      LAYER met5 ;
        RECT 2122.000 105.015 2124.000 129.965 ;
      LAYER met5 ;
        RECT 2125.600 105.015 2130.400 129.965 ;
      LAYER met5 ;
        RECT 2132.000 105.015 2134.000 129.965 ;
        RECT 2137.000 105.015 2261.000 129.965 ;
      LAYER met5 ;
        RECT 2262.600 105.015 2277.400 129.965 ;
      LAYER met5 ;
        RECT 2279.000 105.015 2281.000 129.965 ;
      LAYER met5 ;
        RECT 2282.600 105.015 2287.400 129.965 ;
      LAYER met5 ;
        RECT 2289.000 105.015 2291.000 129.965 ;
        RECT 2294.000 105.015 2298.270 129.965 ;
      LAYER met5 ;
        RECT 2299.870 103.415 2374.130 181.715 ;
      LAYER met5 ;
        RECT 2375.730 175.665 2572.270 180.115 ;
        RECT 2375.730 169.615 2572.270 174.065 ;
        RECT 2375.730 164.765 2572.270 168.015 ;
        RECT 2377.000 163.160 2571.000 163.165 ;
        RECT 2375.730 159.915 2572.270 163.160 ;
        RECT 2375.730 153.865 2572.270 158.315 ;
        RECT 2375.730 143.265 2572.270 152.265 ;
        RECT 2375.730 137.415 2572.270 141.665 ;
        RECT 2375.730 131.565 2572.270 135.815 ;
        RECT 2375.730 105.015 2378.000 129.965 ;
      LAYER met5 ;
        RECT 2379.600 105.015 2394.400 129.965 ;
      LAYER met5 ;
        RECT 2396.000 105.015 2398.000 129.965 ;
      LAYER met5 ;
        RECT 2399.600 105.015 2404.400 129.965 ;
      LAYER met5 ;
        RECT 2406.000 105.015 2408.000 129.965 ;
        RECT 2411.000 105.015 2535.000 129.965 ;
      LAYER met5 ;
        RECT 2536.600 105.015 2551.400 129.965 ;
      LAYER met5 ;
        RECT 2553.000 105.015 2555.000 129.965 ;
      LAYER met5 ;
        RECT 2556.600 105.015 2561.400 129.965 ;
      LAYER met5 ;
        RECT 2563.000 105.015 2565.000 129.965 ;
        RECT 2568.000 105.015 2572.270 129.965 ;
      LAYER met5 ;
        RECT 2573.870 103.415 2648.130 181.715 ;
      LAYER met5 ;
        RECT 2649.730 175.665 2846.270 180.115 ;
        RECT 2649.730 169.615 2846.270 174.065 ;
        RECT 2649.730 164.765 2846.270 168.015 ;
      LAYER met5 ;
        RECT 2847.870 163.165 2917.130 181.715 ;
      LAYER met5 ;
        RECT 2918.730 175.665 3115.270 180.115 ;
        RECT 2918.730 169.615 3115.270 174.065 ;
        RECT 2918.730 164.765 3115.270 168.015 ;
      LAYER met5 ;
        RECT 3116.870 163.165 3186.130 181.715 ;
      LAYER met5 ;
        RECT 3187.730 175.665 3385.270 180.115 ;
      LAYER met5 ;
        RECT 3386.870 175.245 3434.135 181.715 ;
      LAYER met5 ;
        RECT 3435.735 176.845 3444.735 345.000 ;
        RECT 3446.335 198.375 3450.585 501.270 ;
        RECT 3452.185 198.520 3456.435 501.270 ;
        RECT 3458.035 499.000 3482.985 501.270 ;
      LAYER met5 ;
        RECT 3484.585 500.000 3588.000 502.870 ;
      LAYER met5 ;
        RECT 3458.035 494.000 3482.985 496.000 ;
      LAYER met5 ;
        RECT 3458.035 477.600 3482.985 492.400 ;
      LAYER met5 ;
        RECT 3458.035 474.000 3482.985 476.000 ;
      LAYER met5 ;
        RECT 3458.035 457.600 3482.985 472.400 ;
      LAYER met5 ;
        RECT 3458.035 454.000 3482.985 456.000 ;
      LAYER met5 ;
        RECT 3458.035 437.600 3482.985 452.400 ;
      LAYER met5 ;
        RECT 3458.035 434.000 3482.985 436.000 ;
      LAYER met5 ;
        RECT 3458.035 417.600 3482.985 432.400 ;
      LAYER met5 ;
        RECT 3458.035 414.000 3482.985 416.000 ;
      LAYER met5 ;
        RECT 3458.035 397.600 3482.985 412.400 ;
      LAYER met5 ;
        RECT 3458.035 394.000 3482.985 396.000 ;
      LAYER met5 ;
        RECT 3458.035 377.600 3482.985 392.400 ;
      LAYER met5 ;
        RECT 3458.035 374.000 3482.985 376.000 ;
      LAYER met5 ;
        RECT 3458.035 357.600 3482.985 372.400 ;
      LAYER met5 ;
        RECT 3458.035 344.000 3482.985 356.000 ;
        RECT 3458.035 339.000 3482.985 341.000 ;
      LAYER met5 ;
        RECT 3458.035 322.600 3482.985 337.400 ;
      LAYER met5 ;
        RECT 3458.035 319.000 3482.985 321.000 ;
      LAYER met5 ;
        RECT 3458.035 302.600 3482.985 317.400 ;
      LAYER met5 ;
        RECT 3458.035 299.000 3482.985 301.000 ;
      LAYER met5 ;
        RECT 3458.035 282.600 3482.985 297.400 ;
      LAYER met5 ;
        RECT 3458.035 279.000 3482.985 281.000 ;
      LAYER met5 ;
        RECT 3458.035 262.600 3482.985 277.400 ;
      LAYER met5 ;
        RECT 3458.035 259.000 3482.985 261.000 ;
      LAYER met5 ;
        RECT 3458.035 242.600 3482.985 257.400 ;
      LAYER met5 ;
        RECT 3458.035 239.000 3482.985 241.000 ;
      LAYER met5 ;
        RECT 3458.035 222.600 3482.985 237.400 ;
      LAYER met5 ;
        RECT 3458.035 219.000 3482.985 221.000 ;
      LAYER met5 ;
        RECT 3458.035 202.600 3482.985 217.400 ;
      LAYER met5 ;
        RECT 3458.035 197.355 3482.985 201.000 ;
        RECT 3563.785 200.000 3588.000 500.000 ;
      LAYER met5 ;
        RECT 3452.185 196.775 3456.435 196.920 ;
        RECT 3446.335 195.755 3456.435 196.775 ;
        RECT 3484.585 195.755 3588.000 200.000 ;
        RECT 3446.335 175.245 3588.000 195.755 ;
      LAYER met5 ;
        RECT 3187.730 169.615 3385.270 174.065 ;
        RECT 3187.730 164.765 3385.270 168.015 ;
        RECT 2651.000 163.160 2845.000 163.165 ;
      LAYER met5 ;
        RECT 2845.000 163.160 2920.000 163.165 ;
      LAYER met5 ;
        RECT 2920.000 163.160 3114.000 163.165 ;
      LAYER met5 ;
        RECT 3114.000 163.160 3189.000 163.165 ;
      LAYER met5 ;
        RECT 3189.000 163.160 3384.000 163.165 ;
        RECT 2649.730 159.915 2846.270 163.160 ;
        RECT 2649.730 153.865 2846.270 158.315 ;
        RECT 2649.730 143.265 2846.270 152.265 ;
        RECT 2649.730 137.415 2846.270 141.665 ;
        RECT 2649.730 131.565 2846.270 135.815 ;
        RECT 2649.730 105.015 2652.000 129.965 ;
      LAYER met5 ;
        RECT 2653.600 105.015 2668.400 129.965 ;
      LAYER met5 ;
        RECT 2670.000 105.015 2672.000 129.965 ;
      LAYER met5 ;
        RECT 2673.600 105.015 2678.400 129.965 ;
      LAYER met5 ;
        RECT 2680.000 105.015 2682.000 129.965 ;
        RECT 2685.000 105.015 2809.000 129.965 ;
      LAYER met5 ;
        RECT 2810.600 105.015 2825.400 129.965 ;
      LAYER met5 ;
        RECT 2827.000 105.015 2829.000 129.965 ;
      LAYER met5 ;
        RECT 2830.600 105.015 2835.400 129.965 ;
      LAYER met5 ;
        RECT 2837.000 105.015 2839.000 129.965 ;
        RECT 2842.000 105.015 2846.270 129.965 ;
      LAYER met5 ;
        RECT 2847.870 103.415 2917.130 163.160 ;
      LAYER met5 ;
        RECT 2918.730 159.915 3115.270 163.160 ;
        RECT 2918.730 153.865 3115.270 158.315 ;
        RECT 2918.730 143.265 3115.270 152.265 ;
        RECT 2918.730 137.415 3115.270 141.665 ;
        RECT 2918.730 131.565 3115.270 135.815 ;
        RECT 2918.730 105.015 2921.000 129.965 ;
      LAYER met5 ;
        RECT 2922.600 105.015 2937.400 129.965 ;
      LAYER met5 ;
        RECT 2939.000 105.015 2941.000 129.965 ;
      LAYER met5 ;
        RECT 2942.600 105.015 2947.400 129.965 ;
      LAYER met5 ;
        RECT 2949.000 105.015 2951.000 129.965 ;
        RECT 2954.000 105.015 3078.000 129.965 ;
      LAYER met5 ;
        RECT 3079.600 105.015 3094.400 129.965 ;
      LAYER met5 ;
        RECT 3096.000 105.015 3098.000 129.965 ;
      LAYER met5 ;
        RECT 3099.600 105.015 3104.400 129.965 ;
      LAYER met5 ;
        RECT 3106.000 105.015 3108.000 129.965 ;
        RECT 3111.000 105.015 3115.270 129.965 ;
      LAYER met5 ;
        RECT 3116.870 103.415 3186.130 163.160 ;
      LAYER met5 ;
        RECT 3187.730 159.915 3385.270 163.160 ;
        RECT 3187.730 153.865 3385.270 158.315 ;
      LAYER met5 ;
        RECT 3386.870 153.865 3588.000 175.245 ;
      LAYER met5 ;
        RECT 3187.730 143.265 3411.155 152.265 ;
      LAYER met5 ;
        RECT 3412.755 141.665 3588.000 153.865 ;
      LAYER met5 ;
        RECT 3187.730 137.415 3385.270 141.665 ;
        RECT 3187.730 131.565 3385.270 135.815 ;
      LAYER met5 ;
        RECT 3386.870 131.565 3588.000 141.665 ;
      LAYER met5 ;
        RECT 3187.730 105.015 3190.000 129.965 ;
      LAYER met5 ;
        RECT 3191.600 105.015 3206.400 129.965 ;
      LAYER met5 ;
        RECT 3208.000 105.015 3210.000 129.965 ;
      LAYER met5 ;
        RECT 3211.600 105.015 3216.400 129.965 ;
      LAYER met5 ;
        RECT 3218.000 105.015 3220.000 129.965 ;
        RECT 3223.000 105.015 3347.000 129.965 ;
      LAYER met5 ;
        RECT 3348.600 105.015 3363.400 129.965 ;
      LAYER met5 ;
        RECT 3365.000 105.015 3367.000 129.965 ;
      LAYER met5 ;
        RECT 3368.600 105.015 3373.400 129.965 ;
      LAYER met5 ;
        RECT 3375.000 105.015 3377.000 129.965 ;
        RECT 3380.000 105.015 3385.855 129.965 ;
      LAYER met5 ;
        RECT 3387.455 103.415 3588.000 131.565 ;
        RECT 0.000 0.000 200.000 103.415 ;
        RECT 394.000 96.480 469.000 103.415 ;
        RECT 394.000 32.455 399.510 96.480 ;
        RECT 463.550 32.455 469.000 96.480 ;
      LAYER met5 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met5 ;
        RECT 394.000 0.000 469.000 32.455 ;
        RECT 663.000 93.145 738.000 103.415 ;
        RECT 663.000 34.115 681.965 93.145 ;
        RECT 722.350 34.115 738.000 93.145 ;
        RECT 663.000 25.815 738.000 34.115 ;
        RECT 932.000 97.040 1012.000 103.415 ;
        RECT 932.000 31.390 936.600 97.040 ;
        RECT 1002.400 31.390 1012.000 97.040 ;
      LAYER met5 ;
        RECT 469.000 0.000 664.270 24.215 ;
      LAYER met5 ;
        RECT 665.870 0.000 735.130 25.815 ;
      LAYER met5 ;
        RECT 736.730 0.000 932.000 24.215 ;
      LAYER met5 ;
        RECT 932.000 0.000 1012.000 31.390 ;
        RECT 1206.000 99.700 1281.000 103.415 ;
        RECT 1206.000 29.235 1214.730 99.700 ;
        RECT 1272.330 29.235 1281.000 99.700 ;
      LAYER met5 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met5 ;
        RECT 1206.000 0.000 1281.000 29.235 ;
        RECT 1475.000 97.040 1555.000 103.415 ;
        RECT 1475.000 31.390 1479.600 97.040 ;
        RECT 1545.400 31.390 1555.000 97.040 ;
      LAYER met5 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met5 ;
        RECT 1475.000 0.000 1555.000 31.390 ;
        RECT 1749.000 97.040 1829.000 103.415 ;
        RECT 1749.000 31.390 1753.600 97.040 ;
        RECT 1819.400 31.390 1829.000 97.040 ;
      LAYER met5 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met5 ;
        RECT 1749.000 0.000 1829.000 31.390 ;
        RECT 2023.000 97.040 2103.000 103.415 ;
        RECT 2023.000 31.390 2027.600 97.040 ;
        RECT 2093.400 31.390 2103.000 97.040 ;
      LAYER met5 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met5 ;
        RECT 2023.000 0.000 2103.000 31.390 ;
        RECT 2297.000 97.040 2377.000 103.415 ;
        RECT 2297.000 31.390 2301.600 97.040 ;
        RECT 2367.400 31.390 2377.000 97.040 ;
      LAYER met5 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met5 ;
        RECT 2297.000 0.000 2377.000 31.390 ;
        RECT 2571.000 97.040 2651.000 103.415 ;
        RECT 2571.000 31.390 2575.600 97.040 ;
        RECT 2641.400 31.390 2651.000 97.040 ;
      LAYER met5 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met5 ;
        RECT 2571.000 0.000 2651.000 31.390 ;
        RECT 2845.000 96.480 2920.000 103.415 ;
        RECT 2845.000 32.455 2850.510 96.480 ;
        RECT 2914.550 32.455 2920.000 96.480 ;
      LAYER met5 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met5 ;
        RECT 2845.000 0.000 2920.000 32.455 ;
        RECT 3114.000 96.480 3189.000 103.415 ;
        RECT 3114.000 32.455 3119.510 96.480 ;
        RECT 3183.550 32.455 3189.000 96.480 ;
      LAYER met5 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met5 ;
        RECT 3114.000 0.000 3189.000 32.455 ;
      LAYER met5 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met5 ;
        RECT 3384.000 0.000 3588.000 103.415 ;
  END
END chip_io
END LIBRARY

