* NGSPICE file created from sky130_fd_io__top_gpiov2.ext - technology: sky130A

.subckt sky130_fd_io__hvsbt_inv_x1 OUT VPWR VGND VSUBS a_119_118# w_n46_415#
X0 OUT a_119_118# VPWR w_n46_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 OUT a_119_118# VPWR w_n46_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 OUT a_119_118# VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__hvsbt_xor VPWR VGND IN0 IN1 OUT VSUBS w_95_503#
X0 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 a_862_167# a_566_375# OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X2 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X4 VGND a_161_167# a_862_167# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X5 a_510_167# IN0 VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X6 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X7 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X8 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X9 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X10 VGND IN0 a_161_167# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X11 OUT IN1 a_510_167# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X12 a_566_375# IN1 VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X13 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X14 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X15 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X16 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X17 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
.ends

.subckt sky130_fd_io__hvsbt_nor IN0 VSUBS a_66_482# a_66_144# w_0_415# a_295_118#
+ a_239_144#
X0 a_239_482# IN0 a_66_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 a_239_144# a_295_118# a_239_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 a_239_482# IN0 a_66_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 a_66_144# a_295_118# a_239_144# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X4 a_239_144# a_295_118# a_239_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X5 a_239_144# IN0 a_66_144# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__hvsbt_inv_x2 VPWR VGND IN OUT VSUBS w_0_415#
X0 OUT IN VPWR w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 VPWR IN OUT w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 OUT IN VPWR w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X4 VPWR IN OUT w_0_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X5 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__com_ctl_ls_octl VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H HLD_H_N
+ VSUBS a_181_1305# a_992_934# w_n17_1379#
X0 a_957_1391# a_181_1305# a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X1 VSUBS RST_H a_65_861# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X2 a_634_829# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X3 OUT_H a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X4 a_128_1391# a_181_1305# a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X5 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X6 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X7 a_361_1391# HLD_H_N a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X8 a_634_829# a_992_934# a_181_1305# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_724_1391# a_181_1305# a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X10 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X12 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X13 VSUBS IN a_992_934# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X14 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X15 a_181_1305# IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X17 VSUBS a_65_861# a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X18 a_361_1391# a_181_1305# a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X19 VSUBS a_65_861# OUT_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X20 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X21 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X22 a_957_1391# a_181_1305# a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X23 a_65_861# HLD_H_N a_957_1391# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X24 a_361_1391# a_181_1305# a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X25 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X26 a_724_1391# a_181_1305# a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X27 a_130_181# SET_H VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X28 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X29 a_128_1391# a_181_1305# a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X30 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X31 a_65_861# a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
.ends

.subckt sky130_fd_io__hvsbt_nand2 IN1 IN0 OUT VGND VPWR VSUBS w_n42_415#
X0 OUT IN0 VPWR w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 VPWR IN1 OUT w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 OUT IN0 VPWR w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 OUT IN1 a_239_144# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X4 VPWR IN1 OUT w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X5 a_239_144# IN0 VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__hvsbt_xorv2 VPWR VGND IN0 IN1 OUT VSUBS a_742_141# a_566_375#
+ w_95_503#
X0 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 a_862_167# a_742_141# OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X2 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X4 VGND a_161_167# a_862_167# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X5 a_510_167# IN0 VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X6 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X7 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X8 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X9 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X10 VGND IN0 a_161_167# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X11 OUT IN1 a_510_167# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X12 a_566_375# IN1 VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X13 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X14 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X15 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X16 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X17 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_octl DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2] PUEN_2OR1_H
+ DM_H[1] PDEN_H_N[1] PDEN_H_N[0] OD_H SLOW SLOW_H SLOW_H_N HLD_I_H_N VCC_IO VGND
+ VPWR sky130_fd_io__hvsbt_nand2_0/OUT sky130_fd_io__hvsbt_nand2_4/IN1 sky130_fd_io__hvsbt_xorv2_0/a_566_375#
+ m1_n8856_3102# sky130_fd_io__hvsbt_nor_0/IN0 sky130_fd_io__hvsbt_nand2_0/IN0 sky130_fd_io__hvsbt_inv_x2_3/OUT
+ li_n9202_2336# sky130_fd_io__hvsbt_inv_x2_2/OUT sky130_fd_io__hvsbt_nand2_0/VGND
+ sky130_fd_io__hvsbt_nor_0/w_0_415# sky130_fd_io__hvsbt_nand2_0/VPWR sky130_fd_io__hvsbt_xorv2_0/a_742_141#
+
Xsky130_fd_io__hvsbt_inv_x1_4 sky130_fd_io__hvsbt_inv_x2_2/IN VCC_IO VGND VGND li_5323_4140#
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_xor_0 VCC_IO VGND DM_H[2] DM_H[1] sky130_fd_io__hvsbt_xor_0/OUT
+ VGND VCC_IO sky130_fd_io__hvsbt_xor
Xsky130_fd_io__hvsbt_nor_0 sky130_fd_io__hvsbt_nor_0/IN0 VGND sky130_fd_io__hvsbt_nand2_0/VPWR
+ sky130_fd_io__hvsbt_nand2_0/VGND sky130_fd_io__hvsbt_nor_0/w_0_415# li_n9202_2336#
+ sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_inv_x2_0 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_0/IN PDEN_H_N[0]
+ VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_nor_1 DM_H_N[2] VGND VCC_IO VGND VCC_IO DM_H_N[1] sky130_fd_io__hvsbt_nand2_3/IN0
+ sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_inv_x2_1 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_1/IN PDEN_H_N[1]
+ VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__com_ctl_ls_octl_0 VCC_IO VPWR SLOW_H_N SLOW_H SLOW OD_H VGND HLD_I_H_N
+ VGND VPWR m2_5755_2254# VGND sky130_fd_io__com_ctl_ls_octl
Xsky130_fd_io__hvsbt_nor_2 sky130_fd_io__hvsbt_nor_2/IN0 VGND VCC_IO VGND VCC_IO DM_H_N[1]
+ li_5323_4140# sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__hvsbt_nand2_0/IN0
+ sky130_fd_io__hvsbt_nand2_0/OUT sky130_fd_io__hvsbt_nand2_0/VGND sky130_fd_io__hvsbt_nand2_0/VPWR
+ VGND sky130_fd_io__hvsbt_nor_0/w_0_415# sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_1 sky130_fd_io__hvsbt_nand2_3/OUT sky130_fd_io__hvsbt_nand2_2/OUT
+ PUEN_2OR1_H VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x2_2 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_2/IN sky130_fd_io__hvsbt_inv_x2_2/OUT
+ VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_nand2_2 DM_H[0] sky130_fd_io__hvsbt_xor_0/OUT sky130_fd_io__hvsbt_nand2_2/OUT
+ VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x2_3 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_3/IN sky130_fd_io__hvsbt_inv_x2_3/OUT
+ VGND VCC_IO sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_nand2_3 DM_H_N[0] sky130_fd_io__hvsbt_nand2_3/IN0 sky130_fd_io__hvsbt_nand2_3/OUT
+ VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_4 sky130_fd_io__hvsbt_nand2_4/IN1 PUEN_2OR1_H sky130_fd_io__hvsbt_nand2_4/OUT
+ VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_5 DM_H_N[1] DM_H_N[2] sky130_fd_io__hvsbt_nand2_6/IN1 VGND
+ VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_6 sky130_fd_io__hvsbt_nand2_6/IN1 DM_H_N[0] sky130_fd_io__hvsbt_nand2_6/OUT
+ VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_7 DM_H[0] DM_H[1] sky130_fd_io__hvsbt_nand2_7/OUT VGND
+ VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_xorv2_0 VCC_IO VGND DM_H[2] DM_H[0] sky130_fd_io__hvsbt_nor_2/IN0
+ VGND sky130_fd_io__hvsbt_xorv2_0/a_742_141# sky130_fd_io__hvsbt_xorv2_0/a_566_375#
+ VCC_IO sky130_fd_io__hvsbt_xorv2
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x2_0/IN VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_7/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_inv_x2_3/IN VCC_IO VGND VGND sky130_fd_io__hvsbt_inv_x1_3/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_2 sky130_fd_io__hvsbt_inv_x2_1/IN VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_6/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_3 sky130_fd_io__hvsbt_inv_x1_3/OUT VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_4/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__gpio_dat_ls_1v2 IN OUT_H_N RST_H SET_H HLD_H_N VCC_IO VGND OUT_H
+ VPWR_KA
X0 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X1 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X2 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X4 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X5 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X6 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X7 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt w=3e+06u l=250000u
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X10 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X11 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X12 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X13 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X14 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X15 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X16 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X17 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X18 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X19 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X20 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X21 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X22 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X23 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X24 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X25 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X26 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X27 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt w=3e+06u l=250000u
X28 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X29 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X30 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X31 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X32 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X33 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X34 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X35 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X36 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X37 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X38 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X39 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X40 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X41 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X42 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X43 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X44 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X45 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X46 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X47 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X48 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X49 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
.ends

.subckt sky130_fd_io__gpio_dat_lsv2 IN OUT_H_N RST_H SET_H HLD_H_N VCC_IO VGND OUT_H
+ VPWR_KA a_28_14#
X0 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X1 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X2 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X4 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X5 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X6 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X7 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt w=3e+06u l=250000u
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X10 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X11 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X12 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X13 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X14 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X15 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X16 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X17 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X18 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X19 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X20 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X21 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X22 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X23 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X24 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X25 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X26 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X27 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt w=3e+06u l=250000u
X28 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X29 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X30 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X31 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X32 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X33 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X34 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X35 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X36 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X37 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X38 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X39 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X40 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X41 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X42 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X43 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X44 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X45 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X46 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X47 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X48 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X49 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
.ends

.subckt sky130_fd_io__com_cclat PU_DIS_H PD_DIS_H_uq1 VGND OE_H_N DRVLO_H_N_uq5 DRVHI_H_uq5
+ VCC_IO
X0 DRVLO_H_N_uq5 a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X1 a_4762_1193# DRVHI_H_uq5 a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X2 VCC_IO PU_DIS_H a_638_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X3 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X4 a_2361_1095# DRVHI_H_uq5 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X5 VCC_IO a_638_279# a_947_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X6 DRVHI_H_uq5 a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X7 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X8 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X9 a_987_279# DRVLO_H_N_uq5 a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X10 DRVHI_H_uq5 a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X11 a_2361_1095# a_505_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X12 VGND PD_DIS_H_uq1 a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X13 VCC_IO a_2361_1095# DRVLO_H_N_uq5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X14 VGND OE_H_N a_176_279# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X15 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X16 VGND DRVHI_H_uq5 a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X17 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X18 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X19 VCC_IO a_947_1193# DRVHI_H_uq5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X20 VCC_IO a_947_1193# DRVHI_H_uq5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X21 a_505_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X22 a_2361_1095# PD_DIS_H_uq1 a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X23 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X24 a_1628_279# DRVLO_H_N_uq5 a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X25 VGND a_2361_1095# DRVLO_H_N_uq5 VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X26 VGND a_947_1193# DRVHI_H_uq5 VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X27 DRVLO_H_N_uq5 a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X28 a_947_1193# a_638_279# a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X29 DRVHI_H_uq5 a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X30 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X31 a_3417_1193# DRVHI_H_uq5 a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X32 DRVHI_H_uq5 a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X33 a_947_1193# DRVLO_H_N_uq5 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X34 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X35 DRVLO_H_N_uq5 a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X36 VCC_IO a_947_1193# DRVHI_H_uq5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X37 a_4762_1193# DRVHI_H_uq5 a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X38 a_1628_279# a_638_279# a_947_1193# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X39 VGND a_2361_1095# DRVLO_H_N_uq5 VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X40 VGND a_2361_1095# DRVLO_H_N_uq5 VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X41 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X42 DRVLO_H_N_uq5 a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X43 VGND a_947_1193# DRVHI_H_uq5 VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X44 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X45 VCC_IO a_2361_1095# DRVLO_H_N_uq5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X46 a_2361_1095# PD_DIS_H_uq1 a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X47 a_947_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X48 DRVHI_H_uq5 a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X49 DRVLO_H_N_uq5 a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X50 VCC_IO OE_H_N a_176_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X51 a_4762_1193# PD_DIS_H_uq1 a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X52 a_505_1193# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X53 DRVLO_H_N_uq5 a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X54 a_2361_1095# PD_DIS_H_uq1 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X55 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X56 a_4762_1193# PD_DIS_H_uq1 a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X57 DRVHI_H_uq5 a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X58 VGND a_505_1193# a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X59 VCC_IO a_2361_1095# DRVLO_H_N_uq5 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X60 a_3417_1193# DRVHI_H_uq5 a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X61 VGND PU_DIS_H a_638_279# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X62 VGND a_947_1193# DRVHI_H_uq5 VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
.ends

.subckt sky130_fd_io__com_opath_datoev2 OUT OE_N DRVHI_H DRVLO_H_N VCC_IO VGND HLD_I_OVR_H
+ VPWR_KA OE_H OD_H sky130_fd_io__gpio_dat_ls_1v2_0/SET_H li_5565_99# w_5565_99# sky130_fd_io__gpio_dat_ls_1v2_0/OUT_H
+ w_n227_n1072#
Xsky130_fd_io__gpio_dat_ls_1v2_0 OUT sky130_fd_io__com_cclat_0/PU_DIS_H VGND sky130_fd_io__gpio_dat_ls_1v2_0/SET_H
+ HLD_I_OVR_H VCC_IO VGND sky130_fd_io__gpio_dat_ls_1v2_0/OUT_H VPWR_KA sky130_fd_io__gpio_dat_ls_1v2
Xsky130_fd_io__gpio_dat_lsv2_0 OE_N OE_H VGND OD_H HLD_I_OVR_H VCC_IO VGND sky130_fd_io__com_cclat_0/OE_H_N
+ VPWR_KA a_28_1762# sky130_fd_io__gpio_dat_lsv2
Xsky130_fd_io__com_cclat_0 sky130_fd_io__com_cclat_0/PU_DIS_H sky130_fd_io__gpio_dat_ls_1v2_0/OUT_H
+ VGND sky130_fd_io__com_cclat_0/OE_H_N DRVLO_H_N DRVHI_H VCC_IO sky130_fd_io__com_cclat
.ends

.subckt sky130_fd_io__com_pdpredrvr_strong_slowv2 DRVLO_H_N PDEN_H_N VCC_IO VGND_IO
+ PD_H VSUBS w_59_800#
X0 a_125_866# DRVLO_H_N PD_H w_59_800# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X1 a_125_866# PDEN_H_N VCC_IO w_59_800# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X2 PD_H DRVLO_H_N VGND_IO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X3 VCC_IO PDEN_H_N a_125_866# w_59_800# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X4 PD_H DRVLO_H_N a_125_866# w_59_800# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X5 VGND_IO PDEN_H_N PD_H VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
.ends

.subckt sky130_fd_io__com_pdpredrvr_weakv2 DRVLO_H_N PDEN_H_N VGND_IO VCC_IO PD_H
X0 VCC_IO PDEN_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X1 PD_H DRVLO_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X2 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X3 a_73_866# PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X4 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
.ends

.subckt sky130_fd_io__com_pdpredrvr_pbiasv2 EN_H VGND_IO VCC_IO_uq1 PBIAS_uq5 DRVLO_H_N_uq1
+ EN_H_N PDEN_H_N PD_H VSUBS a_16799_2980# a_18190_3078# a_13911_2980# a_12120_4573#
+ a_12434_3172# a_16899_3078#
X0 a_11460_4784# DRVLO_H_N_uq1 VGND_IO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X1 a_12578_4025# PD_H a_12434_3172# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=4e+06u
X2 PBIAS_uq5 PBIAS_uq5 a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R0 PBIAS_uq5 m1_12872_3935# short w=650000u l=10000u
R1 a_13911_2980# m1_15141_3027# short w=230000u l=10000u
X3 a_13911_2980# a_13911_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R2 a_11368_4652# m1_11681_3387# short w=260000u l=10000u
X4 PBIAS_uq5 a_11581_4213# VGND_IO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=1e+06u
X5 VCC_IO_uq1 a_13911_2980# a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X6 a_13911_2980# PBIAS_uq5 PBIAS_uq5 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X7 VGND_IO a_11581_4213# PBIAS_uq5 VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=1e+06u
X8 a_16899_3078# a_16799_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X9 VCC_IO_uq1 a_16799_2980# a_16899_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X10 a_12120_4573# a_12120_4573# a_18190_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X11 a_11581_4213# DRVLO_H_N_uq1 VGND_IO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
R3 a_13911_2980# m1_16797_3553# short w=230000u l=10000u
X12 a_16799_2980# a_18190_3078# a_18190_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R4 m1_16797_3553# a_16899_3078# short w=230000u l=10000u
X13 PBIAS_uq5 PBIAS_uq5 a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X14 VGND_IO PD_H a_12434_3172# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=4e+06u
X15 a_16899_3078# a_16799_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X16 VGND_IO PDEN_H_N a_11460_4784# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X17 VCC_IO_uq1 EN_H_N a_13361_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X18 a_13911_2980# a_13911_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X19 a_13911_2980# PBIAS_uq5 PBIAS_uq5 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X20 a_18190_3078# a_12120_4573# a_12120_4573# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X21 VCC_IO_uq1 a_16799_2980# a_16899_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X22 a_18190_3078# a_12120_4573# a_12120_4573# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X23 a_16799_2980# VGND_IO VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=8e+06u
X24 VCC_IO_uq1 a_13911_2980# a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X25 VCC_IO_uq1 a_13911_2980# a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X26 a_13347_3873# DRVLO_H_N_uq1 VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X27 PBIAS_uq5 PBIAS_uq5 a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X28 VCC_IO_uq1 EN_H PBIAS_uq5 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R5 m1_12872_3935# a_12906_4025# short w=650000u l=10000u
X29 PBIAS_uq5 PBIAS_uq5 a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R6 a_11368_4652# m1_11524_4701# short w=2.5e+06u l=10000u
X30 VGND_IO a_11460_4784# a_11581_4213# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X31 a_13347_3873# DRVLO_H_N_uq1 VGND_IO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X32 a_13911_2980# a_13911_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R7 a_11781_4311# m1_11840_4382# short w=260000u l=10000u
X33 a_13219_3078# DRVLO_H_N_uq1 a_11581_4213# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X34 a_16899_3078# a_16799_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X35 a_16799_2980# a_18190_3078# a_18190_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X36 VGND_IO a_11581_4213# a_12120_4573# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X37 VCC_IO_uq1 a_13347_3873# a_16799_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R8 m1_13288_3471# EN_H_N short w=640000u l=10000u
X38 a_11781_4311# a_11581_4213# VGND_IO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=1e+06u
X39 a_13361_3078# a_11368_4652# a_13219_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X40 VCC_IO_uq1 a_16799_2980# a_16899_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X41 a_18190_3078# a_18190_3078# a_16799_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R9 m1_11840_4382# PBIAS_uq5 short w=260000u l=10000u
X42 VGND_IO a_11581_4213# a_11781_4311# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=1e+06u
X43 VGND_IO EN_H_N a_11581_4213# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X44 a_13911_2980# PBIAS_uq5 PBIAS_uq5 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R10 m1_11681_3387# PD_H short w=260000u l=10000u
X45 VCC_IO_uq1 a_16799_2980# a_16899_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X46 a_12906_4025# a_11581_4213# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=4e+06u
R11 m1_15178_3027# PBIAS_uq5 short w=230000u l=10000u
X47 VCC_IO_uq1 a_13911_2980# a_13911_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X48 a_12120_4573# a_12120_4573# a_18190_3078# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X49 a_16899_3078# a_16799_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R12 a_11368_4652# m1_13251_3471# short w=640000u l=10000u
R13 a_11460_4784# m1_11524_4738# short w=2.5e+06u l=10000u
R14 a_12578_4025# m1_12556_4086# short w=650000u l=10000u
X50 VCC_IO_uq1 DRVLO_H_N_uq1 a_13347_3873# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X51 a_13911_2980# a_13911_2980# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X52 a_18190_3078# a_18190_3078# a_16799_2980# VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X53 PBIAS_uq5 a_13347_3873# VCC_IO_uq1 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
R15 m1_12556_4086# a_11581_4213# short w=650000u l=10000u
X54 a_11460_4784# a_11368_4652# a_11368_4652# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X55 a_13911_2980# PBIAS_uq5 PBIAS_uq5 VCC_IO_uq1 sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_octl_mux SEL_H_N A_H Y_H B_H SEL_H VSUBS w_1191_2415#
+ w_1266_1185#
X0 A_H SEL_H_N Y_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X1 Y_H SEL_H A_H VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X2 B_H SEL_H_N Y_H VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 Y_H SEL_H B_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 DRVLO_H_N PD_I2C_H PDEN_H_N PD_H
+ VCC_IO I2C_MODE_H VGND_IO EN_FAST_N[0] EN_FAST_N[1] w_4658_n980#
X0 a_7724_n1285# DRVLO_H_N PD_I2C_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X1 a_4877_n914# I2C_MODE_H VCC_IO w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X2 PD_H I2C_MODE_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X3 PD_H DRVLO_H_N a_5469_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X4 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X5 a_5781_n914# DRVLO_H_N PD_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X6 a_7449_n1327# PDEN_H_N a_4877_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=4e+06u
X7 a_7449_n1327# PDEN_H_N a_6596_n1327# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=4e+06u
X8 a_6596_n1327# DRVLO_H_N PD_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=4e+06u
X9 VGND_IO DRVLO_H_N PD_I2C_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X10 PD_I2C_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X11 VCC_IO I2C_MODE_H a_4877_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X12 PD_I2C_H DRVLO_H_N a_6596_n885# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=4e+06u
X13 a_5469_n914# DRVLO_H_N PD_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X14 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X15 a_4877_n914# I2C_MODE_H VCC_IO w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X16 VGND_IO PDEN_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X17 a_4877_n914# EN_FAST_N[0] a_5469_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X18 VCC_IO PDEN_H_N a_6596_n885# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=4e+06u
X19 VCC_IO EN_FAST_N[1] a_7724_n1285# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X20 a_5781_n914# EN_FAST_N[1] a_4877_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X21 PD_H DRVLO_H_N a_5781_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X22 PD_I2C_H DRVLO_H_N a_7724_n1285# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X23 PD_I2C_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong_nr3 EN_FAST_N[0] EN_FAST_N[1] I2C_MODE_H
+ PDEN_H_N DRVLO_H_N PD_H VCC_IO VGND_IO
X0 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X1 a_1708_456# DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X3 a_1992_n250# DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=2e+06u
X4 PD_H DRVLO_H_N a_2477_n356# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X6 a_1592_172# PDEN_H_N a_1139_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=2e+06u
X7 PD_H DRVLO_H_N a_1592_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=2e+06u
X8 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X9 PD_H DRVLO_H_N a_1708_456# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X11 a_1708_456# EN_FAST_N[0] a_1139_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 VCC_IO EN_FAST_N[0] a_2168_n356# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 a_2168_n356# DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VCC_IO I2C_MODE_H a_1139_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X15 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X16 a_1139_172# EN_FAST_N[1] a_1708_456# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X17 a_1139_172# I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X18 a_2477_n356# EN_FAST_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 a_1992_n250# PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=4e+06u
X20 VGND_IO PDEN_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong PD_H[3] PD_H[2] VGND VCC_IO DRVLO_H_N
+ SLOW_H PDEN_H_N_uq2 I2C_MODE_H_N PD_H[4] sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ m2_9346_3319# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078# sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5 sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
Xsky130_fd_io__com_pdpredrvr_pbiasv2_0 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H
+ VGND VCC_IO sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5 DRVLO_H_N sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N
+ PDEN_H_N_uq2 PD_H[4] VGND sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ sky130_fd_io__com_pdpredrvr_pbiasv2
Xsky130_fd_io__gpiov2_octl_mux_0 I2C_MODE_H_N sky130_fd_io__gpiov2_octl_mux_0/A_H
+ sky130_fd_io__gpiov2_octl_mux_0/Y_H DRVLO_H_N sky130_fd_io__hvsbt_nand2_1/IN0 VGND
+ VCC_IO VGND sky130_fd_io__gpiov2_octl_mux
Xsky130_fd_io__hvsbt_nand2_0 SLOW_H I2C_MODE_H_N sky130_fd_io__hvsbt_nand2_0/OUT VGND
+ VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_1 SLOW_H sky130_fd_io__hvsbt_nand2_1/IN0 sky130_fd_io__hvsbt_nand2_1/OUT
+ VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__gpiov2_pdpredrvr_strong_nr2_0 DRVLO_H_N PD_H[4] PDEN_H_N_uq2 PD_H[2]
+ VCC_IO sky130_fd_io__hvsbt_inv_x1_1/OUT VGND sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5 VCC_IO sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x1_0/OUT VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_0/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[0]
+ sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] sky130_fd_io__hvsbt_inv_x1_1/OUT
+ PDEN_H_N_uq2 sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VCC_IO VGND sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_inv_x1_1/OUT VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_1/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
R0 m1_9403_1623# m1_9430_1596# short w=260000u l=10000u
X0 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
R1 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[0] m1_9575_2734# short w=260000u l=10000u
X1 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H PDEN_H_N_uq2 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X2 VGND PD_H[4] sky130_fd_io__gpiov2_octl_mux_0/A_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
R2 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] m1_9830_1715# short w=260000u l=10000u
R3 sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5 m1_9427_1780# short w=260000u l=10000u
X3 sky130_fd_io__hvsbt_nand2_1/IN0 I2C_MODE_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X4 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
R4 m1_9427_1780# sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] short w=260000u l=10000u
R5 sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5 m1_9364_1624# short w=260000u l=10000u
R6 m1_9364_1624# m1_9403_1623# short w=260000u l=10000u
R7 m1_9575_2734# VCC_IO short w=260000u l=10000u
R8 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N m1_9430_1559# short w=260000u l=10000u
X5 sky130_fd_io__hvsbt_nand2_1/IN0 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X6 VGND sky130_fd_io__hvsbt_inv_x1_0/OUT sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
R9 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[0] m1_9830_1752# short w=260000u l=10000u
X7 VCC_IO PD_H[4] sky130_fd_io__gpiov2_octl_mux_0/A_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X8 a_8987_763# PDEN_H_N_uq2 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
R10 m1_9599_1482# sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] short w=260000u l=10000u
X9 VCC_IO sky130_fd_io__hvsbt_inv_x1_0/OUT a_8987_763# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X10 sky130_fd_io__hvsbt_nand2_1/IN0 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
R11 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N m1_9562_1482# short w=260000u l=10000u
.ends

.subckt sky130_fd_io__com_pupredrvr_strong_slowv2 PUEN_H DRVHI_H PU_H_N VGND_IO VCC_IO
+ a_93_102#
X0 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X1 VGND_IO PUEN_H a_93_102# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X2 PU_H_N DRVHI_H a_93_102# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X3 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X4 a_93_102# PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X5 a_93_102# DRVHI_H PU_H_N VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X6 VCC_IO PUEN_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X7 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
.ends

.subckt sky130_fd_io__feas_com_pupredrvr_weak DRVHI_H PUEN_H PU_H_N VGND_IO VCC_IO
+ VSUBS w_21_799#
X0 PU_H_N DRVHI_H a_280_102# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X1 VCC_IO DRVHI_H PU_H_N w_21_799# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X2 VCC_IO PUEN_H PU_H_N w_21_799# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X3 PU_H_N DRVHI_H VCC_IO w_21_799# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X4 a_280_102# PUEN_H VGND_IO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
.ends

.subckt sky130_fd_io__feascom_pupredrvr_nbiasv2 EN_H_N EN_H_uq1 VGND_IO_uq2 NBIAS_uq3
+ DRVHI_H PUEN_H VCC_IO PU_H_N_uq1 a_1772_220# a_2874_118# a_2821_220# a_261_220#
X0 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X1 NBIAS_uq3 NBIAS_uq3 a_261_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X2 NBIAS_uq3 EN_H_N VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 NBIAS_uq3 a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X4 VGND_IO_uq2 a_261_220# a_261_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X5 NBIAS_uq3 NBIAS_uq3 a_261_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X6 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X7 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X8 a_1672_194# a_2821_220# a_2821_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X9 VGND_IO_uq2 a_261_220# a_261_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
R0 m1_1014_800# a_1004_990# short w=260000u l=10000u
X10 VCC_IO a_250_1898# a_2874_118# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X11 VGND_IO_uq2 a_1672_194# a_1772_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
R1 a_562_1898# m1_2838_1831# short w=260000u l=10000u
R2 a_620_1263# m1_2838_1794# short w=260000u l=10000u
X12 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X13 VGND_IO_uq2 a_1672_194# a_1772_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
R3 NBIAS_uq3 m1_1409_1332# short w=230000u l=10000u
X14 VGND_IO_uq2 a_207_1014# NBIAS_uq3 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X15 a_2821_220# a_2874_118# a_2874_118# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
R4 a_261_220# m1_1608_646# short w=230000u l=10000u
R5 m1_1046_126# a_261_220# short w=260000u l=10000u
X16 VCC_IO DRVHI_H a_562_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
R6 m1_702_1715# a_620_1263# short w=230000u l=10000u
X17 a_2421_2014# PU_H_N_uq1 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=8e+06u
X18 VCC_IO a_250_1898# NBIAS_uq3 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X19 a_2821_220# a_2821_220# a_1672_194# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
R7 EN_H_uq1 m1_575_1252# short w=260000u l=10000u
R8 m1_612_1252# a_620_1263# short w=260000u l=10000u
R9 m1_1409_1332# a_1507_1397# short w=230000u l=10000u
X20 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X21 a_562_1898# a_620_1263# a_620_1263# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X22 a_261_220# NBIAS_uq3 NBIAS_uq3 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X23 a_261_220# a_261_220# VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X24 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X25 a_261_220# NBIAS_uq3 NBIAS_uq3 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X26 a_250_1898# DRVHI_H a_737_914# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X27 VCC_IO DRVHI_H a_207_1014# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X28 a_583_914# EN_H_uq1 VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X29 a_1772_220# a_1672_194# VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
R10 NBIAS_uq3 m1_1014_800# short w=260000u l=10000u
X30 VCC_IO EN_H_uq1 a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
R11 a_2421_2014# m1_2596_1928# short w=260000u l=10000u
R12 m1_2596_1928# a_250_1898# short w=260000u l=10000u
X31 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X32 a_1772_220# a_1672_194# VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
R13 NBIAS_uq3 m1_1014_127# short w=260000u l=10000u
X33 a_562_1898# PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X34 VGND_IO_uq2 DRVHI_H a_207_1014# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X35 a_2874_118# a_2874_118# a_2821_220# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X36 a_2874_118# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X37 a_737_914# a_620_1263# a_583_914# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X38 NBIAS_uq3 a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X39 VCC_IO a_250_1898# NBIAS_uq3 VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=800000u
X40 a_1672_194# VCC_IO VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=8e+06u
R14 PU_H_N_uq1 m1_702_1715# short w=230000u l=10000u
X41 a_261_220# a_261_220# VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X42 a_207_1014# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X43 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X44 VGND_IO_uq2 a_250_1898# a_1004_990# VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=4e+06u
R15 m1_1608_646# a_1772_220# short w=230000u l=10000u
X45 a_250_1898# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X46 a_1672_194# a_207_1014# VGND_IO_uq2 VGND_IO_uq2 sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2 DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] VGND_IO VCC_IO PU_H_N a_158_632#
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X1 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
X2 a_809_632# EN_FAST[2] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
X3 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
X4 PU_H_N DRVHI_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=4e+06u
X5 VGND_IO EN_FAST[3] a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
R0 a_158_632# a_1008_2434# sky130_fd_pr__res_generic_po w=330000u l=1.1e+07u
R1 a_158_632# m1_1184_866# short w=260000u l=10000u
R2 m1_1184_866# PU_H_N short w=260000u l=10000u
X6 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X7 VGND_IO PUEN_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=4e+06u
R3 PU_H_N a_1008_2434# sky130_fd_pr__res_generic_po w=330000u l=4e+06u
X8 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X12 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X13 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] VGND_IO VCC_IO PU_H_N a_609_606# a_353_606#
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X1 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
X2 a_809_632# a_609_606# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
X3 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
X4 VGND_IO a_353_606# a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=1e+06u
R0 a_158_632# a_1008_2434# sky130_fd_pr__res_generic_po w=330000u l=1.1e+07u
R1 a_158_632# m1_1184_866# short w=260000u l=10000u
X5 VGND_IO PUEN_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=4e+06u
R2 m1_1184_866# PU_H_N short w=260000u l=10000u
X6 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
R3 PU_H_N a_1008_2434# sky130_fd_pr__res_generic_po w=330000u l=4e+06u
X7 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X10 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X11 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X12 PU_H_N DRVHI_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=4e+06u
X13 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends

.subckt sky130_fd_io__gpio_pupredrvr_strongv2 VCC_IO VSUBS DRVHI_H PU_H_N[3] PUEN_H
+ PU_H_N[2] SLOW_H_N sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+
Xsky130_fd_io__feascom_pupredrvr_nbiasv2_0 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_uq1 VSUBS sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ DRVHI_H PUEN_H VCC_IO PU_H_N[2] sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220# sky130_fd_io__feascom_pupredrvr_nbiasv2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] VSUBS VCC_IO PU_H_N[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] VSUBS VCC_IO PU_H_N[2]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a
X0 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N SLOW_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
R0 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_uq1 m1_4740_1326# short w=260000u l=10000u
X1 VSUBS PUEN_H a_483_1179# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
R1 m1_6555_1273# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] short w=650000u l=10000u
X2 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_uq1 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
R2 m1_4777_1326# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] short w=260000u l=10000u
R3 VSUBS m1_6555_1273# short w=650000u l=10000u
R4 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6300_1402# short w=650000u l=10000u
R5 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] m1_6300_1365# short w=650000u l=10000u
R6 m1_6265_477# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] short w=650000u l=10000u
R7 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6265_477# short w=650000u l=10000u
X3 a_483_1179# SLOW_H_N sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
R8 m1_5759_509# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] short w=260000u l=10000u
R9 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_uq1 m1_5722_509# short w=260000u l=10000u
R10 m1_5786_421# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] short w=260000u l=10000u
R11 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6556_1402# short w=650000u l=10000u
R12 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] m1_6556_1365# short w=650000u l=10000u
R13 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3 m1_4655_1468# short w=260000u l=10000u
R14 m1_4655_1468# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] short w=260000u l=10000u
X4 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_uq1 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
R15 VSUBS m1_6266_605# short w=650000u l=10000u
R16 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] m1_6266_568# short w=650000u l=10000u
X5 VCC_IO PUEN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
R17 m1_6299_1273# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] short w=650000u l=10000u
R18 VSUBS m1_6299_1273# short w=650000u l=10000u
R19 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3 m1_5786_421# short w=260000u l=10000u
.ends

.subckt sky130_fd_io__gpiov2_obpredrvr PD_H[3] PD_H[2] PDEN_H_N[1] DRVHI_H DRVLO_H_N_uq2
+ VGND PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] PD_H[1] PD_H[0] PD_H[4] SLOW_H PUEN_H[1]
+ PUEN_H[0] PDEN_H_N[0] VCC_IO SLOW_H_N I2C_MODE_H_N sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102# sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+
Xsky130_fd_io__com_pdpredrvr_strong_slowv2_0 DRVLO_H_N_uq2 PDEN_H_N[1] VCC_IO VGND
+ PD_H[1] VGND VCC_IO sky130_fd_io__com_pdpredrvr_strong_slowv2
Xsky130_fd_io__com_pdpredrvr_weakv2_0 DRVLO_H_N_uq2 PDEN_H_N[0] VGND VCC_IO PD_H[0]
+ sky130_fd_io__com_pdpredrvr_weakv2
Xsky130_fd_io__gpiov2_pdpredrvr_strong_0 PD_H[3] PD_H[2] VGND VCC_IO DRVLO_H_N_uq2
+ SLOW_H PDEN_H_N[1] I2C_MODE_H_N PD_H[4] sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ PUEN_H[1] sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_pdpredrvr_strong
Xsky130_fd_io__com_pupredrvr_strong_slowv2_0 PUEN_H[1] DRVHI_H PU_H_N[1] VGND VCC_IO
+ sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102# sky130_fd_io__com_pupredrvr_strong_slowv2
Xsky130_fd_io__feas_com_pupredrvr_weak_0 DRVHI_H PUEN_H[0] PU_H_N[0] VGND VCC_IO VGND
+ VCC_IO sky130_fd_io__feas_com_pupredrvr_weak
Xsky130_fd_io__gpio_pupredrvr_strongv2_0 VCC_IO VGND DRVHI_H PU_H_N[3] PUEN_H[1] PU_H_N[2]
+ SLOW_H_N sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2
.ends

.subckt sky130_fd_io__gpiov2_octl_dat VPWR VGND VCC_IO VPWR_KA SLOW HLD_I_H_N HLD_I_OVR_H
+ OD_H SLOW_H_N DRVHI_H PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] PD_H[1] PD_H[0] PD_H[4]
+ DRVLO_H_N DM_H_N[2] DM_H_N[0] DM_H[2] DM_H[1] DM_H[0] OUT OE_N DM_H_N[1] PD_H[3]
+ PD_H[2] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__com_opath_datoev2_0/w_5565_99# sky130_fd_io__com_opath_datoev2_0/li_5565_99#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__com_opath_datoev2_0/w_n227_n1072# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+
Xsky130_fd_io__gpiov2_octl_0 DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2] sky130_fd_io__gpiov2_octl_0/PUEN_2OR1_H
+ DM_H[1] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0]
+ OD_H SLOW sky130_fd_io__gpiov2_octl_0/SLOW_H SLOW_H_N HLD_I_H_N VCC_IO VGND VPWR
+ sky130_fd_io__gpiov2_obpredrvr_0/I2C_MODE_H_N VCC_IO a_13335_4479# VCC_IO DM_H[1]
+ DM_H[2] sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[1] DM_H[0] sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[0]
+ VGND VCC_IO VCC_IO a_13335_4479# sky130_fd_io__gpiov2_octl
Xsky130_fd_io__com_opath_datoev2_0 OUT OE_N DRVHI_H DRVLO_H_N VCC_IO VGND HLD_I_OVR_H
+ VPWR_KA sky130_fd_io__com_opath_datoev2_0/OE_H OD_H OD_H sky130_fd_io__com_opath_datoev2_0/li_5565_99#
+ sky130_fd_io__com_opath_datoev2_0/w_5565_99# sky130_fd_io__com_opath_datoev2_0/sky130_fd_io__gpio_dat_ls_1v2_0/OUT_H
+ sky130_fd_io__com_opath_datoev2_0/w_n227_n1072# sky130_fd_io__com_opath_datoev2
Xsky130_fd_io__gpiov2_obpredrvr_0 PD_H[3] PD_H[2] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1]
+ DRVHI_H DRVLO_H_N VGND PU_H_N[3] PU_H_N[2] PU_H_N[1] PU_H_N[0] PD_H[1] PD_H[0] PD_H[4]
+ sky130_fd_io__gpiov2_octl_0/SLOW_H sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[1] sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[0]
+ sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0] VCC_IO SLOW_H_N sky130_fd_io__gpiov2_obpredrvr_0/I2C_MODE_H_N
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_obpredrvr
.ends

.subckt sky130_fd_io__com_pudrvr_strong_slowv2 PU_H_N PAD VSUBS a_356_297# w_122_n30#
+ w_n10_n150#
X0 w_122_n30# PU_H_N PAD w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X1 PAD PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X2 a_356_297# PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X3 w_122_n30# PU_H_N a_356_297# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X4 w_122_n30# PU_H_N PAD w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X5 PAD PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X6 a_356_297# PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X7 w_122_n30# PU_H_N a_356_297# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
.ends

.subckt sky130_fd_io__com_res_weak_bentbigres VSUBS a_n2_6046# a_419_9396# a_419_8146#
+ a_n256_8772# a_419_8054# a_419_6804#
R0 a_419_8146# a_419_9396# sky130_fd_pr__res_generic_po w=800000u l=6e+06u
R1 a_n258_6046# a_n2_6046# sky130_fd_pr__res_generic_po w=800000u l=5e+07u
R2 a_n258_6046# a_n256_8772# sky130_fd_pr__res_generic_po w=800000u l=1.2e+07u
R3 a_419_6804# a_419_8054# sky130_fd_pr__res_generic_po w=800000u l=6e+06u
.ends

.subckt sky130_fd_io__com_res_weak RB RA VSUBS
Xsky130_fd_io__com_res_weak_bentbigres_0 VSUBS RA a_n160_9488# li_n135_8054# li_n135_6820#
+ li_n135_8054# li_n135_6820# sky130_fd_io__com_res_weak_bentbigres
R0 m1_n147_10115# a_n160_10423# short w=660000u l=10000u
R1 m1_n147_8777# a_n160_9488# short w=660000u l=10000u
R2 a_n160_9838# m1_n147_10115# short w=660000u l=10000u
R3 m1_n147_9555# a_n160_9838# short w=660000u l=10000u
R4 li_n135_8054# m1_n147_8777# short w=660000u l=10000u
R5 RB a_517_9818# sky130_fd_pr__res_generic_po w=800000u l=1.5e+06u
R6 a_n160_9488# m1_n147_9555# short w=660000u l=10000u
R7 m1_532_9534# a_517_9818# short w=660000u l=10000u
R8 RB m1_532_9534# short w=660000u l=10000u
R9 a_n160_9488# a_n160_9838# sky130_fd_pr__res_generic_po w=800000u l=1.5e+06u
R10 li_n135_8054# m1_n146_7735# short w=660000u l=10000u
R11 li_n135_6820# m1_n146_7434# short w=660000u l=10000u
R12 a_n160_9838# a_n160_10423# sky130_fd_pr__res_generic_po w=800000u l=1.5e+06u
R13 m1_532_10115# a_n160_10423# short w=660000u l=10000u
R14 a_517_9818# a_n160_10423# sky130_fd_pr__res_generic_po w=800000u l=1.5e+06u
R15 a_517_9818# m1_532_10115# short w=660000u l=10000u
.ends

.subckt sky130_fd_io__pfet_con_diff_wo_abt_270v2 VSUBS a_6833_1380# w_36_314# a_881_1380#
+ a_11793_1380# a_3857_1380# a_13215_1380# a_1873_1380# a_8255_1380# a_10239_1380#
+ a_11231_1380# a_5279_1380# a_6271_1380# a_1001_1552# a_9809_1380# a_3295_1380# a_7825_1380#
+ a_12785_1380# a_1311_1380# a_14135_1380# a_10801_1380# a_4849_1380# a_5841_1380#
+ a_2865_1380# a_9247_1380# a_12223_1380# a_7263_1380# a_4287_1380# a_8817_1380# a_13777_1380#
+ a_2303_1380# w_415_600#
X0 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X1 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X2 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X3 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X4 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X5 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X6 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X7 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X8 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X9 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X10 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X11 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X12 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X13 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X14 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X15 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X16 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X17 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X18 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X19 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X20 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X21 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X22 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X23 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X24 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X25 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X26 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X27 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X28 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X29 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X30 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X31 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X32 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X33 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X34 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X35 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X36 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X37 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X38 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X39 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X40 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X41 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X42 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X43 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X44 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X45 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X46 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X47 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X48 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X49 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X50 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X51 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X52 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X53 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X54 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
X55 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=600000u
.ends

.subckt sky130_fd_io__gpio_pudrvr_strongv2 PU_H_N[3] PU_H_N[2] VCC_IO TIE_HI_ESD VNB
+ PAD VSUBS li_9083_n155# m1_6033_n459# m1_14880_n614# m1_3028_333# a_14575_n157#
+ m1_6658_n459# m1_1330_n459# m1_3421_98#
Xsky130_fd_io__pfet_con_diff_wo_abt_270v2_0 VSUBS PU_H_N[3] VNB PU_H_N[2] m1_11745_1478#
+ PU_H_N[3] m1_13667_1478# PU_H_N[2] m1_8837_1478# m1_10391_1478# m1_11745_1478# PU_H_N[3]
+ PU_H_N[3] PAD m1_10391_1478# PU_H_N[2] PU_H_N[3] PU_H_N[2] PU_H_N[2] m1_14229_1478#
+ m1_10391_1478# PU_H_N[3] PU_H_N[3] PU_H_N[2] m1_8837_1478# m1_11745_1478# PU_H_N[3]
+ PU_H_N[3] m1_8837_1478# m1_14229_1478# PU_H_N[2] VCC_IO sky130_fd_io__pfet_con_diff_wo_abt_270v2
R0 m1_11745_1478# m2_12608_116# short w=650000u l=10000u
R1 TIE_HI_ESD m2_10197_n209# short w=650000u l=10000u
R2 PU_H_N[3] m2_10439_n209# short w=650000u l=10000u
R3 PU_H_N[2] m2_11422_n209# short w=650000u l=10000u
R4 PU_H_N[2] m2_12849_n185# short w=650000u l=10000u
R5 m1_13667_1478# m2_13593_958# short w=650000u l=10000u
R6 TIE_HI_ESD m2_13593_657# short w=650000u l=10000u
R7 m1_8837_1478# m2_10197_92# short w=650000u l=10000u
R8 m1_10391_1478# m2_10945_92# short w=650000u l=10000u
R9 PU_H_N[3] m2_11186_n208# short w=650000u l=10000u
R10 m1_13667_1478# m2_14075_958# short w=650000u l=10000u
R11 m2_14286_658# m1_14229_1478# short w=650000u l=10000u
R12 m2_10673_n208# m1_8837_1478# short w=650000u l=10000u
R13 m2_12365_n184# m1_11745_1478# short w=650000u l=10000u
R14 TIE_HI_ESD m2_14286_658# short w=650000u l=10000u
R15 PU_H_N[2] m2_14075_657# short w=650000u l=10000u
R16 m2_11186_n208# m1_10391_1478# short w=650000u l=10000u
R17 m1_11745_1478# m2_12849_116# short w=650000u l=10000u
R18 TIE_HI_ESD m2_12365_n184# short w=650000u l=10000u
R19 PU_H_N[3] m2_12608_n185# short w=650000u l=10000u
R20 m2_13837_658# m1_13667_1478# short w=650000u l=10000u
R21 TIE_HI_ESD a_14575_n157# sky130_fd_pr__res_generic_po w=500000u l=1.02e+07u
R22 TIE_HI_ESD m2_10945_n209# short w=650000u l=10000u
R23 m1_14229_1478# m2_14532_958# short w=650000u l=10000u
R24 m1_14229_1478# m2_14769_958# short w=650000u l=10000u
R25 m1_8837_1478# m2_10439_92# short w=650000u l=10000u
R26 m1_10391_1478# m2_11422_92# short w=650000u l=10000u
R27 PU_H_N[2] m2_10673_n208# short w=650000u l=10000u
R28 PU_H_N[3] m2_13837_658# short w=650000u l=10000u
R29 PU_H_N[3] m2_14532_657# short w=650000u l=10000u
R30 PU_H_N[2] m2_14769_657# short w=650000u l=10000u
.ends

.subckt sky130_fd_io__nfet_con_diff_wo_abt_270v2 VCC_IO VSSIO PAD VSUBS a_9852_1285#
+ a_2346_1285# a_11836_1285# a_924_1285# a_6876_1285# a_4892_1285# a_1916_1285# a_9290_1285#
+ a_13258_1285# a_8298_1285# a_6314_1285# a_11274_1285# a_3338_1285# a_4330_1285#
+ a_13820_1285# a_8860_1285# a_12828_1285# a_7868_1285# a_1354_1285# a_10844_1285#
+ a_14178_1285# a_5884_1285# a_2908_1285# a_3900_1285# a_7306_1285# a_12266_1285#
+ a_5322_1285# a_10282_1285#
X0 PAD a_3900_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X1 PAD a_5884_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X2 VSSIO a_14178_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X3 VSSIO a_7306_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X4 PAD a_7868_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X5 VSSIO a_13258_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X6 VSSIO a_1354_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X7 PAD a_8860_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X8 PAD a_11836_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X9 VSSIO a_6314_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X10 VSSIO a_8298_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X11 VSSIO a_9290_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X12 VSSIO a_12266_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X13 PAD a_6876_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X14 PAD a_10844_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X15 PAD a_924_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X16 VSSIO a_2346_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X17 PAD a_9852_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X18 PAD a_12828_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X19 VSSIO a_7306_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X20 PAD a_13820_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X21 VSSIO a_13258_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X22 VSSIO a_1354_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X23 PAD a_7868_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X24 PAD a_8860_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X25 PAD a_11836_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X26 VSSIO a_3338_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X27 VSSIO a_4330_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X28 PAD a_1916_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X29 PAD a_4892_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X30 VSSIO a_10282_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X31 PAD a_924_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X32 VSSIO a_2346_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X33 PAD a_9852_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X34 PAD a_12828_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X35 PAD a_13820_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X36 VSSIO a_5322_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X37 PAD a_2908_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X38 PAD a_5884_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X39 VSSIO a_11274_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X40 VSSIO a_14178_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X41 PAD a_3900_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X42 VSSIO a_3338_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X43 VSSIO a_4330_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X44 PAD a_1916_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X45 VSSIO a_10282_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X46 PAD a_4892_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X47 VSSIO a_6314_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X48 VSSIO a_8298_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X49 PAD a_6876_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X50 VSSIO a_9290_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X51 VSSIO a_12266_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X52 PAD a_10844_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X53 VSSIO a_5322_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X54 PAD a_2908_1285# VSSIO VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X55 VSSIO a_11274_1285# PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_pddrvr_strong VCC_IO PD_H[2] PD_H[3] TIE_LO_ESD VGND_IO
+ VSSIO_AMX FORCE_LOVOL_H FORCE_LO_H PAD PD_H_I2C VSUBS m1_9575_2540# m1_4511_2373#
+ m1_225_1760# m1_320_1652# m2_8958_2367# m1_2396_2540#
Xsky130_fd_io__nfet_con_diff_wo_abt_270v2_0 VCC_IO VGND_IO PAD VSUBS PD_H[3] m1_12747_3898#
+ PD_H[3] m1_12747_3898# m1_8232_3898# m1_9769_3898# m1_12747_3898# PD_H[3] m1_785_3898#
+ PD_H[2] m1_8232_3898# PD_H[3] m1_11193_3898# m1_9769_3898# m1_785_3898# PD_H[2]
+ m1_2135_3898# PD_H[2] m1_12747_3898# PD_H[3] m1_785_3898# m1_8232_3898# m1_11193_3898#
+ m1_11193_3898# m1_7657_3898# PD_H_I2C m1_9769_3898# PD_H[3] sky130_fd_io__nfet_con_diff_wo_abt_270v2
R0 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po w=500000u l=1.02e+07u
R1 TIE_LO_ESD m2_1848_1637# short w=650000u l=10000u
R2 TIE_LO_ESD m2_9366_1637# short w=650000u l=10000u
R3 TIE_LO_ESD m2_7664_1637# short w=650000u l=10000u
R4 m1_12747_3898# m2_12763_1938# short w=650000u l=10000u
R5 m1_9769_3898# m2_10846_1938# short w=650000u l=10000u
R6 m1_12747_3898# m2_13193_1938# short w=650000u l=10000u
R7 PD_H[2] m2_12763_1637# short w=650000u l=10000u
R8 TIE_LO_ESD m2_10846_1637# short w=650000u l=10000u
R9 PD_H[3] m2_13193_1637# short w=650000u l=10000u
R10 m1_8232_3898# m2_8506_1938# short w=650000u l=10000u
R11 m1_785_3898# m2_414_1938# short w=650000u l=10000u
R12 m1_7657_3898# m2_6804_1938# short w=650000u l=10000u
R13 m2_7233_1638# m1_7657_3898# short w=650000u l=10000u
R14 PD_H[2] m2_6804_1637# short w=650000u l=10000u
R15 PD_H[2] m2_8506_1637# short w=650000u l=10000u
R16 m2_655_1638# m1_785_3898# short w=650000u l=10000u
R17 TIE_LO_ESD m2_414_1637# short w=650000u l=10000u
R18 PD_H[3] m2_7233_1638# short w=650000u l=10000u
R19 PD_H[3] m2_655_1638# short w=650000u l=10000u
R20 m2_10415_1638# m1_9769_3898# short w=650000u l=10000u
R21 m2_11758_1638# m1_11193_3898# short w=650000u l=10000u
R22 m1_2135_3898# m2_1565_1938# short w=650000u l=10000u
R23 PD_H[3] m2_10415_1638# short w=650000u l=10000u
R24 m2_1260_1638# m1_2135_3898# short w=650000u l=10000u
R25 m1_11193_3898# m2_12189_1938# short w=650000u l=10000u
R26 PD_H[3] m2_11758_1638# short w=650000u l=10000u
R27 PD_H[3] m2_1565_1637# short w=650000u l=10000u
R28 PD_H[2] m2_1260_1638# short w=650000u l=10000u
R29 m1_9769_3898# m2_9986_1938# short w=650000u l=10000u
R30 m2_13622_1638# m1_12747_3898# short w=650000u l=10000u
R31 TIE_LO_ESD m2_12189_1637# short w=650000u l=10000u
R32 PD_H[2] m2_9986_1637# short w=650000u l=10000u
R33 m1_785_3898# m2_897_1938# short w=650000u l=10000u
R34 TIE_LO_ESD m2_13622_1638# short w=650000u l=10000u
R35 PD_H[2] m2_897_1637# short w=650000u l=10000u
R36 m1_11193_3898# m2_11329_1938# short w=650000u l=10000u
R37 m1_2135_3898# m2_1848_1938# short w=650000u l=10000u
R38 m2_8935_1638# m1_8232_3898# short w=650000u l=10000u
R39 PD_H[2] m2_11329_1637# short w=650000u l=10000u
R40 m1_7657_3898# m2_7664_1938# short w=650000u l=10000u
R41 m1_8232_3898# m2_9366_1938# short w=650000u l=10000u
R42 PD_H[3] m2_8935_1638# short w=650000u l=10000u
.ends

.subckt sky130_fd_io__com_pudrvr_weakv2 PU_H_N PAD VSUBS a_756_297# w_n10_n150# w_258_n30#
X0 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X1 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X2 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X3 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X4 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X5 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X6 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X7 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
.ends

.subckt sky130_fd_io__gpio_pddrvr_strong_slowv2 PD_H PAD VSUBS dw_n122_n335# w_254_254#
X0 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X1 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X2 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X3 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
.ends

.subckt sky130_fd_io__res250_sub_small VSUBS a_2142_2# a_10_2#
R0 a_10_2# a_2142_2# sky130_fd_pr__res_generic_po w=2e+06u l=1.007e+07u
.ends

.subckt sky130_fd_io__res250only_small PAD ROUT VSUBS
Xsky130_fd_io__res250_sub_small_0 VSUBS ROUT PAD sky130_fd_io__res250_sub_small
.ends

.subckt sky130_fd_io__gpio_pddrvr_weakv2 PD_H PAD VSUBS dw_n122_84# w_254_254#
X0 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X1 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X2 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X3 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X4 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
X5 w_254_254# PD_H PAD VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=600000u
.ends

.subckt sky130_fd_io__gpio_odrvr_subv2 VGND PD_H[0] PD_H[2] PD_H[1] PD_H[3] VCC_IO
+ PAD TIE_LO_ESD FORCE_HI_H_N FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2]
+ PU_H_N[3] VSSIO_AMX VGND_IO TIE_HI_ESD w_n947_8961# sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614# m3_9047_13425# m2_8191_n10933#
+ li_5884_n9263# m3_4600_13425# sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C m3_6107_13425#
+
Xsky130_fd_io__com_pudrvr_strong_slowv2_0 PU_H_N[1] sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD
+ VGND sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD VCC_IO VGND sky130_fd_io__com_pudrvr_strong_slowv2
Xsky130_fd_io__com_res_weak_0 sky130_fd_io__com_res_weak_0/RB sky130_fd_io__com_res_weak_0/RA
+ VGND sky130_fd_io__com_res_weak
Xsky130_fd_io__gpio_pudrvr_strongv2_0 PU_H_N[3] PU_H_N[2] VCC_IO TIE_HI_ESD VGND PAD
+ VGND sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155# VCC_IO sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ VCC_IO VCC_IO VCC_IO VCC_IO PU_H_N[0] sky130_fd_io__gpio_pudrvr_strongv2
Xsky130_fd_io__gpiov2_pddrvr_strong_0 VCC_IO PD_H[2] PD_H[3] TIE_LO_ESD VGND_IO VCC_IO
+ VCC_IO VCC_IO PAD sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C VGND PD_H[0] m3_4600_13425#
+ sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD sky130_fd_io__com_res_weak_0/RA m3_9047_13425#
+ PD_H[1] sky130_fd_io__gpiov2_pddrvr_strong
Xsky130_fd_io__com_pudrvr_weakv2_0 PU_H_N[0] sky130_fd_io__com_res_weak_0/RA VGND
+ sky130_fd_io__com_res_weak_0/RA VGND VCC_IO sky130_fd_io__com_pudrvr_weakv2
Xsky130_fd_io__gpio_pddrvr_strong_slowv2_0 PD_H[1] sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD
+ VGND VCC_IO m3_4600_13425# sky130_fd_io__gpio_pddrvr_strong_slowv2
Xsky130_fd_io__res250only_small_0 PAD sky130_fd_io__com_res_weak_0/RB VGND sky130_fd_io__res250only_small
Xsky130_fd_io__gpio_pddrvr_weakv2_0 PD_H[0] sky130_fd_io__com_res_weak_0/RA VGND VCC_IO
+ m3_9047_13425# sky130_fd_io__gpio_pddrvr_weakv2
R0 a_10314_7886# sky130_fd_io__com_res_weak_0/RB sky130_fd_pr__res_generic_po w=2e+06u l=2e+06u
R1 a_9612_7886# a_10314_7886# sky130_fd_pr__res_generic_po w=2e+06u l=3e+06u
R2 m1_9882_7996# a_10314_7886# short w=1.32e+06u l=10000u
R3 sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD a_9612_7886# sky130_fd_pr__res_generic_po w=2e+06u l=5e+06u
R4 a_9612_7886# m1_9882_7996# short w=1.32e+06u l=10000u
.ends

.subckt sky130_fd_io__gpio_odrvrv2 VGND PAD PD_H[0] PD_H[1] PD_H[2] PD_H[3] TIE_LO_ESD
+ VCC_IO PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3] TIE_HI_ESD VGND_IO FORCE_HI_H_N FORCE_LO_H
+ FORCE_LOVOL_H VSSIO_AMX sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvr_subv2_0/w_n947_8961# sky130_fd_io__gpio_odrvr_subv2_0/m3_9047_13425#
+ sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933# sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263#
+ sky130_fd_io__gpio_odrvr_subv2_0/m3_4600_13425# sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C
+ a_68_1251# sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425#
Xsky130_fd_io__gpio_odrvr_subv2_0 VGND PD_H[0] PD_H[2] PD_H[1] PD_H[3] VCC_IO PAD
+ TIE_LO_ESD FORCE_HI_H_N FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3]
+ VSSIO_AMX VGND_IO TIE_HI_ESD sky130_fd_io__gpio_odrvr_subv2_0/w_n947_8961# sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_odrvr_subv2_0/m3_9047_13425# sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933#
+ sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263# sky130_fd_io__gpio_odrvr_subv2_0/m3_4600_13425#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425#
+ sky130_fd_io__gpio_odrvr_subv2
.ends

.subckt sky130_fd_io__gpio_opathv2 VGND HLD_I_H_N OD_H SLOW VCC_IO VPWR VPWR_KA PAD
+ TIE_HI_ESD VSSIO_AMX DM_H[0] DM_H[1] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2] HLD_I_OVR_H
+ OE_N OUT TIE_LO_ESD sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/w_n947_8961# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__com_opath_datoev2_0/w_n227_n1072#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ a_168_16482# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ m2_2157_n626# sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] m1_5007_14860# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ m1_4747_14860# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+
Xsky130_fd_io__gpiov2_octl_dat_0 VPWR VGND VCC_IO VPWR_KA SLOW HLD_I_H_N HLD_I_OVR_H
+ OD_H sky130_fd_io__gpiov2_octl_dat_0/SLOW_H_N sky130_fd_io__gpiov2_octl_dat_0/DRVHI_H
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1] sky130_fd_io__gpio_odrvrv2_0/PD_H[0]
+ sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] sky130_fd_io__gpiov2_octl_dat_0/DRVLO_H_N
+ DM_H_N[2] DM_H_N[0] DM_H[2] DM_H[1] DM_H[0] OUT OE_N DM_H_N[1] sky130_fd_io__gpio_odrvrv2_0/PD_H[3]
+ sky130_fd_io__gpio_odrvrv2_0/PD_H[2] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ VGND VGND sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__com_opath_datoev2_0/w_n227_n1072#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ sky130_fd_io__gpiov2_octl_dat
Xsky130_fd_io__gpio_odrvrv2_0 VGND PAD sky130_fd_io__gpio_odrvrv2_0/PD_H[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1]
+ sky130_fd_io__gpio_odrvrv2_0/PD_H[2] sky130_fd_io__gpio_odrvrv2_0/PD_H[3] TIE_LO_ESD
+ VCC_IO sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3] TIE_HI_ESD
+ VGND VSSIO_AMX VSSIO_AMX VSSIO_AMX VSSIO_AMX sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1]
+ sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/w_n947_8961# VGND
+ VGND VGND VGND sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] a_168_16482# VGND sky130_fd_io__gpio_odrvrv2
.ends

.subckt sky130_fd_io__amux_switch_1v2b AMUXBUS_HV PAD_HV_P0 PG_AMX_VDDA_H_N NG_AMX_VPMP_H
+ NG_PAD_VPMP_H PAD_HV_P1 PG_PAD_VDDIOQ_H_N PAD_HV_N0 PAD_HV_N1 VSSD VDDA PAD_HV_N2
+ VDDIO PAD_HV_N3 w_7097_435# w_4005_333#
X0 PAD_HV_N3 NG_PAD_VPMP_H w_7097_435# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X1 PAD_HV_P0 PG_PAD_VDDIOQ_H_N w_4005_333# VDDIO sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X2 AMUXBUS_HV NG_AMX_VPMP_H w_7097_435# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X3 PAD_HV_N1 NG_PAD_VPMP_H w_4005_333# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X4 w_4005_333# NG_PAD_VPMP_H PAD_HV_N0 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X5 AMUXBUS_HV NG_AMX_VPMP_H w_4005_333# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X6 w_7097_435# NG_PAD_VPMP_H PAD_HV_N2 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X7 w_4005_333# NG_PAD_VPMP_H PAD_HV_N0 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X8 w_7097_435# NG_PAD_VPMP_H PAD_HV_N3 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X9 w_4005_333# NG_AMX_VPMP_H AMUXBUS_HV VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X10 AMUXBUS_HV PG_AMX_VDDA_H_N w_4005_333# VDDA sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X11 w_7097_435# NG_PAD_VPMP_H PAD_HV_N2 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X12 w_4005_333# PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X13 PAD_HV_N2 NG_PAD_VPMP_H w_7097_435# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X14 AMUXBUS_HV NG_AMX_VPMP_H w_4005_333# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X15 PAD_HV_N0 NG_PAD_VPMP_H w_4005_333# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X16 AMUXBUS_HV NG_AMX_VPMP_H w_7097_435# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X17 w_7097_435# NG_AMX_VPMP_H AMUXBUS_HV VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X18 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_4005_333# VDDIO sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X19 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_4005_333# VDDIO sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X20 w_7097_435# NG_AMX_VPMP_H AMUXBUS_HV VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X21 AMUXBUS_HV NG_AMX_VPMP_H w_4005_333# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X22 w_4005_333# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X23 w_7097_435# NG_PAD_VPMP_H PAD_HV_N3 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X24 w_4005_333# NG_PAD_VPMP_H PAD_HV_N1 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X25 AMUXBUS_HV PG_AMX_VDDA_H_N w_4005_333# VDDA sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X26 w_7097_435# NG_AMX_VPMP_H AMUXBUS_HV VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X27 w_4005_333# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X28 AMUXBUS_HV NG_AMX_VPMP_H w_7097_435# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X29 PAD_HV_N2 NG_PAD_VPMP_H w_7097_435# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X30 PAD_HV_N3 NG_PAD_VPMP_H w_7097_435# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X31 w_4005_333# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X32 AMUXBUS_HV NG_AMX_VPMP_H w_4005_333# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X33 PAD_HV_N1 NG_PAD_VPMP_H w_4005_333# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X34 w_4005_333# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X35 w_4005_333# NG_AMX_VPMP_H AMUXBUS_HV VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X36 w_4005_333# NG_PAD_VPMP_H PAD_HV_N1 VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X37 w_7097_435# NG_AMX_VPMP_H AMUXBUS_HV VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
X38 w_4005_333# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 w=7e+06u l=500000u
X39 w_4005_333# NG_AMX_VPMP_H AMUXBUS_HV VSSD sky130_fd_pr__nfet_g5v0d10v5 w=7e+06u l=500000u
.ends

.subckt sky130_fd_io__res75only_small PAD ROUT VSUBS
R0 PAD ROUT sky130_fd_pr__res_generic_po w=2e+06u l=3.15e+06u
.ends

.subckt sky130_fd_io__gpiov2_amx_pucsd_inv VSSA VDA Y A VSUBS w_1_293#
X0 VDA A Y w_1_293# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 Y A VSSA VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X3 VDA A Y w_1_293# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X4 Y A VSSA VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X5 VSSA A Y VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X6 Y A VSSA VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X7 VSSA A Y VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X8 Y A VSSA VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X9 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X10 VDA A Y w_1_293# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X11 VSSA A Y VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X12 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X13 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_amx_inv4 A VDA VSSA Y VSUBS w_0_284#
X0 VDA A Y w_0_284# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 Y A VDA w_0_284# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 Y A VSSA VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
X3 VSSA A Y VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr_lshv2hv VPWR_HV IN VGND RST_H HLD_H_N IN_B
+ OUT_H_N a_n988_3146# w_n1543_3062# a_n1424_3030#
X0 a_472_123# IN_B a_n1424_3030# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X1 a_472_123# IN_B a_n1424_3030# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X2 a_472_123# IN a_n988_3146# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 a_n988_3146# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X4 VGND a_n1424_3030# OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X5 VPWR_HV a_n1424_3030# OUT_H_N w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X6 a_n1424_3030# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X7 VGND HLD_H_N a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X8 VPWR_HV a_n988_3146# a_n1424_3030# w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X9 a_n1424_3030# IN_B a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X10 a_n988_3146# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X11 OUT_H_N a_n1424_3030# VPWR_HV w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X12 a_n988_3146# a_n1424_3030# VPWR_HV w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr_ls VPWR_LV RST_H OUT_H_N IN IN_B HLD_H_N OUT_H
+ VGND VPWR_HV a_226_158# a_398_158#
X0 OUT_H RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_226_158# IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X2 a_594_584# VPWR_LV a_226_158# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X3 VPWR_HV OUT_H OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=700000u l=600000u
X4 a_398_158# IN VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X5 VGND IN_B a_226_158# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X6 VGND RST_H OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_398_158# VPWR_LV a_877_584# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X8 a_594_584# HLD_H_N OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_226_158# VPWR_LV a_594_584# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X10 OUT_H_N HLD_H_N a_877_584# VGND sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VGND IN a_398_158# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X12 OUT_H HLD_H_N a_594_584# VGND sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 a_877_584# HLD_H_N OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_877_584# VPWR_LV a_398_158# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X15 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr_lshv2hv2 VPWR_HV IN VGND RST_H HLD_H_N IN_B
+ OUT_H_N a_940_123# a_319_123#
X0 a_472_123# IN_B a_319_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X1 VPWR_HV a_319_123# a_940_123# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X2 a_472_123# IN_B a_319_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 a_472_123# IN a_940_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X4 VPWR_HV a_319_123# OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X5 a_940_123# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X6 VGND a_319_123# OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X7 a_319_123# a_940_123# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X8 a_319_123# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X9 VGND HLD_H_N a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X10 a_319_123# IN_B a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X11 a_940_123# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X12 OUT_H_N a_319_123# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
.ends

.subckt sky130_fd_io__amx_inv1 VSUBS w_0_316# a_119_10# a_66_36# a_219_36# a_66_382#
X0 a_219_36# a_119_10# a_66_382# w_0_316# sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_219_36# a_119_10# a_66_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr VSSD VDDIO_Q VSWITCH VCCD D_B NMIDA_VCCD_N
+ NMIDA_VCCD NGA_PAD_VSWITCH_H_N PD_CSD_VSWITCH_H_N NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H
+ PD_CSD_VSWITCH_H NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N AMUX_EN_VDDA_H_N
+ NMIDA_ON_N PU_ON_N PU_ON AMUX_EN_VDDIO_H AMUXBUSA_ON_N AMUXBUSA_ON AMUX_EN_VSWITCH_H_N
+ PGB_AMX_VDDA_H_N NGA_AMX_VSWITCH_H PD_ON_N VDDA AMUX_EN_VDDA_H AMUX_EN_VSWITCH_H
+ AMUXBUSB_ON PU_CSD_VDDIOQ_H_N AMUXBUSB_ON_N PD_ON PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N
+ PGA_AMX_VDDA_H_N m1_18386_n10924# sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158#
+ m1_17472_n6692# m2_16610_n11154# m1_23054_n9427# sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ m1_18834_n11156# m2_16276_n11768# li_22905_n10879# m1_17800_n11010# m1_16696_n12226#
+ m1_17457_n12126# m1_18272_n10845# sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158#
+ m2_16613_n11563# m1_17795_n11868# sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146#
+ m2_16478_n11164# sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N m1_18395_n10976# m2_16340_n11711#
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123# sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158#
+ m1_16576_n12293# m1_18095_n11662# sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N sky130_fd_io__gpiov2_amx_inv4_4/A
+ m1_23228_n10198# m1_16635_n11564# m1_17387_n10793# m1_17465_n10807# m2_16539_n11240#
+ m2_16539_n11154# m1_17797_n11059# m2_16610_n11236# sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ m1_19972_n11538# m1_17927_n11010# m2_17359_n12074# sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123#
+ m1_19532_n11662# m1_16789_n12170# sky130_fd_io__gpiov2_amx_inv4_2/A sky130_fd_io__gpiov2_amx_inv4_1/A
+ m1_17059_n11489# sky130_fd_io__hvsbt_inv_x2_1/IN m1_18759_n11083# m1_18222_n11662#
+ m2_27137_n11400# m1_22876_n9465# m1_18090_n11624# m1_18005_n10811# m1_18445_n10934#
+ m2_17856_n11844# m2_16473_n11654# m2_17903_n11844# m2_20939_n11919# m2_19572_n11610#
+ m1_17927_n10793# m1_19746_n11489# m1_18775_n11178# sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158#
+ m1_17928_n11059# m1_16691_n12255# sky130_fd_io__gpiov2_amx_pucsd_inv_0/A m1_17392_n6692#
+ m2_16539_n11002# m1_19616_n11489# sky130_fd_io__gpiov2_amx_inv4_5/A m1_18680_n11104#
+ m2_20007_n11486# m1_23401_n11569# m2_17426_n12074# m2_19532_n11610# m1_16633_n11615#
+ m2_20051_n11486# m2_16549_n11563# sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158#
+ m1_19990_n11490#
Xsky130_fd_io__gpiov2_amx_pucsd_inv_0 VSSD VDDIO_Q PU_CSD_VDDIOQ_H_N sky130_fd_io__gpiov2_amx_pucsd_inv_0/A
+ VSSD VDDIO_Q sky130_fd_io__gpiov2_amx_pucsd_inv
Xsky130_fd_io__gpiov2_amx_inv4_0 sky130_fd_io__gpiov2_amx_inv4_1/A VSWITCH VSSD NGB_PAD_VSWITCH_H
+ VSSD VSWITCH sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_1 sky130_fd_io__gpiov2_amx_inv4_1/A VSWITCH VSSD NGB_AMX_VSWITCH_H
+ VSSD VSWITCH sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_2 sky130_fd_io__gpiov2_amx_inv4_2/A VDDIO_Q VSSD PGB_PAD_VDDIOQ_H_N
+ VSSD VDDIO_Q sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_3 sky130_fd_io__gpiov2_amx_inv4_5/A VSWITCH VSSD NGA_PAD_VSWITCH_H
+ VSSD VSWITCH sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_4 sky130_fd_io__gpiov2_amx_inv4_4/A VDDIO_Q VSSD PGA_PAD_VDDIOQ_H_N
+ VSSD VDDIO_Q sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_5 sky130_fd_io__gpiov2_amx_inv4_5/A VSWITCH VSSD NGA_AMX_VSWITCH_H
+ VSSD VSWITCH sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amux_drvr_lshv2hv_0 VDDA sky130_fd_io__gpiov2_amx_inv4_4/A VSSD
+ AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N PGA_AMX_VDDA_H_N
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146# VDDA sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv
Xsky130_fd_io__hvsbt_inv_x2_0 VCCD VSSD NMIDA_ON_N NMIDA_VCCD VSSD VCCD sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_inv_x2_1 VCCD VSSD sky130_fd_io__hvsbt_inv_x2_1/IN D_B VSSD VCCD
+ sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__gpiov2_amux_drvr_ls_0 VCCD AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amx_inv4_1/A
+ AMUXBUSB_ON AMUXBUSB_ON_N AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_0/OUT_H
+ VSSD VSWITCH sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158# sky130_fd_io__gpiov2_amux_drvr_ls_0/a_398_158#
+ sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0 VDDA sky130_fd_io__gpiov2_amx_inv4_2/A
+ VSSD AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ PGB_AMX_VDDA_H_N sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123# sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123#
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv2
Xsky130_fd_io__gpiov2_amux_drvr_ls_1 VCCD AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ AMUXBUSB_ON AMUXBUSB_ON_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amx_inv4_2/A VSSD
+ VDDIO_Q sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158# sky130_fd_io__gpiov2_amux_drvr_ls_1/a_398_158#
+ sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_2 VCCD AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ PD_ON PD_ON_N AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H VSSD VSWITCH
+ sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158# sky130_fd_io__gpiov2_amux_drvr_ls_2/a_398_158#
+ sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_3 VCCD AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amx_inv4_5/A
+ AMUXBUSA_ON AMUXBUSA_ON_N AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_3/OUT_H
+ VSSD VSWITCH sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158# sky130_fd_io__gpiov2_amux_drvr_ls_3/a_398_158#
+ sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_5 VCCD AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_ls_5/OUT_H_N
+ PU_ON PU_ON_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amx_pucsd_inv_0/A VSSD VDDIO_Q
+ sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158# sky130_fd_io__gpiov2_amux_drvr_ls_5/a_398_158#
+ sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_4 VCCD AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N
+ AMUXBUSA_ON AMUXBUSA_ON_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amx_inv4_4/A VSSD
+ VDDIO_Q m1_16788_n13135# m1_16634_n13346# sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__amx_inv1_0 VSSD VSWITCH PD_CSD_VSWITCH_H VSSD PD_CSD_VSWITCH_H_N VSWITCH
+ sky130_fd_io__amx_inv1
Xsky130_fd_io__amx_inv1_1 VSSD VSWITCH NGB_PAD_VSWITCH_H VSSD NGB_PAD_VSWITCH_H_N
+ VSWITCH sky130_fd_io__amx_inv1
Xsky130_fd_io__amx_inv1_2 VSSD VSWITCH NGA_PAD_VSWITCH_H VSSD NGA_PAD_VSWITCH_H_N
+ VSWITCH sky130_fd_io__amx_inv1
Xsky130_fd_io__hvsbt_inv_x1_0 NMIDA_VCCD_N VCCD VSSD VSSD NMIDA_VCCD VCCD sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 D_B VCCD VSSD VSSD D_B VCCD sky130_fd_io__hvsbt_inv_x1
X0 PD_CSD_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 NGB_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X2 PD_CSD_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=2e+06u
X3 NGA_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X4 PD_CSD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X5 VSSD AMUX_EN_VDDA_H_N NGA_AMX_VSWITCH_H VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X6 VSSD VSSD PD_CSD_VSWITCH_H VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 VSWITCH sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N PD_CSD_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=2e+06u
X8 VSSD AMUX_EN_VDDIO_H_N NGB_PAD_VSWITCH_H VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_amux_nand5 OUT VPWR VGND IN1 IN0 IN3 IN2 IN4
X0 a_59_1018# OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 OUT a_59_1018# VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_59_1018# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR IN0 OUT VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X4 a_386_228# IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X5 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X6 a_698_228# IN3 a_542_228# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X7 VPWR OUT a_59_1018# VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X8 a_542_228# IN4 a_386_228# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X9 a_854_228# IN2 a_698_228# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X10 VGND OUT a_59_1018# VGND sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 OUT IN1 a_854_228# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
.ends

.subckt sky130_fd_io__inv_1 VNB VPB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends

.subckt sky130_fd_io__xor2_1 VNB VPB VPWR VGND A B X
X0 a_42_367# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND a_42_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR B a_293_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 X B a_297_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_293_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_125_367# B a_42_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND A a_42_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_297_69# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR A a_125_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_293_367# a_42_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends

.subckt sky130_fd_io__nor2_1 VNB VPB VPWR VGND B Y A
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 Y B a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends

.subckt sky130_fd_io__gpiov2_amux_nand4 OUT VPWR VGND IN1 IN0 IN3 IN2
X0 VPWR IN0 OUT VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 VPWR OUT a_59_1018# VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 VGND a_59_1018# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X4 a_386_228# IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X5 a_698_228# IN2 a_542_228# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X6 a_542_228# IN3 a_386_228# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X7 OUT IN1 a_698_228# VGND sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X8 a_59_1018# OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X9 VGND OUT a_59_1018# VGND sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 OUT a_59_1018# VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
.ends

.subckt sky130_fd_io__nand2_1 VNB VPB VPWR VGND B Y A
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X2 Y A a_117_74# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_117_74# B VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends

.subckt sky130_fd_io__gpiov2_amux_decoder NMIDA_ON_N D_B PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N
+ PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N PD_ON PD_ON_N PU_ON PU_ON_N AMUXBUSB_ON AMUXBUSB_ON_N
+ OUT ANALOG_EN ANALOG_POL ANALOG_SEL AMUXBUSA_ON AMUXBUSA_ON_N VSSD VCCD NGB_PAD_VSWITCH_H
+ NGA_PAD_VSWITCH_H NGA_PAD_VSWITCH_H_N NGB_PAD_VSWITCH_H_N NMIDA_VCCD_N PU_VDDIOQ_H_N
+ PD_VSWITCH_H_N sky130_fd_io__inv_1_14/Y sky130_fd_io__hvsbt_nand2_3/OUT sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_2/Y sky130_fd_io__hvsbt_nand2_0/IN1
+ sky130_fd_io__hvsbt_nand2_1/IN1 sky130_fd_io__xor2_1_0/A sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__inv_1_3/Y sky130_fd_io__nor2_1_2/B sky130_fd_io__nor2_1_1/Y sky130_fd_io__hvsbt_nand2_2/OUT
+ sky130_fd_io__inv_1_7/A sky130_fd_io__inv_1_2/A sky130_fd_io__gpiov2_amux_nand4_0/OUT
+ sky130_fd_io__gpiov2_amux_nand5_1/IN0 sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_nand5_0/IN0
+ sky130_fd_io__xor2_1_0/X
Xsky130_fd_io__gpiov2_amux_nand5_0 sky130_fd_io__inv_1_7/A VCCD VSSD PGA_PAD_VDDIOQ_H_N
+ sky130_fd_io__gpiov2_amux_nand5_0/IN0 NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N NGB_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_nand5
Xsky130_fd_io__gpiov2_amux_nand5_1 sky130_fd_io__inv_1_5/A VCCD VSSD PGA_PAD_VDDIOQ_H_N
+ sky130_fd_io__gpiov2_amux_nand5_1/IN0 NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N NGB_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_nand5
Xsky130_fd_io__inv_1_10 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_11/A ANALOG_POL sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_11 VSSD VCCD VCCD VSSD sky130_fd_io__xor2_1_0/A sky130_fd_io__inv_1_11/A
+ sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nor_0 NGA_PAD_VSWITCH_H VSSD VCCD VSSD VCCD sky130_fd_io__hvsbt_nand2_3/OUT
+ sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nor_1 NGB_PAD_VSWITCH_H VSSD VCCD VSSD VCCD sky130_fd_io__hvsbt_nand2_2/OUT
+ sky130_fd_io__hvsbt_nand2_1/IN1 sky130_fd_io__hvsbt_nor
Xsky130_fd_io__xor2_1_0 VSSD VCCD VCCD VSSD sky130_fd_io__xor2_1_0/A sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__xor2_1_0/X sky130_fd_io__xor2_1
Xsky130_fd_io__inv_1_13 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_13/Y ANALOG_SEL sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_12 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_14 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_14/Y sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__inv_1_14/Y
+ NMIDA_ON_N VSSD VCCD VSSD VCCD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_0 VSSD VCCD VCCD VSSD PD_ON_N PD_ON sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nand2_1 sky130_fd_io__hvsbt_nand2_1/IN1 sky130_fd_io__inv_1_2/Y
+ D_B VSSD VCCD VSSD VCCD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_2 PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N sky130_fd_io__hvsbt_nand2_2/OUT
+ VSSD VCCD VSSD VCCD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_1 VSSD VCCD VCCD VSSD PU_ON_N PU_ON sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_2 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_2/Y sky130_fd_io__inv_1_2/A
+ sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_3 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_3/Y sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nand2_3 PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__hvsbt_nand2_3/OUT
+ VSSD VCCD VSSD VCCD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_4 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_4/Y OUT sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_5 VSSD VCCD VCCD VSSD PU_ON sky130_fd_io__inv_1_5/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_6 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_6/Y ANALOG_EN sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_0 VSSD VCCD VCCD VSSD sky130_fd_io__nor2_1_0/B sky130_fd_io__inv_1_2/A
+ sky130_fd_io__inv_1_6/Y sky130_fd_io__nor2_1
Xsky130_fd_io__gpiov2_amux_nand4_0 sky130_fd_io__gpiov2_amux_nand4_0/OUT VCCD VSSD
+ PU_VDDIOQ_H_N sky130_fd_io__nor2_1_2/Y NMIDA_VCCD_N PD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_nand4
Xsky130_fd_io__inv_1_7 VSSD VCCD VCCD VSSD PD_ON sky130_fd_io__inv_1_7/A sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_2 VSSD VCCD VCCD VSSD sky130_fd_io__nor2_1_2/B sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__inv_1_6/Y sky130_fd_io__nor2_1
Xsky130_fd_io__nor2_1_1 VSSD VCCD VCCD VSSD sky130_fd_io__nor2_1_1/B sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__inv_1_6/Y sky130_fd_io__nor2_1
Xsky130_fd_io__gpiov2_amux_nand4_1 AMUXBUSB_ON_N VCCD VSSD PU_VDDIOQ_H_N sky130_fd_io__inv_1_2/A
+ D_B PD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_nand4
Xsky130_fd_io__nor2_1_3 VSSD VCCD VCCD VSSD sky130_fd_io__nor2_1_3/B sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__inv_1_6/Y sky130_fd_io__nor2_1
Xsky130_fd_io__inv_1_8 VSSD VCCD VCCD VSSD AMUXBUSA_ON AMUXBUSA_ON_N sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_9 VSSD VCCD VCCD VSSD AMUXBUSB_ON AMUXBUSB_ON_N sky130_fd_io__inv_1
Xsky130_fd_io__nand2_1_0 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_12/Y sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__xor2_1_0/X sky130_fd_io__nand2_1
* Xsky130_fd_io__tap_1_0 VSSD VCCD VCCD VSSD sky130_fd_io__tap_1
Xsky130_fd_io__nand2_1_1 VSSD VCCD VCCD VSSD sky130_fd_io__xor2_1_0/X sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__inv_1_13/Y sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_2 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_4/Y sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__inv_1_11/A sky130_fd_io__nand2_1
* Xsky130_fd_io__tap_1_1 VSSD VCCD VCCD VSSD sky130_fd_io__tap_1
* Xsky130_fd_io__tap_1_2 VSSD VCCD VCCD VSSD sky130_fd_io__tap_1
Xsky130_fd_io__nand2_1_3 VSSD VCCD VCCD VSSD sky130_fd_io__inv_1_3/Y sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__xor2_1_0/A sky130_fd_io__nand2_1
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_ls IN_B OUT_H_N OUT_H VPWR_HV VGND HLD_H_N RST_H
+ IN VPWR_LV
X0 VGND HLD_H_N a_209_617# VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X1 a_292_617# VPWR_LV a_331_899# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X2 a_141_899# VPWR_LV a_636_617# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X3 a_636_617# VPWR_LV a_141_899# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X4 a_292_617# VPWR_LV a_331_899# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X5 a_331_899# VPWR_LV a_292_617# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X6 a_292_617# IN a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X7 a_209_617# IN a_292_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X8 a_209_617# HLD_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X9 VGND a_331_899# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X10 a_636_617# VPWR_LV a_141_899# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X11 a_636_617# IN_B a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X12 a_141_899# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X13 VPWR_HV a_141_899# OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_292_617# IN a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X15 a_209_617# IN_B a_636_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X16 a_141_899# VPWR_LV a_636_617# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X17 a_141_899# a_331_899# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 a_331_899# a_141_899# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X19 OUT_H_N a_141_899# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X20 VGND HLD_H_N a_209_617# VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X21 a_331_899# VPWR_LV a_292_617# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X22 OUT_H a_331_899# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X23 a_636_617# IN_B a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X24 a_209_617# IN_B a_636_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X25 a_209_617# HLD_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X26 a_209_617# IN a_292_617# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_inv_1 VNB VPB VPWR VGND OUT IN
X0 OUT IN VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 OUT IN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_lshv2hv IN_B IN RST_H OUT_H_N OUT_H VPWR_HV
+ HLD_H VGND a_3512_651# a_4133_651#
X0 a_3665_651# IN_B a_3512_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X1 a_3665_651# IN_B a_3512_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X2 a_3512_651# IN_B a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 a_4133_651# a_3512_651# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X4 VPWR_HV a_4133_651# OUT_H VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X5 VPWR_HV a_4133_651# a_3512_651# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X6 OUT_H_N a_3512_651# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_3665_651# IN a_4133_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X8 VGND HLD_H a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X9 VGND RST_H a_3512_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X10 a_4133_651# IN a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X11 OUT_H a_4133_651# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X12 a_4133_651# IN a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X13 OUT_H_N a_3512_651# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_lshv2hv2 IN_B IN RST_H OUT_H_N OUT_H VPWR_HV
+ HLD_H VGND VSUBS li_1122_1924# a_391_3019# a_693_2921# a_291_2921# a_425_1501# w_467_555#
X0 OUT_H a_425_665# VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X1 a_391_3019# a_291_2921# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_578_665# IN_B a_693_2921# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 a_578_665# IN a_425_665# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X4 a_425_665# IN a_578_665# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X5 a_391_3019# a_291_2921# a_425_1501# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X6 a_693_2921# a_425_665# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X7 a_693_2921# IN_B a_578_665# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X8 VGND a_693_2921# OUT_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X9 a_693_2921# RST_H VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=500000u
X10 VPWR_HV a_693_2921# OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VPWR_HV a_291_2921# a_391_3019# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 OUT_H a_425_665# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X13 a_578_665# IN a_425_665# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X14 VGND HLD_H a_578_665# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X15 VPWR_HV a_693_2921# a_425_665# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X16 a_693_2921# IN_B a_578_665# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_amux_ls ANALOG_EN HLD_I_H HLD_I_H_N VDDIO_Q VSWITCH AMUX_EN_VSWITCH_H
+ AMUX_EN_VDDA_H_N VSSD AMUX_EN_VSWITCH_H_N ENABLE_VSWITCH_H AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H
+ AMUX_EN_VDDA_H ENABLE_VDDA_H VDDA VCCD sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_3512_651#
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/w_467_555# sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921# sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/li_1122_1924#
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_4133_651#
+ sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N w_1167_10569#
Xsky130_fd_io__gpiov2_amux_ctl_ls_0 sky130_fd_io__gpiov2_amux_ctl_ls_0/IN_B sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N
+ AMUX_EN_VDDIO_H VDDIO_Q VSSD HLD_I_H_N HLD_I_H sky130_fd_io__gpiov2_amux_ctl_ls_0/IN
+ VCCD sky130_fd_io__gpiov2_amux_ctl_ls
Xsky130_fd_io__gpiov2_amux_ctl_inv_1_0 VSSD VCCD VCCD VSSD sky130_fd_io__gpiov2_amux_ctl_ls_0/IN
+ sky130_fd_io__gpiov2_amux_ctl_ls_0/IN_B sky130_fd_io__gpiov2_amux_ctl_inv_1
Xsky130_fd_io__gpiov2_amux_ctl_inv_1_1 VSSD VCCD VCCD VSSD sky130_fd_io__gpiov2_amux_ctl_ls_0/IN_B
+ ANALOG_EN sky130_fd_io__gpiov2_amux_ctl_inv_1
Xsky130_fd_io__gpiov2_amux_ctl_lshv2hv_0 AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ AMUX_EN_VSWITCH_H_N AMUX_EN_VSWITCH_H VSWITCH ENABLE_VSWITCH_H VSSD sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_3512_651#
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_4133_651# sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xsky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0 AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H VDDA ENABLE_VDDA_H VSSD VSSD sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/li_1122_1924#
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921#
+ ENABLE_VDDA_H VSSD sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/w_467_555# sky130_fd_io__gpiov2_amux_ctl_lshv2hv2
* Xsky130_fd_io__tap_1_0 VSSD VCCD VCCD VSSD sky130_fd_io__tap_1
X0 VSWITCH ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H w_1167_10569# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 VSSD ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H VSSD sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X2 sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H ENABLE_VSWITCH_H VSWITCH w_1167_10569# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_logic ANALOG_EN NMIDA_VCCD D_B PD_CSD_VSWITCH_H
+ NGB_AMX_VSWITCH_H NGA_AMX_VSWITCH_H NGB_PAD_VSWITCH_H NGA_PAD_VSWITCH_H PGB_AMX_VDDA_H_N
+ PGA_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N PU_CSD_VDDIOQ_H_N OUT ANALOG_SEL
+ ANALOG_POL VSSD HLD_I_H_N HLD_I_H ENABLE_VSWITCH_H ENABLE_VDDA_H AMUX_EN_VDDIO_H_N
+ AMUX_EN_VDDA_H_N VCCD VDDA VDDIO_Q VSWITCH sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_3/OUT sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_4/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N
+ m1_31532_n4418# sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123#
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N sky130_fd_io__gpiov2_amux_drvr_0/PGB_AMX_VDDA_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_5/A sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON
+ sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_2/OUT
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/A m2_37354_n6053# sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_0/IN1
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/PU_ON sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123#
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_pucsd_inv_0/A sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_0/m2_27137_n11400# sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_2/A
+ w_28088_n3500# sky130_fd_io__gpiov2_amux_drvr_0/PD_ON sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158#
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146#
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158#
+ m1_31532_n4477# sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921#
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158#
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/X
Xsky130_fd_io__gpiov2_amux_drvr_0 VSSD VDDIO_Q VSWITCH VCCD D_B sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N
+ NMIDA_VCCD sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H PD_CSD_VSWITCH_H
+ NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N AMUX_EN_VDDA_H_N sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N sky130_fd_io__gpiov2_amux_drvr_0/PU_ON
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/PGB_AMX_VDDA_H_N NGA_AMX_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N
+ VDDA sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDA_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON PU_CSD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/PD_ON PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N PGA_AMX_VDDA_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934# sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158#
+ VSWITCH sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ D_B sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158#
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146#
+ ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934# sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123#
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158#
+ sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_4/A
+ sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ VSWITCH VSWITCH sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_2/A sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_1/A
+ AMUX_EN_VDDIO_H_N D_B sky130_fd_io__gpiov2_amux_drvr_0/m1_18759_n11083# sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H
+ sky130_fd_io__gpiov2_amux_drvr_0/m2_27137_n11400# NGA_PAD_VSWITCH_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H
+ VSWITCH sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934# sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H VSWITCH AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_pucsd_inv_0/A VSWITCH
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H AMUX_EN_VDDIO_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_5/A sky130_fd_io__gpiov2_amux_drvr_0/m1_18759_n11083#
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158#
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr
Xsky130_fd_io__gpiov2_amux_decoder_0 sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N D_B
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_drvr_0/PD_ON
+ sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N sky130_fd_io__gpiov2_amux_drvr_0/PU_ON
+ sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N OUT ANALOG_EN ANALOG_POL ANALOG_SEL
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ VSSD VCCD NGB_PAD_VSWITCH_H NGA_PAD_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N
+ PU_CSD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_3/OUT sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_2/OUT
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/X sky130_fd_io__gpiov2_amux_decoder
Xsky130_fd_io__gpiov2_amux_ls_0 ANALOG_EN HLD_I_H HLD_I_H_N VDDIO_Q VSWITCH sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ AMUX_EN_VDDA_H_N VSSD sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N ENABLE_VSWITCH_H
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDA_H
+ ENABLE_VDDA_H VDDA VCCD sky130_fd_io__gpiov2_amux_drvr_0/m1_18759_n11083# VSSD sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921#
+ VSWITCH sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934# sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N
+ VSWITCH sky130_fd_io__gpiov2_amux_ls
.ends

.subckt sky130_fd_io__gpiov2_amux PAD AMUXBUS_B AMUXBUS_A VDDIO_Q VSSD VCCD VDDA VSSIO_Q
+ OUT HLD_I_H_N HLD_I_H ENABLE_VSWITCH_H ENABLE_VDDA_H ANALOG_SEL ANALOG_POL ANALOG_EN
+ VSWITCH w_n874_6088# a_14152_3009#
Xsky130_fd_io__amux_switch_1v2b_0 AMUXBUS_A sky130_fd_io__res75only_small_13/ROUT
+ sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H sky130_fd_io__res75only_small_0/ROUT
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__res75only_small_3/ROUT VSSD VDDA sky130_fd_io__res75only_small_10/ROUT
+ VDDIO_Q sky130_fd_io__res75only_small_10/ROUT a_13552_3035# m1_8800_6769# sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__amux_switch_1v2b_1 AMUXBUS_B sky130_fd_io__res75only_small_13/ROUT
+ sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H sky130_fd_io__res75only_small_0/ROUT
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__res75only_small_3/ROUT VSSD VDDA sky130_fd_io__res75only_small_10/ROUT
+ VDDIO_Q sky130_fd_io__res75only_small_10/ROUT a_13975_3415# m1_8800_4647# sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__res75only_small_10 sky130_fd_io__res75only_small_10/PAD sky130_fd_io__res75only_small_10/ROUT
+ VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_11 PAD sky130_fd_io__res75only_small_10/PAD VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_13 PAD sky130_fd_io__res75only_small_13/ROUT VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_12 PAD PAD VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_0 PAD sky130_fd_io__res75only_small_0/ROUT VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 PAD sky130_fd_io__res75only_small_3/PAD VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 PAD PAD VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD sky130_fd_io__res75only_small_3/ROUT
+ VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_4 PAD sky130_fd_io__res75only_small_4/ROUT VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_amux_ctl_logic_0 ANALOG_EN sky130_fd_io__gpiov2_amux_ctl_logic_0/NMIDA_VCCD
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/D_B sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H
+ sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N OUT ANALOG_SEL ANALOG_POL
+ VSSD HLD_I_H_N HLD_I_H ENABLE_VSWITCH_H ENABLE_VDDA_H sky130_fd_io__gpiov2_amux_ctl_logic_0/AMUX_EN_VDDIO_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/AMUX_EN_VDDA_H_N VCCD VDDA VDDIO_Q VSWITCH
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_3/OUT
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H
+ m1_1514_5549# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_4/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N m1_415_8073# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_5/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_2/OUT
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/A
+ VCCD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_0/IN1
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PU_ON m1_515_8136#
+ m1_10523_333# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_pucsd_inv_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N
+ m1_n206_2973# VSSD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_2/A
+ m1_1260_3234# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PD_ON
+ m1_2332_3812# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ m2_405_5685# m1_8066_354# sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N m1_71_5381#
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ m1_n212_3842# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/X
+ sky130_fd_io__gpiov2_amux_ctl_logic
Xsky130_fd_io__res75only_small_5 PAD sky130_fd_io__res75only_small_5/ROUT VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_6 VSSD sky130_fd_io__res75only_small_6/ROUT VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_7 VSSD sky130_fd_io__res75only_small_7/ROUT VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_8 VSSD sky130_fd_io__res75only_small_8/ROUT VSSD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_9 VSSD sky130_fd_io__res75only_small_9/ROUT VSSD sky130_fd_io__res75only_small
X0 VSSD a_14152_3009# m1_8800_6769# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X2 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X3 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_4/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X4 VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N sky130_fd_io__res75only_small_4/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+07u l=500000u
X5 VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+07u l=500000u
X6 VSSD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H m1_8800_4647# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VSSD a_14152_3009# a_13975_3415# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X9 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+07u l=500000u
X10 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X11 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+07u l=500000u
X12 a_13552_3035# sky130_fd_io__gpiov2_amux_ctl_logic_0/NMIDA_VCCD sky130_fd_io__res75only_small_9/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X13 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_4/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X14 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X15 a_13552_3035# a_14152_3009# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 m1_8800_4647# a_14152_3009# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X18 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X19 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X20 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+07u l=500000u
X21 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X22 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X23 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+07u l=500000u
X24 m1_8800_6769# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 sky130_fd_io__res75only_small_8/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/NMIDA_VCCD m1_8800_6769# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X26 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X27 a_13975_3415# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 a_13975_3415# sky130_fd_io__gpiov2_amux_ctl_logic_0/D_B sky130_fd_io__res75only_small_7/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X29 VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+07u l=500000u
X30 m1_8800_4647# sky130_fd_io__gpiov2_amux_ctl_logic_0/D_B sky130_fd_io__res75only_small_6/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X31 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_4/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X32 VSSD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H a_13552_3035# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_ipath_hvls OUT OUT_B MODE_NORMAL_N IN_VCCHIB INB_VCCHIB
+ IN_VDDIO MODE_VCCHIB_N MODE_NORMAL MODE_VCCHIB VDDIO_Q VSSD
X0 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X1 OUT_B IN_VDDIO a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X2 OUT_B IN_VDDIO a_1752_2267# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X4 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X5 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X6 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X7 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X8 VDDIO_Q MODE_VCCHIB_N a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X9 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X10 VDDIO_Q a_621_2778# a_602_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 VDDIO_Q MODE_NORMAL_N a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X12 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X13 a_1175_2172# a_602_2876# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 a_1752_1955# a_1175_2172# OUT_B VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X15 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X16 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X17 OUT_B a_1175_2172# a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X18 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X19 a_1175_2172# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X20 a_2911_2876# MODE_VCCHIB OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X21 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X22 a_2024_2876# IN_VDDIO OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X23 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X24 a_621_2778# MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X25 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X26 a_1290_2876# MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X27 a_621_2778# INB_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X28 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X29 a_1290_2876# a_1175_2172# OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X30 VDDIO_Q MODE_NORMAL a_2911_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X31 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X32 a_621_2778# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X33 a_2024_2876# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X34 a_1930_201# IN_VCCHIB a_602_2876# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X35 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X36 a_1752_2267# MODE_NORMAL VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X37 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X38 VSSD MODE_VCCHIB a_1752_1955# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X39 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X40 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
.ends

.subckt sky130_fd_io__gpiov2_vcchib_in_buf IN_H MODE_VCCHIB_LV_N VCCHIB VSSD OUT OUT_N
X0 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X1 a_538_595# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
X2 a_538_595# a_591_563# a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X3 a_591_563# IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X4 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X5 a_751_595# IN_H a_591_563# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X6 a_446_3055# a_591_563# VSSD VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X7 VCCHIB MODE_VCCHIB_LV_N a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X8 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X9 VSSD IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X10 OUT OUT_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
X11 VSSD a_446_3055# OUT_N VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X12 VSSD MODE_VCCHIB_LV_N a_446_3055# VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X13 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X14 a_612_3332# a_591_563# a_446_3055# VCCHIB sky130_fd_pr__pfet_01v8 w=1e+06u l=250000u
X15 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
X16 a_446_3055# MODE_VCCHIB_LV_N VSSD VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X17 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
X18 a_751_595# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X19 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X20 VSSD a_591_563# a_446_3055# VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X21 a_612_2476# IN_H a_591_563# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=800000u
X22 VCCHIB a_446_3055# OUT_N VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
X23 a_591_563# IN_H a_612_2476# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=800000u
X24 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X25 a_446_3055# a_591_563# a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 w=1e+06u l=250000u
X26 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X27 a_612_2476# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
.ends

.subckt sky130_fd_io__gpiov2_in_buf OUT OUT_N MODE_NORMAL_N_uq1 IN_H IN_VT VTRIP_SEL_H
+ VTRIP_SEL_H_N VDDIO_Q VSSD m1_n467_n748#
Xsky130_fd_io__hvsbt_nor_0 VTRIP_SEL_H VSSD VDDIO_Q VSSD VDDIO_Q MODE_NORMAL_N_uq1
+ li_3458_2405# sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO_Q VSSD VSSD li_3458_2405#
+ VDDIO_Q sky130_fd_io__hvsbt_inv_x1
X0 VDDIO_Q MODE_NORMAL_N_uq1 a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X1 OUT OUT_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X2 VSSD a_36_n802# a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X3 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X4 VDDIO_Q sky130_fd_io__hvsbt_inv_x1_0/OUT a_1761_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X5 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X6 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X7 a_2073_1865# MODE_NORMAL_N_uq1 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X8 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X9 VSSD a_2651_1865# OUT_N VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X10 a_917_1865# IN_H a_36_n802# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=800000u
X11 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X12 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X13 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X14 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=500000u
X15 VDDIO_Q sky130_fd_io__hvsbt_inv_x1_0/OUT a_917_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X16 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X17 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=800000u
X18 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X19 a_1761_1865# sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X20 VSSD VTRIP_SEL_H_N IN_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=1e+06u
X21 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X22 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X23 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X24 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X25 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X26 VSSD MODE_NORMAL_N_uq1 a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X27 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X28 a_2651_1865# a_36_n802# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X29 VDDIO_Q MODE_NORMAL_N_uq1 a_2073_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X30 VSSD IN_VT a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X31 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X32 a_2651_1865# a_36_n802# a_2385_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=500000u
X33 a_2385_1865# MODE_NORMAL_N_uq1 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X34 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X35 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X36 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X37 a_917_1865# sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X38 a_219_1865# MODE_NORMAL_N_uq1 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X39 VDDIO_Q a_2651_1865# OUT_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X40 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=800000u
X41 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=5e+06u l=800000u
X42 a_2651_1865# MODE_NORMAL_N_uq1 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=500000u
X43 a_36_n802# IN_H a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=800000u
.ends

.subckt sky130_fd_io__gpiov2_ipath_lvls IN_VCCHIB IN_VDDIO MODE_NORMAL_LV MODE_NORMAL_LV_N
+ MODE_VCCHIB_LV MODE_VCCHIB_LV_N VCCHIB VSSD OUT OUT_B a_323_2354#
X0 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X1 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X2 a_1504_2754# IN_VCCHIB OUT_B VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X3 OUT_B a_323_2354# a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X4 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X5 VSSD MODE_NORMAL_LV a_316_n17# VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X6 VCCHIB IN_VDDIO a_114_2354# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X7 a_323_2354# a_114_2354# VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
X8 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X9 VCCHIB MODE_VCCHIB_LV_N a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X10 a_114_2354# IN_VDDIO VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 w=5e+06u l=500000u
X11 a_1679_n317# IN_VCCHIB OUT_B VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X12 a_436_2754# a_323_2354# OUT_B VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X13 VSSD MODE_NORMAL_LV a_823_n317# VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X14 OUT_B IN_VCCHIB a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X15 OUT_B a_323_2354# a_823_n317# VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X16 a_1679_n317# MODE_VCCHIB_LV VSSD VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X17 a_436_2754# MODE_NORMAL_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X18 a_323_2354# a_114_2354# VSSD VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X19 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X20 VCCHIB MODE_NORMAL_LV_N a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X21 OUT_B IN_VCCHIB a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X22 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X23 a_1504_2754# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X24 VCCHIB MODE_VCCHIB_LV a_2141_2754# VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X25 VSSD MODE_VCCHIB_LV a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X26 a_2141_2754# MODE_NORMAL_LV OUT_B VCCHIB sky130_fd_pr__pfet_01v8 w=3e+06u l=250000u
X27 a_823_n317# MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
X28 VCCHIB MODE_NORMAL_LV a_114_2354# VCCHIB sky130_fd_pr__pfet_01v8 w=5e+06u l=250000u
X29 a_316_n17# IN_VDDIO a_114_2354# VSSD sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X30 a_823_n317# a_323_2354# OUT_B VSSD sky130_fd_pr__nfet_01v8 w=3e+06u l=250000u
.ends

.subckt sky130_fd_io__gpiov2_inbuf_lvinv_x1 IN VGND VPWR OUT
X0 VPWR IN OUT VPWR sky130_fd_pr__pfet_01v8_hvt w=3e+06u l=250000u
X1 VGND IN OUT VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
.ends

.subckt sky130_fd_io__gpiov2_ibuf_se VTRIP_SEL_H_N VCCHIB ENABLE_VDDIO_LV MODE_NORMAL_N
+ VSSD VDDIO_Q IBUFMUX_OUT IN_VT IN_H VTRIP_SEL_H MODE_VCCHIB_N IBUFMUX_OUT_H sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354#
+ sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
Xsky130_fd_io__gpiov2_ipath_hvls_0 IBUFMUX_OUT_H sky130_fd_io__gpiov2_ipath_hvls_0/OUT_B
+ MODE_NORMAL_N sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N
+ sky130_fd_io__gpiov2_in_buf_0/OUT MODE_VCCHIB_N sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__hvsbt_nand2_0/IN1 VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_hvls
Xsky130_fd_io__gpiov2_vcchib_in_buf_0 IN_H sky130_fd_io__hvsbt_nand2_0/OUT VCCHIB
+ VSSD sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N
+ sky130_fd_io__gpiov2_vcchib_in_buf
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 ENABLE_VDDIO_LV sky130_fd_io__hvsbt_nand2_0/OUT
+ VSSD VCCHIB VSSD VCCHIB sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_1 sky130_fd_io__hvsbt_nand2_1/IN1 ENABLE_VDDIO_LV sky130_fd_io__hvsbt_nand2_1/OUT
+ VSSD VCCHIB VSSD VCCHIB sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__gpiov2_in_buf_0 sky130_fd_io__gpiov2_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT_N
+ MODE_NORMAL_N IN_H IN_VT VTRIP_SEL_H VTRIP_SEL_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
+ sky130_fd_io__gpiov2_in_buf
Xsky130_fd_io__gpiov2_ipath_lvls_0 sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT sky130_fd_io__hvsbt_nand2_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT
+ sky130_fd_io__hvsbt_nand2_0/OUT VCCHIB VSSD IBUFMUX_OUT sky130_fd_io__gpiov2_ipath_lvls_0/OUT_B
+ sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354# sky130_fd_io__gpiov2_ipath_lvls
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_0 sky130_fd_io__hvsbt_nand2_1/OUT VSSD VCCHIB
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_1 sky130_fd_io__hvsbt_nand2_0/OUT VSSD VCCHIB
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_nand2_0/IN1 VDDIO_Q VSSD VSSD MODE_VCCHIB_N
+ VDDIO_Q sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_nand2_1/IN1 VDDIO_Q VSSD VSSD MODE_NORMAL_N
+ VDDIO_Q sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__hvsbt_nand2v2 IN1 IN0 OUT VGND VPWR VSUBS w_n34_415#
X0 OUT IN0 VPWR w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 VPWR IN1 OUT w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 OUT IN0 VPWR w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 OUT IN1 a_239_144# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X4 VPWR IN1 OUT w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X5 a_239_144# IN0 VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_ictl_logic INP_DIS_I_H_N INP_DIS_I_H INP_DIS_H_N DM_H_N[2]
+ DM_H_N[1] DM_H_N[0] IB_MODE_SEL_H_N VDDIO_Q VSSD VTRIP_SEL_H_N MODE_NORMAL_N MODE_VCCHIB_N
+ TRIPSEL_I_H TRIPSEL_I_H_N IB_MODE_SEL_H
Xsky130_fd_io__hvsbt_nand2v2_0 DM_H_N[0] DM_H_N[1] sky130_fd_io__hvsbt_nand2v2_0/OUT
+ VSSD VDDIO_Q VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2v2
Xsky130_fd_io__hvsbt_nor_0 VTRIP_SEL_H_N VSSD VDDIO_Q VSSD VDDIO_Q MODE_NORMAL_N TRIPSEL_I_H
+ sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nand2_0 IB_MODE_SEL_H INP_DIS_I_H_N MODE_VCCHIB_N VSSD VDDIO_Q
+ VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_1 IB_MODE_SEL_H_N INP_DIS_I_H_N MODE_NORMAL_N VSSD VDDIO_Q
+ VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_2 INP_DIS_H_N sky130_fd_io__hvsbt_nand2_3/OUT INP_DIS_I_H
+ VSSD VDDIO_Q VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_3 sky130_fd_io__hvsbt_nand2_3/IN1 DM_H_N[2] sky130_fd_io__hvsbt_nand2_3/OUT
+ VSSD VDDIO_Q VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x1_0 INP_DIS_I_H_N VDDIO_Q VSSD VSSD INP_DIS_I_H VDDIO_Q
+ sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_nand2_3/IN1 VDDIO_Q VSSD VSSD sky130_fd_io__hvsbt_nand2v2_0/OUT
+ VDDIO_Q sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_2 TRIPSEL_I_H_N VDDIO_Q VSSD VSSD TRIPSEL_I_H VDDIO_Q
+ sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__signal_5_sym_hv_local_5term GATE NWELLRING VGND NBODY IN m1_204_67#
R0 NBODY m1_534_67# short w=20000u l=5000u
R1 NWELLRING m1_204_67# short w=20000u l=5000u
X0 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 w=5.4e+06u l=600000u
.ends

.subckt sky130_fd_io__gpiov2_buf_localesd VTRIP_SEL_H OUT_VT VDDIO_Q VSSD OUT_H IN_H
+ w_1005_268#
Xsky130_fd_io__signal_5_sym_hv_local_5term_0 VSSD VDDIO_Q VSSD VSSD OUT_H VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_1 VSSD VDDIO_Q OUT_H VSSD VDDIO_Q VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__res250only_small_0 IN_H OUT_H VSSD sky130_fd_io__res250only_small
X0 OUT_H VTRIP_SEL_H OUT_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=1e+06u
.ends

.subckt sky130_fd_io__gpiov2_ipath ENABLE_VDDIO_LV OUT_H MODE_VCCHIB_N VCCHIB VDDIO_Q
+ VSSD PAD OUT DM_H_N[1] DM_H_N[0] DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H IB_MODE_SEL_H_N
+ VTRIP_SEL_H_N m1_2064_35655#
Xsky130_fd_io__gpiov2_ibuf_se_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VCCHIB
+ ENABLE_VDDIO_LV sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N VSSD VDDIO_Q OUT sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ sky130_fd_io__gpiov2_ibuf_se_0/IN_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H MODE_VCCHIB_N
+ OUT_H m2_15184_37213# PAD sky130_fd_io__gpiov2_ibuf_se
Xsky130_fd_io__gpiov2_ictl_logic_0 sky130_fd_io__gpiov2_ictl_logic_0/INP_DIS_I_H_N
+ sky130_fd_io__gpiov2_ictl_logic_0/INP_DIS_I_H INP_DIS_H_N DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ IB_MODE_SEL_H_N VDDIO_Q VSSD VTRIP_SEL_H_N sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N
+ MODE_VCCHIB_N sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N
+ IB_MODE_SEL_H sky130_fd_io__gpiov2_ictl_logic
Xsky130_fd_io__gpiov2_buf_localesd_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ VDDIO_Q VSSD sky130_fd_io__gpiov2_ibuf_se_0/IN_H PAD VSSD sky130_fd_io__gpiov2_buf_localesd
.ends

.subckt sky130_fd_io__com_ctl_ls_en_1_v2 DM[1] VCC_IO VPB OUT_H_N OUT_H RST_H SET_H
+ VPWR HLD_H_N VSUBS a_1762_n1276# w_1114_n948# w_n17_1379# a_1150_n777#
X0 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X1 VSUBS RST_H a_65_861# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X2 OUT_H a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X3 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X4 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X5 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X6 a_361_1391# HLD_H_N a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X7 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X8 a_634_829# a_992_934# a_1150_n777# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 a_1150_n777# DM[1] a_992_934# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X12 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X13 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X14 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X15 VSUBS a_65_861# a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X16 a_1762_n1276# DM[1] a_992_934# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X17 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X18 VSUBS a_65_861# OUT_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X19 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X20 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X21 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X22 a_65_861# HLD_H_N a_957_1391# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X23 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X24 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X25 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X26 a_634_829# a_992_934# a_1762_n1276# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X27 a_130_181# SET_H VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X28 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X29 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X30 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X31 a_65_861# a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
.ends

.subckt sky130_fd_io__com_ctl_ls_v2 VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N
+ VSUBS w_n17_1379#
X0 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X1 VSUBS RST_H a_65_861# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X2 a_634_829# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X3 OUT_H a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X4 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X5 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X6 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X7 a_361_1391# HLD_H_N a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X8 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X10 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X12 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X13 VSUBS IN a_992_934# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X14 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X15 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X17 VSUBS a_65_861# a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X18 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X19 VSUBS a_65_861# OUT_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X20 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X21 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X22 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X23 a_65_861# HLD_H_N a_957_1391# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X24 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X25 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X26 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X27 a_130_181# SET_H VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X28 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X29 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X30 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X31 a_65_861# a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
.ends

.subckt sky130_fd_io__com_ctl_lsv2 SET_H HLD_H_N VGND OUT_H OUT_H_N RST_H IN VPWR
+ VCC_IO w_4727_n1281# w_5775_333# m1_5613_1428# m1_5675_1428#
X0 a_4933_638# HLD_H_N a_4793_n866# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X1 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X2 a_4944_2840# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X3 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X4 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X5 a_4739_1530# HLD_H_N a_4700_968# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X6 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X7 OUT_H a_4739_1530# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X8 VGND IN a_4944_2496# VGND sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X9 a_4739_1530# a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X10 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X11 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X12 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X13 a_4793_n866# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X14 VCC_IO a_4793_n866# a_4739_1530# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X15 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X16 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X17 VCC_IO a_4739_1530# a_4793_n866# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X19 a_4700_638# VPWR a_4933_638# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X20 a_4944_2840# a_4944_2496# VPWR w_5775_333# sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 OUT_H_N a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X22 VCC_IO a_4793_n866# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X23 VGND a_4739_1530# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X24 VPWR IN a_4944_2496# w_5775_333# sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X26 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X27 a_4793_n866# a_4739_1530# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X28 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X29 VGND SET_H a_4739_1530# VGND sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X30 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X31 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
.ends

.subckt sky130_fd_io__com_ctl_ls_1v2 VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR
+ HLD_H_N VSUBS w_n17_1379#
X0 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X1 VSUBS RST_H a_65_861# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X2 a_634_829# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X3 OUT_H a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X4 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X5 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X6 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X7 a_361_1391# HLD_H_N a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X8 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X10 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X12 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X13 VSUBS IN a_992_934# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X14 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X15 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X17 VSUBS a_65_861# a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X18 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X19 VSUBS a_65_861# OUT_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X20 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X21 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X22 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X23 a_65_861# HLD_H_N a_957_1391# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X24 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X25 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X26 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X27 a_130_181# SET_H VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X28 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X29 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X30 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X31 a_65_861# a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
.ends

.subckt sky130_fd_io__gpiov2_ctl_lsbank VTRIP_SEL_H VTRIP_SEL VTRIP_SEL_H_N INP_DIS
+ INP_DIS_H INP_DIS_H_N DM[0] DM_H[0] DM_H_N[0] DM_H[1] DM_H_N[1] DM[2] DM_H[2] DM_H_N[2]
+ VPWR DM[1] VCC_IO STARTUP_ST_H VGND STARTUP_RST_H HLD_I_H_N OD_I_H IB_MODE_SEL_H_N
+ IB_MODE_SEL_H IB_MODE_SEL VSUBS m1_2266_545# w_15552_2653# sky130_fd_io__com_ctl_lsv2_0/VCC_IO
+ sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
Xsky130_fd_io__com_ctl_ls_en_1_v2_0 DM[1] VCC_IO VPWR DM_H_N[1] DM_H[1] sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H VPWR HLD_I_H_N VSUBS sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ VPWR VGND VPWR sky130_fd_io__com_ctl_ls_en_1_v2
Xsky130_fd_io__com_ctl_ls_v2_0 VCC_IO VPWR DM_H_N[2] DM_H[2] DM[2] sky130_fd_io__com_ctl_ls_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_v2_0/SET_H VPWR HLD_I_H_N VSUBS VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_1 VCC_IO VPWR INP_DIS_H_N INP_DIS_H INP_DIS sky130_fd_io__com_ctl_ls_v2_1/RST_H
+ sky130_fd_io__com_ctl_ls_v2_1/SET_H VPWR HLD_I_H_N VSUBS VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_2 VCC_IO VPWR DM_H_N[0] DM_H[0] DM[0] sky130_fd_io__com_ctl_ls_v2_2/RST_H
+ sky130_fd_io__com_ctl_ls_v2_2/SET_H VPWR HLD_I_H_N VSUBS VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_lsv2_0 sky130_fd_io__com_ctl_lsv2_0/SET_H HLD_I_H_N VSUBS IB_MODE_SEL_H
+ IB_MODE_SEL_H_N sky130_fd_io__com_ctl_lsv2_0/RST_H IB_MODE_SEL VPWR sky130_fd_io__com_ctl_lsv2_0/VCC_IO
+ w_15552_2653# VPWR VSUBS VSUBS sky130_fd_io__com_ctl_lsv2
Xsky130_fd_io__com_ctl_ls_1v2_0 VCC_IO VPWR VTRIP_SEL_H_N VTRIP_SEL_H VTRIP_SEL sky130_fd_io__com_ctl_ls_1v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_1v2_0/SET_H VPWR HLD_I_H_N VSUBS VSUBS sky130_fd_io__com_ctl_ls_1v2
R0 sky130_fd_io__com_ctl_ls_v2_0/SET_H m1_10303_506# short w=260000u l=10000u
R1 OD_I_H m1_10029_412# short w=230000u l=10000u
R2 STARTUP_ST_H m1_5955_333# short w=230000u l=10000u
R3 sky130_fd_io__com_ctl_ls_v2_1/SET_H m1_6421_356# short w=260000u l=10000u
R4 sky130_fd_io__com_ctl_lsv2_0/SET_H m2_15089_329# short w=260000u l=10000u
R5 m2_15027_104# sky130_fd_io__com_ctl_lsv2_0/SET_H short w=260000u l=10000u
R6 VGND m1_2266_320# short w=260000u l=10000u
R7 m2_14799_410# sky130_fd_io__com_ctl_lsv2_0/RST_H short w=260000u l=10000u
R8 m1_5875_412# sky130_fd_io__com_ctl_ls_v2_2/RST_H short w=230000u l=10000u
R9 OD_I_H m2_14799_410# short w=260000u l=10000u
R10 STARTUP_RST_H m1_5875_412# short w=230000u l=10000u
R11 sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H m1_2467_370# short w=230000u l=10000u
R12 m1_10302_320# sky130_fd_io__com_ctl_ls_v2_0/SET_H short w=260000u l=10000u
R13 STARTUP_ST_H m1_6620_334# short w=230000u l=10000u
R14 m1_2553_412# m1_2266_545# short w=230000u l=10000u
R15 OD_I_H m2_14990_104# short w=260000u l=10000u
R16 VSUBS m1_14911_546# short w=260000u l=10000u
R17 sky130_fd_io__com_ctl_ls_v2_2/SET_H m1_6149_506# short w=260000u l=10000u
R18 sky130_fd_io__com_ctl_ls_v2_0/RST_H m1_10109_370# short w=230000u l=10000u
R19 sky130_fd_io__com_ctl_ls_v2_1/RST_H m1_6707_412# short w=230000u l=10000u
R20 m1_6420_507# STARTUP_RST_H short w=260000u l=10000u
R21 sky130_fd_io__com_ctl_ls_1v2_0/RST_H m1_14263_617# short w=230000u l=10000u
R22 sky130_fd_io__com_ctl_ls_1v2_0/SET_H m1_14457_467# short w=260000u l=10000u
R23 sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H m1_2267_506# short w=260000u l=10000u
R24 sky130_fd_io__com_ctl_ls_1v2_0/SET_H m1_14456_624# short w=260000u l=10000u
R25 OD_I_H m1_10303_543# short w=260000u l=10000u
R26 sky130_fd_io__com_ctl_ls_v2_2/RST_H m1_5955_370# short w=230000u l=10000u
R27 m1_6148_320# sky130_fd_io__com_ctl_ls_v2_2/SET_H short w=260000u l=10000u
R28 m2_15089_329# VSUBS short w=260000u l=10000u
R29 m1_2266_320# sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H short w=260000u l=10000u
R30 sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H m1_2553_412# short w=230000u l=10000u
R31 STARTUP_ST_H m1_6421_319# short w=260000u l=10000u
R32 m1_10029_412# sky130_fd_io__com_ctl_ls_v2_0/RST_H short w=230000u l=10000u
R33 m1_6620_334# sky130_fd_io__com_ctl_ls_v2_1/RST_H short w=230000u l=10000u
R34 VGND m1_10302_320# short w=260000u l=10000u
R35 VGND m1_2467_333# short w=230000u l=10000u
R36 STARTUP_RST_H m1_6149_543# short w=260000u l=10000u
R37 m1_14183_362# sky130_fd_io__com_ctl_ls_1v2_0/RST_H short w=230000u l=10000u
R38 sky130_fd_io__com_ctl_lsv2_0/RST_H m1_14911_509# short w=260000u l=10000u
R39 OD_I_H m1_14183_362# short w=230000u l=10000u
R40 VSUBS m1_14263_654# short w=230000u l=10000u
R41 VGND m1_10109_333# short w=230000u l=10000u
R42 m1_2266_545# m1_2267_543# short w=260000u l=10000u
R43 sky130_fd_io__com_ctl_ls_v2_1/SET_H m1_6420_507# short w=260000u l=10000u
R44 m1_14456_624# VSUBS short w=260000u l=10000u
R45 OD_I_H m1_14457_430# short w=260000u l=10000u
R46 m1_6744_412# STARTUP_RST_H short w=230000u l=10000u
R47 STARTUP_ST_H m1_6148_320# short w=260000u l=10000u
.ends

.subckt sky130_fd_io__hvsbt_inv_x8 IN VPWR VGND OUT VSUBS w_n42_416#
X0 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X4 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X5 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X6 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X7 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X8 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X9 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X10 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X11 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X12 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X13 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X14 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X15 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X16 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X17 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X18 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X19 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X20 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X21 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X22 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X23 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__hvsbt_inv_x4 IN OUT VSUBS a_66_482# a_66_144# w_n42_416#
X0 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 OUT IN a_66_144# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X4 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X5 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X6 a_66_144# IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X7 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X8 a_66_144# IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X9 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X10 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X11 OUT IN a_66_144# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__com_ctl_ls VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N
+ VSUBS w_n17_1379#
X0 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X1 VSUBS RST_H a_65_861# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X2 a_634_829# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X3 OUT_H a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X4 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X5 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X6 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X7 a_361_1391# HLD_H_N a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X8 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X10 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X12 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X13 VSUBS IN a_992_934# VSUBS sky130_fd_pr__nfet_01v8 w=1e+06u l=250000u
X14 VSUBS a_634_829# a_128_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X15 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=3e+06u l=600000u
X17 VSUBS a_65_861# a_130_181# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
X18 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X19 VSUBS a_65_861# OUT_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=1e+06u l=600000u
X20 a_128_1391# a_634_829# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X21 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X22 a_957_1391# VPWR a_724_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X23 a_65_861# HLD_H_N a_957_1391# VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X24 a_361_1391# VPWR a_128_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X25 a_724_1391# a_992_934# VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X26 a_724_1391# VPWR a_957_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X27 a_130_181# SET_H VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=3e+06u l=600000u
X28 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X29 a_128_1391# VPWR a_361_1391# VSUBS sky130_fd_pr__nfet_05v0_nvt w=1e+06u l=900000u
X30 VSUBS a_992_934# a_724_1391# VSUBS sky130_fd_pr__nfet_01v8_lvt w=1e+06u l=150000u
X31 a_65_861# a_130_181# VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=1e+06u
.ends

.subckt sky130_fd_io__hvsbt_inv_x8v2 IN VPWR VGND OUT VSUBS w_n42_416#
X0 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X1 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X2 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X3 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X4 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X5 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X6 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X7 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X8 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X9 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X10 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X11 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X12 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X13 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X14 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X15 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X16 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X17 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X18 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X19 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X20 VGND IN OUT VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
X21 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X22 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=600000u
X23 OUT IN VGND VSUBS sky130_fd_pr__nfet_g5v0d10v5 w=700000u l=600000u
.ends

.subckt sky130_fd_io__com_ctl_hldv2 HLD_OVR VCC_IO VGND HLD_I_H_N OD_I_H VPWR HLD_I_H
+ m2_3665_4183# sky130_fd_io__hvsbt_nand2_0/IN0 m1_3684_4201# sky130_fd_io__hvsbt_nand2_0/IN1
+ li_8226_3758# m2_3561_4196#
Xsky130_fd_io__hvsbt_inv_x8_0 sky130_fd_io__hvsbt_inv_x8_0/IN VCC_IO VGND sky130_fd_io__hvsbt_inv_x8_0/OUT
+ VGND VCC_IO sky130_fd_io__hvsbt_inv_x8
Xsky130_fd_io__hvsbt_inv_x4_0 sky130_fd_io__hvsbt_inv_x4_0/IN OD_I_H VGND VCC_IO VGND
+ VCC_IO sky130_fd_io__hvsbt_inv_x4
Xsky130_fd_io__hvsbt_inv_x4_1 sky130_fd_io__hvsbt_nor_0/IN0 sky130_fd_io__hvsbt_inv_x8_0/IN
+ VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_inv_x4
Xsky130_fd_io__hvsbt_nor_0 sky130_fd_io__hvsbt_nor_0/IN0 VGND VCC_IO VGND VCC_IO sky130_fd_io__com_ctl_ls_0/OUT_H
+ li_8312_3766# sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nor_1 OD_I_H VGND VCC_IO VGND VCC_IO li_8312_3766# li_8226_3758#
+ sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__hvsbt_nand2_0/IN0
+ sky130_fd_io__hvsbt_nand2_0/OUT VGND VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__com_ctl_ls_0 VCC_IO VPWR sky130_fd_io__com_ctl_ls_0/OUT_H_N sky130_fd_io__com_ctl_ls_0/OUT_H
+ HLD_OVR sky130_fd_io__hvsbt_inv_x1_0/OUT VGND VPWR sky130_fd_io__hvsbt_nor_0/IN0
+ VGND VGND sky130_fd_io__com_ctl_ls
Xsky130_fd_io__hvsbt_inv_x8v2_0 sky130_fd_io__hvsbt_inv_x8_0/IN VCC_IO VGND sky130_fd_io__hvsbt_inv_x8v2_0/OUT
+ VGND VCC_IO sky130_fd_io__hvsbt_inv_x8v2
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x1_0/OUT VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_0/IN0
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_inv_x4_0/IN VCC_IO VGND VGND sky130_fd_io__hvsbt_inv_x1_0/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_2 sky130_fd_io__hvsbt_nor_0/IN0 VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_0/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
R0 sky130_fd_io__hvsbt_inv_x8v2_0/OUT HLD_I_H_N short w=230000u l=25000u
R1 HLD_I_H sky130_fd_io__hvsbt_inv_x8_0/IN short w=230000u l=10000u
R2 HLD_I_H_N sky130_fd_io__hvsbt_inv_x8_0/OUT short w=230000u l=25000u
.ends

.subckt sky130_fd_io__gpiov2_ctl VTRIP_SEL_H_N DM[0] DM[2] DM_H[0] DM_H[1] HLD_OVR
+ DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2] INP_DIS INP_DIS_H_N VTRIP_SEL_H VTRIP_SEL
+ VPWR HLD_H_N OD_I_H INP_STARTUP_EN_H IB_MODE_SEL_H_N IB_MODE_SEL_H IB_MODE_SEL DM[1]
+ ENABLE_INP_H VCC_IO HLD_I_H_N ENABLE_H VGND HLD_I_OVR_H sky130_fd_io__com_ctl_hldv2_0/HLD_I_H
+ sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ li_18199_5031# li_11745_4176#
Xsky130_fd_io__gpiov2_ctl_lsbank_0 VTRIP_SEL_H VTRIP_SEL VTRIP_SEL_H_N INP_DIS sky130_fd_io__gpiov2_ctl_lsbank_0/INP_DIS_H
+ INP_DIS_H_N DM[0] DM_H[0] DM_H_N[0] DM_H[1] DM_H_N[1] DM[2] DM_H[2] DM_H_N[2] VPWR
+ DM[1] VCC_IO INP_STARTUP_EN_H VGND sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H
+ HLD_I_H_N OD_I_H IB_MODE_SEL_H_N IB_MODE_SEL_H IB_MODE_SEL VGND OD_I_H VCC_IO VCC_IO
+ sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ sky130_fd_io__gpiov2_ctl_lsbank
Xsky130_fd_io__com_ctl_hldv2_0 HLD_OVR VCC_IO VGND HLD_I_H_N OD_I_H VPWR sky130_fd_io__com_ctl_hldv2_0/HLD_I_H
+ OD_I_H ENABLE_H OD_I_H HLD_H_N HLD_I_OVR_H OD_I_H sky130_fd_io__com_ctl_hldv2
Xsky130_fd_io__hvsbt_nor_0 ENABLE_INP_H VGND VCC_IO VGND VCC_IO li_11745_4176# sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H
+ sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nand2_0 ENABLE_INP_H OD_I_H sky130_fd_io__hvsbt_nand2_0/OUT VGND
+ VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x1_0 INP_STARTUP_EN_H VCC_IO VGND VGND sky130_fd_io__hvsbt_nand2_0/OUT
+ VCC_IO sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__top_gpiov2 PAD VSSIO AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO VSWITCH
+ VDDA VCCD VCCHIB VSSIO_Q PAD_A_NOESD_H ANALOG_POL ENABLE_VDDIO IN_H IN ANALOG_EN
+ OUT TIE_HI_ESD PAD_A_ESD_1_H DM[0] DM[1] DM[2] HLD_H_N HLD_OVR INP_DIS ENABLE_VDDA_H
+ VTRIP_SEL OE_N SLOW TIE_LO_ESD PAD_A_ESD_0_H ANALOG_SEL ENABLE_INP_H ENABLE_H IB_MODE_SEL
+ ENABLE_VSWITCH_H
Xsky130_fd_io__gpio_opathv2_0 VSSIO sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N sky130_fd_io__gpiov2_ctl_0/OD_I_H
+ SLOW VDDIO VCCD VCCHIB PAD TIE_HI_ESD VDDA sky130_fd_io__gpiov2_ctl_0/DM_H[0] sky130_fd_io__gpiov2_ctl_0/DM_H[1]
+ sky130_fd_io__gpiov2_ctl_0/DM_H[2] sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] sky130_fd_io__gpiov2_ctl_0/DM_H_N[1]
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H OE_N
+ OUT TIE_LO_ESD li_3334_5352# li_3958_5352# VSSIO li_4745_6400# VSSIO sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS_uq3
+ a_1009_20453# li_5245_3919# li_2678_6400# li_5278_5352# sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N
+ sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] VSSIO sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS_uq5
+ li_3442_6400# li_7636_6398# PAD VSSIO li_3302_6400# li_10974_4971# li_7854_5377#
+ sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ li_9062_7268# sky130_fd_io__gpio_opathv2
Xsky130_fd_io__gpiov2_amux_0 PAD AMUXBUS_B AMUXBUS_A VDDIO_Q VSSIO VCCD VDDA VSSIO_Q
+ OUT sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N sky130_fd_io__gpiov2_amux_0/HLD_I_H ENABLE_VSWITCH_H
+ ENABLE_VDDA_H ANALOG_SEL ANALOG_POL ANALOG_EN sky130_fd_io__gpiov2_amux_0/VSWITCH
+ VSSIO sky130_fd_io__gpiov2_amux_0/HLD_I_H sky130_fd_io__gpiov2_amux
Xsky130_fd_io__res75only_small_0 PAD_A_ESD_1_H sky130_fd_io__res75only_small_1/PAD
+ VSSIO sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 sky130_fd_io__res75only_small_1/PAD PAD VSSIO sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 PAD_A_ESD_0_H sky130_fd_io__res75only_small_3/PAD
+ VSSIO sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD PAD VSSIO sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_ipath_0 ENABLE_VDDIO IN_H sky130_fd_io__gpiov2_ipath_0/MODE_VCCHIB_N
+ VCCHIB VDDIO_Q VSSIO PAD IN sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] sky130_fd_io__gpiov2_ctl_0/DM_H_N[0]
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H
+ sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N
+ VDDIO sky130_fd_io__gpiov2_ipath
* Xsky130_fd_io__overlay_gpiov2_m4_0 AMUXBUS_B VSSIO VSSIO AMUXBUS_A VDDA VSSIO VSSIO_Q
* + VCCHIB VSWITCH VCCD VDDIO VDDIO_Q PAD sky130_fd_io__overlay_gpiov2_m4
Xsky130_fd_io__gpiov2_ctl_0 sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N DM[0] DM[2] sky130_fd_io__gpiov2_ctl_0/DM_H[0]
+ sky130_fd_io__gpiov2_ctl_0/DM_H[1] HLD_OVR sky130_fd_io__gpiov2_ctl_0/DM_H[2] sky130_fd_io__gpiov2_ctl_0/DM_H_N[0]
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] INP_DIS
+ sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H VTRIP_SEL
+ VCCD HLD_H_N sky130_fd_io__gpiov2_ctl_0/OD_I_H sky130_fd_io__gpiov2_ctl_0/INP_STARTUP_EN_H
+ sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H
+ IB_MODE_SEL DM[1] ENABLE_INP_H VDDIO_Q sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N ENABLE_H
+ VSSIO sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H sky130_fd_io__gpiov2_amux_0/HLD_I_H
+ VSSIO PAD ENABLE_H sky130_fd_io__gpiov2_ctl
R0 PAD_A_NOESD_H PAD short w=1.237e+07u l=35000u
R1 PAD_A_NOESD_H PAD short w=1.07e+06u l=35000u
.ends

