magic
tech sky130A
magscale 1 2
timestamp 1606075443
<< error_s >>
rect -282 8620 -266 8678
rect 336 8666 340 8678
rect 348 8632 352 8666
rect -94 8054 -82 8100
rect 185 8074 189 8108
<< nwell >>
rect -7877 8875 -1295 9326
<< pwell >>
rect -7484 8100 -7428 8110
rect -5312 7347 -5094 7557
<< locali >>
rect -7906 9806 -7764 9819
rect -7906 9721 -7890 9806
rect -7778 9721 -7764 9806
rect -7906 8982 -7764 9721
rect -1056 9804 -813 9817
rect -1056 9643 -1011 9804
rect -830 9643 -813 9804
rect -1056 8986 -813 9643
rect -4904 8982 -813 8986
rect -7906 8966 -813 8982
rect -7906 8836 -1020 8966
rect -7912 7919 -7826 8710
rect -4904 8553 -1020 8836
rect -837 8853 -813 8966
rect -837 8732 2882 8853
rect -837 8553 -813 8732
rect -4904 8536 -813 8553
rect -5040 8224 -813 8369
rect -5040 7919 -4727 8224
rect -7912 7851 -4727 7919
rect -7912 7849 -7442 7851
rect -7912 7723 -7899 7849
rect -7661 7723 -7442 7849
rect -7912 7722 -7442 7723
rect -4996 7784 -4727 7851
rect -1831 7919 -813 8224
rect -1831 7784 2913 7919
rect -4996 7722 2913 7784
rect -7912 7674 2913 7722
rect -7912 7344 -7258 7674
rect -6941 7344 -6554 7560
rect -6169 7344 -5782 7560
rect -5397 7546 -5010 7560
rect -5397 7360 -5299 7546
rect -5107 7360 -5010 7546
rect -5397 7344 -5010 7360
rect -4625 7344 -4238 7560
rect -3853 7344 -3466 7560
rect -3081 7344 -2694 7560
rect -2309 7344 -1922 7560
rect -1537 7344 -1150 7560
rect -765 7344 -378 7560
rect 7 7344 394 7560
rect 779 7344 1166 7560
rect 1551 7344 1938 7560
rect 2709 7344 2890 7560
rect -7896 1696 -7713 1912
rect -7328 1696 -6941 1912
rect -6556 1696 -6169 1912
rect -5784 1696 -5397 1912
rect -5012 1696 -4625 1912
rect -4240 1696 -3853 1912
rect -3468 1696 -3081 1912
rect -2696 1696 -2309 1912
rect -1924 1696 -1537 1912
rect -1152 1696 -765 1912
rect -380 1696 7 1912
rect 392 1696 779 1912
rect 1164 1696 1551 1912
rect 1936 1696 2323 1912
rect 2708 1696 2888 1912
<< viali >>
rect -7890 9721 -7778 9806
rect -1011 9643 -830 9804
rect 1277 9385 1323 9591
rect -343 9285 -140 9332
rect 1512 9285 1849 9332
rect 2838 9214 2872 9410
rect -1020 8553 -837 8966
rect -77 8306 181 8365
rect -7899 7723 -7661 7849
rect -7442 7722 -4996 7851
rect -4727 7784 -1831 8224
rect 492 8215 559 8409
rect 703 8251 906 8298
rect 2323 8266 2369 8427
rect -5299 7360 -5107 7546
rect 2255 7129 2393 7561
<< metal1 >>
rect -7907 9806 -814 9817
rect -7907 9721 -7890 9806
rect -7778 9804 -814 9806
rect -7778 9800 -1011 9804
rect -7323 9791 -1011 9800
rect -7323 9732 -6921 9791
rect -7778 9724 -6921 9732
rect -830 9740 -814 9804
rect -663 9783 2894 9809
rect -7778 9721 -1011 9724
rect -7907 9710 -1011 9721
rect -7729 9641 -7571 9658
rect -7729 9569 -7511 9641
rect -7238 9613 -7228 9675
rect -7146 9660 -7129 9675
rect -7146 9616 -5449 9660
rect -5118 9616 -4957 9660
rect -7146 9613 -7129 9616
rect -7729 9555 -7665 9569
rect -7729 9172 -7634 9555
rect -7572 9172 -7511 9569
rect -7426 9319 -7380 9571
rect -7320 9423 -5126 9559
rect -7445 9184 -5410 9319
rect -7729 9099 -7511 9172
rect -7426 9128 -7380 9184
rect -7238 9128 -7228 9137
rect -7729 9085 -7572 9099
rect -7729 9032 -7665 9085
rect -7426 9084 -7228 9128
rect -7238 9075 -7228 9084
rect -7146 9128 -7129 9137
rect -5081 9128 -5003 9616
rect -4954 9189 -4647 9335
rect -7146 9087 -4957 9128
rect -7146 9084 -5025 9087
rect -7146 9075 -7129 9084
rect -4587 9032 -4514 9653
rect -4248 9613 -3988 9659
rect -4461 9167 -4391 9566
rect -7729 8984 -4514 9032
rect -7729 8779 -7665 8984
rect -4450 8875 -4391 9167
rect -7762 8652 -7665 8779
rect -5565 8805 -4391 8875
rect -4248 9173 -4166 9613
rect -3664 9612 -2200 9656
rect -1864 9612 -1710 9656
rect -1037 9643 -1011 9710
rect -830 9643 -813 9740
rect -663 9684 -629 9783
rect 2855 9684 2894 9783
rect -663 9656 2894 9684
rect -3959 9336 -3922 9572
rect -3838 9403 -1876 9564
rect -3981 9176 -2145 9336
rect -4248 9131 -4174 9173
rect -4248 9085 -3989 9131
rect -3959 9128 -3922 9176
rect -1821 9128 -1759 9612
rect -1698 9415 -1410 9560
rect -1698 9221 -1685 9415
rect -4248 9032 -4174 9085
rect -3959 9084 -1708 9128
rect -1335 9032 -1273 9643
rect -4248 8984 -1273 9032
rect -7762 8500 -7684 8652
rect -5565 8605 -5495 8805
rect -4248 8696 -4174 8984
rect -5682 8578 -5672 8605
rect -7762 8104 -7665 8500
rect -7922 7849 -7646 7857
rect -7922 7723 -7899 7849
rect -7661 7723 -7646 7849
rect -7922 7716 -7646 7723
rect -7922 6879 -7814 7716
rect -7602 7475 -7548 8564
rect -7166 8534 -5672 8578
rect -5596 8578 -5495 8605
rect -5180 8605 -4174 8696
rect -5596 8534 -5209 8578
rect -7484 8276 -7313 8503
rect -5565 8483 -5495 8534
rect -7226 8346 -5495 8483
rect -7484 8110 -5387 8276
rect -7484 8100 -7313 8110
rect -7442 7857 -7313 8100
rect -5318 8064 -5254 8534
rect -5180 8480 -5105 8605
rect -1195 8596 -1124 9575
rect -1037 8966 -813 9643
rect 1271 9591 1329 9603
rect 1271 9385 1277 9591
rect 1323 9582 1329 9591
rect 2181 9582 2191 9584
rect 1323 9532 2191 9582
rect 1323 9385 1329 9532
rect 2181 9530 2191 9532
rect 2343 9530 2353 9584
rect 1271 9373 1329 9385
rect 2832 9410 2878 9422
rect -355 9332 392 9338
rect -355 9285 -343 9332
rect -140 9285 392 9332
rect -355 9279 392 9285
rect 572 9332 1861 9338
rect 572 9285 1512 9332
rect 1849 9285 1861 9332
rect 572 9279 1861 9285
rect 2832 9259 2838 9410
rect 2872 9259 2878 9410
rect 2796 9205 2806 9259
rect 2958 9205 2968 9259
rect 2832 9202 2878 9205
rect -5191 8104 -5105 8480
rect -1540 8567 -1122 8596
rect -4780 8350 -1773 8373
rect -4780 8224 -3616 8350
rect -2669 8224 -1773 8350
rect -7166 8020 -5672 8064
rect -5682 7991 -5672 8020
rect -5597 7991 -5587 8064
rect -5362 8020 -5208 8064
rect -4780 7857 -4727 8224
rect -7454 7851 -4727 7857
rect -7454 7722 -7442 7851
rect -4996 7784 -4727 7851
rect -1831 8062 -1773 8224
rect -1540 8154 -1515 8567
rect -1144 8371 -1122 8567
rect -1037 8553 -1020 8966
rect -837 8855 -813 8966
rect -668 9074 2889 9101
rect -668 8980 -641 9074
rect 396 8980 671 9074
rect 2702 8980 2889 9074
rect -668 8948 2889 8980
rect -837 8830 2885 8855
rect -837 8655 -776 8830
rect 373 8655 655 8830
rect 2803 8655 2885 8830
rect -837 8625 2885 8655
rect -837 8553 -813 8625
rect 2569 8624 2885 8625
rect -1037 8525 -813 8553
rect 2317 8427 2375 8439
rect 486 8409 565 8421
rect -1144 8365 193 8371
rect -1144 8306 -77 8365
rect 181 8306 193 8365
rect -1144 8300 193 8306
rect -1144 8154 -1122 8300
rect 482 8215 492 8409
rect 559 8304 569 8409
rect 559 8298 918 8304
rect 559 8251 703 8298
rect 906 8251 918 8298
rect 2317 8266 2323 8427
rect 2369 8365 2375 8427
rect 2369 8296 2560 8365
rect 2725 8296 2735 8365
rect 2369 8266 2375 8296
rect 2317 8254 2375 8266
rect 559 8245 918 8251
rect 559 8215 569 8245
rect 486 8203 565 8215
rect -1540 8131 -1122 8154
rect -1831 7850 2880 8062
rect -1831 7784 -1773 7850
rect -4996 7768 -1773 7784
rect 2274 7791 2769 7801
rect -4996 7722 -1772 7768
rect -7454 7716 -1772 7722
rect 2274 7718 2286 7791
rect 2753 7718 2769 7791
rect 2274 7707 2769 7718
rect 2274 7576 2368 7707
rect 2240 7561 2406 7576
rect -5312 7546 -5094 7557
rect -5312 7475 -5299 7546
rect -7602 7421 -5299 7475
rect -5312 7360 -5299 7421
rect -5107 7360 -5094 7546
rect -5312 7347 -5094 7360
rect 2240 7129 2255 7561
rect 2393 7129 2406 7561
rect 2240 7113 2406 7129
rect 2858 6879 2920 7610
rect -7922 6279 2920 6879
rect -7922 5879 -7814 6279
rect 2858 5879 2920 6279
rect -7922 5279 2920 5879
rect -7922 4879 -7814 5279
rect 2858 4879 2920 5279
rect -7922 4279 2920 4879
rect -7922 3879 -7814 4279
rect 2858 3879 2920 4279
rect -7922 3279 2920 3879
rect -7922 2879 -7814 3279
rect 2858 2879 2920 3279
rect -7922 2279 2920 2879
rect -7922 1630 -7814 2279
rect 2858 1630 2920 2279
rect -7922 1542 2920 1630
<< via1 >>
rect -7887 9732 -7778 9800
rect -7778 9732 -7323 9800
rect -6921 9724 -1011 9791
rect -1011 9724 -854 9791
rect -7228 9613 -7146 9675
rect -7228 9075 -7146 9137
rect -629 9684 2855 9783
rect -5672 8534 -5596 8605
rect 2191 9530 2343 9584
rect 392 9279 572 9338
rect 2806 9214 2838 9259
rect 2838 9214 2872 9259
rect 2872 9214 2958 9259
rect 2806 9205 2958 9214
rect -3616 8224 -2669 8350
rect -5672 7991 -5597 8064
rect -3616 7801 -2669 8224
rect -1515 8154 -1144 8567
rect -641 8980 396 9074
rect 671 8980 2702 9074
rect -776 8655 373 8830
rect 655 8655 2803 8830
rect 492 8215 559 8409
rect 2560 8296 2725 8365
rect 2286 7718 2753 7791
<< metal2 >>
rect -6962 9817 -815 9818
rect -7909 9800 -815 9817
rect -7909 9732 -7887 9800
rect -7323 9792 -815 9800
rect -7909 9635 -7870 9732
rect -7313 9718 -7061 9792
rect -856 9791 -815 9792
rect -854 9724 -815 9791
rect -7313 9635 -7293 9718
rect -7909 9592 -7293 9635
rect -7228 9675 -7146 9685
rect -7228 9603 -7146 9613
rect -7081 9635 -7061 9718
rect -856 9635 -815 9724
rect -663 9783 2894 9809
rect -663 9684 -629 9783
rect 2855 9684 2894 9783
rect -663 9656 2894 9684
rect -7218 9147 -7162 9603
rect -7081 9591 -815 9635
rect 2191 9587 2343 9597
rect 2191 9517 2343 9527
rect 392 9338 572 9348
rect 392 9269 572 9279
rect -7228 9137 -7146 9147
rect -7228 9065 -7146 9075
rect -668 9074 427 9101
rect -668 8980 -641 9074
rect 396 8980 427 9074
rect -668 8948 427 8980
rect -806 8830 408 8855
rect -806 8655 -776 8830
rect 373 8655 408 8830
rect -806 8625 408 8655
rect -5672 8605 -5596 8615
rect -5672 8524 -5596 8534
rect -1540 8567 -1122 8596
rect -5659 8074 -5607 8524
rect -3639 8380 -2649 8399
rect -5672 8064 -5597 8074
rect -5672 7981 -5597 7991
rect -3639 7801 -3616 8380
rect -2669 7801 -2649 8380
rect -1540 8154 -1515 8567
rect -1144 8154 -1122 8567
rect 496 8419 553 9269
rect 2806 9262 2958 9272
rect 2806 9192 2958 9202
rect 641 9074 2720 9101
rect 640 8980 671 9074
rect 2702 8980 2720 9074
rect 641 8948 2720 8980
rect 620 8830 2851 8855
rect 620 8655 655 8830
rect 2803 8655 2851 8830
rect 620 8625 2851 8655
rect 492 8409 559 8419
rect 492 8205 559 8215
rect -1540 8131 -1122 8154
rect -3639 7780 -2649 7801
rect 2274 7801 2484 8625
rect 2551 8296 2560 8365
rect 2725 8296 2810 8365
rect 2962 8296 2971 8365
rect 2274 7791 2769 7801
rect 2274 7718 2286 7791
rect 2753 7718 2769 7791
rect 2274 7707 2769 7718
<< via2 >>
rect -7870 9732 -7323 9792
rect -7323 9732 -7313 9792
rect -7870 9635 -7313 9732
rect -7061 9791 -856 9792
rect -7061 9724 -6921 9791
rect -6921 9724 -856 9791
rect -7061 9635 -856 9724
rect -629 9684 2855 9783
rect 2191 9584 2343 9587
rect 2191 9530 2343 9584
rect 2191 9527 2343 9530
rect -641 8980 396 9074
rect -3616 8350 -2669 8380
rect -3616 8053 -2669 8350
rect -1515 8154 -1144 8567
rect 2806 9259 2958 9262
rect 2806 9205 2958 9259
rect 2806 9202 2958 9205
rect 671 8980 2702 9074
rect 2810 8296 2962 8365
<< metal3 >>
rect -7909 9792 -821 9814
rect -7909 9775 -7870 9792
rect -7313 9775 -7061 9792
rect -7909 9531 -7874 9775
rect -856 9635 -821 9792
rect -663 9783 2894 9809
rect -663 9684 -629 9783
rect 2855 9684 2894 9783
rect -663 9656 2894 9684
rect -874 9531 -821 9635
rect -7909 9496 -821 9531
rect 2181 9587 2348 9595
rect 2181 9527 2191 9587
rect 2343 9527 2484 9587
rect 2181 9522 2348 9527
rect 2424 9447 2484 9527
rect 2424 9387 3396 9447
rect 2796 9262 2963 9270
rect 2796 9202 2806 9262
rect 2958 9202 2963 9262
rect 2796 9197 2963 9202
rect -668 9074 2720 9101
rect -668 8980 -641 9074
rect 2702 8980 2720 9074
rect 2845 9082 2905 9197
rect 2845 9022 3397 9082
rect -668 8948 2720 8980
rect -3836 8808 -2648 8848
rect -3836 8380 -3597 8808
rect -2679 8380 -2648 8808
rect -3836 8053 -3616 8380
rect -2669 8053 -2648 8380
rect -1539 8567 -1122 8596
rect -1539 8154 -1515 8567
rect -1144 8154 -1122 8567
rect 2800 8365 2971 8371
rect 2800 8296 2810 8365
rect 2962 8296 3395 8365
rect 2800 8289 2971 8296
rect -1539 8131 -1122 8154
rect -3836 8025 -2648 8053
rect -3836 7782 -3640 8025
<< via3 >>
rect -7874 9635 -7870 9775
rect -7870 9635 -7313 9775
rect -7313 9635 -7061 9775
rect -7061 9635 -874 9775
rect -629 9684 2855 9783
rect -7874 9531 -874 9635
rect -641 8980 396 9074
rect 396 8980 671 9074
rect 671 8980 2702 9074
rect -3597 8380 -2679 8808
rect -3597 8089 -2679 8380
rect -1515 8154 -1144 8567
<< metal4 >>
rect -7909 9775 -821 9814
rect -7909 9531 -7874 9775
rect -874 9531 -821 9775
rect -7909 9496 -821 9531
rect -706 9783 3233 9822
rect -706 9684 -629 9783
rect 2855 9684 3233 9783
rect -706 9493 3233 9684
rect 2896 9286 3231 9305
rect -7909 9074 2720 9186
rect -7909 8980 -641 9074
rect 2702 8980 2720 9074
rect -7909 8808 2720 8980
rect -7909 8786 -3597 8808
rect -3930 8089 -3597 8786
rect -2679 8786 2720 8808
rect -2679 8089 -2648 8786
rect 2896 8605 2932 9286
rect -1561 8567 2932 8605
rect -1561 8154 -1515 8567
rect -1144 8154 2932 8567
rect -1561 8146 2932 8154
rect 3199 8146 3231 9286
rect -1561 8122 3231 8146
rect -3930 8053 -2648 8089
rect -3930 1582 -3736 8053
<< via4 >>
rect -3597 8089 -2679 8778
rect 2932 8146 3199 9286
<< metal5 >>
rect 2904 9286 3224 9310
rect -3634 8778 -2648 8848
rect -3634 8089 -3597 8778
rect -2679 8089 -2648 8778
rect -3634 8025 -2648 8089
rect -3440 7666 -2648 8025
rect 2904 8146 2932 9286
rect 3199 8146 3224 9286
rect 2904 7773 3224 8146
use sky130_fd_pr__nfet_g5v0d10v5_TGFUGS  sky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0
timestamp 1606063140
transform 1 0 -6432 0 1 8300
box -962 -458 962 458
use sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC  sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1
timestamp 1605994897
transform -1 0 -7576 0 1 8300
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ  sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0
timestamp 1606063140
transform 1 0 -6290 0 1 9372
box -1101 -497 1101 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3
timestamp 1606063140
transform 1 0 -7539 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__nfet_g5v0d10v5_PKVMTM  sky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0
timestamp 1606063140
transform 1 0 -5287 0 1 8301
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_YUHPBG  sky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0
timestamp 1606063140
transform 1 0 -5041 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0
timestamp 1606063140
transform 1 0 -4555 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1
timestamp 1606063140
transform 1 0 -4069 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_YEUEBV  sky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0
timestamp 1606063140
transform 1 0 -2929 0 1 9372
box -992 -497 992 497
use sky130_fd_pr__pfet_g5v0d10v5_YUHPXE  sky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0
timestamp 1606063140
transform 1 0 -1789 0 1 9372
box -338 -497 338 497
use sky130_fd_pr__pfet_g5v0d10v5_3YBPVB  sky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2
timestamp 1606063140
transform 1 0 -1303 0 1 9372
box -338 -497 338 497
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1606075443
transform 1 0 -480 0 1 7935
box -66 -23 1122 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1606075443
transform 1 0 576 0 1 7935
box -66 -23 1986 897
use sky130_fd_sc_hvl__buf_8  sky130_fd_sc_hvl__buf_8_1
timestamp 1606075443
transform 1 0 -470 0 1 8969
box -66 -23 1986 897
use sky130_fd_sc_hvl__fill_4  sky130_fd_sc_hvl__fill_4_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1606075443
transform 1 0 2496 0 1 7935
box -66 -23 450 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1606075443
transform 1 0 1450 0 1 8969
box -66 -23 1506 897
use sky130_fd_pr__res_xhigh_po_0p69_S5N9F3  sky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0
timestamp 1606074388
transform 1 0 -2501 0 1 4629
box -5446 -3098 5446 3098
use sky130_fd_pr__cap_mim_m3_1_N249RX  sky130_fd_pr__cap_mim_m3_1_N249RX_0
timestamp 1605923309
transform -1 0 -650 0 1 4682
box -3186 -3100 3186 3100
use sky130_fd_pr__cap_mim_m3_2_N249RX  sky130_fd_pr__cap_mim_m3_2_N249RX_0
timestamp 1605923309
transform 1 0 -177 0 1 4682
box -3379 -3101 3401 3101
<< labels >>
flabel metal2 520 8895 520 8895 0 FreeSans 320 0 0 0 out
flabel metal4 s -7909 9496 -7874 9814 0 FreeSans 320 0 0 0 vdd3v3
port 0 nsew
flabel metal4 s -7909 8786 -7715 9186 0 FreeSans 320 0 0 0 vss
port 2 nsew
flabel metal3 3022 8296 3395 8365 0 FreeSans 320 0 0 0 porb_h
port 3 nsew
flabel metal4 s 3027 9493 3233 9822 0 FreeSans 320 0 0 0 vdd1v8
port 1 nsew
flabel metal3 3242 9022 3397 9082 0 FreeSans 320 0 0 0 por_l
port 4 nsew
flabel metal3 3241 9387 3396 9447 0 FreeSans 320 0 0 0 porb_l
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 4360 9164
<< end >>
