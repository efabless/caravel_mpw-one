magic
tech sky130A
magscale 1 2
timestamp 1606426375
<< error_p >>
rect -8820 381 -8762 387
rect -8702 381 -8644 387
rect -8584 381 -8526 387
rect -8466 381 -8408 387
rect -8348 381 -8290 387
rect -8230 381 -8172 387
rect -8112 381 -8054 387
rect -7994 381 -7936 387
rect -7876 381 -7818 387
rect -7758 381 -7700 387
rect -7640 381 -7582 387
rect -7522 381 -7464 387
rect -7404 381 -7346 387
rect -7286 381 -7228 387
rect -7168 381 -7110 387
rect -7050 381 -6992 387
rect -6932 381 -6874 387
rect -6814 381 -6756 387
rect -6696 381 -6638 387
rect -6578 381 -6520 387
rect -6460 381 -6402 387
rect -6342 381 -6284 387
rect -6224 381 -6166 387
rect -6106 381 -6048 387
rect -5988 381 -5930 387
rect -5870 381 -5812 387
rect -5752 381 -5694 387
rect -5634 381 -5576 387
rect -5516 381 -5458 387
rect -5398 381 -5340 387
rect -5280 381 -5222 387
rect -5162 381 -5104 387
rect -5044 381 -4986 387
rect -4926 381 -4868 387
rect -4808 381 -4750 387
rect -4690 381 -4632 387
rect -4572 381 -4514 387
rect -4454 381 -4396 387
rect -4336 381 -4278 387
rect -4218 381 -4160 387
rect -4100 381 -4042 387
rect -3982 381 -3924 387
rect -3864 381 -3806 387
rect -3746 381 -3688 387
rect -3628 381 -3570 387
rect -3510 381 -3452 387
rect -3392 381 -3334 387
rect -3274 381 -3216 387
rect -3156 381 -3098 387
rect -3038 381 -2980 387
rect -2920 381 -2862 387
rect -2802 381 -2744 387
rect -2684 381 -2626 387
rect -2566 381 -2508 387
rect -2448 381 -2390 387
rect -2330 381 -2272 387
rect -2212 381 -2154 387
rect -2094 381 -2036 387
rect -1976 381 -1918 387
rect -1858 381 -1800 387
rect -1740 381 -1682 387
rect -1622 381 -1564 387
rect -1504 381 -1446 387
rect -1386 381 -1328 387
rect -1268 381 -1210 387
rect -1150 381 -1092 387
rect -1032 381 -974 387
rect -914 381 -856 387
rect -796 381 -738 387
rect -678 381 -620 387
rect -560 381 -502 387
rect -442 381 -384 387
rect -324 381 -266 387
rect -206 381 -148 387
rect -88 381 -30 387
rect 30 381 88 387
rect 148 381 206 387
rect 266 381 324 387
rect 384 381 442 387
rect 502 381 560 387
rect 620 381 678 387
rect 738 381 796 387
rect 856 381 914 387
rect 974 381 1032 387
rect 1092 381 1150 387
rect 1210 381 1268 387
rect 1328 381 1386 387
rect 1446 381 1504 387
rect 1564 381 1622 387
rect 1682 381 1740 387
rect 1800 381 1858 387
rect 1918 381 1976 387
rect 2036 381 2094 387
rect 2154 381 2212 387
rect 2272 381 2330 387
rect 2390 381 2448 387
rect 2508 381 2566 387
rect 2626 381 2684 387
rect 2744 381 2802 387
rect 2862 381 2920 387
rect 2980 381 3038 387
rect 3098 381 3156 387
rect 3216 381 3274 387
rect 3334 381 3392 387
rect 3452 381 3510 387
rect 3570 381 3628 387
rect 3688 381 3746 387
rect 3806 381 3864 387
rect 3924 381 3982 387
rect 4042 381 4100 387
rect 4160 381 4218 387
rect 4278 381 4336 387
rect 4396 381 4454 387
rect 4514 381 4572 387
rect 4632 381 4690 387
rect 4750 381 4808 387
rect 4868 381 4926 387
rect 4986 381 5044 387
rect 5104 381 5162 387
rect 5222 381 5280 387
rect 5340 381 5398 387
rect 5458 381 5516 387
rect 5576 381 5634 387
rect 5694 381 5752 387
rect 5812 381 5870 387
rect 5930 381 5988 387
rect 6048 381 6106 387
rect 6166 381 6224 387
rect 6284 381 6342 387
rect 6402 381 6460 387
rect 6520 381 6578 387
rect 6638 381 6696 387
rect 6756 381 6814 387
rect 6874 381 6932 387
rect 6992 381 7050 387
rect 7110 381 7168 387
rect 7228 381 7286 387
rect 7346 381 7404 387
rect 7464 381 7522 387
rect 7582 381 7640 387
rect 7700 381 7758 387
rect 7818 381 7876 387
rect 7936 381 7994 387
rect 8054 381 8112 387
rect 8172 381 8230 387
rect 8290 381 8348 387
rect 8408 381 8466 387
rect 8526 381 8584 387
rect 8644 381 8702 387
rect 8762 381 8820 387
rect -8820 347 -8808 381
rect -8702 347 -8690 381
rect -8584 347 -8572 381
rect -8466 347 -8454 381
rect -8348 347 -8336 381
rect -8230 347 -8218 381
rect -8112 347 -8100 381
rect -7994 347 -7982 381
rect -7876 347 -7864 381
rect -7758 347 -7746 381
rect -7640 347 -7628 381
rect -7522 347 -7510 381
rect -7404 347 -7392 381
rect -7286 347 -7274 381
rect -7168 347 -7156 381
rect -7050 347 -7038 381
rect -6932 347 -6920 381
rect -6814 347 -6802 381
rect -6696 347 -6684 381
rect -6578 347 -6566 381
rect -6460 347 -6448 381
rect -6342 347 -6330 381
rect -6224 347 -6212 381
rect -6106 347 -6094 381
rect -5988 347 -5976 381
rect -5870 347 -5858 381
rect -5752 347 -5740 381
rect -5634 347 -5622 381
rect -5516 347 -5504 381
rect -5398 347 -5386 381
rect -5280 347 -5268 381
rect -5162 347 -5150 381
rect -5044 347 -5032 381
rect -4926 347 -4914 381
rect -4808 347 -4796 381
rect -4690 347 -4678 381
rect -4572 347 -4560 381
rect -4454 347 -4442 381
rect -4336 347 -4324 381
rect -4218 347 -4206 381
rect -4100 347 -4088 381
rect -3982 347 -3970 381
rect -3864 347 -3852 381
rect -3746 347 -3734 381
rect -3628 347 -3616 381
rect -3510 347 -3498 381
rect -3392 347 -3380 381
rect -3274 347 -3262 381
rect -3156 347 -3144 381
rect -3038 347 -3026 381
rect -2920 347 -2908 381
rect -2802 347 -2790 381
rect -2684 347 -2672 381
rect -2566 347 -2554 381
rect -2448 347 -2436 381
rect -2330 347 -2318 381
rect -2212 347 -2200 381
rect -2094 347 -2082 381
rect -1976 347 -1964 381
rect -1858 347 -1846 381
rect -1740 347 -1728 381
rect -1622 347 -1610 381
rect -1504 347 -1492 381
rect -1386 347 -1374 381
rect -1268 347 -1256 381
rect -1150 347 -1138 381
rect -1032 347 -1020 381
rect -914 347 -902 381
rect -796 347 -784 381
rect -678 347 -666 381
rect -560 347 -548 381
rect -442 347 -430 381
rect -324 347 -312 381
rect -206 347 -194 381
rect -88 347 -76 381
rect 30 347 42 381
rect 148 347 160 381
rect 266 347 278 381
rect 384 347 396 381
rect 502 347 514 381
rect 620 347 632 381
rect 738 347 750 381
rect 856 347 868 381
rect 974 347 986 381
rect 1092 347 1104 381
rect 1210 347 1222 381
rect 1328 347 1340 381
rect 1446 347 1458 381
rect 1564 347 1576 381
rect 1682 347 1694 381
rect 1800 347 1812 381
rect 1918 347 1930 381
rect 2036 347 2048 381
rect 2154 347 2166 381
rect 2272 347 2284 381
rect 2390 347 2402 381
rect 2508 347 2520 381
rect 2626 347 2638 381
rect 2744 347 2756 381
rect 2862 347 2874 381
rect 2980 347 2992 381
rect 3098 347 3110 381
rect 3216 347 3228 381
rect 3334 347 3346 381
rect 3452 347 3464 381
rect 3570 347 3582 381
rect 3688 347 3700 381
rect 3806 347 3818 381
rect 3924 347 3936 381
rect 4042 347 4054 381
rect 4160 347 4172 381
rect 4278 347 4290 381
rect 4396 347 4408 381
rect 4514 347 4526 381
rect 4632 347 4644 381
rect 4750 347 4762 381
rect 4868 347 4880 381
rect 4986 347 4998 381
rect 5104 347 5116 381
rect 5222 347 5234 381
rect 5340 347 5352 381
rect 5458 347 5470 381
rect 5576 347 5588 381
rect 5694 347 5706 381
rect 5812 347 5824 381
rect 5930 347 5942 381
rect 6048 347 6060 381
rect 6166 347 6178 381
rect 6284 347 6296 381
rect 6402 347 6414 381
rect 6520 347 6532 381
rect 6638 347 6650 381
rect 6756 347 6768 381
rect 6874 347 6886 381
rect 6992 347 7004 381
rect 7110 347 7122 381
rect 7228 347 7240 381
rect 7346 347 7358 381
rect 7464 347 7476 381
rect 7582 347 7594 381
rect 7700 347 7712 381
rect 7818 347 7830 381
rect 7936 347 7948 381
rect 8054 347 8066 381
rect 8172 347 8184 381
rect 8290 347 8302 381
rect 8408 347 8420 381
rect 8526 347 8538 381
rect 8644 347 8656 381
rect 8762 347 8774 381
rect -8820 341 -8762 347
rect -8702 341 -8644 347
rect -8584 341 -8526 347
rect -8466 341 -8408 347
rect -8348 341 -8290 347
rect -8230 341 -8172 347
rect -8112 341 -8054 347
rect -7994 341 -7936 347
rect -7876 341 -7818 347
rect -7758 341 -7700 347
rect -7640 341 -7582 347
rect -7522 341 -7464 347
rect -7404 341 -7346 347
rect -7286 341 -7228 347
rect -7168 341 -7110 347
rect -7050 341 -6992 347
rect -6932 341 -6874 347
rect -6814 341 -6756 347
rect -6696 341 -6638 347
rect -6578 341 -6520 347
rect -6460 341 -6402 347
rect -6342 341 -6284 347
rect -6224 341 -6166 347
rect -6106 341 -6048 347
rect -5988 341 -5930 347
rect -5870 341 -5812 347
rect -5752 341 -5694 347
rect -5634 341 -5576 347
rect -5516 341 -5458 347
rect -5398 341 -5340 347
rect -5280 341 -5222 347
rect -5162 341 -5104 347
rect -5044 341 -4986 347
rect -4926 341 -4868 347
rect -4808 341 -4750 347
rect -4690 341 -4632 347
rect -4572 341 -4514 347
rect -4454 341 -4396 347
rect -4336 341 -4278 347
rect -4218 341 -4160 347
rect -4100 341 -4042 347
rect -3982 341 -3924 347
rect -3864 341 -3806 347
rect -3746 341 -3688 347
rect -3628 341 -3570 347
rect -3510 341 -3452 347
rect -3392 341 -3334 347
rect -3274 341 -3216 347
rect -3156 341 -3098 347
rect -3038 341 -2980 347
rect -2920 341 -2862 347
rect -2802 341 -2744 347
rect -2684 341 -2626 347
rect -2566 341 -2508 347
rect -2448 341 -2390 347
rect -2330 341 -2272 347
rect -2212 341 -2154 347
rect -2094 341 -2036 347
rect -1976 341 -1918 347
rect -1858 341 -1800 347
rect -1740 341 -1682 347
rect -1622 341 -1564 347
rect -1504 341 -1446 347
rect -1386 341 -1328 347
rect -1268 341 -1210 347
rect -1150 341 -1092 347
rect -1032 341 -974 347
rect -914 341 -856 347
rect -796 341 -738 347
rect -678 341 -620 347
rect -560 341 -502 347
rect -442 341 -384 347
rect -324 341 -266 347
rect -206 341 -148 347
rect -88 341 -30 347
rect 30 341 88 347
rect 148 341 206 347
rect 266 341 324 347
rect 384 341 442 347
rect 502 341 560 347
rect 620 341 678 347
rect 738 341 796 347
rect 856 341 914 347
rect 974 341 1032 347
rect 1092 341 1150 347
rect 1210 341 1268 347
rect 1328 341 1386 347
rect 1446 341 1504 347
rect 1564 341 1622 347
rect 1682 341 1740 347
rect 1800 341 1858 347
rect 1918 341 1976 347
rect 2036 341 2094 347
rect 2154 341 2212 347
rect 2272 341 2330 347
rect 2390 341 2448 347
rect 2508 341 2566 347
rect 2626 341 2684 347
rect 2744 341 2802 347
rect 2862 341 2920 347
rect 2980 341 3038 347
rect 3098 341 3156 347
rect 3216 341 3274 347
rect 3334 341 3392 347
rect 3452 341 3510 347
rect 3570 341 3628 347
rect 3688 341 3746 347
rect 3806 341 3864 347
rect 3924 341 3982 347
rect 4042 341 4100 347
rect 4160 341 4218 347
rect 4278 341 4336 347
rect 4396 341 4454 347
rect 4514 341 4572 347
rect 4632 341 4690 347
rect 4750 341 4808 347
rect 4868 341 4926 347
rect 4986 341 5044 347
rect 5104 341 5162 347
rect 5222 341 5280 347
rect 5340 341 5398 347
rect 5458 341 5516 347
rect 5576 341 5634 347
rect 5694 341 5752 347
rect 5812 341 5870 347
rect 5930 341 5988 347
rect 6048 341 6106 347
rect 6166 341 6224 347
rect 6284 341 6342 347
rect 6402 341 6460 347
rect 6520 341 6578 347
rect 6638 341 6696 347
rect 6756 341 6814 347
rect 6874 341 6932 347
rect 6992 341 7050 347
rect 7110 341 7168 347
rect 7228 341 7286 347
rect 7346 341 7404 347
rect 7464 341 7522 347
rect 7582 341 7640 347
rect 7700 341 7758 347
rect 7818 341 7876 347
rect 7936 341 7994 347
rect 8054 341 8112 347
rect 8172 341 8230 347
rect 8290 341 8348 347
rect 8408 341 8466 347
rect 8526 341 8584 347
rect 8644 341 8702 347
rect 8762 341 8820 347
rect -8820 -347 -8762 -341
rect -8702 -347 -8644 -341
rect -8584 -347 -8526 -341
rect -8466 -347 -8408 -341
rect -8348 -347 -8290 -341
rect -8230 -347 -8172 -341
rect -8112 -347 -8054 -341
rect -7994 -347 -7936 -341
rect -7876 -347 -7818 -341
rect -7758 -347 -7700 -341
rect -7640 -347 -7582 -341
rect -7522 -347 -7464 -341
rect -7404 -347 -7346 -341
rect -7286 -347 -7228 -341
rect -7168 -347 -7110 -341
rect -7050 -347 -6992 -341
rect -6932 -347 -6874 -341
rect -6814 -347 -6756 -341
rect -6696 -347 -6638 -341
rect -6578 -347 -6520 -341
rect -6460 -347 -6402 -341
rect -6342 -347 -6284 -341
rect -6224 -347 -6166 -341
rect -6106 -347 -6048 -341
rect -5988 -347 -5930 -341
rect -5870 -347 -5812 -341
rect -5752 -347 -5694 -341
rect -5634 -347 -5576 -341
rect -5516 -347 -5458 -341
rect -5398 -347 -5340 -341
rect -5280 -347 -5222 -341
rect -5162 -347 -5104 -341
rect -5044 -347 -4986 -341
rect -4926 -347 -4868 -341
rect -4808 -347 -4750 -341
rect -4690 -347 -4632 -341
rect -4572 -347 -4514 -341
rect -4454 -347 -4396 -341
rect -4336 -347 -4278 -341
rect -4218 -347 -4160 -341
rect -4100 -347 -4042 -341
rect -3982 -347 -3924 -341
rect -3864 -347 -3806 -341
rect -3746 -347 -3688 -341
rect -3628 -347 -3570 -341
rect -3510 -347 -3452 -341
rect -3392 -347 -3334 -341
rect -3274 -347 -3216 -341
rect -3156 -347 -3098 -341
rect -3038 -347 -2980 -341
rect -2920 -347 -2862 -341
rect -2802 -347 -2744 -341
rect -2684 -347 -2626 -341
rect -2566 -347 -2508 -341
rect -2448 -347 -2390 -341
rect -2330 -347 -2272 -341
rect -2212 -347 -2154 -341
rect -2094 -347 -2036 -341
rect -1976 -347 -1918 -341
rect -1858 -347 -1800 -341
rect -1740 -347 -1682 -341
rect -1622 -347 -1564 -341
rect -1504 -347 -1446 -341
rect -1386 -347 -1328 -341
rect -1268 -347 -1210 -341
rect -1150 -347 -1092 -341
rect -1032 -347 -974 -341
rect -914 -347 -856 -341
rect -796 -347 -738 -341
rect -678 -347 -620 -341
rect -560 -347 -502 -341
rect -442 -347 -384 -341
rect -324 -347 -266 -341
rect -206 -347 -148 -341
rect -88 -347 -30 -341
rect 30 -347 88 -341
rect 148 -347 206 -341
rect 266 -347 324 -341
rect 384 -347 442 -341
rect 502 -347 560 -341
rect 620 -347 678 -341
rect 738 -347 796 -341
rect 856 -347 914 -341
rect 974 -347 1032 -341
rect 1092 -347 1150 -341
rect 1210 -347 1268 -341
rect 1328 -347 1386 -341
rect 1446 -347 1504 -341
rect 1564 -347 1622 -341
rect 1682 -347 1740 -341
rect 1800 -347 1858 -341
rect 1918 -347 1976 -341
rect 2036 -347 2094 -341
rect 2154 -347 2212 -341
rect 2272 -347 2330 -341
rect 2390 -347 2448 -341
rect 2508 -347 2566 -341
rect 2626 -347 2684 -341
rect 2744 -347 2802 -341
rect 2862 -347 2920 -341
rect 2980 -347 3038 -341
rect 3098 -347 3156 -341
rect 3216 -347 3274 -341
rect 3334 -347 3392 -341
rect 3452 -347 3510 -341
rect 3570 -347 3628 -341
rect 3688 -347 3746 -341
rect 3806 -347 3864 -341
rect 3924 -347 3982 -341
rect 4042 -347 4100 -341
rect 4160 -347 4218 -341
rect 4278 -347 4336 -341
rect 4396 -347 4454 -341
rect 4514 -347 4572 -341
rect 4632 -347 4690 -341
rect 4750 -347 4808 -341
rect 4868 -347 4926 -341
rect 4986 -347 5044 -341
rect 5104 -347 5162 -341
rect 5222 -347 5280 -341
rect 5340 -347 5398 -341
rect 5458 -347 5516 -341
rect 5576 -347 5634 -341
rect 5694 -347 5752 -341
rect 5812 -347 5870 -341
rect 5930 -347 5988 -341
rect 6048 -347 6106 -341
rect 6166 -347 6224 -341
rect 6284 -347 6342 -341
rect 6402 -347 6460 -341
rect 6520 -347 6578 -341
rect 6638 -347 6696 -341
rect 6756 -347 6814 -341
rect 6874 -347 6932 -341
rect 6992 -347 7050 -341
rect 7110 -347 7168 -341
rect 7228 -347 7286 -341
rect 7346 -347 7404 -341
rect 7464 -347 7522 -341
rect 7582 -347 7640 -341
rect 7700 -347 7758 -341
rect 7818 -347 7876 -341
rect 7936 -347 7994 -341
rect 8054 -347 8112 -341
rect 8172 -347 8230 -341
rect 8290 -347 8348 -341
rect 8408 -347 8466 -341
rect 8526 -347 8584 -341
rect 8644 -347 8702 -341
rect 8762 -347 8820 -341
rect -8820 -381 -8808 -347
rect -8702 -381 -8690 -347
rect -8584 -381 -8572 -347
rect -8466 -381 -8454 -347
rect -8348 -381 -8336 -347
rect -8230 -381 -8218 -347
rect -8112 -381 -8100 -347
rect -7994 -381 -7982 -347
rect -7876 -381 -7864 -347
rect -7758 -381 -7746 -347
rect -7640 -381 -7628 -347
rect -7522 -381 -7510 -347
rect -7404 -381 -7392 -347
rect -7286 -381 -7274 -347
rect -7168 -381 -7156 -347
rect -7050 -381 -7038 -347
rect -6932 -381 -6920 -347
rect -6814 -381 -6802 -347
rect -6696 -381 -6684 -347
rect -6578 -381 -6566 -347
rect -6460 -381 -6448 -347
rect -6342 -381 -6330 -347
rect -6224 -381 -6212 -347
rect -6106 -381 -6094 -347
rect -5988 -381 -5976 -347
rect -5870 -381 -5858 -347
rect -5752 -381 -5740 -347
rect -5634 -381 -5622 -347
rect -5516 -381 -5504 -347
rect -5398 -381 -5386 -347
rect -5280 -381 -5268 -347
rect -5162 -381 -5150 -347
rect -5044 -381 -5032 -347
rect -4926 -381 -4914 -347
rect -4808 -381 -4796 -347
rect -4690 -381 -4678 -347
rect -4572 -381 -4560 -347
rect -4454 -381 -4442 -347
rect -4336 -381 -4324 -347
rect -4218 -381 -4206 -347
rect -4100 -381 -4088 -347
rect -3982 -381 -3970 -347
rect -3864 -381 -3852 -347
rect -3746 -381 -3734 -347
rect -3628 -381 -3616 -347
rect -3510 -381 -3498 -347
rect -3392 -381 -3380 -347
rect -3274 -381 -3262 -347
rect -3156 -381 -3144 -347
rect -3038 -381 -3026 -347
rect -2920 -381 -2908 -347
rect -2802 -381 -2790 -347
rect -2684 -381 -2672 -347
rect -2566 -381 -2554 -347
rect -2448 -381 -2436 -347
rect -2330 -381 -2318 -347
rect -2212 -381 -2200 -347
rect -2094 -381 -2082 -347
rect -1976 -381 -1964 -347
rect -1858 -381 -1846 -347
rect -1740 -381 -1728 -347
rect -1622 -381 -1610 -347
rect -1504 -381 -1492 -347
rect -1386 -381 -1374 -347
rect -1268 -381 -1256 -347
rect -1150 -381 -1138 -347
rect -1032 -381 -1020 -347
rect -914 -381 -902 -347
rect -796 -381 -784 -347
rect -678 -381 -666 -347
rect -560 -381 -548 -347
rect -442 -381 -430 -347
rect -324 -381 -312 -347
rect -206 -381 -194 -347
rect -88 -381 -76 -347
rect 30 -381 42 -347
rect 148 -381 160 -347
rect 266 -381 278 -347
rect 384 -381 396 -347
rect 502 -381 514 -347
rect 620 -381 632 -347
rect 738 -381 750 -347
rect 856 -381 868 -347
rect 974 -381 986 -347
rect 1092 -381 1104 -347
rect 1210 -381 1222 -347
rect 1328 -381 1340 -347
rect 1446 -381 1458 -347
rect 1564 -381 1576 -347
rect 1682 -381 1694 -347
rect 1800 -381 1812 -347
rect 1918 -381 1930 -347
rect 2036 -381 2048 -347
rect 2154 -381 2166 -347
rect 2272 -381 2284 -347
rect 2390 -381 2402 -347
rect 2508 -381 2520 -347
rect 2626 -381 2638 -347
rect 2744 -381 2756 -347
rect 2862 -381 2874 -347
rect 2980 -381 2992 -347
rect 3098 -381 3110 -347
rect 3216 -381 3228 -347
rect 3334 -381 3346 -347
rect 3452 -381 3464 -347
rect 3570 -381 3582 -347
rect 3688 -381 3700 -347
rect 3806 -381 3818 -347
rect 3924 -381 3936 -347
rect 4042 -381 4054 -347
rect 4160 -381 4172 -347
rect 4278 -381 4290 -347
rect 4396 -381 4408 -347
rect 4514 -381 4526 -347
rect 4632 -381 4644 -347
rect 4750 -381 4762 -347
rect 4868 -381 4880 -347
rect 4986 -381 4998 -347
rect 5104 -381 5116 -347
rect 5222 -381 5234 -347
rect 5340 -381 5352 -347
rect 5458 -381 5470 -347
rect 5576 -381 5588 -347
rect 5694 -381 5706 -347
rect 5812 -381 5824 -347
rect 5930 -381 5942 -347
rect 6048 -381 6060 -347
rect 6166 -381 6178 -347
rect 6284 -381 6296 -347
rect 6402 -381 6414 -347
rect 6520 -381 6532 -347
rect 6638 -381 6650 -347
rect 6756 -381 6768 -347
rect 6874 -381 6886 -347
rect 6992 -381 7004 -347
rect 7110 -381 7122 -347
rect 7228 -381 7240 -347
rect 7346 -381 7358 -347
rect 7464 -381 7476 -347
rect 7582 -381 7594 -347
rect 7700 -381 7712 -347
rect 7818 -381 7830 -347
rect 7936 -381 7948 -347
rect 8054 -381 8066 -347
rect 8172 -381 8184 -347
rect 8290 -381 8302 -347
rect 8408 -381 8420 -347
rect 8526 -381 8538 -347
rect 8644 -381 8656 -347
rect 8762 -381 8774 -347
rect -8820 -387 -8762 -381
rect -8702 -387 -8644 -381
rect -8584 -387 -8526 -381
rect -8466 -387 -8408 -381
rect -8348 -387 -8290 -381
rect -8230 -387 -8172 -381
rect -8112 -387 -8054 -381
rect -7994 -387 -7936 -381
rect -7876 -387 -7818 -381
rect -7758 -387 -7700 -381
rect -7640 -387 -7582 -381
rect -7522 -387 -7464 -381
rect -7404 -387 -7346 -381
rect -7286 -387 -7228 -381
rect -7168 -387 -7110 -381
rect -7050 -387 -6992 -381
rect -6932 -387 -6874 -381
rect -6814 -387 -6756 -381
rect -6696 -387 -6638 -381
rect -6578 -387 -6520 -381
rect -6460 -387 -6402 -381
rect -6342 -387 -6284 -381
rect -6224 -387 -6166 -381
rect -6106 -387 -6048 -381
rect -5988 -387 -5930 -381
rect -5870 -387 -5812 -381
rect -5752 -387 -5694 -381
rect -5634 -387 -5576 -381
rect -5516 -387 -5458 -381
rect -5398 -387 -5340 -381
rect -5280 -387 -5222 -381
rect -5162 -387 -5104 -381
rect -5044 -387 -4986 -381
rect -4926 -387 -4868 -381
rect -4808 -387 -4750 -381
rect -4690 -387 -4632 -381
rect -4572 -387 -4514 -381
rect -4454 -387 -4396 -381
rect -4336 -387 -4278 -381
rect -4218 -387 -4160 -381
rect -4100 -387 -4042 -381
rect -3982 -387 -3924 -381
rect -3864 -387 -3806 -381
rect -3746 -387 -3688 -381
rect -3628 -387 -3570 -381
rect -3510 -387 -3452 -381
rect -3392 -387 -3334 -381
rect -3274 -387 -3216 -381
rect -3156 -387 -3098 -381
rect -3038 -387 -2980 -381
rect -2920 -387 -2862 -381
rect -2802 -387 -2744 -381
rect -2684 -387 -2626 -381
rect -2566 -387 -2508 -381
rect -2448 -387 -2390 -381
rect -2330 -387 -2272 -381
rect -2212 -387 -2154 -381
rect -2094 -387 -2036 -381
rect -1976 -387 -1918 -381
rect -1858 -387 -1800 -381
rect -1740 -387 -1682 -381
rect -1622 -387 -1564 -381
rect -1504 -387 -1446 -381
rect -1386 -387 -1328 -381
rect -1268 -387 -1210 -381
rect -1150 -387 -1092 -381
rect -1032 -387 -974 -381
rect -914 -387 -856 -381
rect -796 -387 -738 -381
rect -678 -387 -620 -381
rect -560 -387 -502 -381
rect -442 -387 -384 -381
rect -324 -387 -266 -381
rect -206 -387 -148 -381
rect -88 -387 -30 -381
rect 30 -387 88 -381
rect 148 -387 206 -381
rect 266 -387 324 -381
rect 384 -387 442 -381
rect 502 -387 560 -381
rect 620 -387 678 -381
rect 738 -387 796 -381
rect 856 -387 914 -381
rect 974 -387 1032 -381
rect 1092 -387 1150 -381
rect 1210 -387 1268 -381
rect 1328 -387 1386 -381
rect 1446 -387 1504 -381
rect 1564 -387 1622 -381
rect 1682 -387 1740 -381
rect 1800 -387 1858 -381
rect 1918 -387 1976 -381
rect 2036 -387 2094 -381
rect 2154 -387 2212 -381
rect 2272 -387 2330 -381
rect 2390 -387 2448 -381
rect 2508 -387 2566 -381
rect 2626 -387 2684 -381
rect 2744 -387 2802 -381
rect 2862 -387 2920 -381
rect 2980 -387 3038 -381
rect 3098 -387 3156 -381
rect 3216 -387 3274 -381
rect 3334 -387 3392 -381
rect 3452 -387 3510 -381
rect 3570 -387 3628 -381
rect 3688 -387 3746 -381
rect 3806 -387 3864 -381
rect 3924 -387 3982 -381
rect 4042 -387 4100 -381
rect 4160 -387 4218 -381
rect 4278 -387 4336 -381
rect 4396 -387 4454 -381
rect 4514 -387 4572 -381
rect 4632 -387 4690 -381
rect 4750 -387 4808 -381
rect 4868 -387 4926 -381
rect 4986 -387 5044 -381
rect 5104 -387 5162 -381
rect 5222 -387 5280 -381
rect 5340 -387 5398 -381
rect 5458 -387 5516 -381
rect 5576 -387 5634 -381
rect 5694 -387 5752 -381
rect 5812 -387 5870 -381
rect 5930 -387 5988 -381
rect 6048 -387 6106 -381
rect 6166 -387 6224 -381
rect 6284 -387 6342 -381
rect 6402 -387 6460 -381
rect 6520 -387 6578 -381
rect 6638 -387 6696 -381
rect 6756 -387 6814 -381
rect 6874 -387 6932 -381
rect 6992 -387 7050 -381
rect 7110 -387 7168 -381
rect 7228 -387 7286 -381
rect 7346 -387 7404 -381
rect 7464 -387 7522 -381
rect 7582 -387 7640 -381
rect 7700 -387 7758 -381
rect 7818 -387 7876 -381
rect 7936 -387 7994 -381
rect 8054 -387 8112 -381
rect 8172 -387 8230 -381
rect 8290 -387 8348 -381
rect 8408 -387 8466 -381
rect 8526 -387 8584 -381
rect 8644 -387 8702 -381
rect 8762 -387 8820 -381
<< nwell >>
rect -9017 -519 9017 519
<< pmos >>
rect -8821 -300 -8761 300
rect -8703 -300 -8643 300
rect -8585 -300 -8525 300
rect -8467 -300 -8407 300
rect -8349 -300 -8289 300
rect -8231 -300 -8171 300
rect -8113 -300 -8053 300
rect -7995 -300 -7935 300
rect -7877 -300 -7817 300
rect -7759 -300 -7699 300
rect -7641 -300 -7581 300
rect -7523 -300 -7463 300
rect -7405 -300 -7345 300
rect -7287 -300 -7227 300
rect -7169 -300 -7109 300
rect -7051 -300 -6991 300
rect -6933 -300 -6873 300
rect -6815 -300 -6755 300
rect -6697 -300 -6637 300
rect -6579 -300 -6519 300
rect -6461 -300 -6401 300
rect -6343 -300 -6283 300
rect -6225 -300 -6165 300
rect -6107 -300 -6047 300
rect -5989 -300 -5929 300
rect -5871 -300 -5811 300
rect -5753 -300 -5693 300
rect -5635 -300 -5575 300
rect -5517 -300 -5457 300
rect -5399 -300 -5339 300
rect -5281 -300 -5221 300
rect -5163 -300 -5103 300
rect -5045 -300 -4985 300
rect -4927 -300 -4867 300
rect -4809 -300 -4749 300
rect -4691 -300 -4631 300
rect -4573 -300 -4513 300
rect -4455 -300 -4395 300
rect -4337 -300 -4277 300
rect -4219 -300 -4159 300
rect -4101 -300 -4041 300
rect -3983 -300 -3923 300
rect -3865 -300 -3805 300
rect -3747 -300 -3687 300
rect -3629 -300 -3569 300
rect -3511 -300 -3451 300
rect -3393 -300 -3333 300
rect -3275 -300 -3215 300
rect -3157 -300 -3097 300
rect -3039 -300 -2979 300
rect -2921 -300 -2861 300
rect -2803 -300 -2743 300
rect -2685 -300 -2625 300
rect -2567 -300 -2507 300
rect -2449 -300 -2389 300
rect -2331 -300 -2271 300
rect -2213 -300 -2153 300
rect -2095 -300 -2035 300
rect -1977 -300 -1917 300
rect -1859 -300 -1799 300
rect -1741 -300 -1681 300
rect -1623 -300 -1563 300
rect -1505 -300 -1445 300
rect -1387 -300 -1327 300
rect -1269 -300 -1209 300
rect -1151 -300 -1091 300
rect -1033 -300 -973 300
rect -915 -300 -855 300
rect -797 -300 -737 300
rect -679 -300 -619 300
rect -561 -300 -501 300
rect -443 -300 -383 300
rect -325 -300 -265 300
rect -207 -300 -147 300
rect -89 -300 -29 300
rect 29 -300 89 300
rect 147 -300 207 300
rect 265 -300 325 300
rect 383 -300 443 300
rect 501 -300 561 300
rect 619 -300 679 300
rect 737 -300 797 300
rect 855 -300 915 300
rect 973 -300 1033 300
rect 1091 -300 1151 300
rect 1209 -300 1269 300
rect 1327 -300 1387 300
rect 1445 -300 1505 300
rect 1563 -300 1623 300
rect 1681 -300 1741 300
rect 1799 -300 1859 300
rect 1917 -300 1977 300
rect 2035 -300 2095 300
rect 2153 -300 2213 300
rect 2271 -300 2331 300
rect 2389 -300 2449 300
rect 2507 -300 2567 300
rect 2625 -300 2685 300
rect 2743 -300 2803 300
rect 2861 -300 2921 300
rect 2979 -300 3039 300
rect 3097 -300 3157 300
rect 3215 -300 3275 300
rect 3333 -300 3393 300
rect 3451 -300 3511 300
rect 3569 -300 3629 300
rect 3687 -300 3747 300
rect 3805 -300 3865 300
rect 3923 -300 3983 300
rect 4041 -300 4101 300
rect 4159 -300 4219 300
rect 4277 -300 4337 300
rect 4395 -300 4455 300
rect 4513 -300 4573 300
rect 4631 -300 4691 300
rect 4749 -300 4809 300
rect 4867 -300 4927 300
rect 4985 -300 5045 300
rect 5103 -300 5163 300
rect 5221 -300 5281 300
rect 5339 -300 5399 300
rect 5457 -300 5517 300
rect 5575 -300 5635 300
rect 5693 -300 5753 300
rect 5811 -300 5871 300
rect 5929 -300 5989 300
rect 6047 -300 6107 300
rect 6165 -300 6225 300
rect 6283 -300 6343 300
rect 6401 -300 6461 300
rect 6519 -300 6579 300
rect 6637 -300 6697 300
rect 6755 -300 6815 300
rect 6873 -300 6933 300
rect 6991 -300 7051 300
rect 7109 -300 7169 300
rect 7227 -300 7287 300
rect 7345 -300 7405 300
rect 7463 -300 7523 300
rect 7581 -300 7641 300
rect 7699 -300 7759 300
rect 7817 -300 7877 300
rect 7935 -300 7995 300
rect 8053 -300 8113 300
rect 8171 -300 8231 300
rect 8289 -300 8349 300
rect 8407 -300 8467 300
rect 8525 -300 8585 300
rect 8643 -300 8703 300
rect 8761 -300 8821 300
<< pdiff >>
rect -8879 288 -8821 300
rect -8879 -288 -8867 288
rect -8833 -288 -8821 288
rect -8879 -300 -8821 -288
rect -8761 288 -8703 300
rect -8761 -288 -8749 288
rect -8715 -288 -8703 288
rect -8761 -300 -8703 -288
rect -8643 288 -8585 300
rect -8643 -288 -8631 288
rect -8597 -288 -8585 288
rect -8643 -300 -8585 -288
rect -8525 288 -8467 300
rect -8525 -288 -8513 288
rect -8479 -288 -8467 288
rect -8525 -300 -8467 -288
rect -8407 288 -8349 300
rect -8407 -288 -8395 288
rect -8361 -288 -8349 288
rect -8407 -300 -8349 -288
rect -8289 288 -8231 300
rect -8289 -288 -8277 288
rect -8243 -288 -8231 288
rect -8289 -300 -8231 -288
rect -8171 288 -8113 300
rect -8171 -288 -8159 288
rect -8125 -288 -8113 288
rect -8171 -300 -8113 -288
rect -8053 288 -7995 300
rect -8053 -288 -8041 288
rect -8007 -288 -7995 288
rect -8053 -300 -7995 -288
rect -7935 288 -7877 300
rect -7935 -288 -7923 288
rect -7889 -288 -7877 288
rect -7935 -300 -7877 -288
rect -7817 288 -7759 300
rect -7817 -288 -7805 288
rect -7771 -288 -7759 288
rect -7817 -300 -7759 -288
rect -7699 288 -7641 300
rect -7699 -288 -7687 288
rect -7653 -288 -7641 288
rect -7699 -300 -7641 -288
rect -7581 288 -7523 300
rect -7581 -288 -7569 288
rect -7535 -288 -7523 288
rect -7581 -300 -7523 -288
rect -7463 288 -7405 300
rect -7463 -288 -7451 288
rect -7417 -288 -7405 288
rect -7463 -300 -7405 -288
rect -7345 288 -7287 300
rect -7345 -288 -7333 288
rect -7299 -288 -7287 288
rect -7345 -300 -7287 -288
rect -7227 288 -7169 300
rect -7227 -288 -7215 288
rect -7181 -288 -7169 288
rect -7227 -300 -7169 -288
rect -7109 288 -7051 300
rect -7109 -288 -7097 288
rect -7063 -288 -7051 288
rect -7109 -300 -7051 -288
rect -6991 288 -6933 300
rect -6991 -288 -6979 288
rect -6945 -288 -6933 288
rect -6991 -300 -6933 -288
rect -6873 288 -6815 300
rect -6873 -288 -6861 288
rect -6827 -288 -6815 288
rect -6873 -300 -6815 -288
rect -6755 288 -6697 300
rect -6755 -288 -6743 288
rect -6709 -288 -6697 288
rect -6755 -300 -6697 -288
rect -6637 288 -6579 300
rect -6637 -288 -6625 288
rect -6591 -288 -6579 288
rect -6637 -300 -6579 -288
rect -6519 288 -6461 300
rect -6519 -288 -6507 288
rect -6473 -288 -6461 288
rect -6519 -300 -6461 -288
rect -6401 288 -6343 300
rect -6401 -288 -6389 288
rect -6355 -288 -6343 288
rect -6401 -300 -6343 -288
rect -6283 288 -6225 300
rect -6283 -288 -6271 288
rect -6237 -288 -6225 288
rect -6283 -300 -6225 -288
rect -6165 288 -6107 300
rect -6165 -288 -6153 288
rect -6119 -288 -6107 288
rect -6165 -300 -6107 -288
rect -6047 288 -5989 300
rect -6047 -288 -6035 288
rect -6001 -288 -5989 288
rect -6047 -300 -5989 -288
rect -5929 288 -5871 300
rect -5929 -288 -5917 288
rect -5883 -288 -5871 288
rect -5929 -300 -5871 -288
rect -5811 288 -5753 300
rect -5811 -288 -5799 288
rect -5765 -288 -5753 288
rect -5811 -300 -5753 -288
rect -5693 288 -5635 300
rect -5693 -288 -5681 288
rect -5647 -288 -5635 288
rect -5693 -300 -5635 -288
rect -5575 288 -5517 300
rect -5575 -288 -5563 288
rect -5529 -288 -5517 288
rect -5575 -300 -5517 -288
rect -5457 288 -5399 300
rect -5457 -288 -5445 288
rect -5411 -288 -5399 288
rect -5457 -300 -5399 -288
rect -5339 288 -5281 300
rect -5339 -288 -5327 288
rect -5293 -288 -5281 288
rect -5339 -300 -5281 -288
rect -5221 288 -5163 300
rect -5221 -288 -5209 288
rect -5175 -288 -5163 288
rect -5221 -300 -5163 -288
rect -5103 288 -5045 300
rect -5103 -288 -5091 288
rect -5057 -288 -5045 288
rect -5103 -300 -5045 -288
rect -4985 288 -4927 300
rect -4985 -288 -4973 288
rect -4939 -288 -4927 288
rect -4985 -300 -4927 -288
rect -4867 288 -4809 300
rect -4867 -288 -4855 288
rect -4821 -288 -4809 288
rect -4867 -300 -4809 -288
rect -4749 288 -4691 300
rect -4749 -288 -4737 288
rect -4703 -288 -4691 288
rect -4749 -300 -4691 -288
rect -4631 288 -4573 300
rect -4631 -288 -4619 288
rect -4585 -288 -4573 288
rect -4631 -300 -4573 -288
rect -4513 288 -4455 300
rect -4513 -288 -4501 288
rect -4467 -288 -4455 288
rect -4513 -300 -4455 -288
rect -4395 288 -4337 300
rect -4395 -288 -4383 288
rect -4349 -288 -4337 288
rect -4395 -300 -4337 -288
rect -4277 288 -4219 300
rect -4277 -288 -4265 288
rect -4231 -288 -4219 288
rect -4277 -300 -4219 -288
rect -4159 288 -4101 300
rect -4159 -288 -4147 288
rect -4113 -288 -4101 288
rect -4159 -300 -4101 -288
rect -4041 288 -3983 300
rect -4041 -288 -4029 288
rect -3995 -288 -3983 288
rect -4041 -300 -3983 -288
rect -3923 288 -3865 300
rect -3923 -288 -3911 288
rect -3877 -288 -3865 288
rect -3923 -300 -3865 -288
rect -3805 288 -3747 300
rect -3805 -288 -3793 288
rect -3759 -288 -3747 288
rect -3805 -300 -3747 -288
rect -3687 288 -3629 300
rect -3687 -288 -3675 288
rect -3641 -288 -3629 288
rect -3687 -300 -3629 -288
rect -3569 288 -3511 300
rect -3569 -288 -3557 288
rect -3523 -288 -3511 288
rect -3569 -300 -3511 -288
rect -3451 288 -3393 300
rect -3451 -288 -3439 288
rect -3405 -288 -3393 288
rect -3451 -300 -3393 -288
rect -3333 288 -3275 300
rect -3333 -288 -3321 288
rect -3287 -288 -3275 288
rect -3333 -300 -3275 -288
rect -3215 288 -3157 300
rect -3215 -288 -3203 288
rect -3169 -288 -3157 288
rect -3215 -300 -3157 -288
rect -3097 288 -3039 300
rect -3097 -288 -3085 288
rect -3051 -288 -3039 288
rect -3097 -300 -3039 -288
rect -2979 288 -2921 300
rect -2979 -288 -2967 288
rect -2933 -288 -2921 288
rect -2979 -300 -2921 -288
rect -2861 288 -2803 300
rect -2861 -288 -2849 288
rect -2815 -288 -2803 288
rect -2861 -300 -2803 -288
rect -2743 288 -2685 300
rect -2743 -288 -2731 288
rect -2697 -288 -2685 288
rect -2743 -300 -2685 -288
rect -2625 288 -2567 300
rect -2625 -288 -2613 288
rect -2579 -288 -2567 288
rect -2625 -300 -2567 -288
rect -2507 288 -2449 300
rect -2507 -288 -2495 288
rect -2461 -288 -2449 288
rect -2507 -300 -2449 -288
rect -2389 288 -2331 300
rect -2389 -288 -2377 288
rect -2343 -288 -2331 288
rect -2389 -300 -2331 -288
rect -2271 288 -2213 300
rect -2271 -288 -2259 288
rect -2225 -288 -2213 288
rect -2271 -300 -2213 -288
rect -2153 288 -2095 300
rect -2153 -288 -2141 288
rect -2107 -288 -2095 288
rect -2153 -300 -2095 -288
rect -2035 288 -1977 300
rect -2035 -288 -2023 288
rect -1989 -288 -1977 288
rect -2035 -300 -1977 -288
rect -1917 288 -1859 300
rect -1917 -288 -1905 288
rect -1871 -288 -1859 288
rect -1917 -300 -1859 -288
rect -1799 288 -1741 300
rect -1799 -288 -1787 288
rect -1753 -288 -1741 288
rect -1799 -300 -1741 -288
rect -1681 288 -1623 300
rect -1681 -288 -1669 288
rect -1635 -288 -1623 288
rect -1681 -300 -1623 -288
rect -1563 288 -1505 300
rect -1563 -288 -1551 288
rect -1517 -288 -1505 288
rect -1563 -300 -1505 -288
rect -1445 288 -1387 300
rect -1445 -288 -1433 288
rect -1399 -288 -1387 288
rect -1445 -300 -1387 -288
rect -1327 288 -1269 300
rect -1327 -288 -1315 288
rect -1281 -288 -1269 288
rect -1327 -300 -1269 -288
rect -1209 288 -1151 300
rect -1209 -288 -1197 288
rect -1163 -288 -1151 288
rect -1209 -300 -1151 -288
rect -1091 288 -1033 300
rect -1091 -288 -1079 288
rect -1045 -288 -1033 288
rect -1091 -300 -1033 -288
rect -973 288 -915 300
rect -973 -288 -961 288
rect -927 -288 -915 288
rect -973 -300 -915 -288
rect -855 288 -797 300
rect -855 -288 -843 288
rect -809 -288 -797 288
rect -855 -300 -797 -288
rect -737 288 -679 300
rect -737 -288 -725 288
rect -691 -288 -679 288
rect -737 -300 -679 -288
rect -619 288 -561 300
rect -619 -288 -607 288
rect -573 -288 -561 288
rect -619 -300 -561 -288
rect -501 288 -443 300
rect -501 -288 -489 288
rect -455 -288 -443 288
rect -501 -300 -443 -288
rect -383 288 -325 300
rect -383 -288 -371 288
rect -337 -288 -325 288
rect -383 -300 -325 -288
rect -265 288 -207 300
rect -265 -288 -253 288
rect -219 -288 -207 288
rect -265 -300 -207 -288
rect -147 288 -89 300
rect -147 -288 -135 288
rect -101 -288 -89 288
rect -147 -300 -89 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 89 288 147 300
rect 89 -288 101 288
rect 135 -288 147 288
rect 89 -300 147 -288
rect 207 288 265 300
rect 207 -288 219 288
rect 253 -288 265 288
rect 207 -300 265 -288
rect 325 288 383 300
rect 325 -288 337 288
rect 371 -288 383 288
rect 325 -300 383 -288
rect 443 288 501 300
rect 443 -288 455 288
rect 489 -288 501 288
rect 443 -300 501 -288
rect 561 288 619 300
rect 561 -288 573 288
rect 607 -288 619 288
rect 561 -300 619 -288
rect 679 288 737 300
rect 679 -288 691 288
rect 725 -288 737 288
rect 679 -300 737 -288
rect 797 288 855 300
rect 797 -288 809 288
rect 843 -288 855 288
rect 797 -300 855 -288
rect 915 288 973 300
rect 915 -288 927 288
rect 961 -288 973 288
rect 915 -300 973 -288
rect 1033 288 1091 300
rect 1033 -288 1045 288
rect 1079 -288 1091 288
rect 1033 -300 1091 -288
rect 1151 288 1209 300
rect 1151 -288 1163 288
rect 1197 -288 1209 288
rect 1151 -300 1209 -288
rect 1269 288 1327 300
rect 1269 -288 1281 288
rect 1315 -288 1327 288
rect 1269 -300 1327 -288
rect 1387 288 1445 300
rect 1387 -288 1399 288
rect 1433 -288 1445 288
rect 1387 -300 1445 -288
rect 1505 288 1563 300
rect 1505 -288 1517 288
rect 1551 -288 1563 288
rect 1505 -300 1563 -288
rect 1623 288 1681 300
rect 1623 -288 1635 288
rect 1669 -288 1681 288
rect 1623 -300 1681 -288
rect 1741 288 1799 300
rect 1741 -288 1753 288
rect 1787 -288 1799 288
rect 1741 -300 1799 -288
rect 1859 288 1917 300
rect 1859 -288 1871 288
rect 1905 -288 1917 288
rect 1859 -300 1917 -288
rect 1977 288 2035 300
rect 1977 -288 1989 288
rect 2023 -288 2035 288
rect 1977 -300 2035 -288
rect 2095 288 2153 300
rect 2095 -288 2107 288
rect 2141 -288 2153 288
rect 2095 -300 2153 -288
rect 2213 288 2271 300
rect 2213 -288 2225 288
rect 2259 -288 2271 288
rect 2213 -300 2271 -288
rect 2331 288 2389 300
rect 2331 -288 2343 288
rect 2377 -288 2389 288
rect 2331 -300 2389 -288
rect 2449 288 2507 300
rect 2449 -288 2461 288
rect 2495 -288 2507 288
rect 2449 -300 2507 -288
rect 2567 288 2625 300
rect 2567 -288 2579 288
rect 2613 -288 2625 288
rect 2567 -300 2625 -288
rect 2685 288 2743 300
rect 2685 -288 2697 288
rect 2731 -288 2743 288
rect 2685 -300 2743 -288
rect 2803 288 2861 300
rect 2803 -288 2815 288
rect 2849 -288 2861 288
rect 2803 -300 2861 -288
rect 2921 288 2979 300
rect 2921 -288 2933 288
rect 2967 -288 2979 288
rect 2921 -300 2979 -288
rect 3039 288 3097 300
rect 3039 -288 3051 288
rect 3085 -288 3097 288
rect 3039 -300 3097 -288
rect 3157 288 3215 300
rect 3157 -288 3169 288
rect 3203 -288 3215 288
rect 3157 -300 3215 -288
rect 3275 288 3333 300
rect 3275 -288 3287 288
rect 3321 -288 3333 288
rect 3275 -300 3333 -288
rect 3393 288 3451 300
rect 3393 -288 3405 288
rect 3439 -288 3451 288
rect 3393 -300 3451 -288
rect 3511 288 3569 300
rect 3511 -288 3523 288
rect 3557 -288 3569 288
rect 3511 -300 3569 -288
rect 3629 288 3687 300
rect 3629 -288 3641 288
rect 3675 -288 3687 288
rect 3629 -300 3687 -288
rect 3747 288 3805 300
rect 3747 -288 3759 288
rect 3793 -288 3805 288
rect 3747 -300 3805 -288
rect 3865 288 3923 300
rect 3865 -288 3877 288
rect 3911 -288 3923 288
rect 3865 -300 3923 -288
rect 3983 288 4041 300
rect 3983 -288 3995 288
rect 4029 -288 4041 288
rect 3983 -300 4041 -288
rect 4101 288 4159 300
rect 4101 -288 4113 288
rect 4147 -288 4159 288
rect 4101 -300 4159 -288
rect 4219 288 4277 300
rect 4219 -288 4231 288
rect 4265 -288 4277 288
rect 4219 -300 4277 -288
rect 4337 288 4395 300
rect 4337 -288 4349 288
rect 4383 -288 4395 288
rect 4337 -300 4395 -288
rect 4455 288 4513 300
rect 4455 -288 4467 288
rect 4501 -288 4513 288
rect 4455 -300 4513 -288
rect 4573 288 4631 300
rect 4573 -288 4585 288
rect 4619 -288 4631 288
rect 4573 -300 4631 -288
rect 4691 288 4749 300
rect 4691 -288 4703 288
rect 4737 -288 4749 288
rect 4691 -300 4749 -288
rect 4809 288 4867 300
rect 4809 -288 4821 288
rect 4855 -288 4867 288
rect 4809 -300 4867 -288
rect 4927 288 4985 300
rect 4927 -288 4939 288
rect 4973 -288 4985 288
rect 4927 -300 4985 -288
rect 5045 288 5103 300
rect 5045 -288 5057 288
rect 5091 -288 5103 288
rect 5045 -300 5103 -288
rect 5163 288 5221 300
rect 5163 -288 5175 288
rect 5209 -288 5221 288
rect 5163 -300 5221 -288
rect 5281 288 5339 300
rect 5281 -288 5293 288
rect 5327 -288 5339 288
rect 5281 -300 5339 -288
rect 5399 288 5457 300
rect 5399 -288 5411 288
rect 5445 -288 5457 288
rect 5399 -300 5457 -288
rect 5517 288 5575 300
rect 5517 -288 5529 288
rect 5563 -288 5575 288
rect 5517 -300 5575 -288
rect 5635 288 5693 300
rect 5635 -288 5647 288
rect 5681 -288 5693 288
rect 5635 -300 5693 -288
rect 5753 288 5811 300
rect 5753 -288 5765 288
rect 5799 -288 5811 288
rect 5753 -300 5811 -288
rect 5871 288 5929 300
rect 5871 -288 5883 288
rect 5917 -288 5929 288
rect 5871 -300 5929 -288
rect 5989 288 6047 300
rect 5989 -288 6001 288
rect 6035 -288 6047 288
rect 5989 -300 6047 -288
rect 6107 288 6165 300
rect 6107 -288 6119 288
rect 6153 -288 6165 288
rect 6107 -300 6165 -288
rect 6225 288 6283 300
rect 6225 -288 6237 288
rect 6271 -288 6283 288
rect 6225 -300 6283 -288
rect 6343 288 6401 300
rect 6343 -288 6355 288
rect 6389 -288 6401 288
rect 6343 -300 6401 -288
rect 6461 288 6519 300
rect 6461 -288 6473 288
rect 6507 -288 6519 288
rect 6461 -300 6519 -288
rect 6579 288 6637 300
rect 6579 -288 6591 288
rect 6625 -288 6637 288
rect 6579 -300 6637 -288
rect 6697 288 6755 300
rect 6697 -288 6709 288
rect 6743 -288 6755 288
rect 6697 -300 6755 -288
rect 6815 288 6873 300
rect 6815 -288 6827 288
rect 6861 -288 6873 288
rect 6815 -300 6873 -288
rect 6933 288 6991 300
rect 6933 -288 6945 288
rect 6979 -288 6991 288
rect 6933 -300 6991 -288
rect 7051 288 7109 300
rect 7051 -288 7063 288
rect 7097 -288 7109 288
rect 7051 -300 7109 -288
rect 7169 288 7227 300
rect 7169 -288 7181 288
rect 7215 -288 7227 288
rect 7169 -300 7227 -288
rect 7287 288 7345 300
rect 7287 -288 7299 288
rect 7333 -288 7345 288
rect 7287 -300 7345 -288
rect 7405 288 7463 300
rect 7405 -288 7417 288
rect 7451 -288 7463 288
rect 7405 -300 7463 -288
rect 7523 288 7581 300
rect 7523 -288 7535 288
rect 7569 -288 7581 288
rect 7523 -300 7581 -288
rect 7641 288 7699 300
rect 7641 -288 7653 288
rect 7687 -288 7699 288
rect 7641 -300 7699 -288
rect 7759 288 7817 300
rect 7759 -288 7771 288
rect 7805 -288 7817 288
rect 7759 -300 7817 -288
rect 7877 288 7935 300
rect 7877 -288 7889 288
rect 7923 -288 7935 288
rect 7877 -300 7935 -288
rect 7995 288 8053 300
rect 7995 -288 8007 288
rect 8041 -288 8053 288
rect 7995 -300 8053 -288
rect 8113 288 8171 300
rect 8113 -288 8125 288
rect 8159 -288 8171 288
rect 8113 -300 8171 -288
rect 8231 288 8289 300
rect 8231 -288 8243 288
rect 8277 -288 8289 288
rect 8231 -300 8289 -288
rect 8349 288 8407 300
rect 8349 -288 8361 288
rect 8395 -288 8407 288
rect 8349 -300 8407 -288
rect 8467 288 8525 300
rect 8467 -288 8479 288
rect 8513 -288 8525 288
rect 8467 -300 8525 -288
rect 8585 288 8643 300
rect 8585 -288 8597 288
rect 8631 -288 8643 288
rect 8585 -300 8643 -288
rect 8703 288 8761 300
rect 8703 -288 8715 288
rect 8749 -288 8761 288
rect 8703 -300 8761 -288
rect 8821 288 8879 300
rect 8821 -288 8833 288
rect 8867 -288 8879 288
rect 8821 -300 8879 -288
<< pdiffc >>
rect -8867 -288 -8833 288
rect -8749 -288 -8715 288
rect -8631 -288 -8597 288
rect -8513 -288 -8479 288
rect -8395 -288 -8361 288
rect -8277 -288 -8243 288
rect -8159 -288 -8125 288
rect -8041 -288 -8007 288
rect -7923 -288 -7889 288
rect -7805 -288 -7771 288
rect -7687 -288 -7653 288
rect -7569 -288 -7535 288
rect -7451 -288 -7417 288
rect -7333 -288 -7299 288
rect -7215 -288 -7181 288
rect -7097 -288 -7063 288
rect -6979 -288 -6945 288
rect -6861 -288 -6827 288
rect -6743 -288 -6709 288
rect -6625 -288 -6591 288
rect -6507 -288 -6473 288
rect -6389 -288 -6355 288
rect -6271 -288 -6237 288
rect -6153 -288 -6119 288
rect -6035 -288 -6001 288
rect -5917 -288 -5883 288
rect -5799 -288 -5765 288
rect -5681 -288 -5647 288
rect -5563 -288 -5529 288
rect -5445 -288 -5411 288
rect -5327 -288 -5293 288
rect -5209 -288 -5175 288
rect -5091 -288 -5057 288
rect -4973 -288 -4939 288
rect -4855 -288 -4821 288
rect -4737 -288 -4703 288
rect -4619 -288 -4585 288
rect -4501 -288 -4467 288
rect -4383 -288 -4349 288
rect -4265 -288 -4231 288
rect -4147 -288 -4113 288
rect -4029 -288 -3995 288
rect -3911 -288 -3877 288
rect -3793 -288 -3759 288
rect -3675 -288 -3641 288
rect -3557 -288 -3523 288
rect -3439 -288 -3405 288
rect -3321 -288 -3287 288
rect -3203 -288 -3169 288
rect -3085 -288 -3051 288
rect -2967 -288 -2933 288
rect -2849 -288 -2815 288
rect -2731 -288 -2697 288
rect -2613 -288 -2579 288
rect -2495 -288 -2461 288
rect -2377 -288 -2343 288
rect -2259 -288 -2225 288
rect -2141 -288 -2107 288
rect -2023 -288 -1989 288
rect -1905 -288 -1871 288
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
rect 1871 -288 1905 288
rect 1989 -288 2023 288
rect 2107 -288 2141 288
rect 2225 -288 2259 288
rect 2343 -288 2377 288
rect 2461 -288 2495 288
rect 2579 -288 2613 288
rect 2697 -288 2731 288
rect 2815 -288 2849 288
rect 2933 -288 2967 288
rect 3051 -288 3085 288
rect 3169 -288 3203 288
rect 3287 -288 3321 288
rect 3405 -288 3439 288
rect 3523 -288 3557 288
rect 3641 -288 3675 288
rect 3759 -288 3793 288
rect 3877 -288 3911 288
rect 3995 -288 4029 288
rect 4113 -288 4147 288
rect 4231 -288 4265 288
rect 4349 -288 4383 288
rect 4467 -288 4501 288
rect 4585 -288 4619 288
rect 4703 -288 4737 288
rect 4821 -288 4855 288
rect 4939 -288 4973 288
rect 5057 -288 5091 288
rect 5175 -288 5209 288
rect 5293 -288 5327 288
rect 5411 -288 5445 288
rect 5529 -288 5563 288
rect 5647 -288 5681 288
rect 5765 -288 5799 288
rect 5883 -288 5917 288
rect 6001 -288 6035 288
rect 6119 -288 6153 288
rect 6237 -288 6271 288
rect 6355 -288 6389 288
rect 6473 -288 6507 288
rect 6591 -288 6625 288
rect 6709 -288 6743 288
rect 6827 -288 6861 288
rect 6945 -288 6979 288
rect 7063 -288 7097 288
rect 7181 -288 7215 288
rect 7299 -288 7333 288
rect 7417 -288 7451 288
rect 7535 -288 7569 288
rect 7653 -288 7687 288
rect 7771 -288 7805 288
rect 7889 -288 7923 288
rect 8007 -288 8041 288
rect 8125 -288 8159 288
rect 8243 -288 8277 288
rect 8361 -288 8395 288
rect 8479 -288 8513 288
rect 8597 -288 8631 288
rect 8715 -288 8749 288
rect 8833 -288 8867 288
<< nsubdiff >>
rect -8981 449 -8885 483
rect 8885 449 8981 483
rect -8981 387 -8947 449
rect 8947 387 8981 449
rect -8981 -449 -8947 -387
rect 8947 -449 8981 -387
rect -8981 -483 -8885 -449
rect 8885 -483 8981 -449
<< nsubdiffcont >>
rect -8885 449 8885 483
rect -8981 -387 -8947 387
rect 8947 -387 8981 387
rect -8885 -483 8885 -449
<< poly >>
rect -8824 381 -8758 397
rect -8824 347 -8808 381
rect -8774 347 -8758 381
rect -8824 331 -8758 347
rect -8706 381 -8640 397
rect -8706 347 -8690 381
rect -8656 347 -8640 381
rect -8706 331 -8640 347
rect -8588 381 -8522 397
rect -8588 347 -8572 381
rect -8538 347 -8522 381
rect -8588 331 -8522 347
rect -8470 381 -8404 397
rect -8470 347 -8454 381
rect -8420 347 -8404 381
rect -8470 331 -8404 347
rect -8352 381 -8286 397
rect -8352 347 -8336 381
rect -8302 347 -8286 381
rect -8352 331 -8286 347
rect -8234 381 -8168 397
rect -8234 347 -8218 381
rect -8184 347 -8168 381
rect -8234 331 -8168 347
rect -8116 381 -8050 397
rect -8116 347 -8100 381
rect -8066 347 -8050 381
rect -8116 331 -8050 347
rect -7998 381 -7932 397
rect -7998 347 -7982 381
rect -7948 347 -7932 381
rect -7998 331 -7932 347
rect -7880 381 -7814 397
rect -7880 347 -7864 381
rect -7830 347 -7814 381
rect -7880 331 -7814 347
rect -7762 381 -7696 397
rect -7762 347 -7746 381
rect -7712 347 -7696 381
rect -7762 331 -7696 347
rect -7644 381 -7578 397
rect -7644 347 -7628 381
rect -7594 347 -7578 381
rect -7644 331 -7578 347
rect -7526 381 -7460 397
rect -7526 347 -7510 381
rect -7476 347 -7460 381
rect -7526 331 -7460 347
rect -7408 381 -7342 397
rect -7408 347 -7392 381
rect -7358 347 -7342 381
rect -7408 331 -7342 347
rect -7290 381 -7224 397
rect -7290 347 -7274 381
rect -7240 347 -7224 381
rect -7290 331 -7224 347
rect -7172 381 -7106 397
rect -7172 347 -7156 381
rect -7122 347 -7106 381
rect -7172 331 -7106 347
rect -7054 381 -6988 397
rect -7054 347 -7038 381
rect -7004 347 -6988 381
rect -7054 331 -6988 347
rect -6936 381 -6870 397
rect -6936 347 -6920 381
rect -6886 347 -6870 381
rect -6936 331 -6870 347
rect -6818 381 -6752 397
rect -6818 347 -6802 381
rect -6768 347 -6752 381
rect -6818 331 -6752 347
rect -6700 381 -6634 397
rect -6700 347 -6684 381
rect -6650 347 -6634 381
rect -6700 331 -6634 347
rect -6582 381 -6516 397
rect -6582 347 -6566 381
rect -6532 347 -6516 381
rect -6582 331 -6516 347
rect -6464 381 -6398 397
rect -6464 347 -6448 381
rect -6414 347 -6398 381
rect -6464 331 -6398 347
rect -6346 381 -6280 397
rect -6346 347 -6330 381
rect -6296 347 -6280 381
rect -6346 331 -6280 347
rect -6228 381 -6162 397
rect -6228 347 -6212 381
rect -6178 347 -6162 381
rect -6228 331 -6162 347
rect -6110 381 -6044 397
rect -6110 347 -6094 381
rect -6060 347 -6044 381
rect -6110 331 -6044 347
rect -5992 381 -5926 397
rect -5992 347 -5976 381
rect -5942 347 -5926 381
rect -5992 331 -5926 347
rect -5874 381 -5808 397
rect -5874 347 -5858 381
rect -5824 347 -5808 381
rect -5874 331 -5808 347
rect -5756 381 -5690 397
rect -5756 347 -5740 381
rect -5706 347 -5690 381
rect -5756 331 -5690 347
rect -5638 381 -5572 397
rect -5638 347 -5622 381
rect -5588 347 -5572 381
rect -5638 331 -5572 347
rect -5520 381 -5454 397
rect -5520 347 -5504 381
rect -5470 347 -5454 381
rect -5520 331 -5454 347
rect -5402 381 -5336 397
rect -5402 347 -5386 381
rect -5352 347 -5336 381
rect -5402 331 -5336 347
rect -5284 381 -5218 397
rect -5284 347 -5268 381
rect -5234 347 -5218 381
rect -5284 331 -5218 347
rect -5166 381 -5100 397
rect -5166 347 -5150 381
rect -5116 347 -5100 381
rect -5166 331 -5100 347
rect -5048 381 -4982 397
rect -5048 347 -5032 381
rect -4998 347 -4982 381
rect -5048 331 -4982 347
rect -4930 381 -4864 397
rect -4930 347 -4914 381
rect -4880 347 -4864 381
rect -4930 331 -4864 347
rect -4812 381 -4746 397
rect -4812 347 -4796 381
rect -4762 347 -4746 381
rect -4812 331 -4746 347
rect -4694 381 -4628 397
rect -4694 347 -4678 381
rect -4644 347 -4628 381
rect -4694 331 -4628 347
rect -4576 381 -4510 397
rect -4576 347 -4560 381
rect -4526 347 -4510 381
rect -4576 331 -4510 347
rect -4458 381 -4392 397
rect -4458 347 -4442 381
rect -4408 347 -4392 381
rect -4458 331 -4392 347
rect -4340 381 -4274 397
rect -4340 347 -4324 381
rect -4290 347 -4274 381
rect -4340 331 -4274 347
rect -4222 381 -4156 397
rect -4222 347 -4206 381
rect -4172 347 -4156 381
rect -4222 331 -4156 347
rect -4104 381 -4038 397
rect -4104 347 -4088 381
rect -4054 347 -4038 381
rect -4104 331 -4038 347
rect -3986 381 -3920 397
rect -3986 347 -3970 381
rect -3936 347 -3920 381
rect -3986 331 -3920 347
rect -3868 381 -3802 397
rect -3868 347 -3852 381
rect -3818 347 -3802 381
rect -3868 331 -3802 347
rect -3750 381 -3684 397
rect -3750 347 -3734 381
rect -3700 347 -3684 381
rect -3750 331 -3684 347
rect -3632 381 -3566 397
rect -3632 347 -3616 381
rect -3582 347 -3566 381
rect -3632 331 -3566 347
rect -3514 381 -3448 397
rect -3514 347 -3498 381
rect -3464 347 -3448 381
rect -3514 331 -3448 347
rect -3396 381 -3330 397
rect -3396 347 -3380 381
rect -3346 347 -3330 381
rect -3396 331 -3330 347
rect -3278 381 -3212 397
rect -3278 347 -3262 381
rect -3228 347 -3212 381
rect -3278 331 -3212 347
rect -3160 381 -3094 397
rect -3160 347 -3144 381
rect -3110 347 -3094 381
rect -3160 331 -3094 347
rect -3042 381 -2976 397
rect -3042 347 -3026 381
rect -2992 347 -2976 381
rect -3042 331 -2976 347
rect -2924 381 -2858 397
rect -2924 347 -2908 381
rect -2874 347 -2858 381
rect -2924 331 -2858 347
rect -2806 381 -2740 397
rect -2806 347 -2790 381
rect -2756 347 -2740 381
rect -2806 331 -2740 347
rect -2688 381 -2622 397
rect -2688 347 -2672 381
rect -2638 347 -2622 381
rect -2688 331 -2622 347
rect -2570 381 -2504 397
rect -2570 347 -2554 381
rect -2520 347 -2504 381
rect -2570 331 -2504 347
rect -2452 381 -2386 397
rect -2452 347 -2436 381
rect -2402 347 -2386 381
rect -2452 331 -2386 347
rect -2334 381 -2268 397
rect -2334 347 -2318 381
rect -2284 347 -2268 381
rect -2334 331 -2268 347
rect -2216 381 -2150 397
rect -2216 347 -2200 381
rect -2166 347 -2150 381
rect -2216 331 -2150 347
rect -2098 381 -2032 397
rect -2098 347 -2082 381
rect -2048 347 -2032 381
rect -2098 331 -2032 347
rect -1980 381 -1914 397
rect -1980 347 -1964 381
rect -1930 347 -1914 381
rect -1980 331 -1914 347
rect -1862 381 -1796 397
rect -1862 347 -1846 381
rect -1812 347 -1796 381
rect -1862 331 -1796 347
rect -1744 381 -1678 397
rect -1744 347 -1728 381
rect -1694 347 -1678 381
rect -1744 331 -1678 347
rect -1626 381 -1560 397
rect -1626 347 -1610 381
rect -1576 347 -1560 381
rect -1626 331 -1560 347
rect -1508 381 -1442 397
rect -1508 347 -1492 381
rect -1458 347 -1442 381
rect -1508 331 -1442 347
rect -1390 381 -1324 397
rect -1390 347 -1374 381
rect -1340 347 -1324 381
rect -1390 331 -1324 347
rect -1272 381 -1206 397
rect -1272 347 -1256 381
rect -1222 347 -1206 381
rect -1272 331 -1206 347
rect -1154 381 -1088 397
rect -1154 347 -1138 381
rect -1104 347 -1088 381
rect -1154 331 -1088 347
rect -1036 381 -970 397
rect -1036 347 -1020 381
rect -986 347 -970 381
rect -1036 331 -970 347
rect -918 381 -852 397
rect -918 347 -902 381
rect -868 347 -852 381
rect -918 331 -852 347
rect -800 381 -734 397
rect -800 347 -784 381
rect -750 347 -734 381
rect -800 331 -734 347
rect -682 381 -616 397
rect -682 347 -666 381
rect -632 347 -616 381
rect -682 331 -616 347
rect -564 381 -498 397
rect -564 347 -548 381
rect -514 347 -498 381
rect -564 331 -498 347
rect -446 381 -380 397
rect -446 347 -430 381
rect -396 347 -380 381
rect -446 331 -380 347
rect -328 381 -262 397
rect -328 347 -312 381
rect -278 347 -262 381
rect -328 331 -262 347
rect -210 381 -144 397
rect -210 347 -194 381
rect -160 347 -144 381
rect -210 331 -144 347
rect -92 381 -26 397
rect -92 347 -76 381
rect -42 347 -26 381
rect -92 331 -26 347
rect 26 381 92 397
rect 26 347 42 381
rect 76 347 92 381
rect 26 331 92 347
rect 144 381 210 397
rect 144 347 160 381
rect 194 347 210 381
rect 144 331 210 347
rect 262 381 328 397
rect 262 347 278 381
rect 312 347 328 381
rect 262 331 328 347
rect 380 381 446 397
rect 380 347 396 381
rect 430 347 446 381
rect 380 331 446 347
rect 498 381 564 397
rect 498 347 514 381
rect 548 347 564 381
rect 498 331 564 347
rect 616 381 682 397
rect 616 347 632 381
rect 666 347 682 381
rect 616 331 682 347
rect 734 381 800 397
rect 734 347 750 381
rect 784 347 800 381
rect 734 331 800 347
rect 852 381 918 397
rect 852 347 868 381
rect 902 347 918 381
rect 852 331 918 347
rect 970 381 1036 397
rect 970 347 986 381
rect 1020 347 1036 381
rect 970 331 1036 347
rect 1088 381 1154 397
rect 1088 347 1104 381
rect 1138 347 1154 381
rect 1088 331 1154 347
rect 1206 381 1272 397
rect 1206 347 1222 381
rect 1256 347 1272 381
rect 1206 331 1272 347
rect 1324 381 1390 397
rect 1324 347 1340 381
rect 1374 347 1390 381
rect 1324 331 1390 347
rect 1442 381 1508 397
rect 1442 347 1458 381
rect 1492 347 1508 381
rect 1442 331 1508 347
rect 1560 381 1626 397
rect 1560 347 1576 381
rect 1610 347 1626 381
rect 1560 331 1626 347
rect 1678 381 1744 397
rect 1678 347 1694 381
rect 1728 347 1744 381
rect 1678 331 1744 347
rect 1796 381 1862 397
rect 1796 347 1812 381
rect 1846 347 1862 381
rect 1796 331 1862 347
rect 1914 381 1980 397
rect 1914 347 1930 381
rect 1964 347 1980 381
rect 1914 331 1980 347
rect 2032 381 2098 397
rect 2032 347 2048 381
rect 2082 347 2098 381
rect 2032 331 2098 347
rect 2150 381 2216 397
rect 2150 347 2166 381
rect 2200 347 2216 381
rect 2150 331 2216 347
rect 2268 381 2334 397
rect 2268 347 2284 381
rect 2318 347 2334 381
rect 2268 331 2334 347
rect 2386 381 2452 397
rect 2386 347 2402 381
rect 2436 347 2452 381
rect 2386 331 2452 347
rect 2504 381 2570 397
rect 2504 347 2520 381
rect 2554 347 2570 381
rect 2504 331 2570 347
rect 2622 381 2688 397
rect 2622 347 2638 381
rect 2672 347 2688 381
rect 2622 331 2688 347
rect 2740 381 2806 397
rect 2740 347 2756 381
rect 2790 347 2806 381
rect 2740 331 2806 347
rect 2858 381 2924 397
rect 2858 347 2874 381
rect 2908 347 2924 381
rect 2858 331 2924 347
rect 2976 381 3042 397
rect 2976 347 2992 381
rect 3026 347 3042 381
rect 2976 331 3042 347
rect 3094 381 3160 397
rect 3094 347 3110 381
rect 3144 347 3160 381
rect 3094 331 3160 347
rect 3212 381 3278 397
rect 3212 347 3228 381
rect 3262 347 3278 381
rect 3212 331 3278 347
rect 3330 381 3396 397
rect 3330 347 3346 381
rect 3380 347 3396 381
rect 3330 331 3396 347
rect 3448 381 3514 397
rect 3448 347 3464 381
rect 3498 347 3514 381
rect 3448 331 3514 347
rect 3566 381 3632 397
rect 3566 347 3582 381
rect 3616 347 3632 381
rect 3566 331 3632 347
rect 3684 381 3750 397
rect 3684 347 3700 381
rect 3734 347 3750 381
rect 3684 331 3750 347
rect 3802 381 3868 397
rect 3802 347 3818 381
rect 3852 347 3868 381
rect 3802 331 3868 347
rect 3920 381 3986 397
rect 3920 347 3936 381
rect 3970 347 3986 381
rect 3920 331 3986 347
rect 4038 381 4104 397
rect 4038 347 4054 381
rect 4088 347 4104 381
rect 4038 331 4104 347
rect 4156 381 4222 397
rect 4156 347 4172 381
rect 4206 347 4222 381
rect 4156 331 4222 347
rect 4274 381 4340 397
rect 4274 347 4290 381
rect 4324 347 4340 381
rect 4274 331 4340 347
rect 4392 381 4458 397
rect 4392 347 4408 381
rect 4442 347 4458 381
rect 4392 331 4458 347
rect 4510 381 4576 397
rect 4510 347 4526 381
rect 4560 347 4576 381
rect 4510 331 4576 347
rect 4628 381 4694 397
rect 4628 347 4644 381
rect 4678 347 4694 381
rect 4628 331 4694 347
rect 4746 381 4812 397
rect 4746 347 4762 381
rect 4796 347 4812 381
rect 4746 331 4812 347
rect 4864 381 4930 397
rect 4864 347 4880 381
rect 4914 347 4930 381
rect 4864 331 4930 347
rect 4982 381 5048 397
rect 4982 347 4998 381
rect 5032 347 5048 381
rect 4982 331 5048 347
rect 5100 381 5166 397
rect 5100 347 5116 381
rect 5150 347 5166 381
rect 5100 331 5166 347
rect 5218 381 5284 397
rect 5218 347 5234 381
rect 5268 347 5284 381
rect 5218 331 5284 347
rect 5336 381 5402 397
rect 5336 347 5352 381
rect 5386 347 5402 381
rect 5336 331 5402 347
rect 5454 381 5520 397
rect 5454 347 5470 381
rect 5504 347 5520 381
rect 5454 331 5520 347
rect 5572 381 5638 397
rect 5572 347 5588 381
rect 5622 347 5638 381
rect 5572 331 5638 347
rect 5690 381 5756 397
rect 5690 347 5706 381
rect 5740 347 5756 381
rect 5690 331 5756 347
rect 5808 381 5874 397
rect 5808 347 5824 381
rect 5858 347 5874 381
rect 5808 331 5874 347
rect 5926 381 5992 397
rect 5926 347 5942 381
rect 5976 347 5992 381
rect 5926 331 5992 347
rect 6044 381 6110 397
rect 6044 347 6060 381
rect 6094 347 6110 381
rect 6044 331 6110 347
rect 6162 381 6228 397
rect 6162 347 6178 381
rect 6212 347 6228 381
rect 6162 331 6228 347
rect 6280 381 6346 397
rect 6280 347 6296 381
rect 6330 347 6346 381
rect 6280 331 6346 347
rect 6398 381 6464 397
rect 6398 347 6414 381
rect 6448 347 6464 381
rect 6398 331 6464 347
rect 6516 381 6582 397
rect 6516 347 6532 381
rect 6566 347 6582 381
rect 6516 331 6582 347
rect 6634 381 6700 397
rect 6634 347 6650 381
rect 6684 347 6700 381
rect 6634 331 6700 347
rect 6752 381 6818 397
rect 6752 347 6768 381
rect 6802 347 6818 381
rect 6752 331 6818 347
rect 6870 381 6936 397
rect 6870 347 6886 381
rect 6920 347 6936 381
rect 6870 331 6936 347
rect 6988 381 7054 397
rect 6988 347 7004 381
rect 7038 347 7054 381
rect 6988 331 7054 347
rect 7106 381 7172 397
rect 7106 347 7122 381
rect 7156 347 7172 381
rect 7106 331 7172 347
rect 7224 381 7290 397
rect 7224 347 7240 381
rect 7274 347 7290 381
rect 7224 331 7290 347
rect 7342 381 7408 397
rect 7342 347 7358 381
rect 7392 347 7408 381
rect 7342 331 7408 347
rect 7460 381 7526 397
rect 7460 347 7476 381
rect 7510 347 7526 381
rect 7460 331 7526 347
rect 7578 381 7644 397
rect 7578 347 7594 381
rect 7628 347 7644 381
rect 7578 331 7644 347
rect 7696 381 7762 397
rect 7696 347 7712 381
rect 7746 347 7762 381
rect 7696 331 7762 347
rect 7814 381 7880 397
rect 7814 347 7830 381
rect 7864 347 7880 381
rect 7814 331 7880 347
rect 7932 381 7998 397
rect 7932 347 7948 381
rect 7982 347 7998 381
rect 7932 331 7998 347
rect 8050 381 8116 397
rect 8050 347 8066 381
rect 8100 347 8116 381
rect 8050 331 8116 347
rect 8168 381 8234 397
rect 8168 347 8184 381
rect 8218 347 8234 381
rect 8168 331 8234 347
rect 8286 381 8352 397
rect 8286 347 8302 381
rect 8336 347 8352 381
rect 8286 331 8352 347
rect 8404 381 8470 397
rect 8404 347 8420 381
rect 8454 347 8470 381
rect 8404 331 8470 347
rect 8522 381 8588 397
rect 8522 347 8538 381
rect 8572 347 8588 381
rect 8522 331 8588 347
rect 8640 381 8706 397
rect 8640 347 8656 381
rect 8690 347 8706 381
rect 8640 331 8706 347
rect 8758 381 8824 397
rect 8758 347 8774 381
rect 8808 347 8824 381
rect 8758 331 8824 347
rect -8821 300 -8761 331
rect -8703 300 -8643 331
rect -8585 300 -8525 331
rect -8467 300 -8407 331
rect -8349 300 -8289 331
rect -8231 300 -8171 331
rect -8113 300 -8053 331
rect -7995 300 -7935 331
rect -7877 300 -7817 331
rect -7759 300 -7699 331
rect -7641 300 -7581 331
rect -7523 300 -7463 331
rect -7405 300 -7345 331
rect -7287 300 -7227 331
rect -7169 300 -7109 331
rect -7051 300 -6991 331
rect -6933 300 -6873 331
rect -6815 300 -6755 331
rect -6697 300 -6637 331
rect -6579 300 -6519 331
rect -6461 300 -6401 331
rect -6343 300 -6283 331
rect -6225 300 -6165 331
rect -6107 300 -6047 331
rect -5989 300 -5929 331
rect -5871 300 -5811 331
rect -5753 300 -5693 331
rect -5635 300 -5575 331
rect -5517 300 -5457 331
rect -5399 300 -5339 331
rect -5281 300 -5221 331
rect -5163 300 -5103 331
rect -5045 300 -4985 331
rect -4927 300 -4867 331
rect -4809 300 -4749 331
rect -4691 300 -4631 331
rect -4573 300 -4513 331
rect -4455 300 -4395 331
rect -4337 300 -4277 331
rect -4219 300 -4159 331
rect -4101 300 -4041 331
rect -3983 300 -3923 331
rect -3865 300 -3805 331
rect -3747 300 -3687 331
rect -3629 300 -3569 331
rect -3511 300 -3451 331
rect -3393 300 -3333 331
rect -3275 300 -3215 331
rect -3157 300 -3097 331
rect -3039 300 -2979 331
rect -2921 300 -2861 331
rect -2803 300 -2743 331
rect -2685 300 -2625 331
rect -2567 300 -2507 331
rect -2449 300 -2389 331
rect -2331 300 -2271 331
rect -2213 300 -2153 331
rect -2095 300 -2035 331
rect -1977 300 -1917 331
rect -1859 300 -1799 331
rect -1741 300 -1681 331
rect -1623 300 -1563 331
rect -1505 300 -1445 331
rect -1387 300 -1327 331
rect -1269 300 -1209 331
rect -1151 300 -1091 331
rect -1033 300 -973 331
rect -915 300 -855 331
rect -797 300 -737 331
rect -679 300 -619 331
rect -561 300 -501 331
rect -443 300 -383 331
rect -325 300 -265 331
rect -207 300 -147 331
rect -89 300 -29 331
rect 29 300 89 331
rect 147 300 207 331
rect 265 300 325 331
rect 383 300 443 331
rect 501 300 561 331
rect 619 300 679 331
rect 737 300 797 331
rect 855 300 915 331
rect 973 300 1033 331
rect 1091 300 1151 331
rect 1209 300 1269 331
rect 1327 300 1387 331
rect 1445 300 1505 331
rect 1563 300 1623 331
rect 1681 300 1741 331
rect 1799 300 1859 331
rect 1917 300 1977 331
rect 2035 300 2095 331
rect 2153 300 2213 331
rect 2271 300 2331 331
rect 2389 300 2449 331
rect 2507 300 2567 331
rect 2625 300 2685 331
rect 2743 300 2803 331
rect 2861 300 2921 331
rect 2979 300 3039 331
rect 3097 300 3157 331
rect 3215 300 3275 331
rect 3333 300 3393 331
rect 3451 300 3511 331
rect 3569 300 3629 331
rect 3687 300 3747 331
rect 3805 300 3865 331
rect 3923 300 3983 331
rect 4041 300 4101 331
rect 4159 300 4219 331
rect 4277 300 4337 331
rect 4395 300 4455 331
rect 4513 300 4573 331
rect 4631 300 4691 331
rect 4749 300 4809 331
rect 4867 300 4927 331
rect 4985 300 5045 331
rect 5103 300 5163 331
rect 5221 300 5281 331
rect 5339 300 5399 331
rect 5457 300 5517 331
rect 5575 300 5635 331
rect 5693 300 5753 331
rect 5811 300 5871 331
rect 5929 300 5989 331
rect 6047 300 6107 331
rect 6165 300 6225 331
rect 6283 300 6343 331
rect 6401 300 6461 331
rect 6519 300 6579 331
rect 6637 300 6697 331
rect 6755 300 6815 331
rect 6873 300 6933 331
rect 6991 300 7051 331
rect 7109 300 7169 331
rect 7227 300 7287 331
rect 7345 300 7405 331
rect 7463 300 7523 331
rect 7581 300 7641 331
rect 7699 300 7759 331
rect 7817 300 7877 331
rect 7935 300 7995 331
rect 8053 300 8113 331
rect 8171 300 8231 331
rect 8289 300 8349 331
rect 8407 300 8467 331
rect 8525 300 8585 331
rect 8643 300 8703 331
rect 8761 300 8821 331
rect -8821 -331 -8761 -300
rect -8703 -331 -8643 -300
rect -8585 -331 -8525 -300
rect -8467 -331 -8407 -300
rect -8349 -331 -8289 -300
rect -8231 -331 -8171 -300
rect -8113 -331 -8053 -300
rect -7995 -331 -7935 -300
rect -7877 -331 -7817 -300
rect -7759 -331 -7699 -300
rect -7641 -331 -7581 -300
rect -7523 -331 -7463 -300
rect -7405 -331 -7345 -300
rect -7287 -331 -7227 -300
rect -7169 -331 -7109 -300
rect -7051 -331 -6991 -300
rect -6933 -331 -6873 -300
rect -6815 -331 -6755 -300
rect -6697 -331 -6637 -300
rect -6579 -331 -6519 -300
rect -6461 -331 -6401 -300
rect -6343 -331 -6283 -300
rect -6225 -331 -6165 -300
rect -6107 -331 -6047 -300
rect -5989 -331 -5929 -300
rect -5871 -331 -5811 -300
rect -5753 -331 -5693 -300
rect -5635 -331 -5575 -300
rect -5517 -331 -5457 -300
rect -5399 -331 -5339 -300
rect -5281 -331 -5221 -300
rect -5163 -331 -5103 -300
rect -5045 -331 -4985 -300
rect -4927 -331 -4867 -300
rect -4809 -331 -4749 -300
rect -4691 -331 -4631 -300
rect -4573 -331 -4513 -300
rect -4455 -331 -4395 -300
rect -4337 -331 -4277 -300
rect -4219 -331 -4159 -300
rect -4101 -331 -4041 -300
rect -3983 -331 -3923 -300
rect -3865 -331 -3805 -300
rect -3747 -331 -3687 -300
rect -3629 -331 -3569 -300
rect -3511 -331 -3451 -300
rect -3393 -331 -3333 -300
rect -3275 -331 -3215 -300
rect -3157 -331 -3097 -300
rect -3039 -331 -2979 -300
rect -2921 -331 -2861 -300
rect -2803 -331 -2743 -300
rect -2685 -331 -2625 -300
rect -2567 -331 -2507 -300
rect -2449 -331 -2389 -300
rect -2331 -331 -2271 -300
rect -2213 -331 -2153 -300
rect -2095 -331 -2035 -300
rect -1977 -331 -1917 -300
rect -1859 -331 -1799 -300
rect -1741 -331 -1681 -300
rect -1623 -331 -1563 -300
rect -1505 -331 -1445 -300
rect -1387 -331 -1327 -300
rect -1269 -331 -1209 -300
rect -1151 -331 -1091 -300
rect -1033 -331 -973 -300
rect -915 -331 -855 -300
rect -797 -331 -737 -300
rect -679 -331 -619 -300
rect -561 -331 -501 -300
rect -443 -331 -383 -300
rect -325 -331 -265 -300
rect -207 -331 -147 -300
rect -89 -331 -29 -300
rect 29 -331 89 -300
rect 147 -331 207 -300
rect 265 -331 325 -300
rect 383 -331 443 -300
rect 501 -331 561 -300
rect 619 -331 679 -300
rect 737 -331 797 -300
rect 855 -331 915 -300
rect 973 -331 1033 -300
rect 1091 -331 1151 -300
rect 1209 -331 1269 -300
rect 1327 -331 1387 -300
rect 1445 -331 1505 -300
rect 1563 -331 1623 -300
rect 1681 -331 1741 -300
rect 1799 -331 1859 -300
rect 1917 -331 1977 -300
rect 2035 -331 2095 -300
rect 2153 -331 2213 -300
rect 2271 -331 2331 -300
rect 2389 -331 2449 -300
rect 2507 -331 2567 -300
rect 2625 -331 2685 -300
rect 2743 -331 2803 -300
rect 2861 -331 2921 -300
rect 2979 -331 3039 -300
rect 3097 -331 3157 -300
rect 3215 -331 3275 -300
rect 3333 -331 3393 -300
rect 3451 -331 3511 -300
rect 3569 -331 3629 -300
rect 3687 -331 3747 -300
rect 3805 -331 3865 -300
rect 3923 -331 3983 -300
rect 4041 -331 4101 -300
rect 4159 -331 4219 -300
rect 4277 -331 4337 -300
rect 4395 -331 4455 -300
rect 4513 -331 4573 -300
rect 4631 -331 4691 -300
rect 4749 -331 4809 -300
rect 4867 -331 4927 -300
rect 4985 -331 5045 -300
rect 5103 -331 5163 -300
rect 5221 -331 5281 -300
rect 5339 -331 5399 -300
rect 5457 -331 5517 -300
rect 5575 -331 5635 -300
rect 5693 -331 5753 -300
rect 5811 -331 5871 -300
rect 5929 -331 5989 -300
rect 6047 -331 6107 -300
rect 6165 -331 6225 -300
rect 6283 -331 6343 -300
rect 6401 -331 6461 -300
rect 6519 -331 6579 -300
rect 6637 -331 6697 -300
rect 6755 -331 6815 -300
rect 6873 -331 6933 -300
rect 6991 -331 7051 -300
rect 7109 -331 7169 -300
rect 7227 -331 7287 -300
rect 7345 -331 7405 -300
rect 7463 -331 7523 -300
rect 7581 -331 7641 -300
rect 7699 -331 7759 -300
rect 7817 -331 7877 -300
rect 7935 -331 7995 -300
rect 8053 -331 8113 -300
rect 8171 -331 8231 -300
rect 8289 -331 8349 -300
rect 8407 -331 8467 -300
rect 8525 -331 8585 -300
rect 8643 -331 8703 -300
rect 8761 -331 8821 -300
rect -8824 -347 -8758 -331
rect -8824 -381 -8808 -347
rect -8774 -381 -8758 -347
rect -8824 -397 -8758 -381
rect -8706 -347 -8640 -331
rect -8706 -381 -8690 -347
rect -8656 -381 -8640 -347
rect -8706 -397 -8640 -381
rect -8588 -347 -8522 -331
rect -8588 -381 -8572 -347
rect -8538 -381 -8522 -347
rect -8588 -397 -8522 -381
rect -8470 -347 -8404 -331
rect -8470 -381 -8454 -347
rect -8420 -381 -8404 -347
rect -8470 -397 -8404 -381
rect -8352 -347 -8286 -331
rect -8352 -381 -8336 -347
rect -8302 -381 -8286 -347
rect -8352 -397 -8286 -381
rect -8234 -347 -8168 -331
rect -8234 -381 -8218 -347
rect -8184 -381 -8168 -347
rect -8234 -397 -8168 -381
rect -8116 -347 -8050 -331
rect -8116 -381 -8100 -347
rect -8066 -381 -8050 -347
rect -8116 -397 -8050 -381
rect -7998 -347 -7932 -331
rect -7998 -381 -7982 -347
rect -7948 -381 -7932 -347
rect -7998 -397 -7932 -381
rect -7880 -347 -7814 -331
rect -7880 -381 -7864 -347
rect -7830 -381 -7814 -347
rect -7880 -397 -7814 -381
rect -7762 -347 -7696 -331
rect -7762 -381 -7746 -347
rect -7712 -381 -7696 -347
rect -7762 -397 -7696 -381
rect -7644 -347 -7578 -331
rect -7644 -381 -7628 -347
rect -7594 -381 -7578 -347
rect -7644 -397 -7578 -381
rect -7526 -347 -7460 -331
rect -7526 -381 -7510 -347
rect -7476 -381 -7460 -347
rect -7526 -397 -7460 -381
rect -7408 -347 -7342 -331
rect -7408 -381 -7392 -347
rect -7358 -381 -7342 -347
rect -7408 -397 -7342 -381
rect -7290 -347 -7224 -331
rect -7290 -381 -7274 -347
rect -7240 -381 -7224 -347
rect -7290 -397 -7224 -381
rect -7172 -347 -7106 -331
rect -7172 -381 -7156 -347
rect -7122 -381 -7106 -347
rect -7172 -397 -7106 -381
rect -7054 -347 -6988 -331
rect -7054 -381 -7038 -347
rect -7004 -381 -6988 -347
rect -7054 -397 -6988 -381
rect -6936 -347 -6870 -331
rect -6936 -381 -6920 -347
rect -6886 -381 -6870 -347
rect -6936 -397 -6870 -381
rect -6818 -347 -6752 -331
rect -6818 -381 -6802 -347
rect -6768 -381 -6752 -347
rect -6818 -397 -6752 -381
rect -6700 -347 -6634 -331
rect -6700 -381 -6684 -347
rect -6650 -381 -6634 -347
rect -6700 -397 -6634 -381
rect -6582 -347 -6516 -331
rect -6582 -381 -6566 -347
rect -6532 -381 -6516 -347
rect -6582 -397 -6516 -381
rect -6464 -347 -6398 -331
rect -6464 -381 -6448 -347
rect -6414 -381 -6398 -347
rect -6464 -397 -6398 -381
rect -6346 -347 -6280 -331
rect -6346 -381 -6330 -347
rect -6296 -381 -6280 -347
rect -6346 -397 -6280 -381
rect -6228 -347 -6162 -331
rect -6228 -381 -6212 -347
rect -6178 -381 -6162 -347
rect -6228 -397 -6162 -381
rect -6110 -347 -6044 -331
rect -6110 -381 -6094 -347
rect -6060 -381 -6044 -347
rect -6110 -397 -6044 -381
rect -5992 -347 -5926 -331
rect -5992 -381 -5976 -347
rect -5942 -381 -5926 -347
rect -5992 -397 -5926 -381
rect -5874 -347 -5808 -331
rect -5874 -381 -5858 -347
rect -5824 -381 -5808 -347
rect -5874 -397 -5808 -381
rect -5756 -347 -5690 -331
rect -5756 -381 -5740 -347
rect -5706 -381 -5690 -347
rect -5756 -397 -5690 -381
rect -5638 -347 -5572 -331
rect -5638 -381 -5622 -347
rect -5588 -381 -5572 -347
rect -5638 -397 -5572 -381
rect -5520 -347 -5454 -331
rect -5520 -381 -5504 -347
rect -5470 -381 -5454 -347
rect -5520 -397 -5454 -381
rect -5402 -347 -5336 -331
rect -5402 -381 -5386 -347
rect -5352 -381 -5336 -347
rect -5402 -397 -5336 -381
rect -5284 -347 -5218 -331
rect -5284 -381 -5268 -347
rect -5234 -381 -5218 -347
rect -5284 -397 -5218 -381
rect -5166 -347 -5100 -331
rect -5166 -381 -5150 -347
rect -5116 -381 -5100 -347
rect -5166 -397 -5100 -381
rect -5048 -347 -4982 -331
rect -5048 -381 -5032 -347
rect -4998 -381 -4982 -347
rect -5048 -397 -4982 -381
rect -4930 -347 -4864 -331
rect -4930 -381 -4914 -347
rect -4880 -381 -4864 -347
rect -4930 -397 -4864 -381
rect -4812 -347 -4746 -331
rect -4812 -381 -4796 -347
rect -4762 -381 -4746 -347
rect -4812 -397 -4746 -381
rect -4694 -347 -4628 -331
rect -4694 -381 -4678 -347
rect -4644 -381 -4628 -347
rect -4694 -397 -4628 -381
rect -4576 -347 -4510 -331
rect -4576 -381 -4560 -347
rect -4526 -381 -4510 -347
rect -4576 -397 -4510 -381
rect -4458 -347 -4392 -331
rect -4458 -381 -4442 -347
rect -4408 -381 -4392 -347
rect -4458 -397 -4392 -381
rect -4340 -347 -4274 -331
rect -4340 -381 -4324 -347
rect -4290 -381 -4274 -347
rect -4340 -397 -4274 -381
rect -4222 -347 -4156 -331
rect -4222 -381 -4206 -347
rect -4172 -381 -4156 -347
rect -4222 -397 -4156 -381
rect -4104 -347 -4038 -331
rect -4104 -381 -4088 -347
rect -4054 -381 -4038 -347
rect -4104 -397 -4038 -381
rect -3986 -347 -3920 -331
rect -3986 -381 -3970 -347
rect -3936 -381 -3920 -347
rect -3986 -397 -3920 -381
rect -3868 -347 -3802 -331
rect -3868 -381 -3852 -347
rect -3818 -381 -3802 -347
rect -3868 -397 -3802 -381
rect -3750 -347 -3684 -331
rect -3750 -381 -3734 -347
rect -3700 -381 -3684 -347
rect -3750 -397 -3684 -381
rect -3632 -347 -3566 -331
rect -3632 -381 -3616 -347
rect -3582 -381 -3566 -347
rect -3632 -397 -3566 -381
rect -3514 -347 -3448 -331
rect -3514 -381 -3498 -347
rect -3464 -381 -3448 -347
rect -3514 -397 -3448 -381
rect -3396 -347 -3330 -331
rect -3396 -381 -3380 -347
rect -3346 -381 -3330 -347
rect -3396 -397 -3330 -381
rect -3278 -347 -3212 -331
rect -3278 -381 -3262 -347
rect -3228 -381 -3212 -347
rect -3278 -397 -3212 -381
rect -3160 -347 -3094 -331
rect -3160 -381 -3144 -347
rect -3110 -381 -3094 -347
rect -3160 -397 -3094 -381
rect -3042 -347 -2976 -331
rect -3042 -381 -3026 -347
rect -2992 -381 -2976 -347
rect -3042 -397 -2976 -381
rect -2924 -347 -2858 -331
rect -2924 -381 -2908 -347
rect -2874 -381 -2858 -347
rect -2924 -397 -2858 -381
rect -2806 -347 -2740 -331
rect -2806 -381 -2790 -347
rect -2756 -381 -2740 -347
rect -2806 -397 -2740 -381
rect -2688 -347 -2622 -331
rect -2688 -381 -2672 -347
rect -2638 -381 -2622 -347
rect -2688 -397 -2622 -381
rect -2570 -347 -2504 -331
rect -2570 -381 -2554 -347
rect -2520 -381 -2504 -347
rect -2570 -397 -2504 -381
rect -2452 -347 -2386 -331
rect -2452 -381 -2436 -347
rect -2402 -381 -2386 -347
rect -2452 -397 -2386 -381
rect -2334 -347 -2268 -331
rect -2334 -381 -2318 -347
rect -2284 -381 -2268 -347
rect -2334 -397 -2268 -381
rect -2216 -347 -2150 -331
rect -2216 -381 -2200 -347
rect -2166 -381 -2150 -347
rect -2216 -397 -2150 -381
rect -2098 -347 -2032 -331
rect -2098 -381 -2082 -347
rect -2048 -381 -2032 -347
rect -2098 -397 -2032 -381
rect -1980 -347 -1914 -331
rect -1980 -381 -1964 -347
rect -1930 -381 -1914 -347
rect -1980 -397 -1914 -381
rect -1862 -347 -1796 -331
rect -1862 -381 -1846 -347
rect -1812 -381 -1796 -347
rect -1862 -397 -1796 -381
rect -1744 -347 -1678 -331
rect -1744 -381 -1728 -347
rect -1694 -381 -1678 -347
rect -1744 -397 -1678 -381
rect -1626 -347 -1560 -331
rect -1626 -381 -1610 -347
rect -1576 -381 -1560 -347
rect -1626 -397 -1560 -381
rect -1508 -347 -1442 -331
rect -1508 -381 -1492 -347
rect -1458 -381 -1442 -347
rect -1508 -397 -1442 -381
rect -1390 -347 -1324 -331
rect -1390 -381 -1374 -347
rect -1340 -381 -1324 -347
rect -1390 -397 -1324 -381
rect -1272 -347 -1206 -331
rect -1272 -381 -1256 -347
rect -1222 -381 -1206 -347
rect -1272 -397 -1206 -381
rect -1154 -347 -1088 -331
rect -1154 -381 -1138 -347
rect -1104 -381 -1088 -347
rect -1154 -397 -1088 -381
rect -1036 -347 -970 -331
rect -1036 -381 -1020 -347
rect -986 -381 -970 -347
rect -1036 -397 -970 -381
rect -918 -347 -852 -331
rect -918 -381 -902 -347
rect -868 -381 -852 -347
rect -918 -397 -852 -381
rect -800 -347 -734 -331
rect -800 -381 -784 -347
rect -750 -381 -734 -347
rect -800 -397 -734 -381
rect -682 -347 -616 -331
rect -682 -381 -666 -347
rect -632 -381 -616 -347
rect -682 -397 -616 -381
rect -564 -347 -498 -331
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -564 -397 -498 -381
rect -446 -347 -380 -331
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -446 -397 -380 -381
rect -328 -347 -262 -331
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -328 -397 -262 -381
rect -210 -347 -144 -331
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -210 -397 -144 -381
rect -92 -347 -26 -331
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect -92 -397 -26 -381
rect 26 -347 92 -331
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 26 -397 92 -381
rect 144 -347 210 -331
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 144 -397 210 -381
rect 262 -347 328 -331
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 262 -397 328 -381
rect 380 -347 446 -331
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 380 -397 446 -381
rect 498 -347 564 -331
rect 498 -381 514 -347
rect 548 -381 564 -347
rect 498 -397 564 -381
rect 616 -347 682 -331
rect 616 -381 632 -347
rect 666 -381 682 -347
rect 616 -397 682 -381
rect 734 -347 800 -331
rect 734 -381 750 -347
rect 784 -381 800 -347
rect 734 -397 800 -381
rect 852 -347 918 -331
rect 852 -381 868 -347
rect 902 -381 918 -347
rect 852 -397 918 -381
rect 970 -347 1036 -331
rect 970 -381 986 -347
rect 1020 -381 1036 -347
rect 970 -397 1036 -381
rect 1088 -347 1154 -331
rect 1088 -381 1104 -347
rect 1138 -381 1154 -347
rect 1088 -397 1154 -381
rect 1206 -347 1272 -331
rect 1206 -381 1222 -347
rect 1256 -381 1272 -347
rect 1206 -397 1272 -381
rect 1324 -347 1390 -331
rect 1324 -381 1340 -347
rect 1374 -381 1390 -347
rect 1324 -397 1390 -381
rect 1442 -347 1508 -331
rect 1442 -381 1458 -347
rect 1492 -381 1508 -347
rect 1442 -397 1508 -381
rect 1560 -347 1626 -331
rect 1560 -381 1576 -347
rect 1610 -381 1626 -347
rect 1560 -397 1626 -381
rect 1678 -347 1744 -331
rect 1678 -381 1694 -347
rect 1728 -381 1744 -347
rect 1678 -397 1744 -381
rect 1796 -347 1862 -331
rect 1796 -381 1812 -347
rect 1846 -381 1862 -347
rect 1796 -397 1862 -381
rect 1914 -347 1980 -331
rect 1914 -381 1930 -347
rect 1964 -381 1980 -347
rect 1914 -397 1980 -381
rect 2032 -347 2098 -331
rect 2032 -381 2048 -347
rect 2082 -381 2098 -347
rect 2032 -397 2098 -381
rect 2150 -347 2216 -331
rect 2150 -381 2166 -347
rect 2200 -381 2216 -347
rect 2150 -397 2216 -381
rect 2268 -347 2334 -331
rect 2268 -381 2284 -347
rect 2318 -381 2334 -347
rect 2268 -397 2334 -381
rect 2386 -347 2452 -331
rect 2386 -381 2402 -347
rect 2436 -381 2452 -347
rect 2386 -397 2452 -381
rect 2504 -347 2570 -331
rect 2504 -381 2520 -347
rect 2554 -381 2570 -347
rect 2504 -397 2570 -381
rect 2622 -347 2688 -331
rect 2622 -381 2638 -347
rect 2672 -381 2688 -347
rect 2622 -397 2688 -381
rect 2740 -347 2806 -331
rect 2740 -381 2756 -347
rect 2790 -381 2806 -347
rect 2740 -397 2806 -381
rect 2858 -347 2924 -331
rect 2858 -381 2874 -347
rect 2908 -381 2924 -347
rect 2858 -397 2924 -381
rect 2976 -347 3042 -331
rect 2976 -381 2992 -347
rect 3026 -381 3042 -347
rect 2976 -397 3042 -381
rect 3094 -347 3160 -331
rect 3094 -381 3110 -347
rect 3144 -381 3160 -347
rect 3094 -397 3160 -381
rect 3212 -347 3278 -331
rect 3212 -381 3228 -347
rect 3262 -381 3278 -347
rect 3212 -397 3278 -381
rect 3330 -347 3396 -331
rect 3330 -381 3346 -347
rect 3380 -381 3396 -347
rect 3330 -397 3396 -381
rect 3448 -347 3514 -331
rect 3448 -381 3464 -347
rect 3498 -381 3514 -347
rect 3448 -397 3514 -381
rect 3566 -347 3632 -331
rect 3566 -381 3582 -347
rect 3616 -381 3632 -347
rect 3566 -397 3632 -381
rect 3684 -347 3750 -331
rect 3684 -381 3700 -347
rect 3734 -381 3750 -347
rect 3684 -397 3750 -381
rect 3802 -347 3868 -331
rect 3802 -381 3818 -347
rect 3852 -381 3868 -347
rect 3802 -397 3868 -381
rect 3920 -347 3986 -331
rect 3920 -381 3936 -347
rect 3970 -381 3986 -347
rect 3920 -397 3986 -381
rect 4038 -347 4104 -331
rect 4038 -381 4054 -347
rect 4088 -381 4104 -347
rect 4038 -397 4104 -381
rect 4156 -347 4222 -331
rect 4156 -381 4172 -347
rect 4206 -381 4222 -347
rect 4156 -397 4222 -381
rect 4274 -347 4340 -331
rect 4274 -381 4290 -347
rect 4324 -381 4340 -347
rect 4274 -397 4340 -381
rect 4392 -347 4458 -331
rect 4392 -381 4408 -347
rect 4442 -381 4458 -347
rect 4392 -397 4458 -381
rect 4510 -347 4576 -331
rect 4510 -381 4526 -347
rect 4560 -381 4576 -347
rect 4510 -397 4576 -381
rect 4628 -347 4694 -331
rect 4628 -381 4644 -347
rect 4678 -381 4694 -347
rect 4628 -397 4694 -381
rect 4746 -347 4812 -331
rect 4746 -381 4762 -347
rect 4796 -381 4812 -347
rect 4746 -397 4812 -381
rect 4864 -347 4930 -331
rect 4864 -381 4880 -347
rect 4914 -381 4930 -347
rect 4864 -397 4930 -381
rect 4982 -347 5048 -331
rect 4982 -381 4998 -347
rect 5032 -381 5048 -347
rect 4982 -397 5048 -381
rect 5100 -347 5166 -331
rect 5100 -381 5116 -347
rect 5150 -381 5166 -347
rect 5100 -397 5166 -381
rect 5218 -347 5284 -331
rect 5218 -381 5234 -347
rect 5268 -381 5284 -347
rect 5218 -397 5284 -381
rect 5336 -347 5402 -331
rect 5336 -381 5352 -347
rect 5386 -381 5402 -347
rect 5336 -397 5402 -381
rect 5454 -347 5520 -331
rect 5454 -381 5470 -347
rect 5504 -381 5520 -347
rect 5454 -397 5520 -381
rect 5572 -347 5638 -331
rect 5572 -381 5588 -347
rect 5622 -381 5638 -347
rect 5572 -397 5638 -381
rect 5690 -347 5756 -331
rect 5690 -381 5706 -347
rect 5740 -381 5756 -347
rect 5690 -397 5756 -381
rect 5808 -347 5874 -331
rect 5808 -381 5824 -347
rect 5858 -381 5874 -347
rect 5808 -397 5874 -381
rect 5926 -347 5992 -331
rect 5926 -381 5942 -347
rect 5976 -381 5992 -347
rect 5926 -397 5992 -381
rect 6044 -347 6110 -331
rect 6044 -381 6060 -347
rect 6094 -381 6110 -347
rect 6044 -397 6110 -381
rect 6162 -347 6228 -331
rect 6162 -381 6178 -347
rect 6212 -381 6228 -347
rect 6162 -397 6228 -381
rect 6280 -347 6346 -331
rect 6280 -381 6296 -347
rect 6330 -381 6346 -347
rect 6280 -397 6346 -381
rect 6398 -347 6464 -331
rect 6398 -381 6414 -347
rect 6448 -381 6464 -347
rect 6398 -397 6464 -381
rect 6516 -347 6582 -331
rect 6516 -381 6532 -347
rect 6566 -381 6582 -347
rect 6516 -397 6582 -381
rect 6634 -347 6700 -331
rect 6634 -381 6650 -347
rect 6684 -381 6700 -347
rect 6634 -397 6700 -381
rect 6752 -347 6818 -331
rect 6752 -381 6768 -347
rect 6802 -381 6818 -347
rect 6752 -397 6818 -381
rect 6870 -347 6936 -331
rect 6870 -381 6886 -347
rect 6920 -381 6936 -347
rect 6870 -397 6936 -381
rect 6988 -347 7054 -331
rect 6988 -381 7004 -347
rect 7038 -381 7054 -347
rect 6988 -397 7054 -381
rect 7106 -347 7172 -331
rect 7106 -381 7122 -347
rect 7156 -381 7172 -347
rect 7106 -397 7172 -381
rect 7224 -347 7290 -331
rect 7224 -381 7240 -347
rect 7274 -381 7290 -347
rect 7224 -397 7290 -381
rect 7342 -347 7408 -331
rect 7342 -381 7358 -347
rect 7392 -381 7408 -347
rect 7342 -397 7408 -381
rect 7460 -347 7526 -331
rect 7460 -381 7476 -347
rect 7510 -381 7526 -347
rect 7460 -397 7526 -381
rect 7578 -347 7644 -331
rect 7578 -381 7594 -347
rect 7628 -381 7644 -347
rect 7578 -397 7644 -381
rect 7696 -347 7762 -331
rect 7696 -381 7712 -347
rect 7746 -381 7762 -347
rect 7696 -397 7762 -381
rect 7814 -347 7880 -331
rect 7814 -381 7830 -347
rect 7864 -381 7880 -347
rect 7814 -397 7880 -381
rect 7932 -347 7998 -331
rect 7932 -381 7948 -347
rect 7982 -381 7998 -347
rect 7932 -397 7998 -381
rect 8050 -347 8116 -331
rect 8050 -381 8066 -347
rect 8100 -381 8116 -347
rect 8050 -397 8116 -381
rect 8168 -347 8234 -331
rect 8168 -381 8184 -347
rect 8218 -381 8234 -347
rect 8168 -397 8234 -381
rect 8286 -347 8352 -331
rect 8286 -381 8302 -347
rect 8336 -381 8352 -347
rect 8286 -397 8352 -381
rect 8404 -347 8470 -331
rect 8404 -381 8420 -347
rect 8454 -381 8470 -347
rect 8404 -397 8470 -381
rect 8522 -347 8588 -331
rect 8522 -381 8538 -347
rect 8572 -381 8588 -347
rect 8522 -397 8588 -381
rect 8640 -347 8706 -331
rect 8640 -381 8656 -347
rect 8690 -381 8706 -347
rect 8640 -397 8706 -381
rect 8758 -347 8824 -331
rect 8758 -381 8774 -347
rect 8808 -381 8824 -347
rect 8758 -397 8824 -381
<< polycont >>
rect -8808 347 -8774 381
rect -8690 347 -8656 381
rect -8572 347 -8538 381
rect -8454 347 -8420 381
rect -8336 347 -8302 381
rect -8218 347 -8184 381
rect -8100 347 -8066 381
rect -7982 347 -7948 381
rect -7864 347 -7830 381
rect -7746 347 -7712 381
rect -7628 347 -7594 381
rect -7510 347 -7476 381
rect -7392 347 -7358 381
rect -7274 347 -7240 381
rect -7156 347 -7122 381
rect -7038 347 -7004 381
rect -6920 347 -6886 381
rect -6802 347 -6768 381
rect -6684 347 -6650 381
rect -6566 347 -6532 381
rect -6448 347 -6414 381
rect -6330 347 -6296 381
rect -6212 347 -6178 381
rect -6094 347 -6060 381
rect -5976 347 -5942 381
rect -5858 347 -5824 381
rect -5740 347 -5706 381
rect -5622 347 -5588 381
rect -5504 347 -5470 381
rect -5386 347 -5352 381
rect -5268 347 -5234 381
rect -5150 347 -5116 381
rect -5032 347 -4998 381
rect -4914 347 -4880 381
rect -4796 347 -4762 381
rect -4678 347 -4644 381
rect -4560 347 -4526 381
rect -4442 347 -4408 381
rect -4324 347 -4290 381
rect -4206 347 -4172 381
rect -4088 347 -4054 381
rect -3970 347 -3936 381
rect -3852 347 -3818 381
rect -3734 347 -3700 381
rect -3616 347 -3582 381
rect -3498 347 -3464 381
rect -3380 347 -3346 381
rect -3262 347 -3228 381
rect -3144 347 -3110 381
rect -3026 347 -2992 381
rect -2908 347 -2874 381
rect -2790 347 -2756 381
rect -2672 347 -2638 381
rect -2554 347 -2520 381
rect -2436 347 -2402 381
rect -2318 347 -2284 381
rect -2200 347 -2166 381
rect -2082 347 -2048 381
rect -1964 347 -1930 381
rect -1846 347 -1812 381
rect -1728 347 -1694 381
rect -1610 347 -1576 381
rect -1492 347 -1458 381
rect -1374 347 -1340 381
rect -1256 347 -1222 381
rect -1138 347 -1104 381
rect -1020 347 -986 381
rect -902 347 -868 381
rect -784 347 -750 381
rect -666 347 -632 381
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect 632 347 666 381
rect 750 347 784 381
rect 868 347 902 381
rect 986 347 1020 381
rect 1104 347 1138 381
rect 1222 347 1256 381
rect 1340 347 1374 381
rect 1458 347 1492 381
rect 1576 347 1610 381
rect 1694 347 1728 381
rect 1812 347 1846 381
rect 1930 347 1964 381
rect 2048 347 2082 381
rect 2166 347 2200 381
rect 2284 347 2318 381
rect 2402 347 2436 381
rect 2520 347 2554 381
rect 2638 347 2672 381
rect 2756 347 2790 381
rect 2874 347 2908 381
rect 2992 347 3026 381
rect 3110 347 3144 381
rect 3228 347 3262 381
rect 3346 347 3380 381
rect 3464 347 3498 381
rect 3582 347 3616 381
rect 3700 347 3734 381
rect 3818 347 3852 381
rect 3936 347 3970 381
rect 4054 347 4088 381
rect 4172 347 4206 381
rect 4290 347 4324 381
rect 4408 347 4442 381
rect 4526 347 4560 381
rect 4644 347 4678 381
rect 4762 347 4796 381
rect 4880 347 4914 381
rect 4998 347 5032 381
rect 5116 347 5150 381
rect 5234 347 5268 381
rect 5352 347 5386 381
rect 5470 347 5504 381
rect 5588 347 5622 381
rect 5706 347 5740 381
rect 5824 347 5858 381
rect 5942 347 5976 381
rect 6060 347 6094 381
rect 6178 347 6212 381
rect 6296 347 6330 381
rect 6414 347 6448 381
rect 6532 347 6566 381
rect 6650 347 6684 381
rect 6768 347 6802 381
rect 6886 347 6920 381
rect 7004 347 7038 381
rect 7122 347 7156 381
rect 7240 347 7274 381
rect 7358 347 7392 381
rect 7476 347 7510 381
rect 7594 347 7628 381
rect 7712 347 7746 381
rect 7830 347 7864 381
rect 7948 347 7982 381
rect 8066 347 8100 381
rect 8184 347 8218 381
rect 8302 347 8336 381
rect 8420 347 8454 381
rect 8538 347 8572 381
rect 8656 347 8690 381
rect 8774 347 8808 381
rect -8808 -381 -8774 -347
rect -8690 -381 -8656 -347
rect -8572 -381 -8538 -347
rect -8454 -381 -8420 -347
rect -8336 -381 -8302 -347
rect -8218 -381 -8184 -347
rect -8100 -381 -8066 -347
rect -7982 -381 -7948 -347
rect -7864 -381 -7830 -347
rect -7746 -381 -7712 -347
rect -7628 -381 -7594 -347
rect -7510 -381 -7476 -347
rect -7392 -381 -7358 -347
rect -7274 -381 -7240 -347
rect -7156 -381 -7122 -347
rect -7038 -381 -7004 -347
rect -6920 -381 -6886 -347
rect -6802 -381 -6768 -347
rect -6684 -381 -6650 -347
rect -6566 -381 -6532 -347
rect -6448 -381 -6414 -347
rect -6330 -381 -6296 -347
rect -6212 -381 -6178 -347
rect -6094 -381 -6060 -347
rect -5976 -381 -5942 -347
rect -5858 -381 -5824 -347
rect -5740 -381 -5706 -347
rect -5622 -381 -5588 -347
rect -5504 -381 -5470 -347
rect -5386 -381 -5352 -347
rect -5268 -381 -5234 -347
rect -5150 -381 -5116 -347
rect -5032 -381 -4998 -347
rect -4914 -381 -4880 -347
rect -4796 -381 -4762 -347
rect -4678 -381 -4644 -347
rect -4560 -381 -4526 -347
rect -4442 -381 -4408 -347
rect -4324 -381 -4290 -347
rect -4206 -381 -4172 -347
rect -4088 -381 -4054 -347
rect -3970 -381 -3936 -347
rect -3852 -381 -3818 -347
rect -3734 -381 -3700 -347
rect -3616 -381 -3582 -347
rect -3498 -381 -3464 -347
rect -3380 -381 -3346 -347
rect -3262 -381 -3228 -347
rect -3144 -381 -3110 -347
rect -3026 -381 -2992 -347
rect -2908 -381 -2874 -347
rect -2790 -381 -2756 -347
rect -2672 -381 -2638 -347
rect -2554 -381 -2520 -347
rect -2436 -381 -2402 -347
rect -2318 -381 -2284 -347
rect -2200 -381 -2166 -347
rect -2082 -381 -2048 -347
rect -1964 -381 -1930 -347
rect -1846 -381 -1812 -347
rect -1728 -381 -1694 -347
rect -1610 -381 -1576 -347
rect -1492 -381 -1458 -347
rect -1374 -381 -1340 -347
rect -1256 -381 -1222 -347
rect -1138 -381 -1104 -347
rect -1020 -381 -986 -347
rect -902 -381 -868 -347
rect -784 -381 -750 -347
rect -666 -381 -632 -347
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect 632 -381 666 -347
rect 750 -381 784 -347
rect 868 -381 902 -347
rect 986 -381 1020 -347
rect 1104 -381 1138 -347
rect 1222 -381 1256 -347
rect 1340 -381 1374 -347
rect 1458 -381 1492 -347
rect 1576 -381 1610 -347
rect 1694 -381 1728 -347
rect 1812 -381 1846 -347
rect 1930 -381 1964 -347
rect 2048 -381 2082 -347
rect 2166 -381 2200 -347
rect 2284 -381 2318 -347
rect 2402 -381 2436 -347
rect 2520 -381 2554 -347
rect 2638 -381 2672 -347
rect 2756 -381 2790 -347
rect 2874 -381 2908 -347
rect 2992 -381 3026 -347
rect 3110 -381 3144 -347
rect 3228 -381 3262 -347
rect 3346 -381 3380 -347
rect 3464 -381 3498 -347
rect 3582 -381 3616 -347
rect 3700 -381 3734 -347
rect 3818 -381 3852 -347
rect 3936 -381 3970 -347
rect 4054 -381 4088 -347
rect 4172 -381 4206 -347
rect 4290 -381 4324 -347
rect 4408 -381 4442 -347
rect 4526 -381 4560 -347
rect 4644 -381 4678 -347
rect 4762 -381 4796 -347
rect 4880 -381 4914 -347
rect 4998 -381 5032 -347
rect 5116 -381 5150 -347
rect 5234 -381 5268 -347
rect 5352 -381 5386 -347
rect 5470 -381 5504 -347
rect 5588 -381 5622 -347
rect 5706 -381 5740 -347
rect 5824 -381 5858 -347
rect 5942 -381 5976 -347
rect 6060 -381 6094 -347
rect 6178 -381 6212 -347
rect 6296 -381 6330 -347
rect 6414 -381 6448 -347
rect 6532 -381 6566 -347
rect 6650 -381 6684 -347
rect 6768 -381 6802 -347
rect 6886 -381 6920 -347
rect 7004 -381 7038 -347
rect 7122 -381 7156 -347
rect 7240 -381 7274 -347
rect 7358 -381 7392 -347
rect 7476 -381 7510 -347
rect 7594 -381 7628 -347
rect 7712 -381 7746 -347
rect 7830 -381 7864 -347
rect 7948 -381 7982 -347
rect 8066 -381 8100 -347
rect 8184 -381 8218 -347
rect 8302 -381 8336 -347
rect 8420 -381 8454 -347
rect 8538 -381 8572 -347
rect 8656 -381 8690 -347
rect 8774 -381 8808 -347
<< locali >>
rect -8981 449 -8885 483
rect 8885 449 8981 483
rect -8981 387 -8947 449
rect 8947 387 8981 449
rect -8824 347 -8808 381
rect -8774 347 -8758 381
rect -8706 347 -8690 381
rect -8656 347 -8640 381
rect -8588 347 -8572 381
rect -8538 347 -8522 381
rect -8470 347 -8454 381
rect -8420 347 -8404 381
rect -8352 347 -8336 381
rect -8302 347 -8286 381
rect -8234 347 -8218 381
rect -8184 347 -8168 381
rect -8116 347 -8100 381
rect -8066 347 -8050 381
rect -7998 347 -7982 381
rect -7948 347 -7932 381
rect -7880 347 -7864 381
rect -7830 347 -7814 381
rect -7762 347 -7746 381
rect -7712 347 -7696 381
rect -7644 347 -7628 381
rect -7594 347 -7578 381
rect -7526 347 -7510 381
rect -7476 347 -7460 381
rect -7408 347 -7392 381
rect -7358 347 -7342 381
rect -7290 347 -7274 381
rect -7240 347 -7224 381
rect -7172 347 -7156 381
rect -7122 347 -7106 381
rect -7054 347 -7038 381
rect -7004 347 -6988 381
rect -6936 347 -6920 381
rect -6886 347 -6870 381
rect -6818 347 -6802 381
rect -6768 347 -6752 381
rect -6700 347 -6684 381
rect -6650 347 -6634 381
rect -6582 347 -6566 381
rect -6532 347 -6516 381
rect -6464 347 -6448 381
rect -6414 347 -6398 381
rect -6346 347 -6330 381
rect -6296 347 -6280 381
rect -6228 347 -6212 381
rect -6178 347 -6162 381
rect -6110 347 -6094 381
rect -6060 347 -6044 381
rect -5992 347 -5976 381
rect -5942 347 -5926 381
rect -5874 347 -5858 381
rect -5824 347 -5808 381
rect -5756 347 -5740 381
rect -5706 347 -5690 381
rect -5638 347 -5622 381
rect -5588 347 -5572 381
rect -5520 347 -5504 381
rect -5470 347 -5454 381
rect -5402 347 -5386 381
rect -5352 347 -5336 381
rect -5284 347 -5268 381
rect -5234 347 -5218 381
rect -5166 347 -5150 381
rect -5116 347 -5100 381
rect -5048 347 -5032 381
rect -4998 347 -4982 381
rect -4930 347 -4914 381
rect -4880 347 -4864 381
rect -4812 347 -4796 381
rect -4762 347 -4746 381
rect -4694 347 -4678 381
rect -4644 347 -4628 381
rect -4576 347 -4560 381
rect -4526 347 -4510 381
rect -4458 347 -4442 381
rect -4408 347 -4392 381
rect -4340 347 -4324 381
rect -4290 347 -4274 381
rect -4222 347 -4206 381
rect -4172 347 -4156 381
rect -4104 347 -4088 381
rect -4054 347 -4038 381
rect -3986 347 -3970 381
rect -3936 347 -3920 381
rect -3868 347 -3852 381
rect -3818 347 -3802 381
rect -3750 347 -3734 381
rect -3700 347 -3684 381
rect -3632 347 -3616 381
rect -3582 347 -3566 381
rect -3514 347 -3498 381
rect -3464 347 -3448 381
rect -3396 347 -3380 381
rect -3346 347 -3330 381
rect -3278 347 -3262 381
rect -3228 347 -3212 381
rect -3160 347 -3144 381
rect -3110 347 -3094 381
rect -3042 347 -3026 381
rect -2992 347 -2976 381
rect -2924 347 -2908 381
rect -2874 347 -2858 381
rect -2806 347 -2790 381
rect -2756 347 -2740 381
rect -2688 347 -2672 381
rect -2638 347 -2622 381
rect -2570 347 -2554 381
rect -2520 347 -2504 381
rect -2452 347 -2436 381
rect -2402 347 -2386 381
rect -2334 347 -2318 381
rect -2284 347 -2268 381
rect -2216 347 -2200 381
rect -2166 347 -2150 381
rect -2098 347 -2082 381
rect -2048 347 -2032 381
rect -1980 347 -1964 381
rect -1930 347 -1914 381
rect -1862 347 -1846 381
rect -1812 347 -1796 381
rect -1744 347 -1728 381
rect -1694 347 -1678 381
rect -1626 347 -1610 381
rect -1576 347 -1560 381
rect -1508 347 -1492 381
rect -1458 347 -1442 381
rect -1390 347 -1374 381
rect -1340 347 -1324 381
rect -1272 347 -1256 381
rect -1222 347 -1206 381
rect -1154 347 -1138 381
rect -1104 347 -1088 381
rect -1036 347 -1020 381
rect -986 347 -970 381
rect -918 347 -902 381
rect -868 347 -852 381
rect -800 347 -784 381
rect -750 347 -734 381
rect -682 347 -666 381
rect -632 347 -616 381
rect -564 347 -548 381
rect -514 347 -498 381
rect -446 347 -430 381
rect -396 347 -380 381
rect -328 347 -312 381
rect -278 347 -262 381
rect -210 347 -194 381
rect -160 347 -144 381
rect -92 347 -76 381
rect -42 347 -26 381
rect 26 347 42 381
rect 76 347 92 381
rect 144 347 160 381
rect 194 347 210 381
rect 262 347 278 381
rect 312 347 328 381
rect 380 347 396 381
rect 430 347 446 381
rect 498 347 514 381
rect 548 347 564 381
rect 616 347 632 381
rect 666 347 682 381
rect 734 347 750 381
rect 784 347 800 381
rect 852 347 868 381
rect 902 347 918 381
rect 970 347 986 381
rect 1020 347 1036 381
rect 1088 347 1104 381
rect 1138 347 1154 381
rect 1206 347 1222 381
rect 1256 347 1272 381
rect 1324 347 1340 381
rect 1374 347 1390 381
rect 1442 347 1458 381
rect 1492 347 1508 381
rect 1560 347 1576 381
rect 1610 347 1626 381
rect 1678 347 1694 381
rect 1728 347 1744 381
rect 1796 347 1812 381
rect 1846 347 1862 381
rect 1914 347 1930 381
rect 1964 347 1980 381
rect 2032 347 2048 381
rect 2082 347 2098 381
rect 2150 347 2166 381
rect 2200 347 2216 381
rect 2268 347 2284 381
rect 2318 347 2334 381
rect 2386 347 2402 381
rect 2436 347 2452 381
rect 2504 347 2520 381
rect 2554 347 2570 381
rect 2622 347 2638 381
rect 2672 347 2688 381
rect 2740 347 2756 381
rect 2790 347 2806 381
rect 2858 347 2874 381
rect 2908 347 2924 381
rect 2976 347 2992 381
rect 3026 347 3042 381
rect 3094 347 3110 381
rect 3144 347 3160 381
rect 3212 347 3228 381
rect 3262 347 3278 381
rect 3330 347 3346 381
rect 3380 347 3396 381
rect 3448 347 3464 381
rect 3498 347 3514 381
rect 3566 347 3582 381
rect 3616 347 3632 381
rect 3684 347 3700 381
rect 3734 347 3750 381
rect 3802 347 3818 381
rect 3852 347 3868 381
rect 3920 347 3936 381
rect 3970 347 3986 381
rect 4038 347 4054 381
rect 4088 347 4104 381
rect 4156 347 4172 381
rect 4206 347 4222 381
rect 4274 347 4290 381
rect 4324 347 4340 381
rect 4392 347 4408 381
rect 4442 347 4458 381
rect 4510 347 4526 381
rect 4560 347 4576 381
rect 4628 347 4644 381
rect 4678 347 4694 381
rect 4746 347 4762 381
rect 4796 347 4812 381
rect 4864 347 4880 381
rect 4914 347 4930 381
rect 4982 347 4998 381
rect 5032 347 5048 381
rect 5100 347 5116 381
rect 5150 347 5166 381
rect 5218 347 5234 381
rect 5268 347 5284 381
rect 5336 347 5352 381
rect 5386 347 5402 381
rect 5454 347 5470 381
rect 5504 347 5520 381
rect 5572 347 5588 381
rect 5622 347 5638 381
rect 5690 347 5706 381
rect 5740 347 5756 381
rect 5808 347 5824 381
rect 5858 347 5874 381
rect 5926 347 5942 381
rect 5976 347 5992 381
rect 6044 347 6060 381
rect 6094 347 6110 381
rect 6162 347 6178 381
rect 6212 347 6228 381
rect 6280 347 6296 381
rect 6330 347 6346 381
rect 6398 347 6414 381
rect 6448 347 6464 381
rect 6516 347 6532 381
rect 6566 347 6582 381
rect 6634 347 6650 381
rect 6684 347 6700 381
rect 6752 347 6768 381
rect 6802 347 6818 381
rect 6870 347 6886 381
rect 6920 347 6936 381
rect 6988 347 7004 381
rect 7038 347 7054 381
rect 7106 347 7122 381
rect 7156 347 7172 381
rect 7224 347 7240 381
rect 7274 347 7290 381
rect 7342 347 7358 381
rect 7392 347 7408 381
rect 7460 347 7476 381
rect 7510 347 7526 381
rect 7578 347 7594 381
rect 7628 347 7644 381
rect 7696 347 7712 381
rect 7746 347 7762 381
rect 7814 347 7830 381
rect 7864 347 7880 381
rect 7932 347 7948 381
rect 7982 347 7998 381
rect 8050 347 8066 381
rect 8100 347 8116 381
rect 8168 347 8184 381
rect 8218 347 8234 381
rect 8286 347 8302 381
rect 8336 347 8352 381
rect 8404 347 8420 381
rect 8454 347 8470 381
rect 8522 347 8538 381
rect 8572 347 8588 381
rect 8640 347 8656 381
rect 8690 347 8706 381
rect 8758 347 8774 381
rect 8808 347 8824 381
rect -8867 288 -8833 304
rect -8867 -304 -8833 -288
rect -8749 288 -8715 304
rect -8749 -304 -8715 -288
rect -8631 288 -8597 304
rect -8631 -304 -8597 -288
rect -8513 288 -8479 304
rect -8513 -304 -8479 -288
rect -8395 288 -8361 304
rect -8395 -304 -8361 -288
rect -8277 288 -8243 304
rect -8277 -304 -8243 -288
rect -8159 288 -8125 304
rect -8159 -304 -8125 -288
rect -8041 288 -8007 304
rect -8041 -304 -8007 -288
rect -7923 288 -7889 304
rect -7923 -304 -7889 -288
rect -7805 288 -7771 304
rect -7805 -304 -7771 -288
rect -7687 288 -7653 304
rect -7687 -304 -7653 -288
rect -7569 288 -7535 304
rect -7569 -304 -7535 -288
rect -7451 288 -7417 304
rect -7451 -304 -7417 -288
rect -7333 288 -7299 304
rect -7333 -304 -7299 -288
rect -7215 288 -7181 304
rect -7215 -304 -7181 -288
rect -7097 288 -7063 304
rect -7097 -304 -7063 -288
rect -6979 288 -6945 304
rect -6979 -304 -6945 -288
rect -6861 288 -6827 304
rect -6861 -304 -6827 -288
rect -6743 288 -6709 304
rect -6743 -304 -6709 -288
rect -6625 288 -6591 304
rect -6625 -304 -6591 -288
rect -6507 288 -6473 304
rect -6507 -304 -6473 -288
rect -6389 288 -6355 304
rect -6389 -304 -6355 -288
rect -6271 288 -6237 304
rect -6271 -304 -6237 -288
rect -6153 288 -6119 304
rect -6153 -304 -6119 -288
rect -6035 288 -6001 304
rect -6035 -304 -6001 -288
rect -5917 288 -5883 304
rect -5917 -304 -5883 -288
rect -5799 288 -5765 304
rect -5799 -304 -5765 -288
rect -5681 288 -5647 304
rect -5681 -304 -5647 -288
rect -5563 288 -5529 304
rect -5563 -304 -5529 -288
rect -5445 288 -5411 304
rect -5445 -304 -5411 -288
rect -5327 288 -5293 304
rect -5327 -304 -5293 -288
rect -5209 288 -5175 304
rect -5209 -304 -5175 -288
rect -5091 288 -5057 304
rect -5091 -304 -5057 -288
rect -4973 288 -4939 304
rect -4973 -304 -4939 -288
rect -4855 288 -4821 304
rect -4855 -304 -4821 -288
rect -4737 288 -4703 304
rect -4737 -304 -4703 -288
rect -4619 288 -4585 304
rect -4619 -304 -4585 -288
rect -4501 288 -4467 304
rect -4501 -304 -4467 -288
rect -4383 288 -4349 304
rect -4383 -304 -4349 -288
rect -4265 288 -4231 304
rect -4265 -304 -4231 -288
rect -4147 288 -4113 304
rect -4147 -304 -4113 -288
rect -4029 288 -3995 304
rect -4029 -304 -3995 -288
rect -3911 288 -3877 304
rect -3911 -304 -3877 -288
rect -3793 288 -3759 304
rect -3793 -304 -3759 -288
rect -3675 288 -3641 304
rect -3675 -304 -3641 -288
rect -3557 288 -3523 304
rect -3557 -304 -3523 -288
rect -3439 288 -3405 304
rect -3439 -304 -3405 -288
rect -3321 288 -3287 304
rect -3321 -304 -3287 -288
rect -3203 288 -3169 304
rect -3203 -304 -3169 -288
rect -3085 288 -3051 304
rect -3085 -304 -3051 -288
rect -2967 288 -2933 304
rect -2967 -304 -2933 -288
rect -2849 288 -2815 304
rect -2849 -304 -2815 -288
rect -2731 288 -2697 304
rect -2731 -304 -2697 -288
rect -2613 288 -2579 304
rect -2613 -304 -2579 -288
rect -2495 288 -2461 304
rect -2495 -304 -2461 -288
rect -2377 288 -2343 304
rect -2377 -304 -2343 -288
rect -2259 288 -2225 304
rect -2259 -304 -2225 -288
rect -2141 288 -2107 304
rect -2141 -304 -2107 -288
rect -2023 288 -1989 304
rect -2023 -304 -1989 -288
rect -1905 288 -1871 304
rect -1905 -304 -1871 -288
rect -1787 288 -1753 304
rect -1787 -304 -1753 -288
rect -1669 288 -1635 304
rect -1669 -304 -1635 -288
rect -1551 288 -1517 304
rect -1551 -304 -1517 -288
rect -1433 288 -1399 304
rect -1433 -304 -1399 -288
rect -1315 288 -1281 304
rect -1315 -304 -1281 -288
rect -1197 288 -1163 304
rect -1197 -304 -1163 -288
rect -1079 288 -1045 304
rect -1079 -304 -1045 -288
rect -961 288 -927 304
rect -961 -304 -927 -288
rect -843 288 -809 304
rect -843 -304 -809 -288
rect -725 288 -691 304
rect -725 -304 -691 -288
rect -607 288 -573 304
rect -607 -304 -573 -288
rect -489 288 -455 304
rect -489 -304 -455 -288
rect -371 288 -337 304
rect -371 -304 -337 -288
rect -253 288 -219 304
rect -253 -304 -219 -288
rect -135 288 -101 304
rect -135 -304 -101 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 101 288 135 304
rect 101 -304 135 -288
rect 219 288 253 304
rect 219 -304 253 -288
rect 337 288 371 304
rect 337 -304 371 -288
rect 455 288 489 304
rect 455 -304 489 -288
rect 573 288 607 304
rect 573 -304 607 -288
rect 691 288 725 304
rect 691 -304 725 -288
rect 809 288 843 304
rect 809 -304 843 -288
rect 927 288 961 304
rect 927 -304 961 -288
rect 1045 288 1079 304
rect 1045 -304 1079 -288
rect 1163 288 1197 304
rect 1163 -304 1197 -288
rect 1281 288 1315 304
rect 1281 -304 1315 -288
rect 1399 288 1433 304
rect 1399 -304 1433 -288
rect 1517 288 1551 304
rect 1517 -304 1551 -288
rect 1635 288 1669 304
rect 1635 -304 1669 -288
rect 1753 288 1787 304
rect 1753 -304 1787 -288
rect 1871 288 1905 304
rect 1871 -304 1905 -288
rect 1989 288 2023 304
rect 1989 -304 2023 -288
rect 2107 288 2141 304
rect 2107 -304 2141 -288
rect 2225 288 2259 304
rect 2225 -304 2259 -288
rect 2343 288 2377 304
rect 2343 -304 2377 -288
rect 2461 288 2495 304
rect 2461 -304 2495 -288
rect 2579 288 2613 304
rect 2579 -304 2613 -288
rect 2697 288 2731 304
rect 2697 -304 2731 -288
rect 2815 288 2849 304
rect 2815 -304 2849 -288
rect 2933 288 2967 304
rect 2933 -304 2967 -288
rect 3051 288 3085 304
rect 3051 -304 3085 -288
rect 3169 288 3203 304
rect 3169 -304 3203 -288
rect 3287 288 3321 304
rect 3287 -304 3321 -288
rect 3405 288 3439 304
rect 3405 -304 3439 -288
rect 3523 288 3557 304
rect 3523 -304 3557 -288
rect 3641 288 3675 304
rect 3641 -304 3675 -288
rect 3759 288 3793 304
rect 3759 -304 3793 -288
rect 3877 288 3911 304
rect 3877 -304 3911 -288
rect 3995 288 4029 304
rect 3995 -304 4029 -288
rect 4113 288 4147 304
rect 4113 -304 4147 -288
rect 4231 288 4265 304
rect 4231 -304 4265 -288
rect 4349 288 4383 304
rect 4349 -304 4383 -288
rect 4467 288 4501 304
rect 4467 -304 4501 -288
rect 4585 288 4619 304
rect 4585 -304 4619 -288
rect 4703 288 4737 304
rect 4703 -304 4737 -288
rect 4821 288 4855 304
rect 4821 -304 4855 -288
rect 4939 288 4973 304
rect 4939 -304 4973 -288
rect 5057 288 5091 304
rect 5057 -304 5091 -288
rect 5175 288 5209 304
rect 5175 -304 5209 -288
rect 5293 288 5327 304
rect 5293 -304 5327 -288
rect 5411 288 5445 304
rect 5411 -304 5445 -288
rect 5529 288 5563 304
rect 5529 -304 5563 -288
rect 5647 288 5681 304
rect 5647 -304 5681 -288
rect 5765 288 5799 304
rect 5765 -304 5799 -288
rect 5883 288 5917 304
rect 5883 -304 5917 -288
rect 6001 288 6035 304
rect 6001 -304 6035 -288
rect 6119 288 6153 304
rect 6119 -304 6153 -288
rect 6237 288 6271 304
rect 6237 -304 6271 -288
rect 6355 288 6389 304
rect 6355 -304 6389 -288
rect 6473 288 6507 304
rect 6473 -304 6507 -288
rect 6591 288 6625 304
rect 6591 -304 6625 -288
rect 6709 288 6743 304
rect 6709 -304 6743 -288
rect 6827 288 6861 304
rect 6827 -304 6861 -288
rect 6945 288 6979 304
rect 6945 -304 6979 -288
rect 7063 288 7097 304
rect 7063 -304 7097 -288
rect 7181 288 7215 304
rect 7181 -304 7215 -288
rect 7299 288 7333 304
rect 7299 -304 7333 -288
rect 7417 288 7451 304
rect 7417 -304 7451 -288
rect 7535 288 7569 304
rect 7535 -304 7569 -288
rect 7653 288 7687 304
rect 7653 -304 7687 -288
rect 7771 288 7805 304
rect 7771 -304 7805 -288
rect 7889 288 7923 304
rect 7889 -304 7923 -288
rect 8007 288 8041 304
rect 8007 -304 8041 -288
rect 8125 288 8159 304
rect 8125 -304 8159 -288
rect 8243 288 8277 304
rect 8243 -304 8277 -288
rect 8361 288 8395 304
rect 8361 -304 8395 -288
rect 8479 288 8513 304
rect 8479 -304 8513 -288
rect 8597 288 8631 304
rect 8597 -304 8631 -288
rect 8715 288 8749 304
rect 8715 -304 8749 -288
rect 8833 288 8867 304
rect 8833 -304 8867 -288
rect -8824 -381 -8808 -347
rect -8774 -381 -8758 -347
rect -8706 -381 -8690 -347
rect -8656 -381 -8640 -347
rect -8588 -381 -8572 -347
rect -8538 -381 -8522 -347
rect -8470 -381 -8454 -347
rect -8420 -381 -8404 -347
rect -8352 -381 -8336 -347
rect -8302 -381 -8286 -347
rect -8234 -381 -8218 -347
rect -8184 -381 -8168 -347
rect -8116 -381 -8100 -347
rect -8066 -381 -8050 -347
rect -7998 -381 -7982 -347
rect -7948 -381 -7932 -347
rect -7880 -381 -7864 -347
rect -7830 -381 -7814 -347
rect -7762 -381 -7746 -347
rect -7712 -381 -7696 -347
rect -7644 -381 -7628 -347
rect -7594 -381 -7578 -347
rect -7526 -381 -7510 -347
rect -7476 -381 -7460 -347
rect -7408 -381 -7392 -347
rect -7358 -381 -7342 -347
rect -7290 -381 -7274 -347
rect -7240 -381 -7224 -347
rect -7172 -381 -7156 -347
rect -7122 -381 -7106 -347
rect -7054 -381 -7038 -347
rect -7004 -381 -6988 -347
rect -6936 -381 -6920 -347
rect -6886 -381 -6870 -347
rect -6818 -381 -6802 -347
rect -6768 -381 -6752 -347
rect -6700 -381 -6684 -347
rect -6650 -381 -6634 -347
rect -6582 -381 -6566 -347
rect -6532 -381 -6516 -347
rect -6464 -381 -6448 -347
rect -6414 -381 -6398 -347
rect -6346 -381 -6330 -347
rect -6296 -381 -6280 -347
rect -6228 -381 -6212 -347
rect -6178 -381 -6162 -347
rect -6110 -381 -6094 -347
rect -6060 -381 -6044 -347
rect -5992 -381 -5976 -347
rect -5942 -381 -5926 -347
rect -5874 -381 -5858 -347
rect -5824 -381 -5808 -347
rect -5756 -381 -5740 -347
rect -5706 -381 -5690 -347
rect -5638 -381 -5622 -347
rect -5588 -381 -5572 -347
rect -5520 -381 -5504 -347
rect -5470 -381 -5454 -347
rect -5402 -381 -5386 -347
rect -5352 -381 -5336 -347
rect -5284 -381 -5268 -347
rect -5234 -381 -5218 -347
rect -5166 -381 -5150 -347
rect -5116 -381 -5100 -347
rect -5048 -381 -5032 -347
rect -4998 -381 -4982 -347
rect -4930 -381 -4914 -347
rect -4880 -381 -4864 -347
rect -4812 -381 -4796 -347
rect -4762 -381 -4746 -347
rect -4694 -381 -4678 -347
rect -4644 -381 -4628 -347
rect -4576 -381 -4560 -347
rect -4526 -381 -4510 -347
rect -4458 -381 -4442 -347
rect -4408 -381 -4392 -347
rect -4340 -381 -4324 -347
rect -4290 -381 -4274 -347
rect -4222 -381 -4206 -347
rect -4172 -381 -4156 -347
rect -4104 -381 -4088 -347
rect -4054 -381 -4038 -347
rect -3986 -381 -3970 -347
rect -3936 -381 -3920 -347
rect -3868 -381 -3852 -347
rect -3818 -381 -3802 -347
rect -3750 -381 -3734 -347
rect -3700 -381 -3684 -347
rect -3632 -381 -3616 -347
rect -3582 -381 -3566 -347
rect -3514 -381 -3498 -347
rect -3464 -381 -3448 -347
rect -3396 -381 -3380 -347
rect -3346 -381 -3330 -347
rect -3278 -381 -3262 -347
rect -3228 -381 -3212 -347
rect -3160 -381 -3144 -347
rect -3110 -381 -3094 -347
rect -3042 -381 -3026 -347
rect -2992 -381 -2976 -347
rect -2924 -381 -2908 -347
rect -2874 -381 -2858 -347
rect -2806 -381 -2790 -347
rect -2756 -381 -2740 -347
rect -2688 -381 -2672 -347
rect -2638 -381 -2622 -347
rect -2570 -381 -2554 -347
rect -2520 -381 -2504 -347
rect -2452 -381 -2436 -347
rect -2402 -381 -2386 -347
rect -2334 -381 -2318 -347
rect -2284 -381 -2268 -347
rect -2216 -381 -2200 -347
rect -2166 -381 -2150 -347
rect -2098 -381 -2082 -347
rect -2048 -381 -2032 -347
rect -1980 -381 -1964 -347
rect -1930 -381 -1914 -347
rect -1862 -381 -1846 -347
rect -1812 -381 -1796 -347
rect -1744 -381 -1728 -347
rect -1694 -381 -1678 -347
rect -1626 -381 -1610 -347
rect -1576 -381 -1560 -347
rect -1508 -381 -1492 -347
rect -1458 -381 -1442 -347
rect -1390 -381 -1374 -347
rect -1340 -381 -1324 -347
rect -1272 -381 -1256 -347
rect -1222 -381 -1206 -347
rect -1154 -381 -1138 -347
rect -1104 -381 -1088 -347
rect -1036 -381 -1020 -347
rect -986 -381 -970 -347
rect -918 -381 -902 -347
rect -868 -381 -852 -347
rect -800 -381 -784 -347
rect -750 -381 -734 -347
rect -682 -381 -666 -347
rect -632 -381 -616 -347
rect -564 -381 -548 -347
rect -514 -381 -498 -347
rect -446 -381 -430 -347
rect -396 -381 -380 -347
rect -328 -381 -312 -347
rect -278 -381 -262 -347
rect -210 -381 -194 -347
rect -160 -381 -144 -347
rect -92 -381 -76 -347
rect -42 -381 -26 -347
rect 26 -381 42 -347
rect 76 -381 92 -347
rect 144 -381 160 -347
rect 194 -381 210 -347
rect 262 -381 278 -347
rect 312 -381 328 -347
rect 380 -381 396 -347
rect 430 -381 446 -347
rect 498 -381 514 -347
rect 548 -381 564 -347
rect 616 -381 632 -347
rect 666 -381 682 -347
rect 734 -381 750 -347
rect 784 -381 800 -347
rect 852 -381 868 -347
rect 902 -381 918 -347
rect 970 -381 986 -347
rect 1020 -381 1036 -347
rect 1088 -381 1104 -347
rect 1138 -381 1154 -347
rect 1206 -381 1222 -347
rect 1256 -381 1272 -347
rect 1324 -381 1340 -347
rect 1374 -381 1390 -347
rect 1442 -381 1458 -347
rect 1492 -381 1508 -347
rect 1560 -381 1576 -347
rect 1610 -381 1626 -347
rect 1678 -381 1694 -347
rect 1728 -381 1744 -347
rect 1796 -381 1812 -347
rect 1846 -381 1862 -347
rect 1914 -381 1930 -347
rect 1964 -381 1980 -347
rect 2032 -381 2048 -347
rect 2082 -381 2098 -347
rect 2150 -381 2166 -347
rect 2200 -381 2216 -347
rect 2268 -381 2284 -347
rect 2318 -381 2334 -347
rect 2386 -381 2402 -347
rect 2436 -381 2452 -347
rect 2504 -381 2520 -347
rect 2554 -381 2570 -347
rect 2622 -381 2638 -347
rect 2672 -381 2688 -347
rect 2740 -381 2756 -347
rect 2790 -381 2806 -347
rect 2858 -381 2874 -347
rect 2908 -381 2924 -347
rect 2976 -381 2992 -347
rect 3026 -381 3042 -347
rect 3094 -381 3110 -347
rect 3144 -381 3160 -347
rect 3212 -381 3228 -347
rect 3262 -381 3278 -347
rect 3330 -381 3346 -347
rect 3380 -381 3396 -347
rect 3448 -381 3464 -347
rect 3498 -381 3514 -347
rect 3566 -381 3582 -347
rect 3616 -381 3632 -347
rect 3684 -381 3700 -347
rect 3734 -381 3750 -347
rect 3802 -381 3818 -347
rect 3852 -381 3868 -347
rect 3920 -381 3936 -347
rect 3970 -381 3986 -347
rect 4038 -381 4054 -347
rect 4088 -381 4104 -347
rect 4156 -381 4172 -347
rect 4206 -381 4222 -347
rect 4274 -381 4290 -347
rect 4324 -381 4340 -347
rect 4392 -381 4408 -347
rect 4442 -381 4458 -347
rect 4510 -381 4526 -347
rect 4560 -381 4576 -347
rect 4628 -381 4644 -347
rect 4678 -381 4694 -347
rect 4746 -381 4762 -347
rect 4796 -381 4812 -347
rect 4864 -381 4880 -347
rect 4914 -381 4930 -347
rect 4982 -381 4998 -347
rect 5032 -381 5048 -347
rect 5100 -381 5116 -347
rect 5150 -381 5166 -347
rect 5218 -381 5234 -347
rect 5268 -381 5284 -347
rect 5336 -381 5352 -347
rect 5386 -381 5402 -347
rect 5454 -381 5470 -347
rect 5504 -381 5520 -347
rect 5572 -381 5588 -347
rect 5622 -381 5638 -347
rect 5690 -381 5706 -347
rect 5740 -381 5756 -347
rect 5808 -381 5824 -347
rect 5858 -381 5874 -347
rect 5926 -381 5942 -347
rect 5976 -381 5992 -347
rect 6044 -381 6060 -347
rect 6094 -381 6110 -347
rect 6162 -381 6178 -347
rect 6212 -381 6228 -347
rect 6280 -381 6296 -347
rect 6330 -381 6346 -347
rect 6398 -381 6414 -347
rect 6448 -381 6464 -347
rect 6516 -381 6532 -347
rect 6566 -381 6582 -347
rect 6634 -381 6650 -347
rect 6684 -381 6700 -347
rect 6752 -381 6768 -347
rect 6802 -381 6818 -347
rect 6870 -381 6886 -347
rect 6920 -381 6936 -347
rect 6988 -381 7004 -347
rect 7038 -381 7054 -347
rect 7106 -381 7122 -347
rect 7156 -381 7172 -347
rect 7224 -381 7240 -347
rect 7274 -381 7290 -347
rect 7342 -381 7358 -347
rect 7392 -381 7408 -347
rect 7460 -381 7476 -347
rect 7510 -381 7526 -347
rect 7578 -381 7594 -347
rect 7628 -381 7644 -347
rect 7696 -381 7712 -347
rect 7746 -381 7762 -347
rect 7814 -381 7830 -347
rect 7864 -381 7880 -347
rect 7932 -381 7948 -347
rect 7982 -381 7998 -347
rect 8050 -381 8066 -347
rect 8100 -381 8116 -347
rect 8168 -381 8184 -347
rect 8218 -381 8234 -347
rect 8286 -381 8302 -347
rect 8336 -381 8352 -347
rect 8404 -381 8420 -347
rect 8454 -381 8470 -347
rect 8522 -381 8538 -347
rect 8572 -381 8588 -347
rect 8640 -381 8656 -347
rect 8690 -381 8706 -347
rect 8758 -381 8774 -347
rect 8808 -381 8824 -347
rect -8981 -449 -8947 -387
rect 8947 -449 8981 -387
rect -8981 -483 -8885 -449
rect 8885 -483 8981 -449
<< viali >>
rect -8808 347 -8774 381
rect -8690 347 -8656 381
rect -8572 347 -8538 381
rect -8454 347 -8420 381
rect -8336 347 -8302 381
rect -8218 347 -8184 381
rect -8100 347 -8066 381
rect -7982 347 -7948 381
rect -7864 347 -7830 381
rect -7746 347 -7712 381
rect -7628 347 -7594 381
rect -7510 347 -7476 381
rect -7392 347 -7358 381
rect -7274 347 -7240 381
rect -7156 347 -7122 381
rect -7038 347 -7004 381
rect -6920 347 -6886 381
rect -6802 347 -6768 381
rect -6684 347 -6650 381
rect -6566 347 -6532 381
rect -6448 347 -6414 381
rect -6330 347 -6296 381
rect -6212 347 -6178 381
rect -6094 347 -6060 381
rect -5976 347 -5942 381
rect -5858 347 -5824 381
rect -5740 347 -5706 381
rect -5622 347 -5588 381
rect -5504 347 -5470 381
rect -5386 347 -5352 381
rect -5268 347 -5234 381
rect -5150 347 -5116 381
rect -5032 347 -4998 381
rect -4914 347 -4880 381
rect -4796 347 -4762 381
rect -4678 347 -4644 381
rect -4560 347 -4526 381
rect -4442 347 -4408 381
rect -4324 347 -4290 381
rect -4206 347 -4172 381
rect -4088 347 -4054 381
rect -3970 347 -3936 381
rect -3852 347 -3818 381
rect -3734 347 -3700 381
rect -3616 347 -3582 381
rect -3498 347 -3464 381
rect -3380 347 -3346 381
rect -3262 347 -3228 381
rect -3144 347 -3110 381
rect -3026 347 -2992 381
rect -2908 347 -2874 381
rect -2790 347 -2756 381
rect -2672 347 -2638 381
rect -2554 347 -2520 381
rect -2436 347 -2402 381
rect -2318 347 -2284 381
rect -2200 347 -2166 381
rect -2082 347 -2048 381
rect -1964 347 -1930 381
rect -1846 347 -1812 381
rect -1728 347 -1694 381
rect -1610 347 -1576 381
rect -1492 347 -1458 381
rect -1374 347 -1340 381
rect -1256 347 -1222 381
rect -1138 347 -1104 381
rect -1020 347 -986 381
rect -902 347 -868 381
rect -784 347 -750 381
rect -666 347 -632 381
rect -548 347 -514 381
rect -430 347 -396 381
rect -312 347 -278 381
rect -194 347 -160 381
rect -76 347 -42 381
rect 42 347 76 381
rect 160 347 194 381
rect 278 347 312 381
rect 396 347 430 381
rect 514 347 548 381
rect 632 347 666 381
rect 750 347 784 381
rect 868 347 902 381
rect 986 347 1020 381
rect 1104 347 1138 381
rect 1222 347 1256 381
rect 1340 347 1374 381
rect 1458 347 1492 381
rect 1576 347 1610 381
rect 1694 347 1728 381
rect 1812 347 1846 381
rect 1930 347 1964 381
rect 2048 347 2082 381
rect 2166 347 2200 381
rect 2284 347 2318 381
rect 2402 347 2436 381
rect 2520 347 2554 381
rect 2638 347 2672 381
rect 2756 347 2790 381
rect 2874 347 2908 381
rect 2992 347 3026 381
rect 3110 347 3144 381
rect 3228 347 3262 381
rect 3346 347 3380 381
rect 3464 347 3498 381
rect 3582 347 3616 381
rect 3700 347 3734 381
rect 3818 347 3852 381
rect 3936 347 3970 381
rect 4054 347 4088 381
rect 4172 347 4206 381
rect 4290 347 4324 381
rect 4408 347 4442 381
rect 4526 347 4560 381
rect 4644 347 4678 381
rect 4762 347 4796 381
rect 4880 347 4914 381
rect 4998 347 5032 381
rect 5116 347 5150 381
rect 5234 347 5268 381
rect 5352 347 5386 381
rect 5470 347 5504 381
rect 5588 347 5622 381
rect 5706 347 5740 381
rect 5824 347 5858 381
rect 5942 347 5976 381
rect 6060 347 6094 381
rect 6178 347 6212 381
rect 6296 347 6330 381
rect 6414 347 6448 381
rect 6532 347 6566 381
rect 6650 347 6684 381
rect 6768 347 6802 381
rect 6886 347 6920 381
rect 7004 347 7038 381
rect 7122 347 7156 381
rect 7240 347 7274 381
rect 7358 347 7392 381
rect 7476 347 7510 381
rect 7594 347 7628 381
rect 7712 347 7746 381
rect 7830 347 7864 381
rect 7948 347 7982 381
rect 8066 347 8100 381
rect 8184 347 8218 381
rect 8302 347 8336 381
rect 8420 347 8454 381
rect 8538 347 8572 381
rect 8656 347 8690 381
rect 8774 347 8808 381
rect -8867 -288 -8833 288
rect -8749 -288 -8715 288
rect -8631 -288 -8597 288
rect -8513 -288 -8479 288
rect -8395 -288 -8361 288
rect -8277 -288 -8243 288
rect -8159 -288 -8125 288
rect -8041 -288 -8007 288
rect -7923 -288 -7889 288
rect -7805 -288 -7771 288
rect -7687 -288 -7653 288
rect -7569 -288 -7535 288
rect -7451 -288 -7417 288
rect -7333 -288 -7299 288
rect -7215 -288 -7181 288
rect -7097 -288 -7063 288
rect -6979 -288 -6945 288
rect -6861 -288 -6827 288
rect -6743 -288 -6709 288
rect -6625 -288 -6591 288
rect -6507 -288 -6473 288
rect -6389 -288 -6355 288
rect -6271 -288 -6237 288
rect -6153 -288 -6119 288
rect -6035 -288 -6001 288
rect -5917 -288 -5883 288
rect -5799 -288 -5765 288
rect -5681 -288 -5647 288
rect -5563 -288 -5529 288
rect -5445 -288 -5411 288
rect -5327 -288 -5293 288
rect -5209 -288 -5175 288
rect -5091 -288 -5057 288
rect -4973 -288 -4939 288
rect -4855 -288 -4821 288
rect -4737 -288 -4703 288
rect -4619 -288 -4585 288
rect -4501 -288 -4467 288
rect -4383 -288 -4349 288
rect -4265 -288 -4231 288
rect -4147 -288 -4113 288
rect -4029 -288 -3995 288
rect -3911 -288 -3877 288
rect -3793 -288 -3759 288
rect -3675 -288 -3641 288
rect -3557 -288 -3523 288
rect -3439 -288 -3405 288
rect -3321 -288 -3287 288
rect -3203 -288 -3169 288
rect -3085 -288 -3051 288
rect -2967 -288 -2933 288
rect -2849 -288 -2815 288
rect -2731 -288 -2697 288
rect -2613 -288 -2579 288
rect -2495 -288 -2461 288
rect -2377 -288 -2343 288
rect -2259 -288 -2225 288
rect -2141 -288 -2107 288
rect -2023 -288 -1989 288
rect -1905 -288 -1871 288
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
rect 1871 -288 1905 288
rect 1989 -288 2023 288
rect 2107 -288 2141 288
rect 2225 -288 2259 288
rect 2343 -288 2377 288
rect 2461 -288 2495 288
rect 2579 -288 2613 288
rect 2697 -288 2731 288
rect 2815 -288 2849 288
rect 2933 -288 2967 288
rect 3051 -288 3085 288
rect 3169 -288 3203 288
rect 3287 -288 3321 288
rect 3405 -288 3439 288
rect 3523 -288 3557 288
rect 3641 -288 3675 288
rect 3759 -288 3793 288
rect 3877 -288 3911 288
rect 3995 -288 4029 288
rect 4113 -288 4147 288
rect 4231 -288 4265 288
rect 4349 -288 4383 288
rect 4467 -288 4501 288
rect 4585 -288 4619 288
rect 4703 -288 4737 288
rect 4821 -288 4855 288
rect 4939 -288 4973 288
rect 5057 -288 5091 288
rect 5175 -288 5209 288
rect 5293 -288 5327 288
rect 5411 -288 5445 288
rect 5529 -288 5563 288
rect 5647 -288 5681 288
rect 5765 -288 5799 288
rect 5883 -288 5917 288
rect 6001 -288 6035 288
rect 6119 -288 6153 288
rect 6237 -288 6271 288
rect 6355 -288 6389 288
rect 6473 -288 6507 288
rect 6591 -288 6625 288
rect 6709 -288 6743 288
rect 6827 -288 6861 288
rect 6945 -288 6979 288
rect 7063 -288 7097 288
rect 7181 -288 7215 288
rect 7299 -288 7333 288
rect 7417 -288 7451 288
rect 7535 -288 7569 288
rect 7653 -288 7687 288
rect 7771 -288 7805 288
rect 7889 -288 7923 288
rect 8007 -288 8041 288
rect 8125 -288 8159 288
rect 8243 -288 8277 288
rect 8361 -288 8395 288
rect 8479 -288 8513 288
rect 8597 -288 8631 288
rect 8715 -288 8749 288
rect 8833 -288 8867 288
rect -8808 -381 -8774 -347
rect -8690 -381 -8656 -347
rect -8572 -381 -8538 -347
rect -8454 -381 -8420 -347
rect -8336 -381 -8302 -347
rect -8218 -381 -8184 -347
rect -8100 -381 -8066 -347
rect -7982 -381 -7948 -347
rect -7864 -381 -7830 -347
rect -7746 -381 -7712 -347
rect -7628 -381 -7594 -347
rect -7510 -381 -7476 -347
rect -7392 -381 -7358 -347
rect -7274 -381 -7240 -347
rect -7156 -381 -7122 -347
rect -7038 -381 -7004 -347
rect -6920 -381 -6886 -347
rect -6802 -381 -6768 -347
rect -6684 -381 -6650 -347
rect -6566 -381 -6532 -347
rect -6448 -381 -6414 -347
rect -6330 -381 -6296 -347
rect -6212 -381 -6178 -347
rect -6094 -381 -6060 -347
rect -5976 -381 -5942 -347
rect -5858 -381 -5824 -347
rect -5740 -381 -5706 -347
rect -5622 -381 -5588 -347
rect -5504 -381 -5470 -347
rect -5386 -381 -5352 -347
rect -5268 -381 -5234 -347
rect -5150 -381 -5116 -347
rect -5032 -381 -4998 -347
rect -4914 -381 -4880 -347
rect -4796 -381 -4762 -347
rect -4678 -381 -4644 -347
rect -4560 -381 -4526 -347
rect -4442 -381 -4408 -347
rect -4324 -381 -4290 -347
rect -4206 -381 -4172 -347
rect -4088 -381 -4054 -347
rect -3970 -381 -3936 -347
rect -3852 -381 -3818 -347
rect -3734 -381 -3700 -347
rect -3616 -381 -3582 -347
rect -3498 -381 -3464 -347
rect -3380 -381 -3346 -347
rect -3262 -381 -3228 -347
rect -3144 -381 -3110 -347
rect -3026 -381 -2992 -347
rect -2908 -381 -2874 -347
rect -2790 -381 -2756 -347
rect -2672 -381 -2638 -347
rect -2554 -381 -2520 -347
rect -2436 -381 -2402 -347
rect -2318 -381 -2284 -347
rect -2200 -381 -2166 -347
rect -2082 -381 -2048 -347
rect -1964 -381 -1930 -347
rect -1846 -381 -1812 -347
rect -1728 -381 -1694 -347
rect -1610 -381 -1576 -347
rect -1492 -381 -1458 -347
rect -1374 -381 -1340 -347
rect -1256 -381 -1222 -347
rect -1138 -381 -1104 -347
rect -1020 -381 -986 -347
rect -902 -381 -868 -347
rect -784 -381 -750 -347
rect -666 -381 -632 -347
rect -548 -381 -514 -347
rect -430 -381 -396 -347
rect -312 -381 -278 -347
rect -194 -381 -160 -347
rect -76 -381 -42 -347
rect 42 -381 76 -347
rect 160 -381 194 -347
rect 278 -381 312 -347
rect 396 -381 430 -347
rect 514 -381 548 -347
rect 632 -381 666 -347
rect 750 -381 784 -347
rect 868 -381 902 -347
rect 986 -381 1020 -347
rect 1104 -381 1138 -347
rect 1222 -381 1256 -347
rect 1340 -381 1374 -347
rect 1458 -381 1492 -347
rect 1576 -381 1610 -347
rect 1694 -381 1728 -347
rect 1812 -381 1846 -347
rect 1930 -381 1964 -347
rect 2048 -381 2082 -347
rect 2166 -381 2200 -347
rect 2284 -381 2318 -347
rect 2402 -381 2436 -347
rect 2520 -381 2554 -347
rect 2638 -381 2672 -347
rect 2756 -381 2790 -347
rect 2874 -381 2908 -347
rect 2992 -381 3026 -347
rect 3110 -381 3144 -347
rect 3228 -381 3262 -347
rect 3346 -381 3380 -347
rect 3464 -381 3498 -347
rect 3582 -381 3616 -347
rect 3700 -381 3734 -347
rect 3818 -381 3852 -347
rect 3936 -381 3970 -347
rect 4054 -381 4088 -347
rect 4172 -381 4206 -347
rect 4290 -381 4324 -347
rect 4408 -381 4442 -347
rect 4526 -381 4560 -347
rect 4644 -381 4678 -347
rect 4762 -381 4796 -347
rect 4880 -381 4914 -347
rect 4998 -381 5032 -347
rect 5116 -381 5150 -347
rect 5234 -381 5268 -347
rect 5352 -381 5386 -347
rect 5470 -381 5504 -347
rect 5588 -381 5622 -347
rect 5706 -381 5740 -347
rect 5824 -381 5858 -347
rect 5942 -381 5976 -347
rect 6060 -381 6094 -347
rect 6178 -381 6212 -347
rect 6296 -381 6330 -347
rect 6414 -381 6448 -347
rect 6532 -381 6566 -347
rect 6650 -381 6684 -347
rect 6768 -381 6802 -347
rect 6886 -381 6920 -347
rect 7004 -381 7038 -347
rect 7122 -381 7156 -347
rect 7240 -381 7274 -347
rect 7358 -381 7392 -347
rect 7476 -381 7510 -347
rect 7594 -381 7628 -347
rect 7712 -381 7746 -347
rect 7830 -381 7864 -347
rect 7948 -381 7982 -347
rect 8066 -381 8100 -347
rect 8184 -381 8218 -347
rect 8302 -381 8336 -347
rect 8420 -381 8454 -347
rect 8538 -381 8572 -347
rect 8656 -381 8690 -347
rect 8774 -381 8808 -347
<< metal1 >>
rect -8820 381 -8762 387
rect -8820 347 -8808 381
rect -8774 347 -8762 381
rect -8820 341 -8762 347
rect -8702 381 -8644 387
rect -8702 347 -8690 381
rect -8656 347 -8644 381
rect -8702 341 -8644 347
rect -8584 381 -8526 387
rect -8584 347 -8572 381
rect -8538 347 -8526 381
rect -8584 341 -8526 347
rect -8466 381 -8408 387
rect -8466 347 -8454 381
rect -8420 347 -8408 381
rect -8466 341 -8408 347
rect -8348 381 -8290 387
rect -8348 347 -8336 381
rect -8302 347 -8290 381
rect -8348 341 -8290 347
rect -8230 381 -8172 387
rect -8230 347 -8218 381
rect -8184 347 -8172 381
rect -8230 341 -8172 347
rect -8112 381 -8054 387
rect -8112 347 -8100 381
rect -8066 347 -8054 381
rect -8112 341 -8054 347
rect -7994 381 -7936 387
rect -7994 347 -7982 381
rect -7948 347 -7936 381
rect -7994 341 -7936 347
rect -7876 381 -7818 387
rect -7876 347 -7864 381
rect -7830 347 -7818 381
rect -7876 341 -7818 347
rect -7758 381 -7700 387
rect -7758 347 -7746 381
rect -7712 347 -7700 381
rect -7758 341 -7700 347
rect -7640 381 -7582 387
rect -7640 347 -7628 381
rect -7594 347 -7582 381
rect -7640 341 -7582 347
rect -7522 381 -7464 387
rect -7522 347 -7510 381
rect -7476 347 -7464 381
rect -7522 341 -7464 347
rect -7404 381 -7346 387
rect -7404 347 -7392 381
rect -7358 347 -7346 381
rect -7404 341 -7346 347
rect -7286 381 -7228 387
rect -7286 347 -7274 381
rect -7240 347 -7228 381
rect -7286 341 -7228 347
rect -7168 381 -7110 387
rect -7168 347 -7156 381
rect -7122 347 -7110 381
rect -7168 341 -7110 347
rect -7050 381 -6992 387
rect -7050 347 -7038 381
rect -7004 347 -6992 381
rect -7050 341 -6992 347
rect -6932 381 -6874 387
rect -6932 347 -6920 381
rect -6886 347 -6874 381
rect -6932 341 -6874 347
rect -6814 381 -6756 387
rect -6814 347 -6802 381
rect -6768 347 -6756 381
rect -6814 341 -6756 347
rect -6696 381 -6638 387
rect -6696 347 -6684 381
rect -6650 347 -6638 381
rect -6696 341 -6638 347
rect -6578 381 -6520 387
rect -6578 347 -6566 381
rect -6532 347 -6520 381
rect -6578 341 -6520 347
rect -6460 381 -6402 387
rect -6460 347 -6448 381
rect -6414 347 -6402 381
rect -6460 341 -6402 347
rect -6342 381 -6284 387
rect -6342 347 -6330 381
rect -6296 347 -6284 381
rect -6342 341 -6284 347
rect -6224 381 -6166 387
rect -6224 347 -6212 381
rect -6178 347 -6166 381
rect -6224 341 -6166 347
rect -6106 381 -6048 387
rect -6106 347 -6094 381
rect -6060 347 -6048 381
rect -6106 341 -6048 347
rect -5988 381 -5930 387
rect -5988 347 -5976 381
rect -5942 347 -5930 381
rect -5988 341 -5930 347
rect -5870 381 -5812 387
rect -5870 347 -5858 381
rect -5824 347 -5812 381
rect -5870 341 -5812 347
rect -5752 381 -5694 387
rect -5752 347 -5740 381
rect -5706 347 -5694 381
rect -5752 341 -5694 347
rect -5634 381 -5576 387
rect -5634 347 -5622 381
rect -5588 347 -5576 381
rect -5634 341 -5576 347
rect -5516 381 -5458 387
rect -5516 347 -5504 381
rect -5470 347 -5458 381
rect -5516 341 -5458 347
rect -5398 381 -5340 387
rect -5398 347 -5386 381
rect -5352 347 -5340 381
rect -5398 341 -5340 347
rect -5280 381 -5222 387
rect -5280 347 -5268 381
rect -5234 347 -5222 381
rect -5280 341 -5222 347
rect -5162 381 -5104 387
rect -5162 347 -5150 381
rect -5116 347 -5104 381
rect -5162 341 -5104 347
rect -5044 381 -4986 387
rect -5044 347 -5032 381
rect -4998 347 -4986 381
rect -5044 341 -4986 347
rect -4926 381 -4868 387
rect -4926 347 -4914 381
rect -4880 347 -4868 381
rect -4926 341 -4868 347
rect -4808 381 -4750 387
rect -4808 347 -4796 381
rect -4762 347 -4750 381
rect -4808 341 -4750 347
rect -4690 381 -4632 387
rect -4690 347 -4678 381
rect -4644 347 -4632 381
rect -4690 341 -4632 347
rect -4572 381 -4514 387
rect -4572 347 -4560 381
rect -4526 347 -4514 381
rect -4572 341 -4514 347
rect -4454 381 -4396 387
rect -4454 347 -4442 381
rect -4408 347 -4396 381
rect -4454 341 -4396 347
rect -4336 381 -4278 387
rect -4336 347 -4324 381
rect -4290 347 -4278 381
rect -4336 341 -4278 347
rect -4218 381 -4160 387
rect -4218 347 -4206 381
rect -4172 347 -4160 381
rect -4218 341 -4160 347
rect -4100 381 -4042 387
rect -4100 347 -4088 381
rect -4054 347 -4042 381
rect -4100 341 -4042 347
rect -3982 381 -3924 387
rect -3982 347 -3970 381
rect -3936 347 -3924 381
rect -3982 341 -3924 347
rect -3864 381 -3806 387
rect -3864 347 -3852 381
rect -3818 347 -3806 381
rect -3864 341 -3806 347
rect -3746 381 -3688 387
rect -3746 347 -3734 381
rect -3700 347 -3688 381
rect -3746 341 -3688 347
rect -3628 381 -3570 387
rect -3628 347 -3616 381
rect -3582 347 -3570 381
rect -3628 341 -3570 347
rect -3510 381 -3452 387
rect -3510 347 -3498 381
rect -3464 347 -3452 381
rect -3510 341 -3452 347
rect -3392 381 -3334 387
rect -3392 347 -3380 381
rect -3346 347 -3334 381
rect -3392 341 -3334 347
rect -3274 381 -3216 387
rect -3274 347 -3262 381
rect -3228 347 -3216 381
rect -3274 341 -3216 347
rect -3156 381 -3098 387
rect -3156 347 -3144 381
rect -3110 347 -3098 381
rect -3156 341 -3098 347
rect -3038 381 -2980 387
rect -3038 347 -3026 381
rect -2992 347 -2980 381
rect -3038 341 -2980 347
rect -2920 381 -2862 387
rect -2920 347 -2908 381
rect -2874 347 -2862 381
rect -2920 341 -2862 347
rect -2802 381 -2744 387
rect -2802 347 -2790 381
rect -2756 347 -2744 381
rect -2802 341 -2744 347
rect -2684 381 -2626 387
rect -2684 347 -2672 381
rect -2638 347 -2626 381
rect -2684 341 -2626 347
rect -2566 381 -2508 387
rect -2566 347 -2554 381
rect -2520 347 -2508 381
rect -2566 341 -2508 347
rect -2448 381 -2390 387
rect -2448 347 -2436 381
rect -2402 347 -2390 381
rect -2448 341 -2390 347
rect -2330 381 -2272 387
rect -2330 347 -2318 381
rect -2284 347 -2272 381
rect -2330 341 -2272 347
rect -2212 381 -2154 387
rect -2212 347 -2200 381
rect -2166 347 -2154 381
rect -2212 341 -2154 347
rect -2094 381 -2036 387
rect -2094 347 -2082 381
rect -2048 347 -2036 381
rect -2094 341 -2036 347
rect -1976 381 -1918 387
rect -1976 347 -1964 381
rect -1930 347 -1918 381
rect -1976 341 -1918 347
rect -1858 381 -1800 387
rect -1858 347 -1846 381
rect -1812 347 -1800 381
rect -1858 341 -1800 347
rect -1740 381 -1682 387
rect -1740 347 -1728 381
rect -1694 347 -1682 381
rect -1740 341 -1682 347
rect -1622 381 -1564 387
rect -1622 347 -1610 381
rect -1576 347 -1564 381
rect -1622 341 -1564 347
rect -1504 381 -1446 387
rect -1504 347 -1492 381
rect -1458 347 -1446 381
rect -1504 341 -1446 347
rect -1386 381 -1328 387
rect -1386 347 -1374 381
rect -1340 347 -1328 381
rect -1386 341 -1328 347
rect -1268 381 -1210 387
rect -1268 347 -1256 381
rect -1222 347 -1210 381
rect -1268 341 -1210 347
rect -1150 381 -1092 387
rect -1150 347 -1138 381
rect -1104 347 -1092 381
rect -1150 341 -1092 347
rect -1032 381 -974 387
rect -1032 347 -1020 381
rect -986 347 -974 381
rect -1032 341 -974 347
rect -914 381 -856 387
rect -914 347 -902 381
rect -868 347 -856 381
rect -914 341 -856 347
rect -796 381 -738 387
rect -796 347 -784 381
rect -750 347 -738 381
rect -796 341 -738 347
rect -678 381 -620 387
rect -678 347 -666 381
rect -632 347 -620 381
rect -678 341 -620 347
rect -560 381 -502 387
rect -560 347 -548 381
rect -514 347 -502 381
rect -560 341 -502 347
rect -442 381 -384 387
rect -442 347 -430 381
rect -396 347 -384 381
rect -442 341 -384 347
rect -324 381 -266 387
rect -324 347 -312 381
rect -278 347 -266 381
rect -324 341 -266 347
rect -206 381 -148 387
rect -206 347 -194 381
rect -160 347 -148 381
rect -206 341 -148 347
rect -88 381 -30 387
rect -88 347 -76 381
rect -42 347 -30 381
rect -88 341 -30 347
rect 30 381 88 387
rect 30 347 42 381
rect 76 347 88 381
rect 30 341 88 347
rect 148 381 206 387
rect 148 347 160 381
rect 194 347 206 381
rect 148 341 206 347
rect 266 381 324 387
rect 266 347 278 381
rect 312 347 324 381
rect 266 341 324 347
rect 384 381 442 387
rect 384 347 396 381
rect 430 347 442 381
rect 384 341 442 347
rect 502 381 560 387
rect 502 347 514 381
rect 548 347 560 381
rect 502 341 560 347
rect 620 381 678 387
rect 620 347 632 381
rect 666 347 678 381
rect 620 341 678 347
rect 738 381 796 387
rect 738 347 750 381
rect 784 347 796 381
rect 738 341 796 347
rect 856 381 914 387
rect 856 347 868 381
rect 902 347 914 381
rect 856 341 914 347
rect 974 381 1032 387
rect 974 347 986 381
rect 1020 347 1032 381
rect 974 341 1032 347
rect 1092 381 1150 387
rect 1092 347 1104 381
rect 1138 347 1150 381
rect 1092 341 1150 347
rect 1210 381 1268 387
rect 1210 347 1222 381
rect 1256 347 1268 381
rect 1210 341 1268 347
rect 1328 381 1386 387
rect 1328 347 1340 381
rect 1374 347 1386 381
rect 1328 341 1386 347
rect 1446 381 1504 387
rect 1446 347 1458 381
rect 1492 347 1504 381
rect 1446 341 1504 347
rect 1564 381 1622 387
rect 1564 347 1576 381
rect 1610 347 1622 381
rect 1564 341 1622 347
rect 1682 381 1740 387
rect 1682 347 1694 381
rect 1728 347 1740 381
rect 1682 341 1740 347
rect 1800 381 1858 387
rect 1800 347 1812 381
rect 1846 347 1858 381
rect 1800 341 1858 347
rect 1918 381 1976 387
rect 1918 347 1930 381
rect 1964 347 1976 381
rect 1918 341 1976 347
rect 2036 381 2094 387
rect 2036 347 2048 381
rect 2082 347 2094 381
rect 2036 341 2094 347
rect 2154 381 2212 387
rect 2154 347 2166 381
rect 2200 347 2212 381
rect 2154 341 2212 347
rect 2272 381 2330 387
rect 2272 347 2284 381
rect 2318 347 2330 381
rect 2272 341 2330 347
rect 2390 381 2448 387
rect 2390 347 2402 381
rect 2436 347 2448 381
rect 2390 341 2448 347
rect 2508 381 2566 387
rect 2508 347 2520 381
rect 2554 347 2566 381
rect 2508 341 2566 347
rect 2626 381 2684 387
rect 2626 347 2638 381
rect 2672 347 2684 381
rect 2626 341 2684 347
rect 2744 381 2802 387
rect 2744 347 2756 381
rect 2790 347 2802 381
rect 2744 341 2802 347
rect 2862 381 2920 387
rect 2862 347 2874 381
rect 2908 347 2920 381
rect 2862 341 2920 347
rect 2980 381 3038 387
rect 2980 347 2992 381
rect 3026 347 3038 381
rect 2980 341 3038 347
rect 3098 381 3156 387
rect 3098 347 3110 381
rect 3144 347 3156 381
rect 3098 341 3156 347
rect 3216 381 3274 387
rect 3216 347 3228 381
rect 3262 347 3274 381
rect 3216 341 3274 347
rect 3334 381 3392 387
rect 3334 347 3346 381
rect 3380 347 3392 381
rect 3334 341 3392 347
rect 3452 381 3510 387
rect 3452 347 3464 381
rect 3498 347 3510 381
rect 3452 341 3510 347
rect 3570 381 3628 387
rect 3570 347 3582 381
rect 3616 347 3628 381
rect 3570 341 3628 347
rect 3688 381 3746 387
rect 3688 347 3700 381
rect 3734 347 3746 381
rect 3688 341 3746 347
rect 3806 381 3864 387
rect 3806 347 3818 381
rect 3852 347 3864 381
rect 3806 341 3864 347
rect 3924 381 3982 387
rect 3924 347 3936 381
rect 3970 347 3982 381
rect 3924 341 3982 347
rect 4042 381 4100 387
rect 4042 347 4054 381
rect 4088 347 4100 381
rect 4042 341 4100 347
rect 4160 381 4218 387
rect 4160 347 4172 381
rect 4206 347 4218 381
rect 4160 341 4218 347
rect 4278 381 4336 387
rect 4278 347 4290 381
rect 4324 347 4336 381
rect 4278 341 4336 347
rect 4396 381 4454 387
rect 4396 347 4408 381
rect 4442 347 4454 381
rect 4396 341 4454 347
rect 4514 381 4572 387
rect 4514 347 4526 381
rect 4560 347 4572 381
rect 4514 341 4572 347
rect 4632 381 4690 387
rect 4632 347 4644 381
rect 4678 347 4690 381
rect 4632 341 4690 347
rect 4750 381 4808 387
rect 4750 347 4762 381
rect 4796 347 4808 381
rect 4750 341 4808 347
rect 4868 381 4926 387
rect 4868 347 4880 381
rect 4914 347 4926 381
rect 4868 341 4926 347
rect 4986 381 5044 387
rect 4986 347 4998 381
rect 5032 347 5044 381
rect 4986 341 5044 347
rect 5104 381 5162 387
rect 5104 347 5116 381
rect 5150 347 5162 381
rect 5104 341 5162 347
rect 5222 381 5280 387
rect 5222 347 5234 381
rect 5268 347 5280 381
rect 5222 341 5280 347
rect 5340 381 5398 387
rect 5340 347 5352 381
rect 5386 347 5398 381
rect 5340 341 5398 347
rect 5458 381 5516 387
rect 5458 347 5470 381
rect 5504 347 5516 381
rect 5458 341 5516 347
rect 5576 381 5634 387
rect 5576 347 5588 381
rect 5622 347 5634 381
rect 5576 341 5634 347
rect 5694 381 5752 387
rect 5694 347 5706 381
rect 5740 347 5752 381
rect 5694 341 5752 347
rect 5812 381 5870 387
rect 5812 347 5824 381
rect 5858 347 5870 381
rect 5812 341 5870 347
rect 5930 381 5988 387
rect 5930 347 5942 381
rect 5976 347 5988 381
rect 5930 341 5988 347
rect 6048 381 6106 387
rect 6048 347 6060 381
rect 6094 347 6106 381
rect 6048 341 6106 347
rect 6166 381 6224 387
rect 6166 347 6178 381
rect 6212 347 6224 381
rect 6166 341 6224 347
rect 6284 381 6342 387
rect 6284 347 6296 381
rect 6330 347 6342 381
rect 6284 341 6342 347
rect 6402 381 6460 387
rect 6402 347 6414 381
rect 6448 347 6460 381
rect 6402 341 6460 347
rect 6520 381 6578 387
rect 6520 347 6532 381
rect 6566 347 6578 381
rect 6520 341 6578 347
rect 6638 381 6696 387
rect 6638 347 6650 381
rect 6684 347 6696 381
rect 6638 341 6696 347
rect 6756 381 6814 387
rect 6756 347 6768 381
rect 6802 347 6814 381
rect 6756 341 6814 347
rect 6874 381 6932 387
rect 6874 347 6886 381
rect 6920 347 6932 381
rect 6874 341 6932 347
rect 6992 381 7050 387
rect 6992 347 7004 381
rect 7038 347 7050 381
rect 6992 341 7050 347
rect 7110 381 7168 387
rect 7110 347 7122 381
rect 7156 347 7168 381
rect 7110 341 7168 347
rect 7228 381 7286 387
rect 7228 347 7240 381
rect 7274 347 7286 381
rect 7228 341 7286 347
rect 7346 381 7404 387
rect 7346 347 7358 381
rect 7392 347 7404 381
rect 7346 341 7404 347
rect 7464 381 7522 387
rect 7464 347 7476 381
rect 7510 347 7522 381
rect 7464 341 7522 347
rect 7582 381 7640 387
rect 7582 347 7594 381
rect 7628 347 7640 381
rect 7582 341 7640 347
rect 7700 381 7758 387
rect 7700 347 7712 381
rect 7746 347 7758 381
rect 7700 341 7758 347
rect 7818 381 7876 387
rect 7818 347 7830 381
rect 7864 347 7876 381
rect 7818 341 7876 347
rect 7936 381 7994 387
rect 7936 347 7948 381
rect 7982 347 7994 381
rect 7936 341 7994 347
rect 8054 381 8112 387
rect 8054 347 8066 381
rect 8100 347 8112 381
rect 8054 341 8112 347
rect 8172 381 8230 387
rect 8172 347 8184 381
rect 8218 347 8230 381
rect 8172 341 8230 347
rect 8290 381 8348 387
rect 8290 347 8302 381
rect 8336 347 8348 381
rect 8290 341 8348 347
rect 8408 381 8466 387
rect 8408 347 8420 381
rect 8454 347 8466 381
rect 8408 341 8466 347
rect 8526 381 8584 387
rect 8526 347 8538 381
rect 8572 347 8584 381
rect 8526 341 8584 347
rect 8644 381 8702 387
rect 8644 347 8656 381
rect 8690 347 8702 381
rect 8644 341 8702 347
rect 8762 381 8820 387
rect 8762 347 8774 381
rect 8808 347 8820 381
rect 8762 341 8820 347
rect -8873 288 -8827 300
rect -8873 -288 -8867 288
rect -8833 -288 -8827 288
rect -8873 -300 -8827 -288
rect -8755 288 -8709 300
rect -8755 -288 -8749 288
rect -8715 -288 -8709 288
rect -8755 -300 -8709 -288
rect -8637 288 -8591 300
rect -8637 -288 -8631 288
rect -8597 -288 -8591 288
rect -8637 -300 -8591 -288
rect -8519 288 -8473 300
rect -8519 -288 -8513 288
rect -8479 -288 -8473 288
rect -8519 -300 -8473 -288
rect -8401 288 -8355 300
rect -8401 -288 -8395 288
rect -8361 -288 -8355 288
rect -8401 -300 -8355 -288
rect -8283 288 -8237 300
rect -8283 -288 -8277 288
rect -8243 -288 -8237 288
rect -8283 -300 -8237 -288
rect -8165 288 -8119 300
rect -8165 -288 -8159 288
rect -8125 -288 -8119 288
rect -8165 -300 -8119 -288
rect -8047 288 -8001 300
rect -8047 -288 -8041 288
rect -8007 -288 -8001 288
rect -8047 -300 -8001 -288
rect -7929 288 -7883 300
rect -7929 -288 -7923 288
rect -7889 -288 -7883 288
rect -7929 -300 -7883 -288
rect -7811 288 -7765 300
rect -7811 -288 -7805 288
rect -7771 -288 -7765 288
rect -7811 -300 -7765 -288
rect -7693 288 -7647 300
rect -7693 -288 -7687 288
rect -7653 -288 -7647 288
rect -7693 -300 -7647 -288
rect -7575 288 -7529 300
rect -7575 -288 -7569 288
rect -7535 -288 -7529 288
rect -7575 -300 -7529 -288
rect -7457 288 -7411 300
rect -7457 -288 -7451 288
rect -7417 -288 -7411 288
rect -7457 -300 -7411 -288
rect -7339 288 -7293 300
rect -7339 -288 -7333 288
rect -7299 -288 -7293 288
rect -7339 -300 -7293 -288
rect -7221 288 -7175 300
rect -7221 -288 -7215 288
rect -7181 -288 -7175 288
rect -7221 -300 -7175 -288
rect -7103 288 -7057 300
rect -7103 -288 -7097 288
rect -7063 -288 -7057 288
rect -7103 -300 -7057 -288
rect -6985 288 -6939 300
rect -6985 -288 -6979 288
rect -6945 -288 -6939 288
rect -6985 -300 -6939 -288
rect -6867 288 -6821 300
rect -6867 -288 -6861 288
rect -6827 -288 -6821 288
rect -6867 -300 -6821 -288
rect -6749 288 -6703 300
rect -6749 -288 -6743 288
rect -6709 -288 -6703 288
rect -6749 -300 -6703 -288
rect -6631 288 -6585 300
rect -6631 -288 -6625 288
rect -6591 -288 -6585 288
rect -6631 -300 -6585 -288
rect -6513 288 -6467 300
rect -6513 -288 -6507 288
rect -6473 -288 -6467 288
rect -6513 -300 -6467 -288
rect -6395 288 -6349 300
rect -6395 -288 -6389 288
rect -6355 -288 -6349 288
rect -6395 -300 -6349 -288
rect -6277 288 -6231 300
rect -6277 -288 -6271 288
rect -6237 -288 -6231 288
rect -6277 -300 -6231 -288
rect -6159 288 -6113 300
rect -6159 -288 -6153 288
rect -6119 -288 -6113 288
rect -6159 -300 -6113 -288
rect -6041 288 -5995 300
rect -6041 -288 -6035 288
rect -6001 -288 -5995 288
rect -6041 -300 -5995 -288
rect -5923 288 -5877 300
rect -5923 -288 -5917 288
rect -5883 -288 -5877 288
rect -5923 -300 -5877 -288
rect -5805 288 -5759 300
rect -5805 -288 -5799 288
rect -5765 -288 -5759 288
rect -5805 -300 -5759 -288
rect -5687 288 -5641 300
rect -5687 -288 -5681 288
rect -5647 -288 -5641 288
rect -5687 -300 -5641 -288
rect -5569 288 -5523 300
rect -5569 -288 -5563 288
rect -5529 -288 -5523 288
rect -5569 -300 -5523 -288
rect -5451 288 -5405 300
rect -5451 -288 -5445 288
rect -5411 -288 -5405 288
rect -5451 -300 -5405 -288
rect -5333 288 -5287 300
rect -5333 -288 -5327 288
rect -5293 -288 -5287 288
rect -5333 -300 -5287 -288
rect -5215 288 -5169 300
rect -5215 -288 -5209 288
rect -5175 -288 -5169 288
rect -5215 -300 -5169 -288
rect -5097 288 -5051 300
rect -5097 -288 -5091 288
rect -5057 -288 -5051 288
rect -5097 -300 -5051 -288
rect -4979 288 -4933 300
rect -4979 -288 -4973 288
rect -4939 -288 -4933 288
rect -4979 -300 -4933 -288
rect -4861 288 -4815 300
rect -4861 -288 -4855 288
rect -4821 -288 -4815 288
rect -4861 -300 -4815 -288
rect -4743 288 -4697 300
rect -4743 -288 -4737 288
rect -4703 -288 -4697 288
rect -4743 -300 -4697 -288
rect -4625 288 -4579 300
rect -4625 -288 -4619 288
rect -4585 -288 -4579 288
rect -4625 -300 -4579 -288
rect -4507 288 -4461 300
rect -4507 -288 -4501 288
rect -4467 -288 -4461 288
rect -4507 -300 -4461 -288
rect -4389 288 -4343 300
rect -4389 -288 -4383 288
rect -4349 -288 -4343 288
rect -4389 -300 -4343 -288
rect -4271 288 -4225 300
rect -4271 -288 -4265 288
rect -4231 -288 -4225 288
rect -4271 -300 -4225 -288
rect -4153 288 -4107 300
rect -4153 -288 -4147 288
rect -4113 -288 -4107 288
rect -4153 -300 -4107 -288
rect -4035 288 -3989 300
rect -4035 -288 -4029 288
rect -3995 -288 -3989 288
rect -4035 -300 -3989 -288
rect -3917 288 -3871 300
rect -3917 -288 -3911 288
rect -3877 -288 -3871 288
rect -3917 -300 -3871 -288
rect -3799 288 -3753 300
rect -3799 -288 -3793 288
rect -3759 -288 -3753 288
rect -3799 -300 -3753 -288
rect -3681 288 -3635 300
rect -3681 -288 -3675 288
rect -3641 -288 -3635 288
rect -3681 -300 -3635 -288
rect -3563 288 -3517 300
rect -3563 -288 -3557 288
rect -3523 -288 -3517 288
rect -3563 -300 -3517 -288
rect -3445 288 -3399 300
rect -3445 -288 -3439 288
rect -3405 -288 -3399 288
rect -3445 -300 -3399 -288
rect -3327 288 -3281 300
rect -3327 -288 -3321 288
rect -3287 -288 -3281 288
rect -3327 -300 -3281 -288
rect -3209 288 -3163 300
rect -3209 -288 -3203 288
rect -3169 -288 -3163 288
rect -3209 -300 -3163 -288
rect -3091 288 -3045 300
rect -3091 -288 -3085 288
rect -3051 -288 -3045 288
rect -3091 -300 -3045 -288
rect -2973 288 -2927 300
rect -2973 -288 -2967 288
rect -2933 -288 -2927 288
rect -2973 -300 -2927 -288
rect -2855 288 -2809 300
rect -2855 -288 -2849 288
rect -2815 -288 -2809 288
rect -2855 -300 -2809 -288
rect -2737 288 -2691 300
rect -2737 -288 -2731 288
rect -2697 -288 -2691 288
rect -2737 -300 -2691 -288
rect -2619 288 -2573 300
rect -2619 -288 -2613 288
rect -2579 -288 -2573 288
rect -2619 -300 -2573 -288
rect -2501 288 -2455 300
rect -2501 -288 -2495 288
rect -2461 -288 -2455 288
rect -2501 -300 -2455 -288
rect -2383 288 -2337 300
rect -2383 -288 -2377 288
rect -2343 -288 -2337 288
rect -2383 -300 -2337 -288
rect -2265 288 -2219 300
rect -2265 -288 -2259 288
rect -2225 -288 -2219 288
rect -2265 -300 -2219 -288
rect -2147 288 -2101 300
rect -2147 -288 -2141 288
rect -2107 -288 -2101 288
rect -2147 -300 -2101 -288
rect -2029 288 -1983 300
rect -2029 -288 -2023 288
rect -1989 -288 -1983 288
rect -2029 -300 -1983 -288
rect -1911 288 -1865 300
rect -1911 -288 -1905 288
rect -1871 -288 -1865 288
rect -1911 -300 -1865 -288
rect -1793 288 -1747 300
rect -1793 -288 -1787 288
rect -1753 -288 -1747 288
rect -1793 -300 -1747 -288
rect -1675 288 -1629 300
rect -1675 -288 -1669 288
rect -1635 -288 -1629 288
rect -1675 -300 -1629 -288
rect -1557 288 -1511 300
rect -1557 -288 -1551 288
rect -1517 -288 -1511 288
rect -1557 -300 -1511 -288
rect -1439 288 -1393 300
rect -1439 -288 -1433 288
rect -1399 -288 -1393 288
rect -1439 -300 -1393 -288
rect -1321 288 -1275 300
rect -1321 -288 -1315 288
rect -1281 -288 -1275 288
rect -1321 -300 -1275 -288
rect -1203 288 -1157 300
rect -1203 -288 -1197 288
rect -1163 -288 -1157 288
rect -1203 -300 -1157 -288
rect -1085 288 -1039 300
rect -1085 -288 -1079 288
rect -1045 -288 -1039 288
rect -1085 -300 -1039 -288
rect -967 288 -921 300
rect -967 -288 -961 288
rect -927 -288 -921 288
rect -967 -300 -921 -288
rect -849 288 -803 300
rect -849 -288 -843 288
rect -809 -288 -803 288
rect -849 -300 -803 -288
rect -731 288 -685 300
rect -731 -288 -725 288
rect -691 -288 -685 288
rect -731 -300 -685 -288
rect -613 288 -567 300
rect -613 -288 -607 288
rect -573 -288 -567 288
rect -613 -300 -567 -288
rect -495 288 -449 300
rect -495 -288 -489 288
rect -455 -288 -449 288
rect -495 -300 -449 -288
rect -377 288 -331 300
rect -377 -288 -371 288
rect -337 -288 -331 288
rect -377 -300 -331 -288
rect -259 288 -213 300
rect -259 -288 -253 288
rect -219 -288 -213 288
rect -259 -300 -213 -288
rect -141 288 -95 300
rect -141 -288 -135 288
rect -101 -288 -95 288
rect -141 -300 -95 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 95 288 141 300
rect 95 -288 101 288
rect 135 -288 141 288
rect 95 -300 141 -288
rect 213 288 259 300
rect 213 -288 219 288
rect 253 -288 259 288
rect 213 -300 259 -288
rect 331 288 377 300
rect 331 -288 337 288
rect 371 -288 377 288
rect 331 -300 377 -288
rect 449 288 495 300
rect 449 -288 455 288
rect 489 -288 495 288
rect 449 -300 495 -288
rect 567 288 613 300
rect 567 -288 573 288
rect 607 -288 613 288
rect 567 -300 613 -288
rect 685 288 731 300
rect 685 -288 691 288
rect 725 -288 731 288
rect 685 -300 731 -288
rect 803 288 849 300
rect 803 -288 809 288
rect 843 -288 849 288
rect 803 -300 849 -288
rect 921 288 967 300
rect 921 -288 927 288
rect 961 -288 967 288
rect 921 -300 967 -288
rect 1039 288 1085 300
rect 1039 -288 1045 288
rect 1079 -288 1085 288
rect 1039 -300 1085 -288
rect 1157 288 1203 300
rect 1157 -288 1163 288
rect 1197 -288 1203 288
rect 1157 -300 1203 -288
rect 1275 288 1321 300
rect 1275 -288 1281 288
rect 1315 -288 1321 288
rect 1275 -300 1321 -288
rect 1393 288 1439 300
rect 1393 -288 1399 288
rect 1433 -288 1439 288
rect 1393 -300 1439 -288
rect 1511 288 1557 300
rect 1511 -288 1517 288
rect 1551 -288 1557 288
rect 1511 -300 1557 -288
rect 1629 288 1675 300
rect 1629 -288 1635 288
rect 1669 -288 1675 288
rect 1629 -300 1675 -288
rect 1747 288 1793 300
rect 1747 -288 1753 288
rect 1787 -288 1793 288
rect 1747 -300 1793 -288
rect 1865 288 1911 300
rect 1865 -288 1871 288
rect 1905 -288 1911 288
rect 1865 -300 1911 -288
rect 1983 288 2029 300
rect 1983 -288 1989 288
rect 2023 -288 2029 288
rect 1983 -300 2029 -288
rect 2101 288 2147 300
rect 2101 -288 2107 288
rect 2141 -288 2147 288
rect 2101 -300 2147 -288
rect 2219 288 2265 300
rect 2219 -288 2225 288
rect 2259 -288 2265 288
rect 2219 -300 2265 -288
rect 2337 288 2383 300
rect 2337 -288 2343 288
rect 2377 -288 2383 288
rect 2337 -300 2383 -288
rect 2455 288 2501 300
rect 2455 -288 2461 288
rect 2495 -288 2501 288
rect 2455 -300 2501 -288
rect 2573 288 2619 300
rect 2573 -288 2579 288
rect 2613 -288 2619 288
rect 2573 -300 2619 -288
rect 2691 288 2737 300
rect 2691 -288 2697 288
rect 2731 -288 2737 288
rect 2691 -300 2737 -288
rect 2809 288 2855 300
rect 2809 -288 2815 288
rect 2849 -288 2855 288
rect 2809 -300 2855 -288
rect 2927 288 2973 300
rect 2927 -288 2933 288
rect 2967 -288 2973 288
rect 2927 -300 2973 -288
rect 3045 288 3091 300
rect 3045 -288 3051 288
rect 3085 -288 3091 288
rect 3045 -300 3091 -288
rect 3163 288 3209 300
rect 3163 -288 3169 288
rect 3203 -288 3209 288
rect 3163 -300 3209 -288
rect 3281 288 3327 300
rect 3281 -288 3287 288
rect 3321 -288 3327 288
rect 3281 -300 3327 -288
rect 3399 288 3445 300
rect 3399 -288 3405 288
rect 3439 -288 3445 288
rect 3399 -300 3445 -288
rect 3517 288 3563 300
rect 3517 -288 3523 288
rect 3557 -288 3563 288
rect 3517 -300 3563 -288
rect 3635 288 3681 300
rect 3635 -288 3641 288
rect 3675 -288 3681 288
rect 3635 -300 3681 -288
rect 3753 288 3799 300
rect 3753 -288 3759 288
rect 3793 -288 3799 288
rect 3753 -300 3799 -288
rect 3871 288 3917 300
rect 3871 -288 3877 288
rect 3911 -288 3917 288
rect 3871 -300 3917 -288
rect 3989 288 4035 300
rect 3989 -288 3995 288
rect 4029 -288 4035 288
rect 3989 -300 4035 -288
rect 4107 288 4153 300
rect 4107 -288 4113 288
rect 4147 -288 4153 288
rect 4107 -300 4153 -288
rect 4225 288 4271 300
rect 4225 -288 4231 288
rect 4265 -288 4271 288
rect 4225 -300 4271 -288
rect 4343 288 4389 300
rect 4343 -288 4349 288
rect 4383 -288 4389 288
rect 4343 -300 4389 -288
rect 4461 288 4507 300
rect 4461 -288 4467 288
rect 4501 -288 4507 288
rect 4461 -300 4507 -288
rect 4579 288 4625 300
rect 4579 -288 4585 288
rect 4619 -288 4625 288
rect 4579 -300 4625 -288
rect 4697 288 4743 300
rect 4697 -288 4703 288
rect 4737 -288 4743 288
rect 4697 -300 4743 -288
rect 4815 288 4861 300
rect 4815 -288 4821 288
rect 4855 -288 4861 288
rect 4815 -300 4861 -288
rect 4933 288 4979 300
rect 4933 -288 4939 288
rect 4973 -288 4979 288
rect 4933 -300 4979 -288
rect 5051 288 5097 300
rect 5051 -288 5057 288
rect 5091 -288 5097 288
rect 5051 -300 5097 -288
rect 5169 288 5215 300
rect 5169 -288 5175 288
rect 5209 -288 5215 288
rect 5169 -300 5215 -288
rect 5287 288 5333 300
rect 5287 -288 5293 288
rect 5327 -288 5333 288
rect 5287 -300 5333 -288
rect 5405 288 5451 300
rect 5405 -288 5411 288
rect 5445 -288 5451 288
rect 5405 -300 5451 -288
rect 5523 288 5569 300
rect 5523 -288 5529 288
rect 5563 -288 5569 288
rect 5523 -300 5569 -288
rect 5641 288 5687 300
rect 5641 -288 5647 288
rect 5681 -288 5687 288
rect 5641 -300 5687 -288
rect 5759 288 5805 300
rect 5759 -288 5765 288
rect 5799 -288 5805 288
rect 5759 -300 5805 -288
rect 5877 288 5923 300
rect 5877 -288 5883 288
rect 5917 -288 5923 288
rect 5877 -300 5923 -288
rect 5995 288 6041 300
rect 5995 -288 6001 288
rect 6035 -288 6041 288
rect 5995 -300 6041 -288
rect 6113 288 6159 300
rect 6113 -288 6119 288
rect 6153 -288 6159 288
rect 6113 -300 6159 -288
rect 6231 288 6277 300
rect 6231 -288 6237 288
rect 6271 -288 6277 288
rect 6231 -300 6277 -288
rect 6349 288 6395 300
rect 6349 -288 6355 288
rect 6389 -288 6395 288
rect 6349 -300 6395 -288
rect 6467 288 6513 300
rect 6467 -288 6473 288
rect 6507 -288 6513 288
rect 6467 -300 6513 -288
rect 6585 288 6631 300
rect 6585 -288 6591 288
rect 6625 -288 6631 288
rect 6585 -300 6631 -288
rect 6703 288 6749 300
rect 6703 -288 6709 288
rect 6743 -288 6749 288
rect 6703 -300 6749 -288
rect 6821 288 6867 300
rect 6821 -288 6827 288
rect 6861 -288 6867 288
rect 6821 -300 6867 -288
rect 6939 288 6985 300
rect 6939 -288 6945 288
rect 6979 -288 6985 288
rect 6939 -300 6985 -288
rect 7057 288 7103 300
rect 7057 -288 7063 288
rect 7097 -288 7103 288
rect 7057 -300 7103 -288
rect 7175 288 7221 300
rect 7175 -288 7181 288
rect 7215 -288 7221 288
rect 7175 -300 7221 -288
rect 7293 288 7339 300
rect 7293 -288 7299 288
rect 7333 -288 7339 288
rect 7293 -300 7339 -288
rect 7411 288 7457 300
rect 7411 -288 7417 288
rect 7451 -288 7457 288
rect 7411 -300 7457 -288
rect 7529 288 7575 300
rect 7529 -288 7535 288
rect 7569 -288 7575 288
rect 7529 -300 7575 -288
rect 7647 288 7693 300
rect 7647 -288 7653 288
rect 7687 -288 7693 288
rect 7647 -300 7693 -288
rect 7765 288 7811 300
rect 7765 -288 7771 288
rect 7805 -288 7811 288
rect 7765 -300 7811 -288
rect 7883 288 7929 300
rect 7883 -288 7889 288
rect 7923 -288 7929 288
rect 7883 -300 7929 -288
rect 8001 288 8047 300
rect 8001 -288 8007 288
rect 8041 -288 8047 288
rect 8001 -300 8047 -288
rect 8119 288 8165 300
rect 8119 -288 8125 288
rect 8159 -288 8165 288
rect 8119 -300 8165 -288
rect 8237 288 8283 300
rect 8237 -288 8243 288
rect 8277 -288 8283 288
rect 8237 -300 8283 -288
rect 8355 288 8401 300
rect 8355 -288 8361 288
rect 8395 -288 8401 288
rect 8355 -300 8401 -288
rect 8473 288 8519 300
rect 8473 -288 8479 288
rect 8513 -288 8519 288
rect 8473 -300 8519 -288
rect 8591 288 8637 300
rect 8591 -288 8597 288
rect 8631 -288 8637 288
rect 8591 -300 8637 -288
rect 8709 288 8755 300
rect 8709 -288 8715 288
rect 8749 -288 8755 288
rect 8709 -300 8755 -288
rect 8827 288 8873 300
rect 8827 -288 8833 288
rect 8867 -288 8873 288
rect 8827 -300 8873 -288
rect -8820 -347 -8762 -341
rect -8820 -381 -8808 -347
rect -8774 -381 -8762 -347
rect -8820 -387 -8762 -381
rect -8702 -347 -8644 -341
rect -8702 -381 -8690 -347
rect -8656 -381 -8644 -347
rect -8702 -387 -8644 -381
rect -8584 -347 -8526 -341
rect -8584 -381 -8572 -347
rect -8538 -381 -8526 -347
rect -8584 -387 -8526 -381
rect -8466 -347 -8408 -341
rect -8466 -381 -8454 -347
rect -8420 -381 -8408 -347
rect -8466 -387 -8408 -381
rect -8348 -347 -8290 -341
rect -8348 -381 -8336 -347
rect -8302 -381 -8290 -347
rect -8348 -387 -8290 -381
rect -8230 -347 -8172 -341
rect -8230 -381 -8218 -347
rect -8184 -381 -8172 -347
rect -8230 -387 -8172 -381
rect -8112 -347 -8054 -341
rect -8112 -381 -8100 -347
rect -8066 -381 -8054 -347
rect -8112 -387 -8054 -381
rect -7994 -347 -7936 -341
rect -7994 -381 -7982 -347
rect -7948 -381 -7936 -347
rect -7994 -387 -7936 -381
rect -7876 -347 -7818 -341
rect -7876 -381 -7864 -347
rect -7830 -381 -7818 -347
rect -7876 -387 -7818 -381
rect -7758 -347 -7700 -341
rect -7758 -381 -7746 -347
rect -7712 -381 -7700 -347
rect -7758 -387 -7700 -381
rect -7640 -347 -7582 -341
rect -7640 -381 -7628 -347
rect -7594 -381 -7582 -347
rect -7640 -387 -7582 -381
rect -7522 -347 -7464 -341
rect -7522 -381 -7510 -347
rect -7476 -381 -7464 -347
rect -7522 -387 -7464 -381
rect -7404 -347 -7346 -341
rect -7404 -381 -7392 -347
rect -7358 -381 -7346 -347
rect -7404 -387 -7346 -381
rect -7286 -347 -7228 -341
rect -7286 -381 -7274 -347
rect -7240 -381 -7228 -347
rect -7286 -387 -7228 -381
rect -7168 -347 -7110 -341
rect -7168 -381 -7156 -347
rect -7122 -381 -7110 -347
rect -7168 -387 -7110 -381
rect -7050 -347 -6992 -341
rect -7050 -381 -7038 -347
rect -7004 -381 -6992 -347
rect -7050 -387 -6992 -381
rect -6932 -347 -6874 -341
rect -6932 -381 -6920 -347
rect -6886 -381 -6874 -347
rect -6932 -387 -6874 -381
rect -6814 -347 -6756 -341
rect -6814 -381 -6802 -347
rect -6768 -381 -6756 -347
rect -6814 -387 -6756 -381
rect -6696 -347 -6638 -341
rect -6696 -381 -6684 -347
rect -6650 -381 -6638 -347
rect -6696 -387 -6638 -381
rect -6578 -347 -6520 -341
rect -6578 -381 -6566 -347
rect -6532 -381 -6520 -347
rect -6578 -387 -6520 -381
rect -6460 -347 -6402 -341
rect -6460 -381 -6448 -347
rect -6414 -381 -6402 -347
rect -6460 -387 -6402 -381
rect -6342 -347 -6284 -341
rect -6342 -381 -6330 -347
rect -6296 -381 -6284 -347
rect -6342 -387 -6284 -381
rect -6224 -347 -6166 -341
rect -6224 -381 -6212 -347
rect -6178 -381 -6166 -347
rect -6224 -387 -6166 -381
rect -6106 -347 -6048 -341
rect -6106 -381 -6094 -347
rect -6060 -381 -6048 -347
rect -6106 -387 -6048 -381
rect -5988 -347 -5930 -341
rect -5988 -381 -5976 -347
rect -5942 -381 -5930 -347
rect -5988 -387 -5930 -381
rect -5870 -347 -5812 -341
rect -5870 -381 -5858 -347
rect -5824 -381 -5812 -347
rect -5870 -387 -5812 -381
rect -5752 -347 -5694 -341
rect -5752 -381 -5740 -347
rect -5706 -381 -5694 -347
rect -5752 -387 -5694 -381
rect -5634 -347 -5576 -341
rect -5634 -381 -5622 -347
rect -5588 -381 -5576 -347
rect -5634 -387 -5576 -381
rect -5516 -347 -5458 -341
rect -5516 -381 -5504 -347
rect -5470 -381 -5458 -347
rect -5516 -387 -5458 -381
rect -5398 -347 -5340 -341
rect -5398 -381 -5386 -347
rect -5352 -381 -5340 -347
rect -5398 -387 -5340 -381
rect -5280 -347 -5222 -341
rect -5280 -381 -5268 -347
rect -5234 -381 -5222 -347
rect -5280 -387 -5222 -381
rect -5162 -347 -5104 -341
rect -5162 -381 -5150 -347
rect -5116 -381 -5104 -347
rect -5162 -387 -5104 -381
rect -5044 -347 -4986 -341
rect -5044 -381 -5032 -347
rect -4998 -381 -4986 -347
rect -5044 -387 -4986 -381
rect -4926 -347 -4868 -341
rect -4926 -381 -4914 -347
rect -4880 -381 -4868 -347
rect -4926 -387 -4868 -381
rect -4808 -347 -4750 -341
rect -4808 -381 -4796 -347
rect -4762 -381 -4750 -347
rect -4808 -387 -4750 -381
rect -4690 -347 -4632 -341
rect -4690 -381 -4678 -347
rect -4644 -381 -4632 -347
rect -4690 -387 -4632 -381
rect -4572 -347 -4514 -341
rect -4572 -381 -4560 -347
rect -4526 -381 -4514 -347
rect -4572 -387 -4514 -381
rect -4454 -347 -4396 -341
rect -4454 -381 -4442 -347
rect -4408 -381 -4396 -347
rect -4454 -387 -4396 -381
rect -4336 -347 -4278 -341
rect -4336 -381 -4324 -347
rect -4290 -381 -4278 -347
rect -4336 -387 -4278 -381
rect -4218 -347 -4160 -341
rect -4218 -381 -4206 -347
rect -4172 -381 -4160 -347
rect -4218 -387 -4160 -381
rect -4100 -347 -4042 -341
rect -4100 -381 -4088 -347
rect -4054 -381 -4042 -347
rect -4100 -387 -4042 -381
rect -3982 -347 -3924 -341
rect -3982 -381 -3970 -347
rect -3936 -381 -3924 -347
rect -3982 -387 -3924 -381
rect -3864 -347 -3806 -341
rect -3864 -381 -3852 -347
rect -3818 -381 -3806 -347
rect -3864 -387 -3806 -381
rect -3746 -347 -3688 -341
rect -3746 -381 -3734 -347
rect -3700 -381 -3688 -347
rect -3746 -387 -3688 -381
rect -3628 -347 -3570 -341
rect -3628 -381 -3616 -347
rect -3582 -381 -3570 -347
rect -3628 -387 -3570 -381
rect -3510 -347 -3452 -341
rect -3510 -381 -3498 -347
rect -3464 -381 -3452 -347
rect -3510 -387 -3452 -381
rect -3392 -347 -3334 -341
rect -3392 -381 -3380 -347
rect -3346 -381 -3334 -347
rect -3392 -387 -3334 -381
rect -3274 -347 -3216 -341
rect -3274 -381 -3262 -347
rect -3228 -381 -3216 -347
rect -3274 -387 -3216 -381
rect -3156 -347 -3098 -341
rect -3156 -381 -3144 -347
rect -3110 -381 -3098 -347
rect -3156 -387 -3098 -381
rect -3038 -347 -2980 -341
rect -3038 -381 -3026 -347
rect -2992 -381 -2980 -347
rect -3038 -387 -2980 -381
rect -2920 -347 -2862 -341
rect -2920 -381 -2908 -347
rect -2874 -381 -2862 -347
rect -2920 -387 -2862 -381
rect -2802 -347 -2744 -341
rect -2802 -381 -2790 -347
rect -2756 -381 -2744 -347
rect -2802 -387 -2744 -381
rect -2684 -347 -2626 -341
rect -2684 -381 -2672 -347
rect -2638 -381 -2626 -347
rect -2684 -387 -2626 -381
rect -2566 -347 -2508 -341
rect -2566 -381 -2554 -347
rect -2520 -381 -2508 -347
rect -2566 -387 -2508 -381
rect -2448 -347 -2390 -341
rect -2448 -381 -2436 -347
rect -2402 -381 -2390 -347
rect -2448 -387 -2390 -381
rect -2330 -347 -2272 -341
rect -2330 -381 -2318 -347
rect -2284 -381 -2272 -347
rect -2330 -387 -2272 -381
rect -2212 -347 -2154 -341
rect -2212 -381 -2200 -347
rect -2166 -381 -2154 -347
rect -2212 -387 -2154 -381
rect -2094 -347 -2036 -341
rect -2094 -381 -2082 -347
rect -2048 -381 -2036 -347
rect -2094 -387 -2036 -381
rect -1976 -347 -1918 -341
rect -1976 -381 -1964 -347
rect -1930 -381 -1918 -347
rect -1976 -387 -1918 -381
rect -1858 -347 -1800 -341
rect -1858 -381 -1846 -347
rect -1812 -381 -1800 -347
rect -1858 -387 -1800 -381
rect -1740 -347 -1682 -341
rect -1740 -381 -1728 -347
rect -1694 -381 -1682 -347
rect -1740 -387 -1682 -381
rect -1622 -347 -1564 -341
rect -1622 -381 -1610 -347
rect -1576 -381 -1564 -347
rect -1622 -387 -1564 -381
rect -1504 -347 -1446 -341
rect -1504 -381 -1492 -347
rect -1458 -381 -1446 -347
rect -1504 -387 -1446 -381
rect -1386 -347 -1328 -341
rect -1386 -381 -1374 -347
rect -1340 -381 -1328 -347
rect -1386 -387 -1328 -381
rect -1268 -347 -1210 -341
rect -1268 -381 -1256 -347
rect -1222 -381 -1210 -347
rect -1268 -387 -1210 -381
rect -1150 -347 -1092 -341
rect -1150 -381 -1138 -347
rect -1104 -381 -1092 -347
rect -1150 -387 -1092 -381
rect -1032 -347 -974 -341
rect -1032 -381 -1020 -347
rect -986 -381 -974 -347
rect -1032 -387 -974 -381
rect -914 -347 -856 -341
rect -914 -381 -902 -347
rect -868 -381 -856 -347
rect -914 -387 -856 -381
rect -796 -347 -738 -341
rect -796 -381 -784 -347
rect -750 -381 -738 -347
rect -796 -387 -738 -381
rect -678 -347 -620 -341
rect -678 -381 -666 -347
rect -632 -381 -620 -347
rect -678 -387 -620 -381
rect -560 -347 -502 -341
rect -560 -381 -548 -347
rect -514 -381 -502 -347
rect -560 -387 -502 -381
rect -442 -347 -384 -341
rect -442 -381 -430 -347
rect -396 -381 -384 -347
rect -442 -387 -384 -381
rect -324 -347 -266 -341
rect -324 -381 -312 -347
rect -278 -381 -266 -347
rect -324 -387 -266 -381
rect -206 -347 -148 -341
rect -206 -381 -194 -347
rect -160 -381 -148 -347
rect -206 -387 -148 -381
rect -88 -347 -30 -341
rect -88 -381 -76 -347
rect -42 -381 -30 -347
rect -88 -387 -30 -381
rect 30 -347 88 -341
rect 30 -381 42 -347
rect 76 -381 88 -347
rect 30 -387 88 -381
rect 148 -347 206 -341
rect 148 -381 160 -347
rect 194 -381 206 -347
rect 148 -387 206 -381
rect 266 -347 324 -341
rect 266 -381 278 -347
rect 312 -381 324 -347
rect 266 -387 324 -381
rect 384 -347 442 -341
rect 384 -381 396 -347
rect 430 -381 442 -347
rect 384 -387 442 -381
rect 502 -347 560 -341
rect 502 -381 514 -347
rect 548 -381 560 -347
rect 502 -387 560 -381
rect 620 -347 678 -341
rect 620 -381 632 -347
rect 666 -381 678 -347
rect 620 -387 678 -381
rect 738 -347 796 -341
rect 738 -381 750 -347
rect 784 -381 796 -347
rect 738 -387 796 -381
rect 856 -347 914 -341
rect 856 -381 868 -347
rect 902 -381 914 -347
rect 856 -387 914 -381
rect 974 -347 1032 -341
rect 974 -381 986 -347
rect 1020 -381 1032 -347
rect 974 -387 1032 -381
rect 1092 -347 1150 -341
rect 1092 -381 1104 -347
rect 1138 -381 1150 -347
rect 1092 -387 1150 -381
rect 1210 -347 1268 -341
rect 1210 -381 1222 -347
rect 1256 -381 1268 -347
rect 1210 -387 1268 -381
rect 1328 -347 1386 -341
rect 1328 -381 1340 -347
rect 1374 -381 1386 -347
rect 1328 -387 1386 -381
rect 1446 -347 1504 -341
rect 1446 -381 1458 -347
rect 1492 -381 1504 -347
rect 1446 -387 1504 -381
rect 1564 -347 1622 -341
rect 1564 -381 1576 -347
rect 1610 -381 1622 -347
rect 1564 -387 1622 -381
rect 1682 -347 1740 -341
rect 1682 -381 1694 -347
rect 1728 -381 1740 -347
rect 1682 -387 1740 -381
rect 1800 -347 1858 -341
rect 1800 -381 1812 -347
rect 1846 -381 1858 -347
rect 1800 -387 1858 -381
rect 1918 -347 1976 -341
rect 1918 -381 1930 -347
rect 1964 -381 1976 -347
rect 1918 -387 1976 -381
rect 2036 -347 2094 -341
rect 2036 -381 2048 -347
rect 2082 -381 2094 -347
rect 2036 -387 2094 -381
rect 2154 -347 2212 -341
rect 2154 -381 2166 -347
rect 2200 -381 2212 -347
rect 2154 -387 2212 -381
rect 2272 -347 2330 -341
rect 2272 -381 2284 -347
rect 2318 -381 2330 -347
rect 2272 -387 2330 -381
rect 2390 -347 2448 -341
rect 2390 -381 2402 -347
rect 2436 -381 2448 -347
rect 2390 -387 2448 -381
rect 2508 -347 2566 -341
rect 2508 -381 2520 -347
rect 2554 -381 2566 -347
rect 2508 -387 2566 -381
rect 2626 -347 2684 -341
rect 2626 -381 2638 -347
rect 2672 -381 2684 -347
rect 2626 -387 2684 -381
rect 2744 -347 2802 -341
rect 2744 -381 2756 -347
rect 2790 -381 2802 -347
rect 2744 -387 2802 -381
rect 2862 -347 2920 -341
rect 2862 -381 2874 -347
rect 2908 -381 2920 -347
rect 2862 -387 2920 -381
rect 2980 -347 3038 -341
rect 2980 -381 2992 -347
rect 3026 -381 3038 -347
rect 2980 -387 3038 -381
rect 3098 -347 3156 -341
rect 3098 -381 3110 -347
rect 3144 -381 3156 -347
rect 3098 -387 3156 -381
rect 3216 -347 3274 -341
rect 3216 -381 3228 -347
rect 3262 -381 3274 -347
rect 3216 -387 3274 -381
rect 3334 -347 3392 -341
rect 3334 -381 3346 -347
rect 3380 -381 3392 -347
rect 3334 -387 3392 -381
rect 3452 -347 3510 -341
rect 3452 -381 3464 -347
rect 3498 -381 3510 -347
rect 3452 -387 3510 -381
rect 3570 -347 3628 -341
rect 3570 -381 3582 -347
rect 3616 -381 3628 -347
rect 3570 -387 3628 -381
rect 3688 -347 3746 -341
rect 3688 -381 3700 -347
rect 3734 -381 3746 -347
rect 3688 -387 3746 -381
rect 3806 -347 3864 -341
rect 3806 -381 3818 -347
rect 3852 -381 3864 -347
rect 3806 -387 3864 -381
rect 3924 -347 3982 -341
rect 3924 -381 3936 -347
rect 3970 -381 3982 -347
rect 3924 -387 3982 -381
rect 4042 -347 4100 -341
rect 4042 -381 4054 -347
rect 4088 -381 4100 -347
rect 4042 -387 4100 -381
rect 4160 -347 4218 -341
rect 4160 -381 4172 -347
rect 4206 -381 4218 -347
rect 4160 -387 4218 -381
rect 4278 -347 4336 -341
rect 4278 -381 4290 -347
rect 4324 -381 4336 -347
rect 4278 -387 4336 -381
rect 4396 -347 4454 -341
rect 4396 -381 4408 -347
rect 4442 -381 4454 -347
rect 4396 -387 4454 -381
rect 4514 -347 4572 -341
rect 4514 -381 4526 -347
rect 4560 -381 4572 -347
rect 4514 -387 4572 -381
rect 4632 -347 4690 -341
rect 4632 -381 4644 -347
rect 4678 -381 4690 -347
rect 4632 -387 4690 -381
rect 4750 -347 4808 -341
rect 4750 -381 4762 -347
rect 4796 -381 4808 -347
rect 4750 -387 4808 -381
rect 4868 -347 4926 -341
rect 4868 -381 4880 -347
rect 4914 -381 4926 -347
rect 4868 -387 4926 -381
rect 4986 -347 5044 -341
rect 4986 -381 4998 -347
rect 5032 -381 5044 -347
rect 4986 -387 5044 -381
rect 5104 -347 5162 -341
rect 5104 -381 5116 -347
rect 5150 -381 5162 -347
rect 5104 -387 5162 -381
rect 5222 -347 5280 -341
rect 5222 -381 5234 -347
rect 5268 -381 5280 -347
rect 5222 -387 5280 -381
rect 5340 -347 5398 -341
rect 5340 -381 5352 -347
rect 5386 -381 5398 -347
rect 5340 -387 5398 -381
rect 5458 -347 5516 -341
rect 5458 -381 5470 -347
rect 5504 -381 5516 -347
rect 5458 -387 5516 -381
rect 5576 -347 5634 -341
rect 5576 -381 5588 -347
rect 5622 -381 5634 -347
rect 5576 -387 5634 -381
rect 5694 -347 5752 -341
rect 5694 -381 5706 -347
rect 5740 -381 5752 -347
rect 5694 -387 5752 -381
rect 5812 -347 5870 -341
rect 5812 -381 5824 -347
rect 5858 -381 5870 -347
rect 5812 -387 5870 -381
rect 5930 -347 5988 -341
rect 5930 -381 5942 -347
rect 5976 -381 5988 -347
rect 5930 -387 5988 -381
rect 6048 -347 6106 -341
rect 6048 -381 6060 -347
rect 6094 -381 6106 -347
rect 6048 -387 6106 -381
rect 6166 -347 6224 -341
rect 6166 -381 6178 -347
rect 6212 -381 6224 -347
rect 6166 -387 6224 -381
rect 6284 -347 6342 -341
rect 6284 -381 6296 -347
rect 6330 -381 6342 -347
rect 6284 -387 6342 -381
rect 6402 -347 6460 -341
rect 6402 -381 6414 -347
rect 6448 -381 6460 -347
rect 6402 -387 6460 -381
rect 6520 -347 6578 -341
rect 6520 -381 6532 -347
rect 6566 -381 6578 -347
rect 6520 -387 6578 -381
rect 6638 -347 6696 -341
rect 6638 -381 6650 -347
rect 6684 -381 6696 -347
rect 6638 -387 6696 -381
rect 6756 -347 6814 -341
rect 6756 -381 6768 -347
rect 6802 -381 6814 -347
rect 6756 -387 6814 -381
rect 6874 -347 6932 -341
rect 6874 -381 6886 -347
rect 6920 -381 6932 -347
rect 6874 -387 6932 -381
rect 6992 -347 7050 -341
rect 6992 -381 7004 -347
rect 7038 -381 7050 -347
rect 6992 -387 7050 -381
rect 7110 -347 7168 -341
rect 7110 -381 7122 -347
rect 7156 -381 7168 -347
rect 7110 -387 7168 -381
rect 7228 -347 7286 -341
rect 7228 -381 7240 -347
rect 7274 -381 7286 -347
rect 7228 -387 7286 -381
rect 7346 -347 7404 -341
rect 7346 -381 7358 -347
rect 7392 -381 7404 -347
rect 7346 -387 7404 -381
rect 7464 -347 7522 -341
rect 7464 -381 7476 -347
rect 7510 -381 7522 -347
rect 7464 -387 7522 -381
rect 7582 -347 7640 -341
rect 7582 -381 7594 -347
rect 7628 -381 7640 -347
rect 7582 -387 7640 -381
rect 7700 -347 7758 -341
rect 7700 -381 7712 -347
rect 7746 -381 7758 -347
rect 7700 -387 7758 -381
rect 7818 -347 7876 -341
rect 7818 -381 7830 -347
rect 7864 -381 7876 -347
rect 7818 -387 7876 -381
rect 7936 -347 7994 -341
rect 7936 -381 7948 -347
rect 7982 -381 7994 -347
rect 7936 -387 7994 -381
rect 8054 -347 8112 -341
rect 8054 -381 8066 -347
rect 8100 -381 8112 -347
rect 8054 -387 8112 -381
rect 8172 -347 8230 -341
rect 8172 -381 8184 -347
rect 8218 -381 8230 -347
rect 8172 -387 8230 -381
rect 8290 -347 8348 -341
rect 8290 -381 8302 -347
rect 8336 -381 8348 -347
rect 8290 -387 8348 -381
rect 8408 -347 8466 -341
rect 8408 -381 8420 -347
rect 8454 -381 8466 -347
rect 8408 -387 8466 -381
rect 8526 -347 8584 -341
rect 8526 -381 8538 -347
rect 8572 -381 8584 -347
rect 8526 -387 8584 -381
rect 8644 -347 8702 -341
rect 8644 -381 8656 -347
rect 8690 -381 8702 -347
rect 8644 -387 8702 -381
rect 8762 -347 8820 -341
rect 8762 -381 8774 -347
rect 8808 -381 8820 -347
rect 8762 -387 8820 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -8964 -466 8964 466
string parameters w 3 l 0.3 m 1 nf 150 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
