VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO storage
  CLASS BLOCK ;
  FOREIGN storage ;
  ORIGIN 0.000 0.000 ;
  SIZE 460.000 BY 960.000 ;
  PIN mgmt_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 440.000 460.000 440.600 ;
    END
  END mgmt_addr[0]
  PIN mgmt_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 446.120 460.000 446.720 ;
    END
  END mgmt_addr[1]
  PIN mgmt_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 452.240 460.000 452.840 ;
    END
  END mgmt_addr[2]
  PIN mgmt_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 458.360 460.000 458.960 ;
    END
  END mgmt_addr[3]
  PIN mgmt_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 464.480 460.000 465.080 ;
    END
  END mgmt_addr[4]
  PIN mgmt_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 470.600 460.000 471.200 ;
    END
  END mgmt_addr[5]
  PIN mgmt_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 476.720 460.000 477.320 ;
    END
  END mgmt_addr[6]
  PIN mgmt_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 482.840 460.000 483.440 ;
    END
  END mgmt_addr[7]
  PIN mgmt_addr_ro[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 488.280 460.000 488.880 ;
    END
  END mgmt_addr_ro[0]
  PIN mgmt_addr_ro[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 494.400 460.000 495.000 ;
    END
  END mgmt_addr_ro[1]
  PIN mgmt_addr_ro[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 500.520 460.000 501.120 ;
    END
  END mgmt_addr_ro[2]
  PIN mgmt_addr_ro[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 506.640 460.000 507.240 ;
    END
  END mgmt_addr_ro[3]
  PIN mgmt_addr_ro[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 512.760 460.000 513.360 ;
    END
  END mgmt_addr_ro[4]
  PIN mgmt_addr_ro[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 518.880 460.000 519.480 ;
    END
  END mgmt_addr_ro[5]
  PIN mgmt_addr_ro[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 525.000 460.000 525.600 ;
    END
  END mgmt_addr_ro[6]
  PIN mgmt_addr_ro[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 531.120 460.000 531.720 ;
    END
  END mgmt_addr_ro[7]
  PIN mgmt_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 433.880 460.000 434.480 ;
    END
  END mgmt_clk
  PIN mgmt_ena[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 2.760 460.000 3.360 ;
    END
  END mgmt_ena[0]
  PIN mgmt_ena[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 731.720 460.000 732.320 ;
    END
  END mgmt_ena[1]
  PIN mgmt_ena_ro
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 8.200 460.000 8.800 ;
    END
  END mgmt_ena_ro
  PIN mgmt_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 44.920 460.000 45.520 ;
    END
  END mgmt_rdata[0]
  PIN mgmt_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 105.440 460.000 106.040 ;
    END
  END mgmt_rdata[10]
  PIN mgmt_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 111.560 460.000 112.160 ;
    END
  END mgmt_rdata[11]
  PIN mgmt_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 117.680 460.000 118.280 ;
    END
  END mgmt_rdata[12]
  PIN mgmt_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 123.800 460.000 124.400 ;
    END
  END mgmt_rdata[13]
  PIN mgmt_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 129.920 460.000 130.520 ;
    END
  END mgmt_rdata[14]
  PIN mgmt_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 136.040 460.000 136.640 ;
    END
  END mgmt_rdata[15]
  PIN mgmt_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 142.160 460.000 142.760 ;
    END
  END mgmt_rdata[16]
  PIN mgmt_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 148.280 460.000 148.880 ;
    END
  END mgmt_rdata[17]
  PIN mgmt_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 154.400 460.000 155.000 ;
    END
  END mgmt_rdata[18]
  PIN mgmt_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 160.520 460.000 161.120 ;
    END
  END mgmt_rdata[19]
  PIN mgmt_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 51.040 460.000 51.640 ;
    END
  END mgmt_rdata[1]
  PIN mgmt_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 166.640 460.000 167.240 ;
    END
  END mgmt_rdata[20]
  PIN mgmt_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 172.760 460.000 173.360 ;
    END
  END mgmt_rdata[21]
  PIN mgmt_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 178.880 460.000 179.480 ;
    END
  END mgmt_rdata[22]
  PIN mgmt_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 185.000 460.000 185.600 ;
    END
  END mgmt_rdata[23]
  PIN mgmt_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 191.120 460.000 191.720 ;
    END
  END mgmt_rdata[24]
  PIN mgmt_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 196.560 460.000 197.160 ;
    END
  END mgmt_rdata[25]
  PIN mgmt_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 202.680 460.000 203.280 ;
    END
  END mgmt_rdata[26]
  PIN mgmt_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 208.800 460.000 209.400 ;
    END
  END mgmt_rdata[27]
  PIN mgmt_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 214.920 460.000 215.520 ;
    END
  END mgmt_rdata[28]
  PIN mgmt_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 221.040 460.000 221.640 ;
    END
  END mgmt_rdata[29]
  PIN mgmt_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 57.160 460.000 57.760 ;
    END
  END mgmt_rdata[2]
  PIN mgmt_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 227.160 460.000 227.760 ;
    END
  END mgmt_rdata[30]
  PIN mgmt_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 233.280 460.000 233.880 ;
    END
  END mgmt_rdata[31]
  PIN mgmt_rdata[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 768.440 460.000 769.040 ;
    END
  END mgmt_rdata[32]
  PIN mgmt_rdata[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 773.880 460.000 774.480 ;
    END
  END mgmt_rdata[33]
  PIN mgmt_rdata[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 780.000 460.000 780.600 ;
    END
  END mgmt_rdata[34]
  PIN mgmt_rdata[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 786.120 460.000 786.720 ;
    END
  END mgmt_rdata[35]
  PIN mgmt_rdata[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 792.240 460.000 792.840 ;
    END
  END mgmt_rdata[36]
  PIN mgmt_rdata[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 798.360 460.000 798.960 ;
    END
  END mgmt_rdata[37]
  PIN mgmt_rdata[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 804.480 460.000 805.080 ;
    END
  END mgmt_rdata[38]
  PIN mgmt_rdata[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 810.600 460.000 811.200 ;
    END
  END mgmt_rdata[39]
  PIN mgmt_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 63.280 460.000 63.880 ;
    END
  END mgmt_rdata[3]
  PIN mgmt_rdata[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 816.720 460.000 817.320 ;
    END
  END mgmt_rdata[40]
  PIN mgmt_rdata[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 822.840 460.000 823.440 ;
    END
  END mgmt_rdata[41]
  PIN mgmt_rdata[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 828.960 460.000 829.560 ;
    END
  END mgmt_rdata[42]
  PIN mgmt_rdata[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 835.080 460.000 835.680 ;
    END
  END mgmt_rdata[43]
  PIN mgmt_rdata[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 841.200 460.000 841.800 ;
    END
  END mgmt_rdata[44]
  PIN mgmt_rdata[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 847.320 460.000 847.920 ;
    END
  END mgmt_rdata[45]
  PIN mgmt_rdata[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 853.440 460.000 854.040 ;
    END
  END mgmt_rdata[46]
  PIN mgmt_rdata[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 859.560 460.000 860.160 ;
    END
  END mgmt_rdata[47]
  PIN mgmt_rdata[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 865.680 460.000 866.280 ;
    END
  END mgmt_rdata[48]
  PIN mgmt_rdata[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 871.120 460.000 871.720 ;
    END
  END mgmt_rdata[49]
  PIN mgmt_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 69.400 460.000 70.000 ;
    END
  END mgmt_rdata[4]
  PIN mgmt_rdata[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 877.240 460.000 877.840 ;
    END
  END mgmt_rdata[50]
  PIN mgmt_rdata[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 883.360 460.000 883.960 ;
    END
  END mgmt_rdata[51]
  PIN mgmt_rdata[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 889.480 460.000 890.080 ;
    END
  END mgmt_rdata[52]
  PIN mgmt_rdata[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 895.600 460.000 896.200 ;
    END
  END mgmt_rdata[53]
  PIN mgmt_rdata[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 901.720 460.000 902.320 ;
    END
  END mgmt_rdata[54]
  PIN mgmt_rdata[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 907.840 460.000 908.440 ;
    END
  END mgmt_rdata[55]
  PIN mgmt_rdata[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 913.960 460.000 914.560 ;
    END
  END mgmt_rdata[56]
  PIN mgmt_rdata[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 920.080 460.000 920.680 ;
    END
  END mgmt_rdata[57]
  PIN mgmt_rdata[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 926.200 460.000 926.800 ;
    END
  END mgmt_rdata[58]
  PIN mgmt_rdata[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 932.320 460.000 932.920 ;
    END
  END mgmt_rdata[59]
  PIN mgmt_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 75.520 460.000 76.120 ;
    END
  END mgmt_rdata[5]
  PIN mgmt_rdata[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 938.440 460.000 939.040 ;
    END
  END mgmt_rdata[60]
  PIN mgmt_rdata[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 944.560 460.000 945.160 ;
    END
  END mgmt_rdata[61]
  PIN mgmt_rdata[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 950.680 460.000 951.280 ;
    END
  END mgmt_rdata[62]
  PIN mgmt_rdata[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 956.800 460.000 957.400 ;
    END
  END mgmt_rdata[63]
  PIN mgmt_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 81.640 460.000 82.240 ;
    END
  END mgmt_rdata[6]
  PIN mgmt_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 87.760 460.000 88.360 ;
    END
  END mgmt_rdata[7]
  PIN mgmt_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 93.880 460.000 94.480 ;
    END
  END mgmt_rdata[8]
  PIN mgmt_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 99.320 460.000 99.920 ;
    END
  END mgmt_rdata[9]
  PIN mgmt_rdata_ro[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 239.400 460.000 240.000 ;
    END
  END mgmt_rdata_ro[0]
  PIN mgmt_rdata_ro[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 299.920 460.000 300.520 ;
    END
  END mgmt_rdata_ro[10]
  PIN mgmt_rdata_ro[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 306.040 460.000 306.640 ;
    END
  END mgmt_rdata_ro[11]
  PIN mgmt_rdata_ro[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 312.160 460.000 312.760 ;
    END
  END mgmt_rdata_ro[12]
  PIN mgmt_rdata_ro[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 318.280 460.000 318.880 ;
    END
  END mgmt_rdata_ro[13]
  PIN mgmt_rdata_ro[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 324.400 460.000 325.000 ;
    END
  END mgmt_rdata_ro[14]
  PIN mgmt_rdata_ro[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 330.520 460.000 331.120 ;
    END
  END mgmt_rdata_ro[15]
  PIN mgmt_rdata_ro[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 336.640 460.000 337.240 ;
    END
  END mgmt_rdata_ro[16]
  PIN mgmt_rdata_ro[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 342.760 460.000 343.360 ;
    END
  END mgmt_rdata_ro[17]
  PIN mgmt_rdata_ro[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 348.880 460.000 349.480 ;
    END
  END mgmt_rdata_ro[18]
  PIN mgmt_rdata_ro[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 355.000 460.000 355.600 ;
    END
  END mgmt_rdata_ro[19]
  PIN mgmt_rdata_ro[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 245.520 460.000 246.120 ;
    END
  END mgmt_rdata_ro[1]
  PIN mgmt_rdata_ro[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 361.120 460.000 361.720 ;
    END
  END mgmt_rdata_ro[20]
  PIN mgmt_rdata_ro[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 367.240 460.000 367.840 ;
    END
  END mgmt_rdata_ro[21]
  PIN mgmt_rdata_ro[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 373.360 460.000 373.960 ;
    END
  END mgmt_rdata_ro[22]
  PIN mgmt_rdata_ro[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 379.480 460.000 380.080 ;
    END
  END mgmt_rdata_ro[23]
  PIN mgmt_rdata_ro[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 385.600 460.000 386.200 ;
    END
  END mgmt_rdata_ro[24]
  PIN mgmt_rdata_ro[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 391.040 460.000 391.640 ;
    END
  END mgmt_rdata_ro[25]
  PIN mgmt_rdata_ro[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 397.160 460.000 397.760 ;
    END
  END mgmt_rdata_ro[26]
  PIN mgmt_rdata_ro[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 403.280 460.000 403.880 ;
    END
  END mgmt_rdata_ro[27]
  PIN mgmt_rdata_ro[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 409.400 460.000 410.000 ;
    END
  END mgmt_rdata_ro[28]
  PIN mgmt_rdata_ro[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 415.520 460.000 416.120 ;
    END
  END mgmt_rdata_ro[29]
  PIN mgmt_rdata_ro[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 251.640 460.000 252.240 ;
    END
  END mgmt_rdata_ro[2]
  PIN mgmt_rdata_ro[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 421.640 460.000 422.240 ;
    END
  END mgmt_rdata_ro[30]
  PIN mgmt_rdata_ro[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 427.760 460.000 428.360 ;
    END
  END mgmt_rdata_ro[31]
  PIN mgmt_rdata_ro[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 257.760 460.000 258.360 ;
    END
  END mgmt_rdata_ro[3]
  PIN mgmt_rdata_ro[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 263.880 460.000 264.480 ;
    END
  END mgmt_rdata_ro[4]
  PIN mgmt_rdata_ro[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 270.000 460.000 270.600 ;
    END
  END mgmt_rdata_ro[5]
  PIN mgmt_rdata_ro[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 276.120 460.000 276.720 ;
    END
  END mgmt_rdata_ro[6]
  PIN mgmt_rdata_ro[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 282.240 460.000 282.840 ;
    END
  END mgmt_rdata_ro[7]
  PIN mgmt_rdata_ro[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 288.360 460.000 288.960 ;
    END
  END mgmt_rdata_ro[8]
  PIN mgmt_rdata_ro[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 293.800 460.000 294.400 ;
    END
  END mgmt_rdata_ro[9]
  PIN mgmt_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 537.240 460.000 537.840 ;
    END
  END mgmt_wdata[0]
  PIN mgmt_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 597.760 460.000 598.360 ;
    END
  END mgmt_wdata[10]
  PIN mgmt_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 603.880 460.000 604.480 ;
    END
  END mgmt_wdata[11]
  PIN mgmt_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 610.000 460.000 610.600 ;
    END
  END mgmt_wdata[12]
  PIN mgmt_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 616.120 460.000 616.720 ;
    END
  END mgmt_wdata[13]
  PIN mgmt_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 622.240 460.000 622.840 ;
    END
  END mgmt_wdata[14]
  PIN mgmt_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 628.360 460.000 628.960 ;
    END
  END mgmt_wdata[15]
  PIN mgmt_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 634.480 460.000 635.080 ;
    END
  END mgmt_wdata[16]
  PIN mgmt_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 640.600 460.000 641.200 ;
    END
  END mgmt_wdata[17]
  PIN mgmt_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 646.720 460.000 647.320 ;
    END
  END mgmt_wdata[18]
  PIN mgmt_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 652.840 460.000 653.440 ;
    END
  END mgmt_wdata[19]
  PIN mgmt_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 543.360 460.000 543.960 ;
    END
  END mgmt_wdata[1]
  PIN mgmt_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 658.960 460.000 659.560 ;
    END
  END mgmt_wdata[20]
  PIN mgmt_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 665.080 460.000 665.680 ;
    END
  END mgmt_wdata[21]
  PIN mgmt_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 671.200 460.000 671.800 ;
    END
  END mgmt_wdata[22]
  PIN mgmt_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 676.640 460.000 677.240 ;
    END
  END mgmt_wdata[23]
  PIN mgmt_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 682.760 460.000 683.360 ;
    END
  END mgmt_wdata[24]
  PIN mgmt_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 688.880 460.000 689.480 ;
    END
  END mgmt_wdata[25]
  PIN mgmt_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 695.000 460.000 695.600 ;
    END
  END mgmt_wdata[26]
  PIN mgmt_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 701.120 460.000 701.720 ;
    END
  END mgmt_wdata[27]
  PIN mgmt_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 707.240 460.000 707.840 ;
    END
  END mgmt_wdata[28]
  PIN mgmt_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 713.360 460.000 713.960 ;
    END
  END mgmt_wdata[29]
  PIN mgmt_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 549.480 460.000 550.080 ;
    END
  END mgmt_wdata[2]
  PIN mgmt_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 719.480 460.000 720.080 ;
    END
  END mgmt_wdata[30]
  PIN mgmt_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 725.600 460.000 726.200 ;
    END
  END mgmt_wdata[31]
  PIN mgmt_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 555.600 460.000 556.200 ;
    END
  END mgmt_wdata[3]
  PIN mgmt_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 561.720 460.000 562.320 ;
    END
  END mgmt_wdata[4]
  PIN mgmt_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 567.840 460.000 568.440 ;
    END
  END mgmt_wdata[5]
  PIN mgmt_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 573.960 460.000 574.560 ;
    END
  END mgmt_wdata[6]
  PIN mgmt_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 579.400 460.000 580.000 ;
    END
  END mgmt_wdata[7]
  PIN mgmt_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 585.520 460.000 586.120 ;
    END
  END mgmt_wdata[8]
  PIN mgmt_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 591.640 460.000 592.240 ;
    END
  END mgmt_wdata[9]
  PIN mgmt_wen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 14.320 460.000 14.920 ;
    END
  END mgmt_wen[0]
  PIN mgmt_wen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 737.840 460.000 738.440 ;
    END
  END mgmt_wen[1]
  PIN mgmt_wen_mask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 20.440 460.000 21.040 ;
    END
  END mgmt_wen_mask[0]
  PIN mgmt_wen_mask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 26.560 460.000 27.160 ;
    END
  END mgmt_wen_mask[1]
  PIN mgmt_wen_mask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 32.680 460.000 33.280 ;
    END
  END mgmt_wen_mask[2]
  PIN mgmt_wen_mask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 38.800 460.000 39.400 ;
    END
  END mgmt_wen_mask[3]
  PIN mgmt_wen_mask[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 743.960 460.000 744.560 ;
    END
  END mgmt_wen_mask[4]
  PIN mgmt_wen_mask[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 750.080 460.000 750.680 ;
    END
  END mgmt_wen_mask[5]
  PIN mgmt_wen_mask[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 756.200 460.000 756.800 ;
    END
  END mgmt_wen_mask[6]
  PIN mgmt_wen_mask[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 456.000 762.320 460.000 762.920 ;
    END
  END mgmt_wen_mask[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 449.720 10.640 451.320 946.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 429.720 10.640 431.320 946.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 946.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 926.490 454.480 928.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 876.490 454.480 878.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 826.490 454.480 828.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 776.490 454.480 778.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 726.490 454.480 728.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 676.490 454.480 678.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 626.490 454.480 628.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 576.490 454.480 578.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 526.490 454.480 528.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 476.490 454.480 478.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 426.490 454.480 428.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 376.490 454.480 378.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 326.490 454.480 328.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 276.490 454.480 278.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 226.490 454.480 228.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 176.490 454.480 178.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 126.490 454.480 128.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 76.490 454.480 78.090 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 454.480 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 439.720 10.640 441.320 946.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 19.720 10.640 21.320 946.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 901.490 454.480 903.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 851.490 454.480 853.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 801.490 454.480 803.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 751.490 454.480 753.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 701.490 454.480 703.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 651.490 454.480 653.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 601.490 454.480 603.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 551.490 454.480 553.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 501.490 454.480 503.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 451.490 454.480 453.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 401.490 454.480 403.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 351.490 454.480 353.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 301.490 454.480 303.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 251.490 454.480 253.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 201.490 454.480 203.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 151.490 454.480 153.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 101.490 454.480 103.090 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 51.490 454.480 53.090 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 5.330 945.145 25.950 946.750 ;
        RECT 5.330 939.705 25.950 942.535 ;
        RECT 5.330 934.265 25.950 937.095 ;
        RECT 5.330 928.825 25.950 931.655 ;
        RECT 5.330 923.385 25.950 926.215 ;
        RECT 5.330 917.945 25.950 920.775 ;
        RECT 5.330 912.505 25.950 915.335 ;
        RECT 5.330 907.065 25.950 909.895 ;
        RECT 5.330 901.625 25.950 904.455 ;
        RECT 5.330 896.185 25.950 899.015 ;
        RECT 5.330 890.745 25.950 893.575 ;
        RECT 5.330 885.305 25.950 888.135 ;
        RECT 5.330 879.865 25.950 882.695 ;
        RECT 5.330 874.425 25.950 877.255 ;
        RECT 5.330 868.985 25.950 871.815 ;
        RECT 5.330 863.545 25.950 866.375 ;
        RECT 5.330 858.105 25.950 860.935 ;
        RECT 5.330 852.665 25.950 855.495 ;
        RECT 5.330 847.225 25.950 850.055 ;
        RECT 5.330 841.785 25.950 844.615 ;
        RECT 5.330 836.345 25.950 839.175 ;
        RECT 5.330 830.905 25.950 833.735 ;
        RECT 5.330 825.465 25.950 828.295 ;
        RECT 5.330 820.025 25.950 822.855 ;
        RECT 5.330 814.585 25.950 817.415 ;
        RECT 5.330 809.145 25.950 811.975 ;
        RECT 5.330 803.705 25.950 806.535 ;
        RECT 5.330 798.265 25.950 801.095 ;
        RECT 5.330 792.825 25.950 795.655 ;
        RECT 5.330 787.385 25.950 790.215 ;
        RECT 5.330 781.945 25.950 784.775 ;
        RECT 5.330 776.505 25.950 779.335 ;
        RECT 5.330 771.065 25.950 773.895 ;
        RECT 5.330 765.625 25.950 768.455 ;
        RECT 5.330 760.185 25.950 763.015 ;
        RECT 5.330 754.745 25.950 757.575 ;
        RECT 5.330 749.305 25.950 752.135 ;
        RECT 5.330 743.865 25.950 746.695 ;
        RECT 5.330 738.425 25.950 741.255 ;
        RECT 5.330 732.985 25.950 735.815 ;
        RECT 5.330 727.545 25.950 730.375 ;
        RECT 5.330 722.105 25.950 724.935 ;
        RECT 5.330 716.665 25.950 719.495 ;
        RECT 5.330 711.225 25.950 714.055 ;
        RECT 5.330 705.785 25.950 708.615 ;
        RECT 5.330 700.345 25.950 703.175 ;
        RECT 5.330 694.905 25.950 697.735 ;
        RECT 5.330 689.465 25.950 692.295 ;
        RECT 5.330 684.025 25.950 686.855 ;
        RECT 5.330 678.585 25.950 681.415 ;
        RECT 5.330 673.145 25.950 675.975 ;
        RECT 5.330 667.705 25.950 670.535 ;
        RECT 5.330 662.265 25.950 665.095 ;
        RECT 5.330 656.825 25.950 659.655 ;
        RECT 5.330 651.385 25.950 654.215 ;
        RECT 5.330 645.945 25.950 648.775 ;
        RECT 5.330 640.505 25.950 643.335 ;
        RECT 5.330 635.065 25.950 637.895 ;
        RECT 5.330 629.625 25.950 632.455 ;
        RECT 5.330 624.185 25.950 627.015 ;
        RECT 5.330 618.745 25.950 621.575 ;
        RECT 5.330 613.305 25.950 616.135 ;
        RECT 5.330 607.865 25.950 610.695 ;
        RECT 5.330 602.425 25.950 605.255 ;
        RECT 5.330 596.985 25.950 599.815 ;
        RECT 5.330 591.545 25.950 594.375 ;
        RECT 5.330 586.105 25.950 588.935 ;
        RECT 5.330 580.665 25.950 583.495 ;
        RECT 5.330 575.225 25.950 578.055 ;
        RECT 5.330 569.785 25.950 572.615 ;
        RECT 5.330 564.345 25.950 567.175 ;
        RECT 5.330 558.905 25.950 561.735 ;
        RECT 5.330 553.465 25.950 556.295 ;
        RECT 5.330 548.025 25.950 550.855 ;
        RECT 5.330 542.585 25.950 545.415 ;
        RECT 5.330 537.145 25.950 539.975 ;
        RECT 5.330 531.705 25.950 534.535 ;
        RECT 5.330 526.265 25.950 529.095 ;
        RECT 5.330 520.825 25.950 523.655 ;
        RECT 5.330 515.385 25.950 518.215 ;
        RECT 5.330 509.945 25.950 512.775 ;
        RECT 5.330 504.505 25.950 507.335 ;
        RECT 5.330 499.065 25.950 501.895 ;
        RECT 5.330 493.625 25.950 496.455 ;
        RECT 5.330 488.185 25.950 491.015 ;
        RECT 5.330 482.745 25.950 485.575 ;
        RECT 5.330 477.305 25.950 480.135 ;
        RECT 5.330 471.865 25.950 474.695 ;
        RECT 5.330 466.425 25.950 469.255 ;
        RECT 5.330 460.985 25.950 463.815 ;
        RECT 5.330 455.545 25.950 458.375 ;
        RECT 5.330 450.105 25.950 452.935 ;
        RECT 5.330 444.665 25.950 447.495 ;
        RECT 5.330 439.225 25.950 442.055 ;
        RECT 5.330 433.785 25.950 436.615 ;
        RECT 5.330 428.345 25.950 431.175 ;
        RECT 5.330 422.905 25.950 425.735 ;
        RECT 5.330 417.465 25.950 420.295 ;
        RECT 5.330 412.025 25.950 414.855 ;
        RECT 5.330 406.585 25.950 409.415 ;
        RECT 5.330 401.145 25.950 403.975 ;
        RECT 5.330 395.705 25.950 398.535 ;
        RECT 5.330 390.265 25.950 393.095 ;
        RECT 5.330 384.825 25.950 387.655 ;
        RECT 5.330 379.385 25.950 382.215 ;
        RECT 5.330 373.945 25.950 376.775 ;
        RECT 5.330 368.505 25.950 371.335 ;
        RECT 5.330 363.065 25.950 365.895 ;
        RECT 5.330 357.625 25.950 360.455 ;
        RECT 5.330 352.185 25.950 355.015 ;
        RECT 5.330 346.745 25.950 349.575 ;
        RECT 5.330 341.305 25.950 344.135 ;
        RECT 5.330 335.865 25.950 338.695 ;
        RECT 5.330 330.425 25.950 333.255 ;
        RECT 5.330 324.985 25.950 327.815 ;
        RECT 5.330 319.545 25.950 322.375 ;
        RECT 5.330 314.105 25.950 316.935 ;
        RECT 5.330 308.665 25.950 311.495 ;
        RECT 5.330 303.225 25.950 306.055 ;
        RECT 5.330 297.785 25.950 300.615 ;
        RECT 5.330 292.345 25.950 295.175 ;
        RECT 5.330 286.905 25.950 289.735 ;
        RECT 5.330 281.465 25.950 284.295 ;
        RECT 5.330 276.025 25.950 278.855 ;
        RECT 5.330 270.585 25.950 273.415 ;
        RECT 5.330 265.145 25.950 267.975 ;
        RECT 5.330 259.705 25.950 262.535 ;
        RECT 5.330 254.265 25.950 257.095 ;
        RECT 5.330 248.825 25.950 251.655 ;
        RECT 5.330 243.385 25.950 246.215 ;
        RECT 5.330 237.945 25.950 240.775 ;
        RECT 5.330 232.505 25.950 235.335 ;
        RECT 5.330 227.065 25.950 229.895 ;
        RECT 5.330 221.625 25.950 224.455 ;
        RECT 5.330 216.185 25.950 219.015 ;
        RECT 5.330 210.745 25.950 213.575 ;
        RECT 5.330 205.305 25.950 208.135 ;
        RECT 5.330 199.865 25.950 202.695 ;
        RECT 5.330 194.425 25.950 197.255 ;
        RECT 5.330 188.985 25.950 191.815 ;
        RECT 5.330 183.545 25.950 186.375 ;
        RECT 5.330 178.105 25.950 180.935 ;
        RECT 5.330 172.665 25.950 175.495 ;
        RECT 5.330 167.225 25.950 170.055 ;
        RECT 5.330 161.785 25.950 164.615 ;
        RECT 5.330 156.345 25.950 159.175 ;
        RECT 5.330 150.905 25.950 153.735 ;
        RECT 5.330 145.465 25.950 148.295 ;
        RECT 5.330 140.025 25.950 142.855 ;
        RECT 5.330 134.585 25.950 137.415 ;
        RECT 5.330 129.145 25.950 131.975 ;
        RECT 5.330 123.705 25.950 126.535 ;
        RECT 5.330 118.265 25.950 121.095 ;
        RECT 5.330 112.825 25.950 115.655 ;
        RECT 5.330 107.385 25.950 110.215 ;
        RECT 5.330 101.945 25.950 104.775 ;
        RECT 5.330 96.505 25.950 99.335 ;
        RECT 5.330 91.065 25.950 93.895 ;
        RECT 5.330 85.625 25.950 88.455 ;
        RECT 5.330 80.185 25.950 83.015 ;
        RECT 5.330 74.745 25.950 77.575 ;
        RECT 5.330 69.305 25.950 72.135 ;
        RECT 5.330 63.865 25.950 66.695 ;
        RECT 5.330 58.425 25.950 61.255 ;
        RECT 5.330 52.985 25.950 55.815 ;
        RECT 5.330 47.545 25.950 50.375 ;
        RECT 5.330 42.105 25.950 44.935 ;
        RECT 5.330 36.665 25.950 39.495 ;
        RECT 5.330 31.225 25.950 34.055 ;
        RECT 5.330 25.785 25.950 28.615 ;
        RECT 5.330 20.345 25.950 23.175 ;
        RECT 5.330 14.905 25.950 17.735 ;
        RECT 5.330 10.690 25.950 12.295 ;
      LAYER li1 ;
        RECT 5.520 6.205 454.480 946.645 ;
      LAYER met1 ;
        RECT 5.520 0.720 454.480 946.800 ;
      LAYER met2 ;
        RECT 9.780 0.690 451.260 951.165 ;
      LAYER met3 ;
        RECT 9.720 956.400 455.600 957.260 ;
        RECT 9.720 951.680 456.000 956.400 ;
        RECT 9.720 950.280 455.600 951.680 ;
        RECT 9.720 945.560 456.000 950.280 ;
        RECT 9.720 944.160 455.600 945.560 ;
        RECT 9.720 939.440 456.000 944.160 ;
        RECT 9.720 938.040 455.600 939.440 ;
        RECT 9.720 933.320 456.000 938.040 ;
        RECT 9.720 931.920 455.600 933.320 ;
        RECT 9.720 927.200 456.000 931.920 ;
        RECT 9.720 925.800 455.600 927.200 ;
        RECT 9.720 921.080 456.000 925.800 ;
        RECT 9.720 919.680 455.600 921.080 ;
        RECT 9.720 914.960 456.000 919.680 ;
        RECT 9.720 913.560 455.600 914.960 ;
        RECT 9.720 908.840 456.000 913.560 ;
        RECT 9.720 907.440 455.600 908.840 ;
        RECT 9.720 902.720 456.000 907.440 ;
        RECT 9.720 901.320 455.600 902.720 ;
        RECT 9.720 896.600 456.000 901.320 ;
        RECT 9.720 895.200 455.600 896.600 ;
        RECT 9.720 890.480 456.000 895.200 ;
        RECT 9.720 889.080 455.600 890.480 ;
        RECT 9.720 884.360 456.000 889.080 ;
        RECT 9.720 882.960 455.600 884.360 ;
        RECT 9.720 878.240 456.000 882.960 ;
        RECT 9.720 876.840 455.600 878.240 ;
        RECT 9.720 872.120 456.000 876.840 ;
        RECT 9.720 870.720 455.600 872.120 ;
        RECT 9.720 866.680 456.000 870.720 ;
        RECT 9.720 865.280 455.600 866.680 ;
        RECT 9.720 860.560 456.000 865.280 ;
        RECT 9.720 859.160 455.600 860.560 ;
        RECT 9.720 854.440 456.000 859.160 ;
        RECT 9.720 853.040 455.600 854.440 ;
        RECT 9.720 848.320 456.000 853.040 ;
        RECT 9.720 846.920 455.600 848.320 ;
        RECT 9.720 842.200 456.000 846.920 ;
        RECT 9.720 840.800 455.600 842.200 ;
        RECT 9.720 836.080 456.000 840.800 ;
        RECT 9.720 834.680 455.600 836.080 ;
        RECT 9.720 829.960 456.000 834.680 ;
        RECT 9.720 828.560 455.600 829.960 ;
        RECT 9.720 823.840 456.000 828.560 ;
        RECT 9.720 822.440 455.600 823.840 ;
        RECT 9.720 817.720 456.000 822.440 ;
        RECT 9.720 816.320 455.600 817.720 ;
        RECT 9.720 811.600 456.000 816.320 ;
        RECT 9.720 810.200 455.600 811.600 ;
        RECT 9.720 805.480 456.000 810.200 ;
        RECT 9.720 804.080 455.600 805.480 ;
        RECT 9.720 799.360 456.000 804.080 ;
        RECT 9.720 797.960 455.600 799.360 ;
        RECT 9.720 793.240 456.000 797.960 ;
        RECT 9.720 791.840 455.600 793.240 ;
        RECT 9.720 787.120 456.000 791.840 ;
        RECT 9.720 785.720 455.600 787.120 ;
        RECT 9.720 781.000 456.000 785.720 ;
        RECT 9.720 779.600 455.600 781.000 ;
        RECT 9.720 774.880 456.000 779.600 ;
        RECT 9.720 773.480 455.600 774.880 ;
        RECT 9.720 769.440 456.000 773.480 ;
        RECT 9.720 768.040 455.600 769.440 ;
        RECT 9.720 763.320 456.000 768.040 ;
        RECT 9.720 761.920 455.600 763.320 ;
        RECT 9.720 757.200 456.000 761.920 ;
        RECT 9.720 755.800 455.600 757.200 ;
        RECT 9.720 751.080 456.000 755.800 ;
        RECT 9.720 749.680 455.600 751.080 ;
        RECT 9.720 744.960 456.000 749.680 ;
        RECT 9.720 743.560 455.600 744.960 ;
        RECT 9.720 738.840 456.000 743.560 ;
        RECT 9.720 737.440 455.600 738.840 ;
        RECT 9.720 732.720 456.000 737.440 ;
        RECT 9.720 731.320 455.600 732.720 ;
        RECT 9.720 726.600 456.000 731.320 ;
        RECT 9.720 725.200 455.600 726.600 ;
        RECT 9.720 720.480 456.000 725.200 ;
        RECT 9.720 719.080 455.600 720.480 ;
        RECT 9.720 714.360 456.000 719.080 ;
        RECT 9.720 712.960 455.600 714.360 ;
        RECT 9.720 708.240 456.000 712.960 ;
        RECT 9.720 706.840 455.600 708.240 ;
        RECT 9.720 702.120 456.000 706.840 ;
        RECT 9.720 700.720 455.600 702.120 ;
        RECT 9.720 696.000 456.000 700.720 ;
        RECT 9.720 694.600 455.600 696.000 ;
        RECT 9.720 689.880 456.000 694.600 ;
        RECT 9.720 688.480 455.600 689.880 ;
        RECT 9.720 683.760 456.000 688.480 ;
        RECT 9.720 682.360 455.600 683.760 ;
        RECT 9.720 677.640 456.000 682.360 ;
        RECT 9.720 676.240 455.600 677.640 ;
        RECT 9.720 672.200 456.000 676.240 ;
        RECT 9.720 670.800 455.600 672.200 ;
        RECT 9.720 666.080 456.000 670.800 ;
        RECT 9.720 664.680 455.600 666.080 ;
        RECT 9.720 659.960 456.000 664.680 ;
        RECT 9.720 658.560 455.600 659.960 ;
        RECT 9.720 653.840 456.000 658.560 ;
        RECT 9.720 652.440 455.600 653.840 ;
        RECT 9.720 647.720 456.000 652.440 ;
        RECT 9.720 646.320 455.600 647.720 ;
        RECT 9.720 641.600 456.000 646.320 ;
        RECT 9.720 640.200 455.600 641.600 ;
        RECT 9.720 635.480 456.000 640.200 ;
        RECT 9.720 634.080 455.600 635.480 ;
        RECT 9.720 629.360 456.000 634.080 ;
        RECT 9.720 627.960 455.600 629.360 ;
        RECT 9.720 623.240 456.000 627.960 ;
        RECT 9.720 621.840 455.600 623.240 ;
        RECT 9.720 617.120 456.000 621.840 ;
        RECT 9.720 615.720 455.600 617.120 ;
        RECT 9.720 611.000 456.000 615.720 ;
        RECT 9.720 609.600 455.600 611.000 ;
        RECT 9.720 604.880 456.000 609.600 ;
        RECT 9.720 603.480 455.600 604.880 ;
        RECT 9.720 598.760 456.000 603.480 ;
        RECT 9.720 597.360 455.600 598.760 ;
        RECT 9.720 592.640 456.000 597.360 ;
        RECT 9.720 591.240 455.600 592.640 ;
        RECT 9.720 586.520 456.000 591.240 ;
        RECT 9.720 585.120 455.600 586.520 ;
        RECT 9.720 580.400 456.000 585.120 ;
        RECT 9.720 579.000 455.600 580.400 ;
        RECT 9.720 574.960 456.000 579.000 ;
        RECT 9.720 573.560 455.600 574.960 ;
        RECT 9.720 568.840 456.000 573.560 ;
        RECT 9.720 567.440 455.600 568.840 ;
        RECT 9.720 562.720 456.000 567.440 ;
        RECT 9.720 561.320 455.600 562.720 ;
        RECT 9.720 556.600 456.000 561.320 ;
        RECT 9.720 555.200 455.600 556.600 ;
        RECT 9.720 550.480 456.000 555.200 ;
        RECT 9.720 549.080 455.600 550.480 ;
        RECT 9.720 544.360 456.000 549.080 ;
        RECT 9.720 542.960 455.600 544.360 ;
        RECT 9.720 538.240 456.000 542.960 ;
        RECT 9.720 536.840 455.600 538.240 ;
        RECT 9.720 532.120 456.000 536.840 ;
        RECT 9.720 530.720 455.600 532.120 ;
        RECT 9.720 526.000 456.000 530.720 ;
        RECT 9.720 524.600 455.600 526.000 ;
        RECT 9.720 519.880 456.000 524.600 ;
        RECT 9.720 518.480 455.600 519.880 ;
        RECT 9.720 513.760 456.000 518.480 ;
        RECT 9.720 512.360 455.600 513.760 ;
        RECT 9.720 507.640 456.000 512.360 ;
        RECT 9.720 506.240 455.600 507.640 ;
        RECT 9.720 501.520 456.000 506.240 ;
        RECT 9.720 500.120 455.600 501.520 ;
        RECT 9.720 495.400 456.000 500.120 ;
        RECT 9.720 494.000 455.600 495.400 ;
        RECT 9.720 489.280 456.000 494.000 ;
        RECT 9.720 487.880 455.600 489.280 ;
        RECT 9.720 483.840 456.000 487.880 ;
        RECT 9.720 482.440 455.600 483.840 ;
        RECT 9.720 477.720 456.000 482.440 ;
        RECT 9.720 476.320 455.600 477.720 ;
        RECT 9.720 471.600 456.000 476.320 ;
        RECT 9.720 470.200 455.600 471.600 ;
        RECT 9.720 465.480 456.000 470.200 ;
        RECT 9.720 464.080 455.600 465.480 ;
        RECT 9.720 459.360 456.000 464.080 ;
        RECT 9.720 457.960 455.600 459.360 ;
        RECT 9.720 453.240 456.000 457.960 ;
        RECT 9.720 451.840 455.600 453.240 ;
        RECT 9.720 447.120 456.000 451.840 ;
        RECT 9.720 445.720 455.600 447.120 ;
        RECT 9.720 441.000 456.000 445.720 ;
        RECT 9.720 439.600 455.600 441.000 ;
        RECT 9.720 434.880 456.000 439.600 ;
        RECT 9.720 433.480 455.600 434.880 ;
        RECT 9.720 428.760 456.000 433.480 ;
        RECT 9.720 427.360 455.600 428.760 ;
        RECT 9.720 422.640 456.000 427.360 ;
        RECT 9.720 421.240 455.600 422.640 ;
        RECT 9.720 416.520 456.000 421.240 ;
        RECT 9.720 415.120 455.600 416.520 ;
        RECT 9.720 410.400 456.000 415.120 ;
        RECT 9.720 409.000 455.600 410.400 ;
        RECT 9.720 404.280 456.000 409.000 ;
        RECT 9.720 402.880 455.600 404.280 ;
        RECT 9.720 398.160 456.000 402.880 ;
        RECT 9.720 396.760 455.600 398.160 ;
        RECT 9.720 392.040 456.000 396.760 ;
        RECT 9.720 390.640 455.600 392.040 ;
        RECT 9.720 386.600 456.000 390.640 ;
        RECT 9.720 385.200 455.600 386.600 ;
        RECT 9.720 380.480 456.000 385.200 ;
        RECT 9.720 379.080 455.600 380.480 ;
        RECT 9.720 374.360 456.000 379.080 ;
        RECT 9.720 372.960 455.600 374.360 ;
        RECT 9.720 368.240 456.000 372.960 ;
        RECT 9.720 366.840 455.600 368.240 ;
        RECT 9.720 362.120 456.000 366.840 ;
        RECT 9.720 360.720 455.600 362.120 ;
        RECT 9.720 356.000 456.000 360.720 ;
        RECT 9.720 354.600 455.600 356.000 ;
        RECT 9.720 349.880 456.000 354.600 ;
        RECT 9.720 348.480 455.600 349.880 ;
        RECT 9.720 343.760 456.000 348.480 ;
        RECT 9.720 342.360 455.600 343.760 ;
        RECT 9.720 337.640 456.000 342.360 ;
        RECT 9.720 336.240 455.600 337.640 ;
        RECT 9.720 331.520 456.000 336.240 ;
        RECT 9.720 330.120 455.600 331.520 ;
        RECT 9.720 325.400 456.000 330.120 ;
        RECT 9.720 324.000 455.600 325.400 ;
        RECT 9.720 319.280 456.000 324.000 ;
        RECT 9.720 317.880 455.600 319.280 ;
        RECT 9.720 313.160 456.000 317.880 ;
        RECT 9.720 311.760 455.600 313.160 ;
        RECT 9.720 307.040 456.000 311.760 ;
        RECT 9.720 305.640 455.600 307.040 ;
        RECT 9.720 300.920 456.000 305.640 ;
        RECT 9.720 299.520 455.600 300.920 ;
        RECT 9.720 294.800 456.000 299.520 ;
        RECT 9.720 293.400 455.600 294.800 ;
        RECT 9.720 289.360 456.000 293.400 ;
        RECT 9.720 287.960 455.600 289.360 ;
        RECT 9.720 283.240 456.000 287.960 ;
        RECT 9.720 281.840 455.600 283.240 ;
        RECT 9.720 277.120 456.000 281.840 ;
        RECT 9.720 275.720 455.600 277.120 ;
        RECT 9.720 271.000 456.000 275.720 ;
        RECT 9.720 269.600 455.600 271.000 ;
        RECT 9.720 264.880 456.000 269.600 ;
        RECT 9.720 263.480 455.600 264.880 ;
        RECT 9.720 258.760 456.000 263.480 ;
        RECT 9.720 257.360 455.600 258.760 ;
        RECT 9.720 252.640 456.000 257.360 ;
        RECT 9.720 251.240 455.600 252.640 ;
        RECT 9.720 246.520 456.000 251.240 ;
        RECT 9.720 245.120 455.600 246.520 ;
        RECT 9.720 240.400 456.000 245.120 ;
        RECT 9.720 239.000 455.600 240.400 ;
        RECT 9.720 234.280 456.000 239.000 ;
        RECT 9.720 232.880 455.600 234.280 ;
        RECT 9.720 228.160 456.000 232.880 ;
        RECT 9.720 226.760 455.600 228.160 ;
        RECT 9.720 222.040 456.000 226.760 ;
        RECT 9.720 220.640 455.600 222.040 ;
        RECT 9.720 215.920 456.000 220.640 ;
        RECT 9.720 214.520 455.600 215.920 ;
        RECT 9.720 209.800 456.000 214.520 ;
        RECT 9.720 208.400 455.600 209.800 ;
        RECT 9.720 203.680 456.000 208.400 ;
        RECT 9.720 202.280 455.600 203.680 ;
        RECT 9.720 197.560 456.000 202.280 ;
        RECT 9.720 196.160 455.600 197.560 ;
        RECT 9.720 192.120 456.000 196.160 ;
        RECT 9.720 190.720 455.600 192.120 ;
        RECT 9.720 186.000 456.000 190.720 ;
        RECT 9.720 184.600 455.600 186.000 ;
        RECT 9.720 179.880 456.000 184.600 ;
        RECT 9.720 178.480 455.600 179.880 ;
        RECT 9.720 173.760 456.000 178.480 ;
        RECT 9.720 172.360 455.600 173.760 ;
        RECT 9.720 167.640 456.000 172.360 ;
        RECT 9.720 166.240 455.600 167.640 ;
        RECT 9.720 161.520 456.000 166.240 ;
        RECT 9.720 160.120 455.600 161.520 ;
        RECT 9.720 155.400 456.000 160.120 ;
        RECT 9.720 154.000 455.600 155.400 ;
        RECT 9.720 149.280 456.000 154.000 ;
        RECT 9.720 147.880 455.600 149.280 ;
        RECT 9.720 143.160 456.000 147.880 ;
        RECT 9.720 141.760 455.600 143.160 ;
        RECT 9.720 137.040 456.000 141.760 ;
        RECT 9.720 135.640 455.600 137.040 ;
        RECT 9.720 130.920 456.000 135.640 ;
        RECT 9.720 129.520 455.600 130.920 ;
        RECT 9.720 124.800 456.000 129.520 ;
        RECT 9.720 123.400 455.600 124.800 ;
        RECT 9.720 118.680 456.000 123.400 ;
        RECT 9.720 117.280 455.600 118.680 ;
        RECT 9.720 112.560 456.000 117.280 ;
        RECT 9.720 111.160 455.600 112.560 ;
        RECT 9.720 106.440 456.000 111.160 ;
        RECT 9.720 105.040 455.600 106.440 ;
        RECT 9.720 100.320 456.000 105.040 ;
        RECT 9.720 98.920 455.600 100.320 ;
        RECT 9.720 94.880 456.000 98.920 ;
        RECT 9.720 93.480 455.600 94.880 ;
        RECT 9.720 88.760 456.000 93.480 ;
        RECT 9.720 87.360 455.600 88.760 ;
        RECT 9.720 82.640 456.000 87.360 ;
        RECT 9.720 81.240 455.600 82.640 ;
        RECT 9.720 76.520 456.000 81.240 ;
        RECT 9.720 75.120 455.600 76.520 ;
        RECT 9.720 70.400 456.000 75.120 ;
        RECT 9.720 69.000 455.600 70.400 ;
        RECT 9.720 64.280 456.000 69.000 ;
        RECT 9.720 62.880 455.600 64.280 ;
        RECT 9.720 58.160 456.000 62.880 ;
        RECT 9.720 56.760 455.600 58.160 ;
        RECT 9.720 52.040 456.000 56.760 ;
        RECT 9.720 50.640 455.600 52.040 ;
        RECT 9.720 45.920 456.000 50.640 ;
        RECT 9.720 44.520 455.600 45.920 ;
        RECT 9.720 39.800 456.000 44.520 ;
        RECT 9.720 38.400 455.600 39.800 ;
        RECT 9.720 33.680 456.000 38.400 ;
        RECT 9.720 32.280 455.600 33.680 ;
        RECT 9.720 27.560 456.000 32.280 ;
        RECT 9.720 26.160 455.600 27.560 ;
        RECT 9.720 21.440 456.000 26.160 ;
        RECT 9.720 20.040 455.600 21.440 ;
        RECT 9.720 15.320 456.000 20.040 ;
        RECT 9.720 13.920 455.600 15.320 ;
        RECT 9.720 9.200 456.000 13.920 ;
        RECT 9.720 7.800 455.600 9.200 ;
        RECT 9.720 3.760 456.000 7.800 ;
        RECT 9.720 2.360 455.600 3.760 ;
        RECT 9.720 0.855 456.000 2.360 ;
      LAYER met4 ;
        RECT 21.950 947.200 438.970 957.265 ;
        RECT 21.950 10.240 429.320 947.200 ;
        RECT 431.720 10.240 438.970 947.200 ;
        RECT 21.950 0.855 438.970 10.240 ;
      LAYER met5 ;
        RECT 21.740 479.690 439.180 488.700 ;
        RECT 21.740 454.690 439.180 474.890 ;
        RECT 21.740 429.690 439.180 449.890 ;
        RECT 21.740 404.690 439.180 424.890 ;
        RECT 21.740 379.690 439.180 399.890 ;
        RECT 21.740 354.690 439.180 374.890 ;
        RECT 21.740 329.690 439.180 349.890 ;
        RECT 21.740 304.690 439.180 324.890 ;
        RECT 21.740 279.690 439.180 299.890 ;
        RECT 21.740 254.690 439.180 274.890 ;
        RECT 21.740 229.690 439.180 249.890 ;
        RECT 21.740 204.690 439.180 224.890 ;
        RECT 21.740 179.690 439.180 199.890 ;
        RECT 21.740 154.690 439.180 174.890 ;
        RECT 21.740 129.690 439.180 149.890 ;
        RECT 21.740 104.690 439.180 124.890 ;
        RECT 21.740 79.690 439.180 99.890 ;
        RECT 21.740 54.690 439.180 74.890 ;
        RECT 21.740 29.690 439.180 49.890 ;
        RECT 21.740 14.500 439.180 24.890 ;
  END
END storage
END LIBRARY

