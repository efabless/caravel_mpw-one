magic
tech sky130A
magscale 1 2
timestamp 1625001917
<< metal1 >>
rect 261328 1006411 261334 1006463
rect 261386 1006451 261392 1006463
rect 276592 1006451 276598 1006463
rect 261386 1006423 276598 1006451
rect 261386 1006411 261392 1006423
rect 276592 1006411 276598 1006423
rect 276650 1006411 276656 1006463
rect 92848 1006115 92854 1006167
rect 92906 1006155 92912 1006167
rect 102448 1006155 102454 1006167
rect 92906 1006127 102454 1006155
rect 92906 1006115 92912 1006127
rect 102448 1006115 102454 1006127
rect 102506 1006115 102512 1006167
rect 356368 1006041 356374 1006093
rect 356426 1006081 356432 1006093
rect 371632 1006081 371638 1006093
rect 356426 1006053 371638 1006081
rect 356426 1006041 356432 1006053
rect 371632 1006041 371638 1006053
rect 371690 1006041 371696 1006093
rect 558160 1006041 558166 1006093
rect 558218 1006081 558224 1006093
rect 574672 1006081 574678 1006093
rect 558218 1006053 574678 1006081
rect 558218 1006041 558224 1006053
rect 574672 1006041 574678 1006053
rect 574730 1006041 574736 1006093
rect 357904 1005967 357910 1006019
rect 357962 1006007 357968 1006019
rect 377296 1006007 377302 1006019
rect 357962 1005979 377302 1006007
rect 357962 1005967 357968 1005979
rect 377296 1005967 377302 1005979
rect 377354 1005967 377360 1006019
rect 358768 1005893 358774 1005945
rect 358826 1005933 358832 1005945
rect 378832 1005933 378838 1005945
rect 358826 1005905 378838 1005933
rect 358826 1005893 358832 1005905
rect 378832 1005893 378838 1005905
rect 378890 1005893 378896 1005945
rect 425680 1005893 425686 1005945
rect 425738 1005933 425744 1005945
rect 471664 1005933 471670 1005945
rect 425738 1005905 471670 1005933
rect 425738 1005893 425744 1005905
rect 471664 1005893 471670 1005905
rect 471722 1005893 471728 1005945
rect 92560 1005819 92566 1005871
rect 92618 1005859 92624 1005871
rect 101008 1005859 101014 1005871
rect 92618 1005831 101014 1005859
rect 92618 1005819 92624 1005831
rect 101008 1005819 101014 1005831
rect 101066 1005819 101072 1005871
rect 262288 1005819 262294 1005871
rect 262346 1005859 262352 1005871
rect 276496 1005859 276502 1005871
rect 262346 1005831 276502 1005859
rect 262346 1005819 262352 1005831
rect 276496 1005819 276502 1005831
rect 276554 1005819 276560 1005871
rect 359344 1005819 359350 1005871
rect 359402 1005859 359408 1005871
rect 380080 1005859 380086 1005871
rect 359402 1005831 380086 1005859
rect 359402 1005819 359408 1005831
rect 380080 1005819 380086 1005831
rect 380138 1005819 380144 1005871
rect 429712 1005819 429718 1005871
rect 429770 1005859 429776 1005871
rect 466480 1005859 466486 1005871
rect 429770 1005831 466486 1005859
rect 429770 1005819 429776 1005831
rect 466480 1005819 466486 1005831
rect 466538 1005819 466544 1005871
rect 551632 1005819 551638 1005871
rect 551690 1005859 551696 1005871
rect 571600 1005859 571606 1005871
rect 551690 1005831 571606 1005859
rect 551690 1005819 551696 1005831
rect 571600 1005819 571606 1005831
rect 571658 1005819 571664 1005871
rect 428272 1005745 428278 1005797
rect 428330 1005785 428336 1005797
rect 460816 1005785 460822 1005797
rect 428330 1005757 460822 1005785
rect 428330 1005745 428336 1005757
rect 460816 1005745 460822 1005757
rect 460874 1005745 460880 1005797
rect 502288 1005745 502294 1005797
rect 502346 1005785 502352 1005797
rect 518512 1005785 518518 1005797
rect 502346 1005757 518518 1005785
rect 502346 1005745 502352 1005757
rect 518512 1005745 518518 1005757
rect 518570 1005745 518576 1005797
rect 553648 1005745 553654 1005797
rect 553706 1005785 553712 1005797
rect 571312 1005785 571318 1005797
rect 553706 1005757 571318 1005785
rect 553706 1005745 553712 1005757
rect 571312 1005745 571318 1005757
rect 571370 1005745 571376 1005797
rect 361840 1005671 361846 1005723
rect 361898 1005711 361904 1005723
rect 383632 1005711 383638 1005723
rect 361898 1005683 383638 1005711
rect 361898 1005671 361904 1005683
rect 383632 1005671 383638 1005683
rect 383690 1005671 383696 1005723
rect 428656 1005671 428662 1005723
rect 428714 1005711 428720 1005723
rect 469264 1005711 469270 1005723
rect 428714 1005683 469270 1005711
rect 428714 1005671 428720 1005683
rect 469264 1005671 469270 1005683
rect 469322 1005671 469328 1005723
rect 501712 1005671 501718 1005723
rect 501770 1005711 501776 1005723
rect 523984 1005711 523990 1005723
rect 501770 1005683 523990 1005711
rect 501770 1005671 501776 1005683
rect 523984 1005671 523990 1005683
rect 524042 1005671 524048 1005723
rect 554608 1005671 554614 1005723
rect 554666 1005711 554672 1005723
rect 573040 1005711 573046 1005723
rect 554666 1005683 573046 1005711
rect 554666 1005671 554672 1005683
rect 573040 1005671 573046 1005683
rect 573098 1005671 573104 1005723
rect 92944 1005597 92950 1005649
rect 93002 1005637 93008 1005649
rect 109936 1005637 109942 1005649
rect 93002 1005609 109942 1005637
rect 93002 1005597 93008 1005609
rect 109936 1005597 109942 1005609
rect 109994 1005597 110000 1005649
rect 358288 1005597 358294 1005649
rect 358346 1005637 358352 1005649
rect 379984 1005637 379990 1005649
rect 358346 1005609 379990 1005637
rect 358346 1005597 358352 1005609
rect 379984 1005597 379990 1005609
rect 380042 1005597 380048 1005649
rect 426736 1005597 426742 1005649
rect 426794 1005637 426800 1005649
rect 472048 1005637 472054 1005649
rect 426794 1005609 472054 1005637
rect 426794 1005597 426800 1005609
rect 472048 1005597 472054 1005609
rect 472106 1005597 472112 1005649
rect 554032 1005597 554038 1005649
rect 554090 1005637 554096 1005649
rect 572944 1005637 572950 1005649
rect 554090 1005609 572950 1005637
rect 554090 1005597 554096 1005609
rect 572944 1005597 572950 1005609
rect 573002 1005597 573008 1005649
rect 94096 1005523 94102 1005575
rect 94154 1005563 94160 1005575
rect 110512 1005563 110518 1005575
rect 94154 1005535 110518 1005563
rect 94154 1005523 94160 1005535
rect 110512 1005523 110518 1005535
rect 110570 1005523 110576 1005575
rect 158512 1005523 158518 1005575
rect 158570 1005563 158576 1005575
rect 172912 1005563 172918 1005575
rect 158570 1005535 172918 1005563
rect 158570 1005523 158576 1005535
rect 172912 1005523 172918 1005535
rect 172970 1005523 172976 1005575
rect 356752 1005523 356758 1005575
rect 356810 1005563 356816 1005575
rect 371536 1005563 371542 1005575
rect 356810 1005535 371542 1005563
rect 356810 1005523 356816 1005535
rect 371536 1005523 371542 1005535
rect 371594 1005523 371600 1005575
rect 425296 1005523 425302 1005575
rect 425354 1005563 425360 1005575
rect 471856 1005563 471862 1005575
rect 425354 1005535 471862 1005563
rect 425354 1005523 425360 1005535
rect 471856 1005523 471862 1005535
rect 471914 1005523 471920 1005575
rect 502672 1005523 502678 1005575
rect 502730 1005563 502736 1005575
rect 502730 1005535 518366 1005563
rect 502730 1005523 502736 1005535
rect 92656 1005449 92662 1005501
rect 92714 1005489 92720 1005501
rect 102064 1005489 102070 1005501
rect 92714 1005461 102070 1005489
rect 92714 1005449 92720 1005461
rect 102064 1005449 102070 1005461
rect 102122 1005449 102128 1005501
rect 151120 1005449 151126 1005501
rect 151178 1005489 151184 1005501
rect 161392 1005489 161398 1005501
rect 151178 1005461 161398 1005489
rect 151178 1005449 151184 1005461
rect 161392 1005449 161398 1005461
rect 161450 1005449 161456 1005501
rect 197200 1005449 197206 1005501
rect 197258 1005489 197264 1005501
rect 207376 1005489 207382 1005501
rect 197258 1005461 207382 1005489
rect 197258 1005449 197264 1005461
rect 207376 1005449 207382 1005461
rect 207434 1005449 207440 1005501
rect 357136 1005449 357142 1005501
rect 357194 1005489 357200 1005501
rect 372016 1005489 372022 1005501
rect 357194 1005461 372022 1005489
rect 357194 1005449 357200 1005461
rect 372016 1005449 372022 1005461
rect 372074 1005449 372080 1005501
rect 423760 1005449 423766 1005501
rect 423818 1005489 423824 1005501
rect 471760 1005489 471766 1005501
rect 423818 1005461 471766 1005489
rect 423818 1005449 423824 1005461
rect 471760 1005449 471766 1005461
rect 471818 1005449 471824 1005501
rect 500752 1005449 500758 1005501
rect 500810 1005489 500816 1005501
rect 509680 1005489 509686 1005501
rect 500810 1005461 509686 1005489
rect 500810 1005449 500816 1005461
rect 509680 1005449 509686 1005461
rect 509738 1005449 509744 1005501
rect 518338 1005489 518366 1005535
rect 518416 1005489 518422 1005501
rect 518338 1005461 518422 1005489
rect 518416 1005449 518422 1005461
rect 518474 1005449 518480 1005501
rect 555184 1005449 555190 1005501
rect 555242 1005489 555248 1005501
rect 571984 1005489 571990 1005501
rect 555242 1005461 571990 1005489
rect 555242 1005449 555248 1005461
rect 571984 1005449 571990 1005461
rect 572042 1005449 572048 1005501
rect 152656 1005375 152662 1005427
rect 152714 1005415 152720 1005427
rect 161872 1005415 161878 1005427
rect 152714 1005387 161878 1005415
rect 152714 1005375 152720 1005387
rect 161872 1005375 161878 1005387
rect 161930 1005375 161936 1005427
rect 361264 1005375 361270 1005427
rect 361322 1005415 361328 1005427
rect 374992 1005415 374998 1005427
rect 361322 1005387 374998 1005415
rect 361322 1005375 361328 1005387
rect 374992 1005375 374998 1005387
rect 375050 1005375 375056 1005427
rect 424720 1005375 424726 1005427
rect 424778 1005415 424784 1005427
rect 472144 1005415 472150 1005427
rect 424778 1005387 472150 1005415
rect 424778 1005375 424784 1005387
rect 472144 1005375 472150 1005387
rect 472202 1005375 472208 1005427
rect 503728 1005375 503734 1005427
rect 503786 1005415 503792 1005427
rect 520528 1005415 520534 1005427
rect 503786 1005387 520534 1005415
rect 503786 1005375 503792 1005387
rect 520528 1005375 520534 1005387
rect 520586 1005375 520592 1005427
rect 107056 1005301 107062 1005353
rect 107114 1005341 107120 1005353
rect 124624 1005341 124630 1005353
rect 107114 1005313 124630 1005341
rect 107114 1005301 107120 1005313
rect 124624 1005301 124630 1005313
rect 124682 1005301 124688 1005353
rect 159472 1005301 159478 1005353
rect 159530 1005341 159536 1005353
rect 172816 1005341 172822 1005353
rect 159530 1005313 172822 1005341
rect 159530 1005301 159536 1005313
rect 172816 1005301 172822 1005313
rect 172874 1005301 172880 1005353
rect 210832 1005301 210838 1005353
rect 210890 1005341 210896 1005353
rect 227344 1005341 227350 1005353
rect 210890 1005313 227350 1005341
rect 210890 1005301 210896 1005313
rect 227344 1005301 227350 1005313
rect 227402 1005301 227408 1005353
rect 316432 1005301 316438 1005353
rect 316490 1005341 316496 1005353
rect 331216 1005341 331222 1005353
rect 316490 1005313 331222 1005341
rect 316490 1005301 316496 1005313
rect 331216 1005301 331222 1005313
rect 331274 1005301 331280 1005353
rect 360880 1005301 360886 1005353
rect 360938 1005341 360944 1005353
rect 374512 1005341 374518 1005353
rect 360938 1005313 374518 1005341
rect 360938 1005301 360944 1005313
rect 374512 1005301 374518 1005313
rect 374570 1005301 374576 1005353
rect 424144 1005301 424150 1005353
rect 424202 1005341 424208 1005353
rect 471952 1005341 471958 1005353
rect 424202 1005313 471958 1005341
rect 424202 1005301 424208 1005313
rect 471952 1005301 471958 1005313
rect 472010 1005301 472016 1005353
rect 505264 1005301 505270 1005353
rect 505322 1005341 505328 1005353
rect 520336 1005341 520342 1005353
rect 505322 1005313 520342 1005341
rect 505322 1005301 505328 1005313
rect 520336 1005301 520342 1005313
rect 520394 1005301 520400 1005353
rect 552592 1005301 552598 1005353
rect 552650 1005341 552656 1005353
rect 561520 1005341 561526 1005353
rect 552650 1005313 561526 1005341
rect 552650 1005301 552656 1005313
rect 561520 1005301 561526 1005313
rect 561578 1005301 561584 1005353
rect 161488 1005227 161494 1005279
rect 161546 1005267 161552 1005279
rect 169936 1005267 169942 1005279
rect 161546 1005239 169942 1005267
rect 161546 1005227 161552 1005239
rect 169936 1005227 169942 1005239
rect 169994 1005227 170000 1005279
rect 201616 1005227 201622 1005279
rect 201674 1005267 201680 1005279
rect 212848 1005267 212854 1005279
rect 201674 1005239 212854 1005267
rect 201674 1005227 201680 1005239
rect 212848 1005227 212854 1005239
rect 212906 1005227 212912 1005279
rect 313840 1005227 313846 1005279
rect 313898 1005267 313904 1005279
rect 329680 1005267 329686 1005279
rect 313898 1005239 329686 1005267
rect 313898 1005227 313904 1005239
rect 329680 1005227 329686 1005239
rect 329738 1005227 329744 1005279
rect 362320 1005227 362326 1005279
rect 362378 1005267 362384 1005279
rect 374608 1005267 374614 1005279
rect 362378 1005239 374614 1005267
rect 362378 1005227 362384 1005239
rect 374608 1005227 374614 1005239
rect 374666 1005227 374672 1005279
rect 426160 1005227 426166 1005279
rect 426218 1005267 426224 1005279
rect 472240 1005267 472246 1005279
rect 426218 1005239 472246 1005267
rect 426218 1005227 426224 1005239
rect 472240 1005227 472246 1005239
rect 472298 1005227 472304 1005279
rect 503248 1005227 503254 1005279
rect 503306 1005267 503312 1005279
rect 521296 1005267 521302 1005279
rect 503306 1005239 521302 1005267
rect 503306 1005227 503312 1005239
rect 521296 1005227 521302 1005239
rect 521354 1005227 521360 1005279
rect 552208 1005227 552214 1005279
rect 552266 1005267 552272 1005279
rect 561040 1005267 561046 1005279
rect 552266 1005239 561046 1005267
rect 552266 1005227 552272 1005239
rect 561040 1005227 561046 1005239
rect 561098 1005227 561104 1005279
rect 98032 1005153 98038 1005205
rect 98090 1005193 98096 1005205
rect 105424 1005193 105430 1005205
rect 98090 1005165 105430 1005193
rect 98090 1005153 98096 1005165
rect 105424 1005153 105430 1005165
rect 105482 1005153 105488 1005205
rect 108016 1005153 108022 1005205
rect 108074 1005193 108080 1005205
rect 126640 1005193 126646 1005205
rect 108074 1005165 126646 1005193
rect 108074 1005153 108080 1005165
rect 126640 1005153 126646 1005165
rect 126698 1005153 126704 1005205
rect 160912 1005153 160918 1005205
rect 160970 1005193 160976 1005205
rect 166958 1005193 166964 1005205
rect 160970 1005165 166964 1005193
rect 160970 1005153 160976 1005165
rect 166958 1005153 166964 1005165
rect 167016 1005153 167022 1005205
rect 209872 1005153 209878 1005205
rect 209930 1005193 209936 1005205
rect 225424 1005193 225430 1005205
rect 209930 1005165 225430 1005193
rect 209930 1005153 209936 1005165
rect 225424 1005153 225430 1005165
rect 225482 1005153 225488 1005205
rect 298480 1005153 298486 1005205
rect 298538 1005193 298544 1005205
rect 308272 1005193 308278 1005205
rect 298538 1005165 308278 1005193
rect 298538 1005153 298544 1005165
rect 308272 1005153 308278 1005165
rect 308330 1005153 308336 1005205
rect 312880 1005153 312886 1005205
rect 312938 1005193 312944 1005205
rect 329776 1005193 329782 1005205
rect 312938 1005165 329782 1005193
rect 312938 1005153 312944 1005165
rect 329776 1005153 329782 1005165
rect 329834 1005153 329840 1005205
rect 362800 1005153 362806 1005205
rect 362858 1005193 362864 1005205
rect 374416 1005193 374422 1005205
rect 362858 1005165 374422 1005193
rect 362858 1005153 362864 1005165
rect 374416 1005153 374422 1005165
rect 374474 1005153 374480 1005205
rect 501136 1005153 501142 1005205
rect 501194 1005193 501200 1005205
rect 501194 1005165 506654 1005193
rect 501194 1005153 501200 1005165
rect 506626 1005119 506654 1005165
rect 506704 1005153 506710 1005205
rect 506762 1005193 506768 1005205
rect 506762 1005165 518414 1005193
rect 506762 1005153 506768 1005165
rect 509776 1005119 509782 1005131
rect 506626 1005091 509782 1005119
rect 509776 1005079 509782 1005091
rect 509834 1005079 509840 1005131
rect 518386 1005119 518414 1005165
rect 552976 1005153 552982 1005205
rect 553034 1005193 553040 1005205
rect 553034 1005165 561566 1005193
rect 553034 1005153 553040 1005165
rect 521488 1005119 521494 1005131
rect 518386 1005091 521494 1005119
rect 521488 1005079 521494 1005091
rect 521546 1005079 521552 1005131
rect 561538 1005119 561566 1005165
rect 564304 1005119 564310 1005131
rect 561538 1005091 564310 1005119
rect 564304 1005079 564310 1005091
rect 564362 1005079 564368 1005131
rect 372016 1005005 372022 1005057
rect 372074 1005045 372080 1005057
rect 380176 1005045 380182 1005057
rect 372074 1005017 380182 1005045
rect 372074 1005005 372080 1005017
rect 380176 1005005 380182 1005017
rect 380234 1005005 380240 1005057
rect 371536 1004931 371542 1004983
rect 371594 1004971 371600 1004983
rect 380368 1004971 380374 1004983
rect 371594 1004943 380374 1004971
rect 371594 1004931 371600 1004943
rect 380368 1004931 380374 1004943
rect 380426 1004931 380432 1004983
rect 371632 1004857 371638 1004909
rect 371690 1004897 371696 1004909
rect 380464 1004897 380470 1004909
rect 371690 1004869 380470 1004897
rect 371690 1004857 371696 1004869
rect 380464 1004857 380470 1004869
rect 380522 1004857 380528 1004909
rect 143824 1004783 143830 1004835
rect 143882 1004823 143888 1004835
rect 156976 1004823 156982 1004835
rect 143882 1004795 156982 1004823
rect 143882 1004783 143888 1004795
rect 156976 1004783 156982 1004795
rect 157034 1004783 157040 1004835
rect 520336 1002711 520342 1002763
rect 520394 1002751 520400 1002763
rect 521584 1002751 521590 1002763
rect 520394 1002723 521590 1002751
rect 520394 1002711 520400 1002723
rect 521584 1002711 521590 1002723
rect 521642 1002711 521648 1002763
rect 299536 1002637 299542 1002689
rect 299594 1002677 299600 1002689
rect 306736 1002677 306742 1002689
rect 299594 1002649 306742 1002677
rect 299594 1002637 299600 1002649
rect 306736 1002637 306742 1002649
rect 306794 1002637 306800 1002689
rect 299728 1002563 299734 1002615
rect 299786 1002603 299792 1002615
rect 307312 1002603 307318 1002615
rect 299786 1002575 307318 1002603
rect 299786 1002563 299792 1002575
rect 307312 1002563 307318 1002575
rect 307370 1002563 307376 1002615
rect 300112 1002489 300118 1002541
rect 300170 1002529 300176 1002541
rect 307888 1002529 307894 1002541
rect 300170 1002501 307894 1002529
rect 300170 1002489 300176 1002501
rect 307888 1002489 307894 1002501
rect 307946 1002489 307952 1002541
rect 97840 1002415 97846 1002467
rect 97898 1002455 97904 1002467
rect 103024 1002455 103030 1002467
rect 97898 1002427 103030 1002455
rect 97898 1002415 97904 1002427
rect 103024 1002415 103030 1002427
rect 103082 1002415 103088 1002467
rect 246928 1002415 246934 1002467
rect 246986 1002455 246992 1002467
rect 255280 1002455 255286 1002467
rect 246986 1002427 255286 1002455
rect 246986 1002415 246992 1002427
rect 255280 1002415 255286 1002427
rect 255338 1002415 255344 1002467
rect 299632 1002415 299638 1002467
rect 299690 1002455 299696 1002467
rect 305296 1002455 305302 1002467
rect 299690 1002427 305302 1002455
rect 299690 1002415 299696 1002427
rect 305296 1002415 305302 1002427
rect 305354 1002415 305360 1002467
rect 95056 1002341 95062 1002393
rect 95114 1002381 95120 1002393
rect 101488 1002381 101494 1002393
rect 95114 1002353 101494 1002381
rect 95114 1002341 95120 1002353
rect 101488 1002341 101494 1002353
rect 101546 1002341 101552 1002393
rect 246544 1002341 246550 1002393
rect 246602 1002381 246608 1002393
rect 253648 1002381 253654 1002393
rect 246602 1002353 253654 1002381
rect 246602 1002341 246608 1002353
rect 253648 1002341 253654 1002353
rect 253706 1002341 253712 1002393
rect 300016 1002341 300022 1002393
rect 300074 1002381 300080 1002393
rect 306352 1002381 306358 1002393
rect 300074 1002353 306358 1002381
rect 300074 1002341 300080 1002353
rect 306352 1002341 306358 1002353
rect 306410 1002341 306416 1002393
rect 561040 1002341 561046 1002393
rect 561098 1002381 561104 1002393
rect 564400 1002381 564406 1002393
rect 561098 1002353 564406 1002381
rect 561098 1002341 561104 1002353
rect 564400 1002341 564406 1002353
rect 564458 1002341 564464 1002393
rect 100528 1002267 100534 1002319
rect 100586 1002307 100592 1002319
rect 103600 1002307 103606 1002319
rect 100586 1002279 103606 1002307
rect 100586 1002267 100592 1002279
rect 103600 1002267 103606 1002279
rect 103658 1002267 103664 1002319
rect 143920 1002267 143926 1002319
rect 143978 1002307 143984 1002319
rect 153040 1002307 153046 1002319
rect 143978 1002279 153046 1002307
rect 143978 1002267 143984 1002279
rect 153040 1002267 153046 1002279
rect 153098 1002267 153104 1002319
rect 246832 1002267 246838 1002319
rect 246890 1002307 246896 1002319
rect 254224 1002307 254230 1002319
rect 246890 1002279 254230 1002307
rect 246890 1002267 246896 1002279
rect 254224 1002267 254230 1002279
rect 254282 1002267 254288 1002319
rect 299824 1002267 299830 1002319
rect 299882 1002307 299888 1002319
rect 305776 1002307 305782 1002319
rect 299882 1002279 305782 1002307
rect 299882 1002267 299888 1002279
rect 305776 1002267 305782 1002279
rect 305834 1002267 305840 1002319
rect 505648 1002267 505654 1002319
rect 505706 1002307 505712 1002319
rect 521392 1002307 521398 1002319
rect 505706 1002279 521398 1002307
rect 505706 1002267 505712 1002279
rect 521392 1002267 521398 1002279
rect 521450 1002267 521456 1002319
rect 558544 1002267 558550 1002319
rect 558602 1002307 558608 1002319
rect 567376 1002307 567382 1002319
rect 558602 1002279 567382 1002307
rect 558602 1002267 558608 1002279
rect 567376 1002267 567382 1002279
rect 567434 1002267 567440 1002319
rect 509680 1002193 509686 1002245
rect 509738 1002233 509744 1002245
rect 515824 1002233 515830 1002245
rect 509738 1002205 515830 1002233
rect 509738 1002193 509744 1002205
rect 515824 1002193 515830 1002205
rect 515882 1002193 515888 1002245
rect 374416 1000935 374422 1000987
rect 374474 1000975 374480 1000987
rect 383440 1000975 383446 1000987
rect 374474 1000947 383446 1000975
rect 374474 1000935 374480 1000947
rect 383440 1000935 383446 1000947
rect 383498 1000935 383504 1000987
rect 430192 1000935 430198 1000987
rect 430250 1000975 430256 1000987
rect 472624 1000975 472630 1000987
rect 430250 1000947 472630 1000975
rect 430250 1000935 430256 1000947
rect 472624 1000935 472630 1000947
rect 472682 1000935 472688 1000987
rect 374992 1000861 374998 1000913
rect 375050 1000901 375056 1000913
rect 383344 1000901 383350 1000913
rect 375050 1000873 383350 1000901
rect 375050 1000861 375056 1000873
rect 383344 1000861 383350 1000873
rect 383402 1000861 383408 1000913
rect 429232 1000861 429238 1000913
rect 429290 1000901 429296 1000913
rect 472528 1000901 472534 1000913
rect 429290 1000873 472534 1000901
rect 429290 1000861 429296 1000873
rect 472528 1000861 472534 1000873
rect 472586 1000861 472592 1000913
rect 195184 1000787 195190 1000839
rect 195242 1000827 195248 1000839
rect 208432 1000827 208438 1000839
rect 195242 1000799 208438 1000827
rect 195242 1000787 195248 1000799
rect 208432 1000787 208438 1000799
rect 208490 1000787 208496 1000839
rect 359728 1000787 359734 1000839
rect 359786 1000827 359792 1000839
rect 383536 1000827 383542 1000839
rect 359786 1000799 383542 1000827
rect 359786 1000787 359792 1000799
rect 383536 1000787 383542 1000799
rect 383594 1000787 383600 1000839
rect 427120 1000787 427126 1000839
rect 427178 1000827 427184 1000839
rect 472624 1000827 472630 1000839
rect 427178 1000799 472630 1000827
rect 427178 1000787 427184 1000799
rect 472624 1000787 472630 1000799
rect 472682 1000787 472688 1000839
rect 507184 1000787 507190 1000839
rect 507242 1000827 507248 1000839
rect 517856 1000827 517862 1000839
rect 507242 1000799 517862 1000827
rect 507242 1000787 507248 1000799
rect 517856 1000787 517862 1000799
rect 517914 1000787 517920 1000839
rect 506224 1000639 506230 1000691
rect 506282 1000679 506288 1000691
rect 518080 1000679 518086 1000691
rect 506282 1000651 518086 1000679
rect 506282 1000639 506288 1000651
rect 518080 1000639 518086 1000651
rect 518138 1000639 518144 1000691
rect 298232 1000121 298238 1000173
rect 298290 1000161 298296 1000173
rect 299632 1000161 299638 1000173
rect 298290 1000133 299638 1000161
rect 298290 1000121 298296 1000133
rect 299632 1000121 299638 1000133
rect 299690 1000121 299696 1000173
rect 92464 999677 92470 999729
rect 92522 999717 92528 999729
rect 95056 999717 95062 999729
rect 92522 999689 95062 999717
rect 92522 999677 92528 999689
rect 95056 999677 95062 999689
rect 95114 999677 95120 999729
rect 590704 999677 590710 999729
rect 590762 999717 590768 999729
rect 625552 999717 625558 999729
rect 590762 999689 625558 999717
rect 590762 999677 590768 999689
rect 625552 999677 625558 999689
rect 625610 999677 625616 999729
rect 609040 999603 609046 999655
rect 609098 999643 609104 999655
rect 625840 999643 625846 999655
rect 609098 999615 625846 999643
rect 609098 999603 609104 999615
rect 625840 999603 625846 999615
rect 625898 999603 625904 999655
rect 246640 999529 246646 999581
rect 246698 999569 246704 999581
rect 259792 999569 259798 999581
rect 246698 999541 259798 999569
rect 246698 999529 246704 999541
rect 259792 999529 259798 999541
rect 259850 999529 259856 999581
rect 298136 999529 298142 999581
rect 298194 999569 298200 999581
rect 311440 999569 311446 999581
rect 298194 999541 311446 999569
rect 298194 999529 298200 999541
rect 311440 999529 311446 999541
rect 311498 999529 311504 999581
rect 540304 999529 540310 999581
rect 540362 999569 540368 999581
rect 572848 999569 572854 999581
rect 540362 999541 572854 999569
rect 540362 999529 540368 999541
rect 572848 999529 572854 999541
rect 572906 999529 572912 999581
rect 590608 999529 590614 999581
rect 590666 999569 590672 999581
rect 625744 999569 625750 999581
rect 590666 999541 625750 999569
rect 590666 999529 590672 999541
rect 625744 999529 625750 999541
rect 625802 999529 625808 999581
rect 92292 999475 92298 999527
rect 92350 999495 92356 999527
rect 100528 999495 100534 999507
rect 92350 999475 100534 999495
rect 92307 999467 100534 999475
rect 100528 999455 100534 999467
rect 100586 999455 100592 999507
rect 247024 999455 247030 999507
rect 247082 999495 247088 999507
rect 256624 999495 256630 999507
rect 247082 999467 256630 999495
rect 247082 999455 247088 999467
rect 256624 999455 256630 999467
rect 256682 999455 256688 999507
rect 298328 999455 298334 999507
rect 298386 999495 298392 999507
rect 299824 999495 299830 999507
rect 298386 999467 299830 999495
rect 298386 999455 298392 999467
rect 299824 999455 299830 999467
rect 299882 999455 299888 999507
rect 380176 999455 380182 999507
rect 380234 999495 380240 999507
rect 382864 999495 382870 999507
rect 380234 999467 382870 999495
rect 380234 999455 380240 999467
rect 382864 999455 382870 999467
rect 382922 999455 382928 999507
rect 469264 999455 469270 999507
rect 469322 999495 469328 999507
rect 472432 999495 472438 999507
rect 469322 999467 472438 999495
rect 469322 999455 469328 999467
rect 472432 999455 472438 999467
rect 472490 999455 472496 999507
rect 504208 999455 504214 999507
rect 504266 999495 504272 999507
rect 518080 999495 518086 999507
rect 504266 999467 518086 999495
rect 504266 999455 504272 999467
rect 518080 999455 518086 999467
rect 518138 999455 518144 999507
rect 561616 999455 561622 999507
rect 561674 999495 561680 999507
rect 574864 999495 574870 999507
rect 561674 999467 574870 999495
rect 561674 999455 561680 999467
rect 574864 999455 574870 999467
rect 574922 999455 574928 999507
rect 590512 999455 590518 999507
rect 590570 999495 590576 999507
rect 625648 999495 625654 999507
rect 590570 999467 625654 999495
rect 590570 999455 590576 999467
rect 625648 999455 625654 999467
rect 625706 999455 625712 999507
rect 92368 999381 92374 999433
rect 92426 999421 92432 999433
rect 98032 999421 98038 999433
rect 92426 999393 98038 999421
rect 92426 999381 92432 999393
rect 98032 999381 98038 999393
rect 98090 999381 98096 999433
rect 143728 999381 143734 999433
rect 143786 999421 143792 999433
rect 154960 999421 154966 999433
rect 143786 999393 154966 999421
rect 143786 999381 143792 999393
rect 154960 999381 154966 999393
rect 155018 999381 155024 999433
rect 195088 999381 195094 999433
rect 195146 999421 195152 999433
rect 206320 999421 206326 999433
rect 195146 999393 206326 999421
rect 195146 999381 195152 999393
rect 206320 999381 206326 999393
rect 206378 999381 206384 999433
rect 246544 999381 246550 999433
rect 246602 999421 246608 999433
rect 257776 999421 257782 999433
rect 246602 999393 257782 999421
rect 246602 999381 246608 999393
rect 257776 999381 257782 999393
rect 257834 999381 257840 999433
rect 298136 999381 298142 999433
rect 298194 999421 298200 999433
rect 309328 999421 309334 999433
rect 298194 999393 309334 999421
rect 298194 999381 298200 999393
rect 309328 999381 309334 999393
rect 309386 999381 309392 999433
rect 380272 999381 380278 999433
rect 380330 999421 380336 999433
rect 382960 999421 382966 999433
rect 380330 999393 382966 999421
rect 380330 999381 380336 999393
rect 382960 999381 382966 999393
rect 383018 999381 383024 999433
rect 399916 999381 399922 999433
rect 399974 999421 399980 999433
rect 446512 999421 446518 999433
rect 399974 999393 446518 999421
rect 399974 999381 399980 999393
rect 446512 999381 446518 999393
rect 446570 999381 446576 999433
rect 460816 999381 460822 999433
rect 460874 999421 460880 999433
rect 469360 999421 469366 999433
rect 460874 999393 469366 999421
rect 460874 999381 460880 999393
rect 469360 999381 469366 999393
rect 469418 999381 469424 999433
rect 509776 999381 509782 999433
rect 509834 999421 509840 999433
rect 517744 999421 517750 999433
rect 509834 999393 517750 999421
rect 509834 999381 509840 999393
rect 517744 999381 517750 999393
rect 517802 999381 517808 999433
rect 564304 999381 564310 999433
rect 564362 999421 564368 999433
rect 564362 999393 570254 999421
rect 564362 999381 564368 999393
rect 570226 999347 570254 999393
rect 573136 999347 573142 999359
rect 570226 999319 573142 999347
rect 573136 999307 573142 999319
rect 573194 999307 573200 999359
rect 564496 998123 564502 998175
rect 564554 998163 564560 998175
rect 573232 998163 573238 998175
rect 564554 998135 573238 998163
rect 564554 998123 564560 998135
rect 573232 998123 573238 998135
rect 573290 998123 573296 998175
rect 92752 997901 92758 997953
rect 92810 997941 92816 997953
rect 106000 997941 106006 997953
rect 92810 997913 106006 997941
rect 92810 997901 92816 997913
rect 106000 997901 106006 997913
rect 106058 997901 106064 997953
rect 567376 997679 567382 997731
rect 567434 997719 567440 997731
rect 590512 997719 590518 997731
rect 567434 997691 590518 997719
rect 567434 997679 567440 997691
rect 590512 997679 590518 997691
rect 590570 997679 590576 997731
rect 555568 997605 555574 997657
rect 555626 997645 555632 997657
rect 625840 997645 625846 997657
rect 555626 997617 625846 997645
rect 555626 997605 555632 997617
rect 625840 997605 625846 997617
rect 625898 997605 625904 997657
rect 571984 997531 571990 997583
rect 572042 997571 572048 997583
rect 609040 997571 609046 997583
rect 572042 997543 609046 997571
rect 572042 997531 572048 997543
rect 609040 997531 609046 997543
rect 609098 997531 609104 997583
rect 557584 997457 557590 997509
rect 557642 997497 557648 997509
rect 590608 997497 590614 997509
rect 557642 997469 590614 997497
rect 557642 997457 557648 997469
rect 590608 997457 590614 997469
rect 590666 997457 590672 997509
rect 574864 997383 574870 997435
rect 574922 997423 574928 997435
rect 590704 997423 590710 997435
rect 574922 997395 590710 997423
rect 574922 997383 574928 997395
rect 590704 997383 590710 997395
rect 590762 997383 590768 997435
rect 377296 997087 377302 997139
rect 377354 997127 377360 997139
rect 382672 997127 382678 997139
rect 377354 997099 382678 997127
rect 377354 997087 377360 997099
rect 382672 997087 382678 997099
rect 382730 997087 382736 997139
rect 246736 996495 246742 996547
rect 246794 996535 246800 996547
rect 256240 996535 256246 996547
rect 246794 996507 256246 996535
rect 246794 996495 246800 996507
rect 256240 996495 256246 996507
rect 256298 996495 256304 996547
rect 299440 996495 299446 996547
rect 299498 996535 299504 996547
rect 309808 996535 309814 996547
rect 299498 996507 309814 996535
rect 299498 996495 299504 996507
rect 309808 996495 309814 996507
rect 309866 996495 309872 996547
rect 378832 996495 378838 996547
rect 378890 996535 378896 996547
rect 382768 996535 382774 996547
rect 378890 996507 382774 996535
rect 378890 996495 378896 996507
rect 382768 996495 382774 996507
rect 382826 996495 382832 996547
rect 572848 996495 572854 996547
rect 572906 996535 572912 996547
rect 576304 996535 576310 996547
rect 572906 996507 576310 996535
rect 572906 996495 572912 996507
rect 576304 996495 576310 996507
rect 576362 996495 576368 996547
rect 146896 996273 146902 996325
rect 146954 996313 146960 996325
rect 154384 996313 154390 996325
rect 146954 996285 154390 996313
rect 146954 996273 146960 996285
rect 154384 996273 154390 996285
rect 154442 996273 154448 996325
rect 108496 996199 108502 996251
rect 108554 996239 108560 996251
rect 112432 996239 112438 996251
rect 108554 996211 112438 996239
rect 108554 996199 108560 996211
rect 112432 996199 112438 996211
rect 112490 996199 112496 996251
rect 149680 996199 149686 996251
rect 149738 996239 149744 996251
rect 153424 996239 153430 996251
rect 149738 996211 153430 996239
rect 149738 996199 149744 996211
rect 153424 996199 153430 996211
rect 153482 996199 153488 996251
rect 159952 996239 159958 996251
rect 155506 996211 159958 996239
rect 115216 996125 115222 996177
rect 115274 996165 115280 996177
rect 155506 996165 155534 996211
rect 159952 996199 159958 996211
rect 160010 996199 160016 996251
rect 201520 996199 201526 996251
rect 201578 996239 201584 996251
rect 204880 996239 204886 996251
rect 201578 996211 204886 996239
rect 201578 996199 201584 996211
rect 204880 996199 204886 996211
rect 204938 996199 204944 996251
rect 115274 996137 155534 996165
rect 115274 996125 115280 996137
rect 166960 996125 166966 996177
rect 167018 996165 167024 996177
rect 211408 996165 211414 996177
rect 167018 996137 211414 996165
rect 167018 996125 167024 996137
rect 211408 996125 211414 996137
rect 211466 996125 211472 996177
rect 216016 996125 216022 996177
rect 216074 996165 216080 996177
rect 262768 996165 262774 996177
rect 216074 996137 262774 996165
rect 216074 996125 216080 996137
rect 262768 996125 262774 996137
rect 262826 996125 262832 996177
rect 276496 996125 276502 996177
rect 276554 996165 276560 996177
rect 314224 996165 314230 996177
rect 276554 996137 314230 996165
rect 276554 996125 276560 996137
rect 314224 996125 314230 996137
rect 314282 996165 314288 996177
rect 321616 996165 321622 996177
rect 314282 996137 321622 996165
rect 314282 996125 314288 996137
rect 321616 996125 321622 996137
rect 321674 996125 321680 996177
rect 374416 996125 374422 996177
rect 374474 996165 374480 996177
rect 432784 996165 432790 996177
rect 374474 996137 432790 996165
rect 374474 996125 374480 996137
rect 432784 996125 432790 996137
rect 432842 996125 432848 996177
rect 440656 996125 440662 996177
rect 440714 996165 440720 996177
rect 509776 996165 509782 996177
rect 440714 996137 509782 996165
rect 440714 996125 440720 996137
rect 509776 996125 509782 996137
rect 509834 996125 509840 996177
rect 510736 996125 510742 996177
rect 510794 996165 510800 996177
rect 515728 996165 515734 996177
rect 510794 996137 515734 996165
rect 510794 996125 510800 996137
rect 515728 996125 515734 996137
rect 515786 996125 515792 996177
rect 126640 996051 126646 996103
rect 126698 996091 126704 996103
rect 126698 996063 155534 996091
rect 126698 996051 126704 996063
rect 124624 995977 124630 996029
rect 124682 996017 124688 996029
rect 124682 995989 126734 996017
rect 124682 995977 124688 995989
rect 92752 995943 92758 995955
rect 78658 995915 92758 995943
rect 78658 995807 78686 995915
rect 92752 995903 92758 995915
rect 92810 995903 92816 995955
rect 100528 995869 100534 995881
rect 82306 995841 100534 995869
rect 82306 995807 82334 995841
rect 100528 995829 100534 995841
rect 100586 995829 100592 995881
rect 126706 995869 126734 995989
rect 146800 995977 146806 996029
rect 146858 996017 146864 996029
rect 152368 996017 152374 996029
rect 146858 995989 152374 996017
rect 146858 995977 146864 995989
rect 152368 995977 152374 995989
rect 152426 995977 152432 996029
rect 146704 995903 146710 995955
rect 146762 995943 146768 995955
rect 151984 995943 151990 995955
rect 146762 995915 151990 995943
rect 146762 995903 146768 995915
rect 151984 995903 151990 995915
rect 152042 995903 152048 995955
rect 155506 995943 155534 996063
rect 158896 996051 158902 996103
rect 158954 996091 158960 996103
rect 164272 996091 164278 996103
rect 158954 996063 164278 996091
rect 158954 996051 158960 996063
rect 164272 996051 164278 996063
rect 164330 996051 164336 996103
rect 172816 996051 172822 996103
rect 172874 996091 172880 996103
rect 210832 996091 210838 996103
rect 172874 996063 210838 996091
rect 172874 996051 172880 996063
rect 210832 996051 210838 996063
rect 210890 996051 210896 996103
rect 212752 996051 212758 996103
rect 212810 996091 212816 996103
rect 216112 996091 216118 996103
rect 212810 996063 216118 996091
rect 212810 996051 212816 996063
rect 216112 996051 216118 996063
rect 216170 996051 216176 996103
rect 227344 996051 227350 996103
rect 227402 996091 227408 996103
rect 227402 996063 247694 996091
rect 227402 996051 227408 996063
rect 172912 995977 172918 996029
rect 172970 996017 172976 996029
rect 172970 995989 210206 996017
rect 172970 995977 172976 995989
rect 159664 995943 159670 995955
rect 155506 995915 159670 995943
rect 159664 995903 159670 995915
rect 159722 995943 159728 995955
rect 164176 995943 164182 995955
rect 159722 995915 164182 995943
rect 159722 995903 159728 995915
rect 164176 995903 164182 995915
rect 164234 995903 164240 995955
rect 198736 995903 198742 995955
rect 198794 995943 198800 995955
rect 205936 995943 205942 995955
rect 198794 995915 205942 995943
rect 198794 995903 198800 995915
rect 205936 995903 205942 995915
rect 205994 995903 206000 995955
rect 210178 995881 210206 995989
rect 210850 995943 210878 996051
rect 247666 996017 247694 996063
rect 263728 996051 263734 996103
rect 263786 996091 263792 996103
rect 313840 996091 313846 996103
rect 263786 996063 313846 996091
rect 263786 996051 263792 996063
rect 313840 996051 313846 996063
rect 313898 996051 313904 996103
rect 366736 996051 366742 996103
rect 366794 996091 366800 996103
rect 371632 996091 371638 996103
rect 366794 996063 371638 996091
rect 366794 996051 366800 996063
rect 371632 996051 371638 996063
rect 371690 996051 371696 996103
rect 434128 996051 434134 996103
rect 434186 996091 434192 996103
rect 437776 996091 437782 996103
rect 434186 996063 437782 996091
rect 434186 996051 434192 996063
rect 437776 996051 437782 996063
rect 437834 996051 437840 996103
rect 512656 996051 512662 996103
rect 512714 996091 512720 996103
rect 561136 996091 561142 996103
rect 512714 996063 561142 996091
rect 512714 996051 512720 996063
rect 561136 996051 561142 996063
rect 561194 996051 561200 996103
rect 561904 996051 561910 996103
rect 561962 996091 561968 996103
rect 569968 996091 569974 996103
rect 561962 996063 569974 996091
rect 561962 996051 561968 996063
rect 569968 996051 569974 996063
rect 570026 996051 570032 996103
rect 262480 996017 262486 996029
rect 247666 995989 262486 996017
rect 262480 995977 262486 995989
rect 262538 996017 262544 996029
rect 268048 996017 268054 996029
rect 262538 995989 268054 996017
rect 262538 995977 262544 995989
rect 268048 995977 268054 995989
rect 268106 995977 268112 996029
rect 276592 995977 276598 996029
rect 276650 996017 276656 996029
rect 313072 996017 313078 996029
rect 276650 995989 313078 996017
rect 276650 995977 276656 995989
rect 313072 995977 313078 995989
rect 313130 996017 313136 996029
rect 317200 996017 317206 996029
rect 313130 995989 317206 996017
rect 313130 995977 313136 995989
rect 317200 995977 317206 995989
rect 317258 995977 317264 996029
rect 366256 995977 366262 996029
rect 366314 996017 366320 996029
rect 371728 996017 371734 996029
rect 366314 995989 371734 996017
rect 366314 995977 366320 995989
rect 371728 995977 371734 995989
rect 371786 995977 371792 996029
rect 382672 995977 382678 996029
rect 382730 996017 382736 996029
rect 382730 995989 393086 996017
rect 382730 995977 382736 995989
rect 216592 995943 216598 995955
rect 210850 995915 216598 995943
rect 216592 995903 216598 995915
rect 216650 995903 216656 995955
rect 225424 995903 225430 995955
rect 225482 995943 225488 995955
rect 261520 995943 261526 995955
rect 225482 995915 261526 995943
rect 225482 995903 225488 995915
rect 261520 995903 261526 995915
rect 261578 995943 261584 995955
rect 265168 995943 265174 995955
rect 261578 995915 265174 995943
rect 261578 995903 261584 995915
rect 265168 995903 265174 995915
rect 265226 995903 265232 995955
rect 382960 995903 382966 995955
rect 383018 995943 383024 995955
rect 383018 995915 387902 995943
rect 383018 995903 383024 995915
rect 158896 995869 158902 995881
rect 126706 995841 158902 995869
rect 158896 995829 158902 995841
rect 158954 995829 158960 995881
rect 203920 995869 203926 995881
rect 188866 995841 203926 995869
rect 188866 995807 188894 995841
rect 203920 995829 203926 995841
rect 203978 995829 203984 995881
rect 210160 995829 210166 995881
rect 210218 995869 210224 995881
rect 213136 995869 213142 995881
rect 210218 995841 213142 995869
rect 210218 995829 210224 995841
rect 213136 995829 213142 995841
rect 213194 995829 213200 995881
rect 246448 995869 246454 995881
rect 240898 995841 246454 995869
rect 240898 995807 240926 995841
rect 246448 995829 246454 995841
rect 246506 995829 246512 995881
rect 298232 995869 298238 995881
rect 296626 995841 298238 995869
rect 78640 995755 78646 995807
rect 78698 995755 78704 995807
rect 82288 995755 82294 995807
rect 82346 995755 82352 995807
rect 86224 995755 86230 995807
rect 86282 995795 86288 995807
rect 94960 995795 94966 995807
rect 86282 995767 94966 995795
rect 86282 995755 86288 995767
rect 94960 995755 94966 995767
rect 95018 995755 95024 995807
rect 142960 995755 142966 995807
rect 143018 995795 143024 995807
rect 143728 995795 143734 995807
rect 143018 995767 143734 995795
rect 143018 995755 143024 995767
rect 143728 995755 143734 995767
rect 143786 995755 143792 995807
rect 146704 995755 146710 995807
rect 146762 995795 146768 995807
rect 154000 995795 154006 995807
rect 146762 995767 154006 995795
rect 146762 995755 146768 995767
rect 154000 995755 154006 995767
rect 154058 995755 154064 995807
rect 188848 995755 188854 995807
rect 188906 995755 188912 995807
rect 189424 995755 189430 995807
rect 189482 995795 189488 995807
rect 202288 995795 202294 995807
rect 189482 995767 202294 995795
rect 189482 995755 189488 995767
rect 202288 995755 202294 995767
rect 202346 995755 202352 995807
rect 240880 995755 240886 995807
rect 240938 995755 240944 995807
rect 245680 995755 245686 995807
rect 245738 995795 245744 995807
rect 246544 995795 246550 995807
rect 245738 995767 246550 995795
rect 245738 995755 245744 995767
rect 246544 995755 246550 995767
rect 246602 995755 246608 995807
rect 292528 995755 292534 995807
rect 292586 995795 292592 995807
rect 296626 995795 296654 995841
rect 298232 995829 298238 995841
rect 298290 995829 298296 995881
rect 383440 995829 383446 995881
rect 383498 995869 383504 995881
rect 383498 995841 386078 995869
rect 383498 995829 383504 995841
rect 386050 995807 386078 995841
rect 292586 995767 296654 995795
rect 292586 995755 292592 995767
rect 297328 995755 297334 995807
rect 297386 995795 297392 995807
rect 298136 995795 298142 995807
rect 297386 995767 298142 995795
rect 297386 995755 297392 995767
rect 298136 995755 298142 995767
rect 298194 995755 298200 995807
rect 383632 995755 383638 995807
rect 383690 995795 383696 995807
rect 384400 995795 384406 995807
rect 383690 995767 384406 995795
rect 383690 995755 383696 995767
rect 384400 995755 384406 995767
rect 384458 995755 384464 995807
rect 386032 995755 386038 995807
rect 386090 995755 386096 995807
rect 387874 995795 387902 995915
rect 393058 995807 393086 995989
rect 433552 995977 433558 996029
rect 433610 996017 433616 996029
rect 437872 996017 437878 996029
rect 433610 995989 437878 996017
rect 433610 995977 433616 995989
rect 437872 995977 437878 995989
rect 437930 995977 437936 996029
rect 511120 995977 511126 996029
rect 511178 996017 511184 996029
rect 515632 996017 515638 996029
rect 511178 995989 515638 996017
rect 511178 995977 511184 995989
rect 515632 995977 515638 995989
rect 515690 995977 515696 996029
rect 471760 995903 471766 995955
rect 471818 995943 471824 995955
rect 471818 995915 478094 995943
rect 471818 995903 471824 995915
rect 472240 995829 472246 995881
rect 472298 995869 472304 995881
rect 472298 995841 477758 995869
rect 472298 995829 472304 995841
rect 477730 995807 477758 995841
rect 388048 995795 388054 995807
rect 387874 995767 388054 995795
rect 388048 995755 388054 995767
rect 388106 995755 388112 995807
rect 393040 995755 393046 995807
rect 393098 995755 393104 995807
rect 396592 995755 396598 995807
rect 396650 995795 396656 995807
rect 399856 995795 399862 995807
rect 396650 995767 399862 995795
rect 396650 995755 396656 995767
rect 399856 995755 399862 995767
rect 399914 995755 399920 995807
rect 472624 995755 472630 995807
rect 472682 995795 472688 995807
rect 474064 995795 474070 995807
rect 472682 995767 474070 995795
rect 472682 995755 472688 995767
rect 474064 995755 474070 995767
rect 474122 995755 474128 995807
rect 477712 995755 477718 995807
rect 477770 995755 477776 995807
rect 478066 995795 478094 995915
rect 523696 995903 523702 995955
rect 523754 995943 523760 995955
rect 523754 995915 529118 995943
rect 523754 995903 523760 995915
rect 523888 995829 523894 995881
rect 523946 995869 523952 995881
rect 523946 995841 526142 995869
rect 523946 995829 523952 995841
rect 526114 995807 526142 995841
rect 529090 995807 529118 995915
rect 625552 995903 625558 995955
rect 625610 995943 625616 995955
rect 625610 995915 634622 995943
rect 625610 995903 625616 995915
rect 625648 995829 625654 995881
rect 625706 995869 625712 995881
rect 625706 995841 627902 995869
rect 625706 995829 625712 995841
rect 627874 995807 627902 995841
rect 634594 995807 634622 995915
rect 482704 995795 482710 995807
rect 478066 995767 482710 995795
rect 482704 995755 482710 995767
rect 482762 995755 482768 995807
rect 524080 995755 524086 995807
rect 524138 995795 524144 995807
rect 525328 995795 525334 995807
rect 524138 995767 525334 995795
rect 524138 995755 524144 995767
rect 525328 995755 525334 995767
rect 525386 995755 525392 995807
rect 526096 995755 526102 995807
rect 526154 995755 526160 995807
rect 529072 995755 529078 995807
rect 529130 995755 529136 995807
rect 537136 995755 537142 995807
rect 537194 995795 537200 995807
rect 540304 995795 540310 995807
rect 537194 995767 540310 995795
rect 537194 995755 537200 995767
rect 540304 995755 540310 995767
rect 540362 995755 540368 995807
rect 625840 995755 625846 995807
rect 625898 995795 625904 995807
rect 627088 995795 627094 995807
rect 625898 995767 627094 995795
rect 625898 995755 625904 995767
rect 627088 995755 627094 995767
rect 627146 995755 627152 995807
rect 627856 995755 627862 995807
rect 627914 995755 627920 995807
rect 634576 995755 634582 995807
rect 634634 995755 634640 995807
rect 91504 995681 91510 995733
rect 91562 995721 91568 995733
rect 92272 995721 92278 995733
rect 91562 995693 92278 995721
rect 91562 995681 91568 995693
rect 92272 995681 92278 995693
rect 92330 995681 92336 995733
rect 141040 995681 141046 995733
rect 141098 995721 141104 995733
rect 143824 995721 143830 995733
rect 141098 995693 143830 995721
rect 141098 995681 141104 995693
rect 143824 995681 143830 995693
rect 143882 995681 143888 995733
rect 194416 995681 194422 995733
rect 194474 995721 194480 995733
rect 195088 995721 195094 995733
rect 194474 995693 195094 995721
rect 194474 995681 194480 995693
rect 195088 995681 195094 995693
rect 195146 995681 195152 995733
rect 243952 995681 243958 995733
rect 244010 995721 244016 995733
rect 246640 995721 246646 995733
rect 244010 995693 246646 995721
rect 244010 995681 244016 995693
rect 246640 995681 246646 995693
rect 246698 995681 246704 995733
rect 295408 995681 295414 995733
rect 295466 995721 295472 995733
rect 298040 995721 298046 995733
rect 295466 995693 298046 995721
rect 295466 995681 295472 995693
rect 298040 995681 298046 995693
rect 298098 995681 298104 995733
rect 383536 995681 383542 995733
rect 383594 995721 383600 995733
rect 384976 995721 384982 995733
rect 383594 995693 384982 995721
rect 383594 995681 383600 995693
rect 384976 995681 384982 995693
rect 385034 995681 385040 995733
rect 472528 995681 472534 995733
rect 472586 995721 472592 995733
rect 473296 995721 473302 995733
rect 472586 995693 473302 995721
rect 472586 995681 472592 995693
rect 473296 995681 473302 995693
rect 473354 995681 473360 995733
rect 523984 995681 523990 995733
rect 524042 995721 524048 995733
rect 524752 995721 524758 995733
rect 524042 995693 524758 995721
rect 524042 995681 524048 995693
rect 524752 995681 524758 995693
rect 524810 995681 524816 995733
rect 625744 995681 625750 995733
rect 625802 995721 625808 995733
rect 626512 995721 626518 995733
rect 625802 995693 626518 995721
rect 625802 995681 625808 995693
rect 626512 995681 626518 995693
rect 626570 995681 626576 995733
rect 89776 995607 89782 995659
rect 89834 995647 89840 995659
rect 92368 995647 92374 995659
rect 89834 995619 92374 995647
rect 89834 995607 89840 995619
rect 92368 995607 92374 995619
rect 92426 995607 92432 995659
rect 139312 995607 139318 995659
rect 139370 995647 139376 995659
rect 143920 995647 143926 995659
rect 139370 995619 143926 995647
rect 139370 995607 139376 995619
rect 143920 995607 143926 995619
rect 143978 995607 143984 995659
rect 192496 995607 192502 995659
rect 192554 995647 192560 995659
rect 195184 995647 195190 995659
rect 192554 995619 195190 995647
rect 192554 995607 192560 995619
rect 195184 995607 195190 995619
rect 195242 995607 195248 995659
rect 235792 995607 235798 995659
rect 235850 995647 235856 995659
rect 246736 995647 246742 995659
rect 235850 995619 246742 995647
rect 235850 995607 235856 995619
rect 246736 995607 246742 995619
rect 246794 995607 246800 995659
rect 290608 995607 290614 995659
rect 290666 995647 290672 995659
rect 299440 995647 299446 995659
rect 290666 995619 299446 995647
rect 290666 995607 290672 995619
rect 299440 995607 299446 995619
rect 299498 995607 299504 995659
rect 383344 995607 383350 995659
rect 383402 995647 383408 995659
rect 387472 995647 387478 995659
rect 383402 995619 387478 995647
rect 383402 995607 383408 995619
rect 387472 995607 387478 995619
rect 387530 995607 387536 995659
rect 472720 995607 472726 995659
rect 472778 995647 472784 995659
rect 474640 995647 474646 995659
rect 472778 995619 474646 995647
rect 472778 995607 472784 995619
rect 474640 995607 474646 995619
rect 474698 995607 474704 995659
rect 523792 995607 523798 995659
rect 523850 995647 523856 995659
rect 529744 995647 529750 995659
rect 523850 995619 529750 995647
rect 523850 995607 523856 995619
rect 529744 995607 529750 995619
rect 529802 995607 529808 995659
rect 625936 995607 625942 995659
rect 625994 995647 626000 995659
rect 630160 995647 630166 995659
rect 625994 995619 630166 995647
rect 625994 995607 626000 995619
rect 630160 995607 630166 995619
rect 630218 995607 630224 995659
rect 85360 995533 85366 995585
rect 85418 995573 85424 995585
rect 94960 995573 94966 995585
rect 85418 995545 94966 995573
rect 85418 995533 85424 995545
rect 94960 995533 94966 995545
rect 95018 995533 95024 995585
rect 236464 995533 236470 995585
rect 236522 995573 236528 995585
rect 254800 995573 254806 995585
rect 236522 995545 254806 995573
rect 236522 995533 236528 995545
rect 254800 995533 254806 995545
rect 254858 995533 254864 995585
rect 291184 995533 291190 995585
rect 291242 995573 291248 995585
rect 298328 995573 298334 995585
rect 291242 995545 298334 995573
rect 291242 995533 291248 995545
rect 298328 995533 298334 995545
rect 298386 995533 298392 995585
rect 382864 995533 382870 995585
rect 382922 995573 382928 995585
rect 389392 995573 389398 995585
rect 382922 995545 389398 995573
rect 382922 995533 382928 995545
rect 389392 995533 389398 995545
rect 389450 995533 389456 995585
rect 472048 995533 472054 995585
rect 472106 995573 472112 995585
rect 476944 995573 476950 995585
rect 472106 995545 476950 995573
rect 472106 995533 472112 995545
rect 476944 995533 476950 995545
rect 477002 995533 477008 995585
rect 480976 995573 480982 995585
rect 478066 995545 480982 995573
rect 87856 995459 87862 995511
rect 87914 995499 87920 995511
rect 92464 995499 92470 995511
rect 87914 995471 92470 995499
rect 87914 995459 87920 995471
rect 92464 995459 92470 995471
rect 92522 995459 92528 995511
rect 183760 995459 183766 995511
rect 183818 995499 183824 995511
rect 205264 995499 205270 995511
rect 183818 995471 205270 995499
rect 183818 995459 183824 995471
rect 205264 995459 205270 995471
rect 205322 995459 205328 995511
rect 239536 995459 239542 995511
rect 239594 995499 239600 995511
rect 246832 995499 246838 995511
rect 239594 995471 246838 995499
rect 239594 995459 239600 995471
rect 246832 995459 246838 995471
rect 246890 995459 246896 995511
rect 287920 995459 287926 995511
rect 287978 995499 287984 995511
rect 300016 995499 300022 995511
rect 287978 995471 300022 995499
rect 287978 995459 287984 995471
rect 300016 995459 300022 995471
rect 300074 995459 300080 995511
rect 380368 995459 380374 995511
rect 380426 995499 380432 995511
rect 392368 995499 392374 995511
rect 380426 995471 392374 995499
rect 380426 995459 380432 995471
rect 392368 995459 392374 995471
rect 392426 995459 392432 995511
rect 472432 995459 472438 995511
rect 472490 995499 472496 995511
rect 476368 995499 476374 995511
rect 472490 995471 476374 995499
rect 472490 995459 472496 995471
rect 476368 995459 476374 995471
rect 476426 995459 476432 995511
rect 380464 995385 380470 995437
rect 380522 995425 380528 995437
rect 393712 995425 393718 995437
rect 380522 995397 393718 995425
rect 380522 995385 380528 995397
rect 393712 995385 393718 995397
rect 393770 995385 393776 995437
rect 469360 995385 469366 995437
rect 469418 995425 469424 995437
rect 478066 995425 478094 995545
rect 480976 995533 480982 995545
rect 481034 995533 481040 995585
rect 523600 995533 523606 995585
rect 523658 995573 523664 995585
rect 528400 995573 528406 995585
rect 523658 995545 528406 995573
rect 523658 995533 523664 995545
rect 528400 995533 528406 995545
rect 528458 995533 528464 995585
rect 469418 995397 478094 995425
rect 469418 995385 469424 995397
rect 140368 995089 140374 995141
rect 140426 995129 140432 995141
rect 140426 995101 155534 995129
rect 140426 995089 140432 995101
rect 155506 995055 155534 995101
rect 186928 995055 186934 995067
rect 155506 995027 186934 995055
rect 186928 995015 186934 995027
rect 186986 995015 186992 995067
rect 517744 994127 517750 994179
rect 517802 994167 517808 994179
rect 532816 994167 532822 994179
rect 517802 994139 532822 994167
rect 517802 994127 517808 994139
rect 532816 994127 532822 994139
rect 532874 994127 532880 994179
rect 515824 993979 515830 994031
rect 515882 994019 515888 994031
rect 534352 994019 534358 994031
rect 515882 993991 534358 994019
rect 515882 993979 515888 993991
rect 534352 993979 534358 993991
rect 534410 993979 534416 994031
rect 571312 993905 571318 993957
rect 571370 993945 571376 993957
rect 635248 993945 635254 993957
rect 571370 993917 635254 993945
rect 571370 993905 571376 993917
rect 635248 993905 635254 993917
rect 635306 993905 635312 993957
rect 129328 993831 129334 993883
rect 129386 993871 129392 993883
rect 146896 993871 146902 993883
rect 129386 993843 146902 993871
rect 129386 993831 129392 993843
rect 146896 993831 146902 993843
rect 146954 993831 146960 993883
rect 180496 993831 180502 993883
rect 180554 993871 180560 993883
rect 198736 993871 198742 993883
rect 180554 993843 198742 993871
rect 180554 993831 180560 993843
rect 198736 993831 198742 993843
rect 198794 993831 198800 993883
rect 77680 993757 77686 993809
rect 77738 993797 77744 993809
rect 97840 993797 97846 993809
rect 77738 993769 97846 993797
rect 77738 993757 77744 993769
rect 97840 993757 97846 993769
rect 97898 993757 97904 993809
rect 131824 993757 131830 993809
rect 131882 993797 131888 993809
rect 156208 993797 156214 993809
rect 131882 993769 156214 993797
rect 131882 993757 131888 993769
rect 156208 993757 156214 993769
rect 156266 993757 156272 993809
rect 179824 993757 179830 993809
rect 179882 993797 179888 993809
rect 207856 993797 207862 993809
rect 179882 993769 207862 993797
rect 179882 993757 179888 993769
rect 207856 993757 207862 993769
rect 207914 993757 207920 993809
rect 561616 993757 561622 993809
rect 561674 993797 561680 993809
rect 634288 993797 634294 993809
rect 561674 993769 634294 993797
rect 561674 993757 561680 993769
rect 634288 993757 634294 993769
rect 634346 993757 634352 993809
rect 77296 993683 77302 993735
rect 77354 993723 77360 993735
rect 103600 993723 103606 993735
rect 77354 993695 103606 993723
rect 77354 993683 77360 993695
rect 103600 993683 103606 993695
rect 103658 993683 103664 993735
rect 128464 993683 128470 993735
rect 128522 993723 128528 993735
rect 156496 993723 156502 993735
rect 128522 993695 156502 993723
rect 128522 993683 128528 993695
rect 156496 993683 156502 993695
rect 156554 993683 156560 993735
rect 181360 993683 181366 993735
rect 181418 993723 181424 993735
rect 209104 993723 209110 993735
rect 181418 993695 209110 993723
rect 181418 993683 181424 993695
rect 209104 993683 209110 993695
rect 209162 993683 209168 993735
rect 232528 993683 232534 993735
rect 232586 993723 232592 993735
rect 260368 993723 260374 993735
rect 232586 993695 260374 993723
rect 232586 993683 232592 993695
rect 260368 993683 260374 993695
rect 260426 993683 260432 993735
rect 360016 993683 360022 993735
rect 360074 993723 360080 993735
rect 398800 993723 398806 993735
rect 360074 993695 398806 993723
rect 360074 993683 360080 993695
rect 398800 993683 398806 993695
rect 398858 993683 398864 993735
rect 427408 993683 427414 993735
rect 427466 993723 427472 993735
rect 487792 993723 487798 993735
rect 427466 993695 487798 993723
rect 427466 993683 427472 993695
rect 487792 993683 487798 993695
rect 487850 993683 487856 993735
rect 504400 993683 504406 993735
rect 504458 993723 504464 993735
rect 538960 993723 538966 993735
rect 504458 993695 538966 993723
rect 504458 993683 504464 993695
rect 538960 993683 538966 993695
rect 539018 993683 539024 993735
rect 555952 993683 555958 993735
rect 556010 993723 556016 993735
rect 641008 993723 641014 993735
rect 556010 993695 641014 993723
rect 556010 993683 556016 993695
rect 641008 993683 641014 993695
rect 641066 993683 641072 993735
rect 362896 993165 362902 993217
rect 362954 993205 362960 993217
rect 430864 993205 430870 993217
rect 362954 993177 430870 993205
rect 362954 993165 362960 993177
rect 430864 993165 430870 993177
rect 430922 993165 430928 993217
rect 363856 993091 363862 993143
rect 363914 993131 363920 993143
rect 431824 993131 431830 993143
rect 363914 993103 431830 993131
rect 363914 993091 363920 993103
rect 431824 993091 431830 993103
rect 431882 993091 431888 993143
rect 434896 993091 434902 993143
rect 434954 993131 434960 993143
rect 507856 993131 507862 993143
rect 434954 993103 507862 993131
rect 434954 993091 434960 993103
rect 507856 993091 507862 993103
rect 507914 993091 507920 993143
rect 559120 993131 559126 993143
rect 512674 993103 559126 993131
rect 431248 993017 431254 993069
rect 431306 993057 431312 993069
rect 508816 993057 508822 993069
rect 431306 993029 508822 993057
rect 431306 993017 431312 993029
rect 508816 993017 508822 993029
rect 508874 993017 508880 993069
rect 430192 992943 430198 992995
rect 430250 992983 430256 992995
rect 434896 992983 434902 992995
rect 430250 992955 434902 992983
rect 430250 992943 430256 992955
rect 434896 992943 434902 992955
rect 434954 992943 434960 992995
rect 507280 992943 507286 992995
rect 507338 992983 507344 992995
rect 512674 992983 512702 993103
rect 559120 993091 559126 993103
rect 559178 993091 559184 993143
rect 560176 993057 560182 993069
rect 507338 992955 512702 992983
rect 518386 993029 560182 993057
rect 507338 992943 507344 992955
rect 508432 992869 508438 992921
rect 508490 992909 508496 992921
rect 518386 992909 518414 993029
rect 560176 993017 560182 993029
rect 560234 993017 560240 993069
rect 508490 992881 518414 992909
rect 508490 992869 508496 992881
rect 331216 992573 331222 992625
rect 331274 992613 331280 992625
rect 332560 992613 332566 992625
rect 331274 992585 332566 992613
rect 331274 992573 331280 992585
rect 332560 992573 332566 992585
rect 332618 992573 332624 992625
rect 105808 990649 105814 990701
rect 105866 990689 105872 990701
rect 109552 990689 109558 990701
rect 105866 990661 109558 990689
rect 105866 990649 105872 990661
rect 109552 990649 109558 990661
rect 109610 990649 109616 990701
rect 373936 990649 373942 990701
rect 373994 990689 374000 990701
rect 381616 990689 381622 990701
rect 373994 990661 381622 990689
rect 373994 990649 374000 990661
rect 381616 990649 381622 990661
rect 381674 990649 381680 990701
rect 89584 989983 89590 990035
rect 89642 990023 89648 990035
rect 94096 990023 94102 990035
rect 89642 989995 94102 990023
rect 89642 989983 89648 989995
rect 94096 989983 94102 989995
rect 94154 989983 94160 990035
rect 569776 989761 569782 989813
rect 569834 989801 569840 989813
rect 592432 989801 592438 989813
rect 569834 989773 592438 989801
rect 569834 989761 569840 989773
rect 592432 989761 592438 989773
rect 592490 989761 592496 989813
rect 138256 989687 138262 989739
rect 138314 989727 138320 989739
rect 151120 989727 151126 989739
rect 138314 989699 151126 989727
rect 138314 989687 138320 989699
rect 151120 989687 151126 989699
rect 151178 989687 151184 989739
rect 371632 989687 371638 989739
rect 371690 989727 371696 989739
rect 397840 989727 397846 989739
rect 371690 989699 397846 989727
rect 371690 989687 371696 989699
rect 397840 989687 397846 989699
rect 397898 989687 397904 989739
rect 437776 989687 437782 989739
rect 437834 989727 437840 989739
rect 462736 989727 462742 989739
rect 437834 989699 462742 989727
rect 437834 989687 437840 989699
rect 462736 989687 462742 989699
rect 462794 989687 462800 989739
rect 515632 989687 515638 989739
rect 515690 989727 515696 989739
rect 527632 989727 527638 989739
rect 515690 989699 527638 989727
rect 515690 989687 515696 989699
rect 527632 989687 527638 989699
rect 527690 989687 527696 989739
rect 569872 989687 569878 989739
rect 569930 989727 569936 989739
rect 608752 989727 608758 989739
rect 569930 989699 608758 989727
rect 569930 989687 569936 989699
rect 608752 989687 608758 989699
rect 608810 989687 608816 989739
rect 371536 989613 371542 989665
rect 371594 989653 371600 989665
rect 414064 989653 414070 989665
rect 371594 989625 414070 989653
rect 371594 989613 371600 989625
rect 414064 989613 414070 989625
rect 414122 989613 414128 989665
rect 437968 989613 437974 989665
rect 438026 989653 438032 989665
rect 478960 989653 478966 989665
rect 438026 989625 478966 989653
rect 438026 989613 438032 989625
rect 478960 989613 478966 989625
rect 479018 989613 479024 989665
rect 491824 989613 491830 989665
rect 491882 989653 491888 989665
rect 511408 989653 511414 989665
rect 491882 989625 511414 989653
rect 491882 989613 491888 989625
rect 511408 989613 511414 989625
rect 511466 989613 511472 989665
rect 515536 989613 515542 989665
rect 515594 989653 515600 989665
rect 543760 989653 543766 989665
rect 515594 989625 543766 989653
rect 515594 989613 515600 989625
rect 543760 989613 543766 989625
rect 543818 989613 543824 989665
rect 569968 989613 569974 989665
rect 570026 989653 570032 989665
rect 624976 989653 624982 989665
rect 570026 989625 624982 989653
rect 570026 989613 570032 989625
rect 624976 989613 624982 989625
rect 625034 989613 625040 989665
rect 319696 989539 319702 989591
rect 319754 989579 319760 989591
rect 365392 989579 365398 989591
rect 319754 989551 365398 989579
rect 319754 989539 319760 989551
rect 365392 989539 365398 989551
rect 365450 989539 365456 989591
rect 371728 989539 371734 989591
rect 371786 989579 371792 989591
rect 430288 989579 430294 989591
rect 371786 989551 430294 989579
rect 371786 989539 371792 989551
rect 430288 989539 430294 989551
rect 430346 989539 430352 989591
rect 437872 989539 437878 989591
rect 437930 989579 437936 989591
rect 495184 989579 495190 989591
rect 437930 989551 495190 989579
rect 437930 989539 437936 989551
rect 495184 989539 495190 989551
rect 495242 989539 495248 989591
rect 515728 989539 515734 989591
rect 515786 989579 515792 989591
rect 560080 989579 560086 989591
rect 515786 989551 560086 989579
rect 515786 989539 515792 989551
rect 560080 989539 560086 989551
rect 560138 989539 560144 989591
rect 567184 989539 567190 989591
rect 567242 989579 567248 989591
rect 660880 989579 660886 989591
rect 567242 989551 660886 989579
rect 567242 989539 567248 989551
rect 660880 989539 660886 989551
rect 660938 989539 660944 989591
rect 216112 989465 216118 989517
rect 216170 989505 216176 989517
rect 235600 989505 235606 989517
rect 216170 989477 235606 989505
rect 216170 989465 216176 989477
rect 235600 989465 235606 989477
rect 235658 989465 235664 989517
rect 267952 989465 267958 989517
rect 268010 989505 268016 989517
rect 300496 989505 300502 989517
rect 268010 989477 300502 989505
rect 268010 989465 268016 989477
rect 300496 989465 300502 989477
rect 300554 989465 300560 989517
rect 319600 989465 319606 989517
rect 319658 989505 319664 989517
rect 349168 989505 349174 989517
rect 319658 989477 349174 989505
rect 319658 989465 319664 989477
rect 349168 989465 349174 989477
rect 349226 989465 349232 989517
rect 351280 989465 351286 989517
rect 351338 989505 351344 989517
rect 649552 989505 649558 989517
rect 351338 989477 649558 989505
rect 351338 989465 351344 989477
rect 649552 989465 649558 989477
rect 649610 989465 649616 989517
rect 110320 989391 110326 989443
rect 110378 989431 110384 989443
rect 122032 989431 122038 989443
rect 110378 989403 122038 989431
rect 110378 989391 110384 989403
rect 122032 989391 122038 989403
rect 122090 989391 122096 989443
rect 270736 989391 270742 989443
rect 270794 989431 270800 989443
rect 284272 989431 284278 989443
rect 270794 989403 284278 989431
rect 270794 989391 270800 989403
rect 284272 989391 284278 989403
rect 284330 989391 284336 989443
rect 305296 989391 305302 989443
rect 305354 989431 305360 989443
rect 649648 989431 649654 989443
rect 305354 989403 649654 989431
rect 305354 989391 305360 989403
rect 649648 989391 649654 989403
rect 649706 989391 649712 989443
rect 73456 989317 73462 989369
rect 73514 989357 73520 989369
rect 92944 989357 92950 989369
rect 73514 989329 92950 989357
rect 73514 989317 73520 989329
rect 92944 989317 92950 989329
rect 93002 989317 93008 989369
rect 265168 989317 265174 989369
rect 265226 989357 265232 989369
rect 658000 989357 658006 989369
rect 265226 989329 658006 989357
rect 265226 989317 265232 989329
rect 658000 989317 658006 989329
rect 658058 989317 658064 989369
rect 45040 989243 45046 989295
rect 45098 989283 45104 989295
rect 108592 989283 108598 989295
rect 45098 989255 108598 989283
rect 45098 989243 45104 989255
rect 108592 989243 108598 989255
rect 108650 989243 108656 989295
rect 250480 989243 250486 989295
rect 250538 989283 250544 989295
rect 649744 989283 649750 989295
rect 250538 989255 649750 989283
rect 250538 989243 250544 989255
rect 649744 989243 649750 989255
rect 649802 989243 649808 989295
rect 152656 989169 152662 989221
rect 152714 989209 152720 989221
rect 154480 989209 154486 989221
rect 152714 989181 154486 989209
rect 152714 989169 152720 989181
rect 154480 989169 154486 989181
rect 154538 989169 154544 989221
rect 201616 988799 201622 988851
rect 201674 988839 201680 988851
rect 203152 988839 203158 988851
rect 201674 988811 203158 988839
rect 201674 988799 201680 988811
rect 203152 988799 203158 988811
rect 203210 988799 203216 988851
rect 329680 987763 329686 987815
rect 329738 987803 329744 987815
rect 650896 987803 650902 987815
rect 329738 987775 650902 987803
rect 329738 987763 329744 987775
rect 650896 987763 650902 987775
rect 650954 987763 650960 987815
rect 329776 987689 329782 987741
rect 329834 987729 329840 987741
rect 650992 987729 650998 987741
rect 329834 987701 650998 987729
rect 329834 987689 329840 987701
rect 650992 987689 650998 987701
rect 651050 987689 651056 987741
rect 44656 987615 44662 987667
rect 44714 987655 44720 987667
rect 364432 987655 364438 987667
rect 44714 987627 364438 987655
rect 44714 987615 44720 987627
rect 364432 987615 364438 987627
rect 364490 987615 364496 987667
rect 44560 987541 44566 987593
rect 44618 987581 44624 987593
rect 363472 987581 363478 987593
rect 44618 987553 363478 987581
rect 44618 987541 44624 987553
rect 363472 987541 363478 987553
rect 363530 987541 363536 987593
rect 44848 987467 44854 987519
rect 44906 987507 44912 987519
rect 363856 987507 363862 987519
rect 44906 987479 363862 987507
rect 44906 987467 44912 987479
rect 363856 987467 363862 987479
rect 363914 987467 363920 987519
rect 44752 987393 44758 987445
rect 44810 987433 44816 987445
rect 362896 987433 362902 987445
rect 44810 987405 362902 987433
rect 44810 987393 44816 987405
rect 362896 987393 362902 987405
rect 362954 987393 362960 987445
rect 417520 987393 417526 987445
rect 417578 987433 417584 987445
rect 649456 987433 649462 987445
rect 417578 987405 649462 987433
rect 417578 987393 417584 987405
rect 649456 987393 649462 987405
rect 649514 987393 649520 987445
rect 321616 987319 321622 987371
rect 321674 987359 321680 987371
rect 652240 987359 652246 987371
rect 321674 987331 652246 987359
rect 321674 987319 321680 987331
rect 652240 987319 652246 987331
rect 652298 987319 652304 987371
rect 317200 987245 317206 987297
rect 317258 987285 317264 987297
rect 652432 987285 652438 987297
rect 317258 987257 652438 987285
rect 317258 987245 317264 987257
rect 652432 987245 652438 987257
rect 652490 987245 652496 987297
rect 268048 987171 268054 987223
rect 268106 987211 268112 987223
rect 658096 987211 658102 987223
rect 268106 987183 658102 987211
rect 268106 987171 268112 987183
rect 658096 987171 658102 987183
rect 658154 987171 658160 987223
rect 45136 987097 45142 987149
rect 45194 987137 45200 987149
rect 431248 987137 431254 987149
rect 45194 987109 431254 987137
rect 45194 987097 45200 987109
rect 431248 987097 431254 987109
rect 431306 987097 431312 987149
rect 44944 987023 44950 987075
rect 45002 987063 45008 987075
rect 430192 987063 430198 987075
rect 45002 987035 430198 987063
rect 45002 987023 45008 987035
rect 430192 987023 430198 987035
rect 430250 987023 430256 987075
rect 495280 987023 495286 987075
rect 495338 987063 495344 987075
rect 649360 987063 649366 987075
rect 495338 987035 649366 987063
rect 495338 987023 495344 987035
rect 649360 987023 649366 987035
rect 649418 987023 649424 987075
rect 216592 986949 216598 987001
rect 216650 986989 216656 987001
rect 658192 986989 658198 987001
rect 216650 986961 658198 986989
rect 216650 986949 216656 986961
rect 658192 986949 658198 986961
rect 658250 986949 658256 987001
rect 213136 986875 213142 986927
rect 213194 986915 213200 986927
rect 658384 986915 658390 986927
rect 213194 986887 658390 986915
rect 213194 986875 213200 986887
rect 658384 986875 658390 986887
rect 658442 986875 658448 986927
rect 198640 986801 198646 986853
rect 198698 986841 198704 986853
rect 649840 986841 649846 986853
rect 198698 986813 649846 986841
rect 198698 986801 198704 986813
rect 649840 986801 649846 986813
rect 649898 986801 649904 986853
rect 45232 986727 45238 986779
rect 45290 986767 45296 986779
rect 507280 986767 507286 986779
rect 45290 986739 507286 986767
rect 45290 986727 45296 986739
rect 507280 986727 507286 986739
rect 507338 986727 507344 986779
rect 45328 986653 45334 986705
rect 45386 986693 45392 986705
rect 508432 986693 508438 986705
rect 45386 986665 508438 986693
rect 45386 986653 45392 986665
rect 508432 986653 508438 986665
rect 508490 986653 508496 986705
rect 571600 986653 571606 986705
rect 571658 986693 571664 986705
rect 653776 986693 653782 986705
rect 571658 986665 653782 986693
rect 571658 986653 571664 986665
rect 653776 986653 653782 986665
rect 653834 986653 653840 986705
rect 164176 986579 164182 986631
rect 164234 986619 164240 986631
rect 655120 986619 655126 986631
rect 164234 986591 655126 986619
rect 164234 986579 164240 986591
rect 655120 986579 655126 986591
rect 655178 986579 655184 986631
rect 146608 986505 146614 986557
rect 146666 986545 146672 986557
rect 649936 986545 649942 986557
rect 146666 986517 649942 986545
rect 146666 986505 146672 986517
rect 649936 986505 649942 986517
rect 649994 986505 650000 986557
rect 62032 986431 62038 986483
rect 62090 986471 62096 986483
rect 112336 986471 112342 986483
rect 62090 986443 112342 986471
rect 62090 986431 62096 986443
rect 112336 986431 112342 986443
rect 112394 986471 112400 986483
rect 669616 986471 669622 986483
rect 112394 986443 669622 986471
rect 112394 986431 112400 986443
rect 669616 986431 669622 986443
rect 669674 986431 669680 986483
rect 62128 986357 62134 986409
rect 62186 986397 62192 986409
rect 112432 986397 112438 986409
rect 62186 986369 112438 986397
rect 62186 986357 62192 986369
rect 112432 986357 112438 986369
rect 112490 986397 112496 986409
rect 669808 986397 669814 986409
rect 112490 986369 669814 986397
rect 112490 986357 112496 986369
rect 669808 986357 669814 986369
rect 669866 986357 669872 986409
rect 565456 985025 565462 985077
rect 565514 985065 565520 985077
rect 566032 985065 566038 985077
rect 565514 985037 566038 985065
rect 565514 985025 565520 985037
rect 566032 985025 566038 985037
rect 566090 985065 566096 985077
rect 669712 985065 669718 985077
rect 566090 985037 669718 985065
rect 566090 985025 566096 985037
rect 669712 985025 669718 985037
rect 669770 985025 669776 985077
rect 565840 984951 565846 985003
rect 565898 984991 565904 985003
rect 566320 984991 566326 985003
rect 565898 984963 566326 984991
rect 565898 984951 565904 984963
rect 566320 984951 566326 984963
rect 566378 984991 566384 985003
rect 669904 984991 669910 985003
rect 566378 984963 669910 984991
rect 566378 984951 566384 984963
rect 669904 984951 669910 984963
rect 669962 984951 669968 985003
rect 164272 983693 164278 983745
rect 164330 983733 164336 983745
rect 660976 983733 660982 983745
rect 164330 983705 660982 983733
rect 164330 983693 164336 983705
rect 660976 983693 660982 983705
rect 661034 983693 661040 983745
rect 61936 983619 61942 983671
rect 61994 983659 62000 983671
rect 566320 983659 566326 983671
rect 61994 983631 566326 983659
rect 61994 983619 62000 983631
rect 566320 983619 566326 983631
rect 566378 983619 566384 983671
rect 61840 983545 61846 983597
rect 61898 983585 61904 983597
rect 565456 983585 565462 983597
rect 61898 983557 565462 983585
rect 61898 983545 61904 983557
rect 565456 983545 565462 983557
rect 565514 983545 565520 983597
rect 94864 983471 94870 983523
rect 94922 983511 94928 983523
rect 650032 983511 650038 983523
rect 94922 983483 650038 983511
rect 94922 983471 94928 983483
rect 650032 983471 650038 983483
rect 650090 983471 650096 983523
rect 65104 983397 65110 983449
rect 65162 983437 65168 983449
rect 652624 983437 652630 983449
rect 65162 983409 652630 983437
rect 65162 983397 65168 983409
rect 652624 983397 652630 983409
rect 652682 983397 652688 983449
rect 63376 983323 63382 983375
rect 63434 983363 63440 983375
rect 652912 983363 652918 983375
rect 63434 983335 652918 983363
rect 63434 983323 63440 983335
rect 652912 983323 652918 983335
rect 652970 983323 652976 983375
rect 63184 983249 63190 983301
rect 63242 983289 63248 983301
rect 652528 983289 652534 983301
rect 63242 983261 652534 983289
rect 63242 983249 63248 983261
rect 652528 983249 652534 983261
rect 652586 983249 652592 983301
rect 62896 983175 62902 983227
rect 62954 983215 62960 983227
rect 652816 983215 652822 983227
rect 62954 983187 652822 983215
rect 62954 983175 62960 983187
rect 652816 983175 652822 983187
rect 652874 983175 652880 983227
rect 63088 983101 63094 983153
rect 63146 983141 63152 983153
rect 653008 983141 653014 983153
rect 63146 983113 653014 983141
rect 63146 983101 63152 983113
rect 653008 983101 653014 983113
rect 653066 983101 653072 983153
rect 60976 983027 60982 983079
rect 61034 983067 61040 983079
rect 655408 983067 655414 983079
rect 61034 983039 655414 983067
rect 61034 983027 61040 983039
rect 655408 983027 655414 983039
rect 655466 983027 655472 983079
rect 63280 982953 63286 983005
rect 63338 982993 63344 983005
rect 655312 982993 655318 983005
rect 63338 982965 655318 982993
rect 63338 982953 63344 982965
rect 655312 982953 655318 982965
rect 655370 982953 655376 983005
rect 57616 982879 57622 982931
rect 57674 982919 57680 982931
rect 652720 982919 652726 982931
rect 57674 982891 652726 982919
rect 57674 982879 57680 982891
rect 652720 982879 652726 982891
rect 652778 982879 652784 982931
rect 48976 982805 48982 982857
rect 49034 982845 49040 982857
rect 652336 982845 652342 982857
rect 49034 982817 652342 982845
rect 49034 982805 49040 982817
rect 652336 982805 652342 982817
rect 652394 982805 652400 982857
rect 58192 979253 58198 979305
rect 58250 979293 58256 979305
rect 63184 979293 63190 979305
rect 58250 979265 63190 979293
rect 58250 979253 58256 979265
rect 63184 979253 63190 979265
rect 63242 979253 63248 979305
rect 55408 979179 55414 979231
rect 55466 979219 55472 979231
rect 60976 979219 60982 979231
rect 55466 979191 60982 979219
rect 55466 979179 55472 979191
rect 60976 979179 60982 979191
rect 61034 979179 61040 979231
rect 52048 977699 52054 977751
rect 52106 977739 52112 977751
rect 63088 977739 63094 977751
rect 52106 977711 63094 977739
rect 52106 977699 52112 977711
rect 63088 977699 63094 977711
rect 63146 977699 63152 977751
rect 58864 976441 58870 976493
rect 58922 976481 58928 976493
rect 63280 976481 63286 976493
rect 58922 976453 63286 976481
rect 58922 976441 58928 976453
rect 63280 976441 63286 976453
rect 63338 976441 63344 976493
rect 58960 976367 58966 976419
rect 59018 976407 59024 976419
rect 65104 976407 65110 976419
rect 59018 976379 65110 976407
rect 59018 976367 59024 976379
rect 65104 976367 65110 976379
rect 65162 976367 65168 976419
rect 51952 974887 51958 974939
rect 52010 974927 52016 974939
rect 62896 974927 62902 974939
rect 52010 974899 62902 974927
rect 52010 974887 52016 974899
rect 62896 974887 62902 974899
rect 62954 974887 62960 974939
rect 56272 973555 56278 973607
rect 56330 973595 56336 973607
rect 58192 973595 58198 973607
rect 56330 973567 58198 973595
rect 56330 973555 56336 973567
rect 58192 973555 58198 973567
rect 58250 973555 58256 973607
rect 51856 973481 51862 973533
rect 51914 973521 51920 973533
rect 58960 973521 58966 973533
rect 51914 973493 58966 973521
rect 51914 973481 51920 973493
rect 58960 973481 58966 973493
rect 59018 973481 59024 973533
rect 63376 973521 63382 973533
rect 60514 973493 63382 973521
rect 56080 973407 56086 973459
rect 56138 973447 56144 973459
rect 60514 973447 60542 973493
rect 63376 973481 63382 973493
rect 63434 973481 63440 973533
rect 56138 973419 60542 973447
rect 56138 973407 56144 973419
rect 45616 972001 45622 972053
rect 45674 972041 45680 972053
rect 48880 972041 48886 972053
rect 45674 972013 48886 972041
rect 45674 972001 45680 972013
rect 48880 972001 48886 972013
rect 48938 972001 48944 972053
rect 42352 970669 42358 970721
rect 42410 970709 42416 970721
rect 59536 970709 59542 970721
rect 42410 970681 59542 970709
rect 42410 970669 42416 970681
rect 59536 970669 59542 970681
rect 59594 970669 59600 970721
rect 52048 970635 52054 970647
rect 46114 970607 52054 970635
rect 44368 970521 44374 970573
rect 44426 970561 44432 970573
rect 46114 970561 46142 970607
rect 52048 970595 52054 970607
rect 52106 970595 52112 970647
rect 44426 970533 46142 970561
rect 44426 970521 44432 970533
rect 48976 969189 48982 969241
rect 49034 969229 49040 969241
rect 57520 969229 57526 969241
rect 49034 969201 57526 969229
rect 49034 969189 49040 969201
rect 57520 969189 57526 969201
rect 57578 969189 57584 969241
rect 50320 969115 50326 969167
rect 50378 969155 50384 969167
rect 58864 969155 58870 969167
rect 50378 969127 58870 969155
rect 50378 969115 50384 969127
rect 58864 969115 58870 969127
rect 58922 969115 58928 969167
rect 46672 968449 46678 968501
rect 46730 968489 46736 968501
rect 51952 968489 51958 968501
rect 46730 968461 51958 968489
rect 46730 968449 46736 968461
rect 51952 968449 51958 968461
rect 52010 968449 52016 968501
rect 45520 967709 45526 967761
rect 45578 967749 45584 967761
rect 51856 967749 51862 967761
rect 45578 967721 51862 967749
rect 45578 967709 45584 967721
rect 51856 967709 51862 967721
rect 51914 967709 51920 967761
rect 42160 967265 42166 967317
rect 42218 967305 42224 967317
rect 42352 967305 42358 967317
rect 42218 967277 42358 967305
rect 42218 967265 42224 967277
rect 42352 967265 42358 967277
rect 42410 967265 42416 967317
rect 44272 966081 44278 966133
rect 44330 966121 44336 966133
rect 46672 966121 46678 966133
rect 44330 966093 46678 966121
rect 44330 966081 44336 966093
rect 46672 966081 46678 966093
rect 46730 966081 46736 966133
rect 46000 964971 46006 965023
rect 46058 965011 46064 965023
rect 55408 965011 55414 965023
rect 46058 964983 55414 965011
rect 46058 964971 46064 964983
rect 55408 964971 55414 964983
rect 55466 964971 55472 965023
rect 51856 964897 51862 964949
rect 51914 964937 51920 964949
rect 56272 964937 56278 964949
rect 51914 964909 56278 964937
rect 51914 964897 51920 964909
rect 56272 964897 56278 964909
rect 56330 964897 56336 964949
rect 48976 964863 48982 964875
rect 46114 964835 48982 964863
rect 45712 964749 45718 964801
rect 45770 964789 45776 964801
rect 46114 964789 46142 964835
rect 48976 964823 48982 964835
rect 49034 964823 49040 964875
rect 52432 964823 52438 964875
rect 52490 964863 52496 964875
rect 56080 964863 56086 964875
rect 52490 964835 56086 964863
rect 52490 964823 52496 964835
rect 56080 964823 56086 964835
rect 56138 964823 56144 964875
rect 45770 964761 46142 964789
rect 45770 964749 45776 964761
rect 47536 961937 47542 961989
rect 47594 961977 47600 961989
rect 59536 961977 59542 961989
rect 47594 961949 59542 961977
rect 47594 961937 47600 961949
rect 59536 961937 59542 961949
rect 59594 961937 59600 961989
rect 674704 961271 674710 961323
rect 674762 961311 674768 961323
rect 675376 961311 675382 961323
rect 674762 961283 675382 961311
rect 674762 961271 674768 961283
rect 675376 961271 675382 961283
rect 675434 961271 675440 961323
rect 655600 959125 655606 959177
rect 655658 959165 655664 959177
rect 674800 959165 674806 959177
rect 655658 959137 674806 959165
rect 655658 959125 655664 959137
rect 674800 959125 674806 959137
rect 674858 959125 674864 959177
rect 45904 959051 45910 959103
rect 45962 959091 45968 959103
rect 50320 959091 50326 959103
rect 45962 959063 50326 959091
rect 45962 959051 45968 959063
rect 50320 959051 50326 959063
rect 50378 959051 50384 959103
rect 674800 955425 674806 955477
rect 674858 955465 674864 955477
rect 675376 955465 675382 955477
rect 674858 955437 675382 955465
rect 674858 955425 674864 955437
rect 675376 955425 675382 955437
rect 675434 955425 675440 955477
rect 48976 953279 48982 953331
rect 49034 953319 49040 953331
rect 52432 953319 52438 953331
rect 49034 953291 52438 953319
rect 49034 953279 49040 953291
rect 52432 953279 52438 953291
rect 52490 953279 52496 953331
rect 47440 951873 47446 951925
rect 47498 951913 47504 951925
rect 51760 951913 51766 951925
rect 47498 951885 51766 951913
rect 47498 951873 47504 951885
rect 51760 951873 51766 951885
rect 51818 951873 51824 951925
rect 38800 950393 38806 950445
rect 38858 950433 38864 950445
rect 42352 950433 42358 950445
rect 38858 950405 42358 950433
rect 38858 950393 38864 950405
rect 42352 950393 42358 950405
rect 42410 950393 42416 950445
rect 34480 947507 34486 947559
rect 34538 947547 34544 947559
rect 59536 947547 59542 947559
rect 34538 947519 59542 947547
rect 34538 947507 34544 947519
rect 59536 947507 59542 947519
rect 59594 947507 59600 947559
rect 44464 945805 44470 945857
rect 44522 945845 44528 945857
rect 48976 945845 48982 945857
rect 44522 945817 48982 945845
rect 44522 945805 44528 945817
rect 48976 945805 48982 945817
rect 49034 945805 49040 945857
rect 41776 943807 41782 943859
rect 41834 943847 41840 943859
rect 47536 943847 47542 943859
rect 41834 943819 47542 943847
rect 41834 943807 41840 943819
rect 47536 943807 47542 943819
rect 47594 943807 47600 943859
rect 41584 943585 41590 943637
rect 41642 943625 41648 943637
rect 45040 943625 45046 943637
rect 41642 943597 45046 943625
rect 41642 943585 41648 943597
rect 45040 943585 45046 943597
rect 45098 943585 45104 943637
rect 40240 941735 40246 941787
rect 40298 941775 40304 941787
rect 62128 941775 62134 941787
rect 40298 941747 62134 941775
rect 40298 941735 40304 941747
rect 62128 941735 62134 941747
rect 62186 941735 62192 941787
rect 660880 939737 660886 939789
rect 660938 939777 660944 939789
rect 676048 939777 676054 939789
rect 660938 939749 676054 939777
rect 660938 939737 660944 939749
rect 676048 939737 676054 939749
rect 676106 939737 676112 939789
rect 655696 939367 655702 939419
rect 655754 939407 655760 939419
rect 676240 939407 676246 939419
rect 655754 939379 676246 939407
rect 655754 939367 655760 939379
rect 676240 939367 676246 939379
rect 676298 939367 676304 939419
rect 655504 939219 655510 939271
rect 655562 939259 655568 939271
rect 676144 939259 676150 939271
rect 655562 939231 676150 939259
rect 655562 939219 655568 939231
rect 676144 939219 676150 939231
rect 676202 939219 676208 939271
rect 670768 939145 670774 939197
rect 670826 939185 670832 939197
rect 676048 939185 676054 939197
rect 670826 939157 676054 939185
rect 670826 939145 670832 939157
rect 676048 939145 676054 939157
rect 676106 939145 676112 939197
rect 655216 939071 655222 939123
rect 655274 939111 655280 939123
rect 676336 939111 676342 939123
rect 655274 939083 676342 939111
rect 655274 939071 655280 939083
rect 676336 939071 676342 939083
rect 676394 939071 676400 939123
rect 41584 938923 41590 938975
rect 41642 938963 41648 938975
rect 62032 938963 62038 938975
rect 41642 938935 62038 938963
rect 41642 938923 41648 938935
rect 62032 938923 62038 938935
rect 62090 938923 62096 938975
rect 39760 938849 39766 938901
rect 39818 938889 39824 938901
rect 59536 938889 59542 938901
rect 39818 938861 59542 938889
rect 39818 938849 39824 938861
rect 59536 938849 59542 938861
rect 59594 938849 59600 938901
rect 669904 938849 669910 938901
rect 669962 938889 669968 938901
rect 676240 938889 676246 938901
rect 669962 938861 676246 938889
rect 669962 938849 669968 938861
rect 676240 938849 676246 938861
rect 676298 938849 676304 938901
rect 670864 938035 670870 938087
rect 670922 938075 670928 938087
rect 676240 938075 676246 938087
rect 670922 938047 676246 938075
rect 670922 938035 670928 938047
rect 676240 938035 676246 938047
rect 676298 938035 676304 938087
rect 669712 937739 669718 937791
rect 669770 937779 669776 937791
rect 676048 937779 676054 937791
rect 669770 937751 676054 937779
rect 669770 937739 669776 937751
rect 676048 937739 676054 937751
rect 676106 937739 676112 937791
rect 670960 937147 670966 937199
rect 671018 937187 671024 937199
rect 676048 937187 676054 937199
rect 671018 937159 676054 937187
rect 671018 937147 671024 937159
rect 676048 937147 676054 937159
rect 676106 937147 676112 937199
rect 41584 932115 41590 932167
rect 41642 932155 41648 932167
rect 45040 932155 45046 932167
rect 41642 932127 45046 932155
rect 41642 932115 41648 932127
rect 45040 932115 45046 932127
rect 45098 932115 45104 932167
rect 660880 927379 660886 927431
rect 660938 927419 660944 927431
rect 679792 927419 679798 927431
rect 660938 927391 679798 927419
rect 660938 927379 660944 927391
rect 679792 927379 679798 927391
rect 679850 927379 679856 927431
rect 43120 921607 43126 921659
rect 43178 921647 43184 921659
rect 58576 921647 58582 921659
rect 43178 921619 58582 921647
rect 43178 921607 43184 921619
rect 58576 921607 58582 921619
rect 58634 921607 58640 921659
rect 656368 921607 656374 921659
rect 656426 921647 656432 921659
rect 666640 921647 666646 921659
rect 656426 921619 666646 921647
rect 656426 921607 656432 921619
rect 666640 921607 666646 921619
rect 666698 921607 666704 921659
rect 50416 910063 50422 910115
rect 50474 910103 50480 910115
rect 59536 910103 59542 910115
rect 50474 910075 59542 910103
rect 50474 910063 50480 910075
rect 59536 910063 59542 910075
rect 59594 910063 59600 910115
rect 654448 908731 654454 908783
rect 654506 908771 654512 908783
rect 661072 908771 661078 908783
rect 654506 908743 661078 908771
rect 654506 908731 654512 908743
rect 661072 908731 661078 908743
rect 661130 908731 661136 908783
rect 47632 895707 47638 895759
rect 47690 895747 47696 895759
rect 59536 895747 59542 895759
rect 47690 895719 59542 895747
rect 47690 895707 47696 895719
rect 59536 895707 59542 895719
rect 59594 895707 59600 895759
rect 654448 895707 654454 895759
rect 654506 895747 654512 895759
rect 672592 895747 672598 895759
rect 654506 895719 672598 895747
rect 654506 895707 654512 895719
rect 672592 895707 672598 895719
rect 672650 895707 672656 895759
rect 53392 884163 53398 884215
rect 53450 884203 53456 884215
rect 58000 884203 58006 884215
rect 53450 884175 58006 884203
rect 53450 884163 53456 884175
rect 58000 884163 58006 884175
rect 58058 884163 58064 884215
rect 673744 876541 673750 876593
rect 673802 876581 673808 876593
rect 675376 876581 675382 876593
rect 673802 876553 675382 876581
rect 673802 876541 673808 876553
rect 675376 876541 675382 876553
rect 675434 876541 675440 876593
rect 673552 873433 673558 873485
rect 673610 873473 673616 873485
rect 675376 873473 675382 873485
rect 673610 873445 675382 873473
rect 673610 873433 673616 873445
rect 675376 873433 675382 873445
rect 675434 873433 675440 873485
rect 673840 872619 673846 872671
rect 673898 872659 673904 872671
rect 675376 872659 675382 872671
rect 673898 872631 675382 872659
rect 673898 872619 673904 872631
rect 675376 872619 675382 872631
rect 675434 872619 675440 872671
rect 672784 872101 672790 872153
rect 672842 872141 672848 872153
rect 675472 872141 675478 872153
rect 672842 872113 675478 872141
rect 672842 872101 672848 872113
rect 675472 872101 675478 872113
rect 675530 872101 675536 872153
rect 656560 871139 656566 871191
rect 656618 871179 656624 871191
rect 674704 871179 674710 871191
rect 656618 871151 674710 871179
rect 656618 871139 656624 871151
rect 674704 871139 674710 871151
rect 674762 871139 674768 871191
rect 47536 869807 47542 869859
rect 47594 869847 47600 869859
rect 59536 869847 59542 869859
rect 47594 869819 59542 869847
rect 47594 869807 47600 869819
rect 59536 869807 59542 869819
rect 59594 869807 59600 869859
rect 654448 869289 654454 869341
rect 654506 869329 654512 869341
rect 663760 869329 663766 869341
rect 654506 869301 663766 869329
rect 654506 869289 654512 869301
rect 663760 869289 663766 869301
rect 663818 869289 663824 869341
rect 673456 869141 673462 869193
rect 673514 869181 673520 869193
rect 675472 869181 675478 869193
rect 673514 869153 675478 869181
rect 673514 869141 673520 869153
rect 675472 869141 675478 869153
rect 675530 869141 675536 869193
rect 674608 868327 674614 868379
rect 674666 868367 674672 868379
rect 675376 868367 675382 868379
rect 674666 868339 675382 868367
rect 674666 868327 674672 868339
rect 675376 868327 675382 868339
rect 675434 868327 675440 868379
rect 673360 867809 673366 867861
rect 673418 867849 673424 867861
rect 675376 867849 675382 867861
rect 673418 867821 675382 867849
rect 673418 867809 673424 867821
rect 675376 867809 675382 867821
rect 675434 867809 675440 867861
rect 669520 866921 669526 866973
rect 669578 866961 669584 866973
rect 675202 866961 675208 866973
rect 669578 866933 675208 866961
rect 669578 866921 669584 866933
rect 675202 866921 675208 866933
rect 675260 866921 675266 866973
rect 674224 866477 674230 866529
rect 674282 866517 674288 866529
rect 675376 866517 675382 866529
rect 674282 866489 675382 866517
rect 674282 866477 674288 866489
rect 675376 866477 675382 866489
rect 675434 866477 675440 866529
rect 674704 866255 674710 866307
rect 674762 866295 674768 866307
rect 675376 866295 675382 866307
rect 674762 866267 675382 866295
rect 674762 866255 674768 866267
rect 675376 866255 675382 866267
rect 675434 866255 675440 866307
rect 53200 858263 53206 858315
rect 53258 858303 53264 858315
rect 58384 858303 58390 858315
rect 53258 858275 58390 858303
rect 53258 858263 53264 858275
rect 58384 858263 58390 858275
rect 58442 858263 58448 858315
rect 654448 855377 654454 855429
rect 654506 855417 654512 855429
rect 672496 855417 672502 855429
rect 654506 855389 672502 855417
rect 654506 855377 654512 855389
rect 672496 855377 672502 855389
rect 672554 855377 672560 855429
rect 53296 843833 53302 843885
rect 53354 843873 53360 843885
rect 59536 843873 59542 843885
rect 53354 843845 59542 843873
rect 53354 843833 53360 843845
rect 59536 843833 59542 843845
rect 59594 843833 59600 843885
rect 654448 840947 654454 840999
rect 654506 840987 654512 840999
rect 666736 840987 666742 840999
rect 654506 840959 666742 840987
rect 654506 840947 654512 840959
rect 666736 840947 666742 840959
rect 666794 840947 666800 840999
rect 50512 832363 50518 832415
rect 50570 832403 50576 832415
rect 59536 832403 59542 832415
rect 50570 832375 59542 832403
rect 50570 832363 50576 832375
rect 59536 832363 59542 832375
rect 59594 832363 59600 832415
rect 654736 829477 654742 829529
rect 654794 829517 654800 829529
rect 661264 829517 661270 829529
rect 654794 829489 661270 829517
rect 654794 829477 654800 829489
rect 661264 829477 661270 829489
rect 661322 829477 661328 829529
rect 41680 823705 41686 823757
rect 41738 823745 41744 823757
rect 62032 823745 62038 823757
rect 41738 823717 62038 823745
rect 41738 823705 41744 823717
rect 62032 823705 62038 823717
rect 62090 823705 62096 823757
rect 39952 820819 39958 820871
rect 40010 820859 40016 820871
rect 41680 820859 41686 820871
rect 40010 820831 41686 820859
rect 40010 820819 40016 820831
rect 41680 820819 41686 820831
rect 41738 820819 41744 820871
rect 41584 819265 41590 819317
rect 41642 819305 41648 819317
rect 47632 819305 47638 819317
rect 41642 819277 47638 819305
rect 41642 819265 41648 819277
rect 47632 819265 47638 819277
rect 47690 819265 47696 819317
rect 41776 818525 41782 818577
rect 41834 818565 41840 818577
rect 53392 818565 53398 818577
rect 41834 818537 53398 818565
rect 41834 818525 41840 818537
rect 53392 818525 53398 818537
rect 53450 818525 53456 818577
rect 41776 818007 41782 818059
rect 41834 818047 41840 818059
rect 50416 818047 50422 818059
rect 41834 818019 50422 818047
rect 41834 818007 41840 818019
rect 50416 818007 50422 818019
rect 50474 818007 50480 818059
rect 50320 817933 50326 817985
rect 50378 817973 50384 817985
rect 59536 817973 59542 817985
rect 50378 817945 59542 817973
rect 50378 817933 50384 817945
rect 59536 817933 59542 817945
rect 59594 817933 59600 817985
rect 41776 816971 41782 817023
rect 41834 817011 41840 817023
rect 43216 817011 43222 817023
rect 41834 816983 43222 817011
rect 41834 816971 41840 816983
rect 43216 816971 43222 816983
rect 43274 816971 43280 817023
rect 655504 815047 655510 815099
rect 655562 815087 655568 815099
rect 661168 815087 661174 815099
rect 655562 815059 661174 815087
rect 655562 815047 655568 815059
rect 661168 815047 661174 815059
rect 661226 815047 661232 815099
rect 41584 812679 41590 812731
rect 41642 812719 41648 812731
rect 43024 812719 43030 812731
rect 41642 812691 43030 812719
rect 41642 812679 41648 812691
rect 43024 812679 43030 812691
rect 43082 812679 43088 812731
rect 41776 812235 41782 812287
rect 41834 812275 41840 812287
rect 42640 812275 42646 812287
rect 41834 812247 42646 812275
rect 41834 812235 41840 812247
rect 42640 812235 42646 812247
rect 42698 812235 42704 812287
rect 42064 810089 42070 810141
rect 42122 810129 42128 810141
rect 43024 810129 43030 810141
rect 42122 810101 43030 810129
rect 42122 810089 42128 810101
rect 43024 810089 43030 810101
rect 43082 810089 43088 810141
rect 41584 806759 41590 806811
rect 41642 806799 41648 806811
rect 42736 806799 42742 806811
rect 41642 806771 42742 806799
rect 41642 806759 41648 806771
rect 42736 806759 42742 806771
rect 42794 806759 42800 806811
rect 47632 806463 47638 806515
rect 47690 806503 47696 806515
rect 59536 806503 59542 806515
rect 47690 806475 59542 806503
rect 47690 806463 47696 806475
rect 59536 806463 59542 806475
rect 59594 806463 59600 806515
rect 41584 806389 41590 806441
rect 41642 806429 41648 806441
rect 45424 806429 45430 806441
rect 41642 806401 45430 806429
rect 41642 806389 41648 806401
rect 45424 806389 45430 806401
rect 45482 806389 45488 806441
rect 42352 802023 42358 802075
rect 42410 802063 42416 802075
rect 42832 802063 42838 802075
rect 42410 802035 42838 802063
rect 42410 802023 42416 802035
rect 42832 802023 42838 802035
rect 42890 802023 42896 802075
rect 654448 800617 654454 800669
rect 654506 800657 654512 800669
rect 670000 800657 670006 800669
rect 654506 800629 670006 800657
rect 654506 800617 654512 800629
rect 670000 800617 670006 800629
rect 670058 800617 670064 800669
rect 41488 800469 41494 800521
rect 41546 800509 41552 800521
rect 43504 800509 43510 800521
rect 41546 800481 43510 800509
rect 41546 800469 41552 800481
rect 43504 800469 43510 800481
rect 43562 800469 43568 800521
rect 42064 800247 42070 800299
rect 42122 800287 42128 800299
rect 43408 800287 43414 800299
rect 42122 800259 43414 800287
rect 42122 800247 42128 800259
rect 43408 800247 43414 800259
rect 43466 800247 43472 800299
rect 41872 800173 41878 800225
rect 41930 800173 41936 800225
rect 42160 800173 42166 800225
rect 42218 800213 42224 800225
rect 43312 800213 43318 800225
rect 42218 800185 43318 800213
rect 42218 800173 42224 800185
rect 43312 800173 43318 800185
rect 43370 800173 43376 800225
rect 41890 800003 41918 800173
rect 41872 799951 41878 800003
rect 41930 799951 41936 800003
rect 42160 798101 42166 798153
rect 42218 798141 42224 798153
rect 42640 798141 42646 798153
rect 42218 798113 42646 798141
rect 42218 798101 42224 798113
rect 42640 798101 42646 798113
rect 42698 798101 42704 798153
rect 653008 797805 653014 797857
rect 653066 797845 653072 797857
rect 653066 797817 656606 797845
rect 653066 797805 653072 797817
rect 656578 797771 656606 797817
rect 657904 797771 657910 797783
rect 656578 797743 657910 797771
rect 657904 797731 657910 797743
rect 657962 797731 657968 797783
rect 42064 797287 42070 797339
rect 42122 797327 42128 797339
rect 43120 797327 43126 797339
rect 42122 797299 43126 797327
rect 42122 797287 42128 797299
rect 43120 797287 43126 797299
rect 43178 797287 43184 797339
rect 43216 797287 43222 797339
rect 43274 797287 43280 797339
rect 43234 797117 43262 797287
rect 43216 797065 43222 797117
rect 43274 797065 43280 797117
rect 42160 794993 42166 795045
rect 42218 795033 42224 795045
rect 42736 795033 42742 795045
rect 42218 795005 42742 795033
rect 42218 794993 42224 795005
rect 42736 794993 42742 795005
rect 42794 794993 42800 795045
rect 42736 794845 42742 794897
rect 42794 794885 42800 794897
rect 43120 794885 43126 794897
rect 42794 794857 43126 794885
rect 42794 794845 42800 794857
rect 43120 794845 43126 794857
rect 43178 794845 43184 794897
rect 43120 794697 43126 794749
rect 43178 794737 43184 794749
rect 43408 794737 43414 794749
rect 43178 794709 43414 794737
rect 43178 794697 43184 794709
rect 43408 794697 43414 794709
rect 43466 794697 43472 794749
rect 42160 793809 42166 793861
rect 42218 793849 42224 793861
rect 42448 793849 42454 793861
rect 42218 793821 42454 793849
rect 42218 793809 42224 793821
rect 42448 793809 42454 793821
rect 42506 793809 42512 793861
rect 42160 793143 42166 793195
rect 42218 793183 42224 793195
rect 42832 793183 42838 793195
rect 42218 793155 42838 793183
rect 42218 793143 42224 793155
rect 42832 793143 42838 793155
rect 42890 793143 42896 793195
rect 42832 792995 42838 793047
rect 42890 793035 42896 793047
rect 43120 793035 43126 793047
rect 42890 793007 43126 793035
rect 42890 792995 42896 793007
rect 43120 792995 43126 793007
rect 43178 792995 43184 793047
rect 43120 792847 43126 792899
rect 43178 792887 43184 792899
rect 43504 792887 43510 792899
rect 43178 792859 43510 792887
rect 43178 792847 43184 792859
rect 43504 792847 43510 792859
rect 43562 792847 43568 792899
rect 47824 792033 47830 792085
rect 47882 792073 47888 792085
rect 59536 792073 59542 792085
rect 47882 792045 59542 792073
rect 47882 792033 47888 792045
rect 59536 792033 59542 792045
rect 59594 792033 59600 792085
rect 42160 790627 42166 790679
rect 42218 790667 42224 790679
rect 42736 790667 42742 790679
rect 42218 790639 42742 790667
rect 42218 790627 42224 790639
rect 42736 790627 42742 790639
rect 42794 790627 42800 790679
rect 42160 789887 42166 789939
rect 42218 789927 42224 789939
rect 43120 789927 43126 789939
rect 42218 789899 43126 789927
rect 42218 789887 42224 789899
rect 43120 789887 43126 789899
rect 43178 789887 43184 789939
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 42832 789483 42838 789495
rect 42218 789455 42838 789483
rect 42218 789443 42224 789455
rect 42832 789443 42838 789455
rect 42890 789443 42896 789495
rect 655600 789147 655606 789199
rect 655658 789187 655664 789199
rect 663856 789187 663862 789199
rect 655658 789159 663862 789187
rect 655658 789147 655664 789159
rect 663856 789147 663862 789159
rect 663914 789147 663920 789199
rect 652912 789073 652918 789125
rect 652970 789113 652976 789125
rect 655504 789113 655510 789125
rect 652970 789085 655510 789113
rect 652970 789073 652976 789085
rect 655504 789073 655510 789085
rect 655562 789073 655568 789125
rect 657904 789073 657910 789125
rect 657962 789113 657968 789125
rect 662320 789113 662326 789125
rect 657962 789085 662326 789113
rect 657962 789073 657968 789085
rect 662320 789073 662326 789085
rect 662378 789073 662384 789125
rect 42160 788777 42166 788829
rect 42218 788817 42224 788829
rect 42928 788817 42934 788829
rect 42218 788789 42934 788817
rect 42218 788777 42224 788789
rect 42928 788777 42934 788789
rect 42986 788777 42992 788829
rect 673264 787297 673270 787349
rect 673322 787337 673328 787349
rect 675472 787337 675478 787349
rect 673322 787309 675478 787337
rect 673322 787297 673328 787309
rect 675472 787297 675478 787309
rect 675530 787297 675536 787349
rect 42160 787001 42166 787053
rect 42218 787041 42224 787053
rect 43024 787041 43030 787053
rect 42218 787013 43030 787041
rect 42218 787001 42224 787013
rect 43024 787001 43030 787013
rect 43082 787001 43088 787053
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42736 786449 42742 786461
rect 42218 786421 42742 786449
rect 42218 786409 42224 786421
rect 42736 786409 42742 786421
rect 42794 786409 42800 786461
rect 42064 785743 42070 785795
rect 42122 785783 42128 785795
rect 42448 785783 42454 785795
rect 42122 785755 42454 785783
rect 42122 785743 42128 785755
rect 42448 785743 42454 785755
rect 42506 785743 42512 785795
rect 42160 784559 42166 784611
rect 42218 784599 42224 784611
rect 45520 784599 45526 784611
rect 42218 784571 45526 784599
rect 42218 784559 42224 784571
rect 45520 784559 45526 784571
rect 45578 784559 45584 784611
rect 42064 784263 42070 784315
rect 42122 784303 42128 784315
rect 45712 784303 45718 784315
rect 42122 784275 45718 784303
rect 42122 784263 42128 784275
rect 45712 784263 45718 784275
rect 45770 784263 45776 784315
rect 673168 784263 673174 784315
rect 673226 784303 673232 784315
rect 675472 784303 675478 784315
rect 673226 784275 675478 784303
rect 673226 784263 673232 784275
rect 675472 784263 675478 784275
rect 675530 784263 675536 784315
rect 662320 783671 662326 783723
rect 662378 783711 662384 783723
rect 666832 783711 666838 783723
rect 662378 783683 666838 783711
rect 662378 783671 662384 783683
rect 666832 783671 666838 783683
rect 666890 783671 666896 783723
rect 673072 783449 673078 783501
rect 673130 783489 673136 783501
rect 675376 783489 675382 783501
rect 673130 783461 675382 783489
rect 673130 783449 673136 783461
rect 675376 783449 675382 783461
rect 675434 783449 675440 783501
rect 661264 783301 661270 783353
rect 661322 783341 661328 783353
rect 674704 783341 674710 783353
rect 661322 783313 674710 783341
rect 661322 783301 661328 783313
rect 674704 783301 674710 783313
rect 674762 783301 674768 783353
rect 672976 782931 672982 782983
rect 673034 782971 673040 782983
rect 675472 782971 675478 782983
rect 673034 782943 675478 782971
rect 673034 782931 673040 782943
rect 675472 782931 675478 782943
rect 675530 782931 675536 782983
rect 673648 779897 673654 779949
rect 673706 779937 673712 779949
rect 675376 779937 675382 779949
rect 673706 779909 675382 779937
rect 673706 779897 673712 779909
rect 675376 779897 675382 779909
rect 675434 779897 675440 779949
rect 672880 778565 672886 778617
rect 672938 778605 672944 778617
rect 675376 778605 675382 778617
rect 672938 778577 675382 778605
rect 672938 778565 672944 778577
rect 675376 778565 675382 778577
rect 675434 778565 675440 778617
rect 53392 777603 53398 777655
rect 53450 777643 53456 777655
rect 59536 777643 59542 777655
rect 53450 777615 59542 777643
rect 53450 777603 53456 777615
rect 59536 777603 59542 777615
rect 59594 777603 59600 777655
rect 674704 777011 674710 777063
rect 674762 777051 674768 777063
rect 675376 777051 675382 777063
rect 674762 777023 675382 777051
rect 674762 777011 674768 777023
rect 675376 777011 675382 777023
rect 675434 777011 675440 777063
rect 41584 776049 41590 776101
rect 41642 776089 41648 776101
rect 53296 776089 53302 776101
rect 41642 776061 53302 776089
rect 41642 776049 41648 776061
rect 53296 776049 53302 776061
rect 53354 776049 53360 776101
rect 41776 775309 41782 775361
rect 41834 775349 41840 775361
rect 50512 775349 50518 775361
rect 41834 775321 50518 775349
rect 41834 775309 41840 775321
rect 50512 775309 50518 775321
rect 50570 775309 50576 775361
rect 41776 774791 41782 774843
rect 41834 774831 41840 774843
rect 53200 774831 53206 774843
rect 41834 774803 53206 774831
rect 41834 774791 41840 774803
rect 53200 774791 53206 774803
rect 53258 774791 53264 774843
rect 41584 774569 41590 774621
rect 41642 774609 41648 774621
rect 43216 774609 43222 774621
rect 41642 774581 43222 774609
rect 41642 774569 41648 774581
rect 43216 774569 43222 774581
rect 43274 774569 43280 774621
rect 41584 773607 41590 773659
rect 41642 773647 41648 773659
rect 43216 773647 43222 773659
rect 41642 773619 43222 773647
rect 41642 773607 41648 773619
rect 43216 773607 43222 773619
rect 43274 773607 43280 773659
rect 41776 769981 41782 770033
rect 41834 770021 41840 770033
rect 42928 770021 42934 770033
rect 41834 769993 42934 770021
rect 41834 769981 41840 769993
rect 42928 769981 42934 769993
rect 42986 769981 42992 770033
rect 41776 769463 41782 769515
rect 41834 769503 41840 769515
rect 43024 769503 43030 769515
rect 41834 769475 43030 769503
rect 41834 769463 41840 769475
rect 43024 769463 43030 769475
rect 43082 769463 43088 769515
rect 41872 766355 41878 766407
rect 41930 766395 41936 766407
rect 43120 766395 43126 766407
rect 41930 766367 43126 766395
rect 41930 766355 41936 766367
rect 43120 766355 43126 766367
rect 43178 766355 43184 766407
rect 41584 766059 41590 766111
rect 41642 766099 41648 766111
rect 42832 766099 42838 766111
rect 41642 766071 42838 766099
rect 41642 766059 41648 766071
rect 42832 766059 42838 766071
rect 42890 766059 42896 766111
rect 53200 766059 53206 766111
rect 53258 766099 53264 766111
rect 59536 766099 59542 766111
rect 53258 766071 59542 766099
rect 53258 766059 53264 766071
rect 59536 766059 59542 766071
rect 59594 766059 59600 766111
rect 41584 763247 41590 763299
rect 41642 763287 41648 763299
rect 45520 763287 45526 763299
rect 41642 763259 45526 763287
rect 41642 763247 41648 763259
rect 45520 763247 45526 763259
rect 45578 763247 45584 763299
rect 654448 763247 654454 763299
rect 654506 763287 654512 763299
rect 672400 763287 672406 763299
rect 654506 763259 672406 763287
rect 654506 763247 654512 763259
rect 672400 763247 672406 763259
rect 672458 763247 672464 763299
rect 661072 762877 661078 762929
rect 661130 762917 661136 762929
rect 676048 762917 676054 762929
rect 661130 762889 676054 762917
rect 661130 762877 661136 762889
rect 676048 762877 676054 762889
rect 676106 762877 676112 762929
rect 666640 762285 666646 762337
rect 666698 762325 666704 762337
rect 676048 762325 676054 762337
rect 666698 762297 676054 762325
rect 666698 762285 666704 762297
rect 676048 762285 676054 762297
rect 676106 762285 676112 762337
rect 672592 761989 672598 762041
rect 672650 762029 672656 762041
rect 676240 762029 676246 762041
rect 672650 762001 676246 762029
rect 672650 761989 672656 762001
rect 676240 761989 676246 762001
rect 676298 761989 676304 762041
rect 655504 761767 655510 761819
rect 655562 761807 655568 761819
rect 666352 761807 666358 761819
rect 655562 761779 666358 761807
rect 655562 761767 655568 761779
rect 666352 761767 666358 761779
rect 666410 761767 666416 761819
rect 670768 761545 670774 761597
rect 670826 761585 670832 761597
rect 676240 761585 676246 761597
rect 670826 761557 676246 761585
rect 670826 761545 670832 761557
rect 676240 761545 676246 761557
rect 676298 761545 676304 761597
rect 672592 760583 672598 760635
rect 672650 760623 672656 760635
rect 676240 760623 676246 760635
rect 672650 760595 676246 760623
rect 672650 760583 672656 760595
rect 676240 760583 676246 760595
rect 676298 760583 676304 760635
rect 670864 760287 670870 760339
rect 670922 760327 670928 760339
rect 676048 760327 676054 760339
rect 670922 760299 676054 760327
rect 670922 760287 670928 760299
rect 676048 760287 676054 760299
rect 676106 760287 676112 760339
rect 670672 759843 670678 759895
rect 670730 759883 670736 759895
rect 676048 759883 676054 759895
rect 670730 759855 676054 759883
rect 670730 759843 670736 759855
rect 676048 759843 676054 759855
rect 676106 759843 676112 759895
rect 670960 759325 670966 759377
rect 671018 759365 671024 759377
rect 676048 759365 676054 759377
rect 671018 759337 676054 759365
rect 671018 759325 671024 759337
rect 676048 759325 676054 759337
rect 676106 759325 676112 759377
rect 666352 758807 666358 758859
rect 666410 758847 666416 758859
rect 670768 758847 670774 758859
rect 666410 758819 670774 758847
rect 666410 758807 666416 758819
rect 670768 758807 670774 758819
rect 670826 758847 670832 758859
rect 676048 758847 676054 758859
rect 670826 758819 676054 758847
rect 670826 758807 670832 758819
rect 676048 758807 676054 758819
rect 676106 758807 676112 758859
rect 669712 757549 669718 757601
rect 669770 757589 669776 757601
rect 670864 757589 670870 757601
rect 669770 757561 670870 757589
rect 669770 757549 669776 757561
rect 670864 757549 670870 757561
rect 670922 757549 670928 757601
rect 42064 757475 42070 757527
rect 42122 757515 42128 757527
rect 42122 757487 42590 757515
rect 42122 757475 42128 757487
rect 40432 757401 40438 757453
rect 40490 757441 40496 757453
rect 42448 757441 42454 757453
rect 40490 757413 42454 757441
rect 40490 757401 40496 757413
rect 42448 757401 42454 757413
rect 42506 757401 42512 757453
rect 42562 757441 42590 757487
rect 43120 757475 43126 757527
rect 43178 757515 43184 757527
rect 43600 757515 43606 757527
rect 43178 757487 43606 757515
rect 43178 757475 43184 757487
rect 43600 757475 43606 757487
rect 43658 757475 43664 757527
rect 43696 757475 43702 757527
rect 43754 757515 43760 757527
rect 47536 757515 47542 757527
rect 43754 757487 47542 757515
rect 43754 757475 43760 757487
rect 47536 757475 47542 757487
rect 47594 757475 47600 757527
rect 669904 757475 669910 757527
rect 669962 757515 669968 757527
rect 670960 757515 670966 757527
rect 669962 757487 670966 757515
rect 669962 757475 669968 757487
rect 670960 757475 670966 757487
rect 671018 757475 671024 757527
rect 45808 757441 45814 757453
rect 42562 757413 45814 757441
rect 45808 757401 45814 757413
rect 45866 757401 45872 757453
rect 40336 757327 40342 757379
rect 40394 757367 40400 757379
rect 40394 757339 41498 757367
rect 40394 757327 40400 757339
rect 41470 756775 41498 757339
rect 41548 757327 41554 757379
rect 41606 757367 41612 757379
rect 43120 757367 43126 757379
rect 41606 757339 43126 757367
rect 41606 757327 41612 757339
rect 43120 757327 43126 757339
rect 43178 757327 43184 757379
rect 41680 757253 41686 757305
rect 41738 757293 41744 757305
rect 42832 757293 42838 757305
rect 41738 757265 42838 757293
rect 41738 757253 41744 757265
rect 42832 757253 42838 757265
rect 42890 757253 42896 757305
rect 43024 757253 43030 757305
rect 43082 757293 43088 757305
rect 43504 757293 43510 757305
rect 43082 757265 43510 757293
rect 43082 757253 43088 757265
rect 43504 757253 43510 757265
rect 43562 757253 43568 757305
rect 42160 757179 42166 757231
rect 42218 757219 42224 757231
rect 43408 757219 43414 757231
rect 42218 757191 43414 757219
rect 42218 757179 42224 757191
rect 43408 757179 43414 757191
rect 43466 757179 43472 757231
rect 41968 757105 41974 757157
rect 42026 757145 42032 757157
rect 43312 757145 43318 757157
rect 42026 757117 43318 757145
rect 42026 757105 42032 757117
rect 43312 757105 43318 757117
rect 43370 757105 43376 757157
rect 41776 757031 41782 757083
rect 41834 757071 41840 757083
rect 43024 757071 43030 757083
rect 41834 757043 43030 757071
rect 41834 757031 41840 757043
rect 43024 757031 43030 757043
rect 43082 757031 43088 757083
rect 41872 756957 41878 757009
rect 41930 756997 41936 757009
rect 42928 756997 42934 757009
rect 41930 756969 42934 756997
rect 41930 756957 41936 756969
rect 42928 756957 42934 756969
rect 42986 756957 42992 757009
rect 41872 756775 41878 756787
rect 41470 756747 41878 756775
rect 41872 756735 41878 756747
rect 41930 756735 41936 756787
rect 42160 755477 42166 755529
rect 42218 755517 42224 755529
rect 42448 755517 42454 755529
rect 42218 755489 42454 755517
rect 42218 755477 42224 755489
rect 42448 755477 42454 755489
rect 42506 755477 42512 755529
rect 673744 755403 673750 755455
rect 673802 755443 673808 755455
rect 676048 755443 676054 755455
rect 673802 755415 676054 755443
rect 673802 755403 673808 755415
rect 676048 755403 676054 755415
rect 676106 755403 676112 755455
rect 42160 755221 42166 755233
rect 42082 755193 42166 755221
rect 42082 754937 42110 755193
rect 42160 755181 42166 755193
rect 42218 755181 42224 755233
rect 673552 755033 673558 755085
rect 673610 755073 673616 755085
rect 676240 755073 676246 755085
rect 673610 755045 676246 755073
rect 673610 755033 673616 755045
rect 676240 755033 676246 755045
rect 676298 755033 676304 755085
rect 42064 754885 42070 754937
rect 42122 754885 42128 754937
rect 673840 754293 673846 754345
rect 673898 754333 673904 754345
rect 676048 754333 676054 754345
rect 673898 754305 676054 754333
rect 673898 754293 673904 754305
rect 676048 754293 676054 754305
rect 676106 754293 676112 754345
rect 42160 754071 42166 754123
rect 42218 754111 42224 754123
rect 43696 754111 43702 754123
rect 42218 754083 43702 754111
rect 42218 754071 42224 754083
rect 43696 754071 43702 754083
rect 43754 754071 43760 754123
rect 42064 753035 42070 753087
rect 42122 753075 42128 753087
rect 42832 753075 42838 753087
rect 42122 753047 42838 753075
rect 42122 753035 42128 753047
rect 42832 753035 42838 753047
rect 42890 753035 42896 753087
rect 42832 752887 42838 752939
rect 42890 752927 42896 752939
rect 43312 752927 43318 752939
rect 42890 752899 43318 752927
rect 42890 752887 42896 752899
rect 43312 752887 43318 752899
rect 43370 752887 43376 752939
rect 672784 752813 672790 752865
rect 672842 752853 672848 752865
rect 676048 752853 676054 752865
rect 672842 752825 676054 752853
rect 672842 752813 672848 752825
rect 676048 752813 676054 752825
rect 676106 752813 676112 752865
rect 673456 752369 673462 752421
rect 673514 752409 673520 752421
rect 676048 752409 676054 752421
rect 673514 752381 676054 752409
rect 673514 752369 673520 752381
rect 676048 752369 676054 752381
rect 676106 752369 676112 752421
rect 673360 751851 673366 751903
rect 673418 751891 673424 751903
rect 676048 751891 676054 751903
rect 673418 751863 676054 751891
rect 673418 751851 673424 751863
rect 676048 751851 676054 751863
rect 676106 751851 676112 751903
rect 42064 751777 42070 751829
rect 42122 751817 42128 751829
rect 42928 751817 42934 751829
rect 42122 751789 42934 751817
rect 42122 751777 42128 751789
rect 42928 751777 42934 751789
rect 42986 751777 42992 751829
rect 47728 751703 47734 751755
rect 47786 751743 47792 751755
rect 59536 751743 59542 751755
rect 47786 751715 59542 751743
rect 47786 751703 47792 751715
rect 59536 751703 59542 751715
rect 59594 751703 59600 751755
rect 652528 751703 652534 751755
rect 652586 751743 652592 751755
rect 655504 751743 655510 751755
rect 652586 751715 655510 751743
rect 652586 751703 652592 751715
rect 655504 751703 655510 751715
rect 655562 751703 655568 751755
rect 42928 751629 42934 751681
rect 42986 751669 42992 751681
rect 43408 751669 43414 751681
rect 42986 751641 43414 751669
rect 42986 751629 42992 751641
rect 43408 751629 43414 751641
rect 43466 751629 43472 751681
rect 42160 750593 42166 750645
rect 42218 750633 42224 750645
rect 43120 750633 43126 750645
rect 42218 750605 43126 750633
rect 42218 750593 42224 750605
rect 43120 750593 43126 750605
rect 43178 750593 43184 750645
rect 43120 750445 43126 750497
rect 43178 750485 43184 750497
rect 43504 750485 43510 750497
rect 43178 750457 43510 750485
rect 43178 750445 43184 750457
rect 43504 750445 43510 750457
rect 43562 750445 43568 750497
rect 42064 749927 42070 749979
rect 42122 749967 42128 749979
rect 43024 749967 43030 749979
rect 42122 749939 43030 749967
rect 42122 749927 42128 749939
rect 43024 749927 43030 749939
rect 43082 749927 43088 749979
rect 654448 748891 654454 748943
rect 654506 748931 654512 748943
rect 666640 748931 666646 748943
rect 654506 748903 666646 748931
rect 654506 748891 654512 748903
rect 666640 748891 666646 748903
rect 666698 748891 666704 748943
rect 658288 748817 658294 748869
rect 658346 748857 658352 748869
rect 679792 748857 679798 748869
rect 658346 748829 679798 748857
rect 658346 748817 658352 748829
rect 679792 748817 679798 748829
rect 679850 748817 679856 748869
rect 42160 746893 42166 746945
rect 42218 746933 42224 746945
rect 42832 746933 42838 746945
rect 42218 746905 42838 746933
rect 42218 746893 42224 746905
rect 42832 746893 42838 746905
rect 42890 746893 42896 746945
rect 42064 746819 42070 746871
rect 42122 746859 42128 746871
rect 42928 746859 42934 746871
rect 42122 746831 42934 746859
rect 42122 746819 42128 746831
rect 42928 746819 42934 746831
rect 42986 746819 42992 746871
rect 42064 746079 42070 746131
rect 42122 746119 42128 746131
rect 43600 746119 43606 746131
rect 42122 746091 43606 746119
rect 42122 746079 42128 746091
rect 43600 746079 43606 746091
rect 43658 746079 43664 746131
rect 42160 745635 42166 745687
rect 42218 745675 42224 745687
rect 43120 745675 43126 745687
rect 42218 745647 43126 745675
rect 42218 745635 42224 745647
rect 43120 745635 43126 745647
rect 43178 745635 43184 745687
rect 42160 743711 42166 743763
rect 42218 743751 42224 743763
rect 43024 743751 43030 743763
rect 42218 743723 43030 743751
rect 42218 743711 42224 743723
rect 43024 743711 43030 743723
rect 43082 743711 43088 743763
rect 42064 743193 42070 743245
rect 42122 743233 42128 743245
rect 42640 743233 42646 743245
rect 42122 743205 42646 743233
rect 42122 743193 42128 743205
rect 42640 743193 42646 743205
rect 42698 743193 42704 743245
rect 42160 742379 42166 742431
rect 42218 742419 42224 742431
rect 42736 742419 42742 742431
rect 42218 742391 42742 742419
rect 42218 742379 42224 742391
rect 42736 742379 42742 742391
rect 42794 742379 42800 742431
rect 42064 741343 42070 741395
rect 42122 741383 42128 741395
rect 45616 741383 45622 741395
rect 42122 741355 45622 741383
rect 42122 741343 42128 741355
rect 45616 741343 45622 741355
rect 45674 741343 45680 741395
rect 41680 741121 41686 741173
rect 41738 741161 41744 741173
rect 44272 741161 44278 741173
rect 41738 741133 44278 741161
rect 41738 741121 41744 741133
rect 44272 741121 44278 741133
rect 44330 741121 44336 741173
rect 47920 740159 47926 740211
rect 47978 740199 47984 740211
rect 58576 740199 58582 740211
rect 47978 740171 58582 740199
rect 47978 740159 47984 740171
rect 58576 740159 58582 740171
rect 58634 740159 58640 740211
rect 673840 739123 673846 739175
rect 673898 739163 673904 739175
rect 675472 739163 675478 739175
rect 673898 739135 675478 739163
rect 673898 739123 673904 739135
rect 675472 739123 675478 739135
rect 675530 739123 675536 739175
rect 655216 738679 655222 738731
rect 655274 738719 655280 738731
rect 674704 738719 674710 738731
rect 655274 738691 674710 738719
rect 655274 738679 655280 738691
rect 674704 738679 674710 738691
rect 674762 738679 674768 738731
rect 673456 738457 673462 738509
rect 673514 738497 673520 738509
rect 675376 738497 675382 738509
rect 673514 738469 675382 738497
rect 673514 738457 673520 738469
rect 675376 738457 675382 738469
rect 675434 738457 675440 738509
rect 673360 737865 673366 737917
rect 673418 737905 673424 737917
rect 675376 737905 675382 737917
rect 673418 737877 675382 737905
rect 673418 737865 673424 737877
rect 675376 737865 675382 737877
rect 675434 737865 675440 737917
rect 654448 735867 654454 735919
rect 654506 735907 654512 735919
rect 661264 735907 661270 735919
rect 654506 735879 661270 735907
rect 654506 735867 654512 735879
rect 661264 735867 661270 735879
rect 661322 735867 661328 735919
rect 673744 734905 673750 734957
rect 673802 734945 673808 734957
rect 675376 734945 675382 734957
rect 673802 734917 675382 734945
rect 673802 734905 673808 734917
rect 675376 734905 675382 734917
rect 675434 734905 675440 734957
rect 672784 733573 672790 733625
rect 672842 733613 672848 733625
rect 675472 733613 675478 733625
rect 672842 733585 675478 733613
rect 672842 733573 672848 733585
rect 675472 733573 675478 733585
rect 675530 733573 675536 733625
rect 41584 732833 41590 732885
rect 41642 732873 41648 732885
rect 47824 732873 47830 732885
rect 41642 732845 47830 732873
rect 41642 732833 41648 732845
rect 47824 732833 47830 732845
rect 47882 732833 47888 732885
rect 672688 732315 672694 732367
rect 672746 732355 672752 732367
rect 675472 732355 675478 732367
rect 672746 732327 675478 732355
rect 672746 732315 672752 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 41776 732093 41782 732145
rect 41834 732133 41840 732145
rect 53392 732133 53398 732145
rect 41834 732105 53398 732133
rect 41834 732093 41840 732105
rect 53392 732093 53398 732105
rect 53450 732093 53456 732145
rect 674704 732019 674710 732071
rect 674762 732059 674768 732071
rect 675376 732059 675382 732071
rect 674762 732031 675382 732059
rect 674762 732019 674768 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 655504 731871 655510 731923
rect 655562 731911 655568 731923
rect 658864 731911 658870 731923
rect 655562 731883 658870 731911
rect 655562 731871 655568 731883
rect 658864 731871 658870 731883
rect 658922 731871 658928 731923
rect 41584 731797 41590 731849
rect 41642 731837 41648 731849
rect 47632 731837 47638 731849
rect 41642 731809 47638 731837
rect 41642 731797 41648 731809
rect 47632 731797 47638 731809
rect 47690 731797 47696 731849
rect 41584 731353 41590 731405
rect 41642 731393 41648 731405
rect 43216 731393 43222 731405
rect 41642 731365 43222 731393
rect 41642 731353 41648 731365
rect 43216 731353 43222 731365
rect 43274 731353 43280 731405
rect 666832 731205 666838 731257
rect 666890 731245 666896 731257
rect 670096 731245 670102 731257
rect 666890 731217 670102 731245
rect 666890 731205 666896 731217
rect 670096 731205 670102 731217
rect 670154 731205 670160 731257
rect 674320 730465 674326 730517
rect 674378 730505 674384 730517
rect 675472 730505 675478 730517
rect 674378 730477 675478 730505
rect 674378 730465 674384 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 41584 730391 41590 730443
rect 41642 730431 41648 730443
rect 43216 730431 43222 730443
rect 41642 730403 43222 730431
rect 41642 730391 41648 730403
rect 43216 730391 43222 730403
rect 43274 730391 43280 730443
rect 674512 728615 674518 728667
rect 674570 728655 674576 728667
rect 675472 728655 675478 728667
rect 674570 728627 675478 728655
rect 674570 728615 674576 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 658864 728541 658870 728593
rect 658922 728581 658928 728593
rect 662128 728581 662134 728593
rect 658922 728553 662134 728581
rect 658922 728541 658928 728553
rect 662128 728541 662134 728553
rect 662186 728541 662192 728593
rect 50512 725803 50518 725855
rect 50570 725843 50576 725855
rect 59152 725843 59158 725855
rect 50570 725815 59158 725843
rect 50570 725803 50576 725815
rect 59152 725803 59158 725815
rect 59210 725803 59216 725855
rect 41776 723287 41782 723339
rect 41834 723327 41840 723339
rect 42928 723327 42934 723339
rect 41834 723299 42934 723327
rect 41834 723287 41840 723299
rect 42928 723287 42934 723299
rect 42986 723287 42992 723339
rect 41776 723139 41782 723191
rect 41834 723179 41840 723191
rect 43024 723179 43030 723191
rect 41834 723151 43030 723179
rect 41834 723139 41840 723151
rect 43024 723139 43030 723151
rect 43082 723139 43088 723191
rect 41584 722991 41590 723043
rect 41642 723031 41648 723043
rect 42832 723031 42838 723043
rect 41642 723003 42838 723031
rect 41642 722991 41648 723003
rect 42832 722991 42838 723003
rect 42890 722991 42896 723043
rect 672592 722917 672598 722969
rect 672650 722957 672656 722969
rect 679696 722957 679702 722969
rect 672650 722929 679702 722957
rect 672650 722917 672656 722929
rect 679696 722917 679702 722929
rect 679754 722917 679760 722969
rect 662128 720919 662134 720971
rect 662186 720959 662192 720971
rect 663376 720959 663382 720971
rect 662186 720931 663382 720959
rect 662186 720919 662192 720931
rect 663376 720919 663382 720931
rect 663434 720919 663440 720971
rect 41776 720179 41782 720231
rect 41834 720219 41840 720231
rect 45616 720219 45622 720231
rect 41834 720191 45622 720219
rect 41834 720179 41840 720191
rect 45616 720179 45622 720191
rect 45674 720179 45680 720231
rect 41584 720105 41590 720157
rect 41642 720145 41648 720157
rect 43120 720145 43126 720157
rect 41642 720117 43126 720145
rect 41642 720105 41648 720117
rect 43120 720105 43126 720117
rect 43178 720105 43184 720157
rect 672496 718033 672502 718085
rect 672554 718073 672560 718085
rect 676240 718073 676246 718085
rect 672554 718045 676246 718073
rect 672554 718033 672560 718045
rect 676240 718033 676246 718045
rect 676298 718033 676304 718085
rect 663760 717293 663766 717345
rect 663818 717333 663824 717345
rect 676048 717333 676054 717345
rect 663818 717305 676054 717333
rect 663818 717293 663824 717305
rect 676048 717293 676054 717305
rect 676106 717293 676112 717345
rect 663376 717145 663382 717197
rect 663434 717185 663440 717197
rect 670384 717185 670390 717197
rect 663434 717157 670390 717185
rect 663434 717145 663440 717157
rect 670384 717145 670390 717157
rect 670442 717145 670448 717197
rect 666736 716997 666742 717049
rect 666794 717037 666800 717049
rect 676240 717037 676246 717049
rect 666794 717009 676246 717037
rect 666794 716997 666800 717009
rect 676240 716997 676246 717009
rect 676298 716997 676304 717049
rect 652528 715665 652534 715717
rect 652586 715705 652592 715717
rect 670672 715705 670678 715717
rect 652586 715677 670678 715705
rect 652586 715665 652592 715677
rect 670672 715665 670678 715677
rect 670730 715665 670736 715717
rect 670672 715295 670678 715347
rect 670730 715335 670736 715347
rect 676048 715335 676054 715347
rect 670730 715307 676054 715335
rect 670730 715295 670736 715307
rect 676048 715295 676054 715307
rect 676106 715295 676112 715347
rect 670096 714851 670102 714903
rect 670154 714891 670160 714903
rect 670960 714891 670966 714903
rect 670154 714863 670966 714891
rect 670154 714851 670160 714863
rect 670960 714851 670966 714863
rect 671018 714891 671024 714903
rect 676048 714891 676054 714903
rect 671018 714863 676054 714891
rect 671018 714851 671024 714863
rect 676048 714851 676054 714863
rect 676106 714851 676112 714903
rect 43696 714333 43702 714385
rect 43754 714373 43760 714385
rect 50320 714373 50326 714385
rect 43754 714345 50326 714373
rect 43754 714333 43760 714345
rect 50320 714333 50326 714345
rect 50378 714333 50384 714385
rect 670768 714333 670774 714385
rect 670826 714373 670832 714385
rect 676048 714373 676054 714385
rect 670826 714345 676054 714373
rect 670826 714333 670832 714345
rect 676048 714333 676054 714345
rect 676106 714333 676112 714385
rect 47536 714259 47542 714311
rect 47594 714299 47600 714311
rect 59536 714299 59542 714311
rect 47594 714271 59542 714299
rect 47594 714259 47600 714271
rect 59536 714259 59542 714271
rect 59594 714259 59600 714311
rect 41488 714049 41494 714101
rect 41546 714077 41552 714101
rect 43600 714077 43606 714089
rect 41546 714049 43606 714077
rect 43600 714037 43606 714049
rect 43658 714037 43664 714089
rect 41872 713815 41878 713867
rect 41930 713815 41936 713867
rect 42064 713815 42070 713867
rect 42122 713855 42128 713867
rect 43408 713855 43414 713867
rect 42122 713827 43414 713855
rect 42122 713815 42128 713827
rect 43408 713815 43414 713827
rect 43466 713815 43472 713867
rect 41890 713571 41918 713815
rect 670384 713741 670390 713793
rect 670442 713781 670448 713793
rect 670864 713781 670870 713793
rect 670442 713753 670870 713781
rect 670442 713741 670448 713753
rect 670864 713741 670870 713753
rect 670922 713781 670928 713793
rect 676048 713781 676054 713793
rect 670922 713753 676054 713781
rect 670922 713741 670928 713753
rect 676048 713741 676054 713753
rect 676106 713741 676112 713793
rect 41872 713519 41878 713571
rect 41930 713519 41936 713571
rect 42448 713223 42454 713275
rect 42506 713263 42512 713275
rect 43504 713263 43510 713275
rect 42506 713235 43510 713263
rect 42506 713223 42512 713235
rect 43504 713223 43510 713235
rect 43562 713223 43568 713275
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 43696 710895 43702 710907
rect 42218 710867 43702 710895
rect 42218 710855 42224 710867
rect 43696 710855 43702 710867
rect 43754 710855 43760 710907
rect 673264 710411 673270 710463
rect 673322 710451 673328 710463
rect 676048 710451 676054 710463
rect 673322 710423 676054 710451
rect 673322 710411 673328 710423
rect 676048 710411 676054 710423
rect 676106 710411 676112 710463
rect 654448 710263 654454 710315
rect 654506 710303 654512 710315
rect 663760 710303 663766 710315
rect 654506 710275 663766 710303
rect 654506 710263 654512 710275
rect 663760 710263 663766 710275
rect 663818 710263 663824 710315
rect 673168 710041 673174 710093
rect 673226 710081 673232 710093
rect 676240 710081 676246 710093
rect 673226 710053 676246 710081
rect 673226 710041 673232 710053
rect 676240 710041 676246 710053
rect 676298 710041 676304 710093
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 42928 709933 42934 709945
rect 42218 709905 42934 709933
rect 42218 709893 42224 709905
rect 42928 709893 42934 709905
rect 42986 709893 42992 709945
rect 673072 709301 673078 709353
rect 673130 709341 673136 709353
rect 676048 709341 676054 709353
rect 673130 709313 676054 709341
rect 673130 709301 673136 709313
rect 676048 709301 676054 709313
rect 676106 709301 676112 709353
rect 42064 708561 42070 708613
rect 42122 708601 42128 708613
rect 43504 708601 43510 708613
rect 42122 708573 43510 708601
rect 42122 708561 42128 708573
rect 43504 708561 43510 708573
rect 43562 708561 43568 708613
rect 42160 708043 42166 708095
rect 42218 708083 42224 708095
rect 43024 708083 43030 708095
rect 42218 708055 43030 708083
rect 42218 708043 42224 708055
rect 43024 708043 43030 708055
rect 43082 708043 43088 708095
rect 672976 707969 672982 708021
rect 673034 708009 673040 708021
rect 676240 708009 676246 708021
rect 673034 707981 676246 708009
rect 673034 707969 673040 707981
rect 676240 707969 676246 707981
rect 676298 707969 676304 708021
rect 43024 707895 43030 707947
rect 43082 707935 43088 707947
rect 43408 707935 43414 707947
rect 43082 707907 43414 707935
rect 43082 707895 43088 707907
rect 43408 707895 43414 707907
rect 43466 707895 43472 707947
rect 42160 707377 42166 707429
rect 42218 707417 42224 707429
rect 43120 707417 43126 707429
rect 42218 707389 43126 707417
rect 42218 707377 42224 707389
rect 43120 707377 43126 707389
rect 43178 707377 43184 707429
rect 673648 707377 673654 707429
rect 673706 707417 673712 707429
rect 676048 707417 676054 707429
rect 673706 707389 676054 707417
rect 673706 707377 673712 707389
rect 676048 707377 676054 707389
rect 676106 707377 676112 707429
rect 672880 706859 672886 706911
rect 672938 706899 672944 706911
rect 676048 706899 676054 706911
rect 672938 706871 676054 706899
rect 672938 706859 672944 706871
rect 676048 706859 676054 706871
rect 676106 706859 676112 706911
rect 42160 706563 42166 706615
rect 42218 706603 42224 706615
rect 43024 706603 43030 706615
rect 42218 706575 43030 706603
rect 42218 706563 42224 706575
rect 43024 706563 43030 706575
rect 43082 706563 43088 706615
rect 43024 706415 43030 706467
rect 43082 706455 43088 706467
rect 43600 706455 43606 706467
rect 43082 706427 43606 706455
rect 43082 706415 43088 706427
rect 43600 706415 43606 706427
rect 43658 706415 43664 706467
rect 42256 704787 42262 704839
rect 42314 704827 42320 704839
rect 42448 704827 42454 704839
rect 42314 704799 42454 704827
rect 42314 704787 42320 704799
rect 42448 704787 42454 704799
rect 42506 704787 42512 704839
rect 42256 703677 42262 703729
rect 42314 703717 42320 703729
rect 42928 703717 42934 703729
rect 42314 703689 42934 703717
rect 42314 703677 42320 703689
rect 42928 703677 42934 703689
rect 42986 703677 42992 703729
rect 42064 703529 42070 703581
rect 42122 703569 42128 703581
rect 42832 703569 42838 703581
rect 42122 703541 42838 703569
rect 42122 703529 42128 703541
rect 42832 703529 42838 703541
rect 42890 703529 42896 703581
rect 658480 702715 658486 702767
rect 658538 702755 658544 702767
rect 679984 702755 679990 702767
rect 658538 702727 679990 702755
rect 658538 702715 658544 702727
rect 679984 702715 679990 702727
rect 680042 702715 680048 702767
rect 42160 702271 42166 702323
rect 42218 702311 42224 702323
rect 43024 702311 43030 702323
rect 42218 702283 43030 702311
rect 42218 702271 42224 702283
rect 43024 702271 43030 702283
rect 43082 702271 43088 702323
rect 42064 700347 42070 700399
rect 42122 700387 42128 700399
rect 43120 700387 43126 700399
rect 42122 700359 43126 700387
rect 42122 700347 42128 700359
rect 43120 700347 43126 700359
rect 43178 700347 43184 700399
rect 42160 700051 42166 700103
rect 42218 700091 42224 700103
rect 42832 700091 42838 700103
rect 42218 700063 42838 700091
rect 42218 700051 42224 700063
rect 42832 700051 42838 700063
rect 42890 700051 42896 700103
rect 47632 699829 47638 699881
rect 47690 699869 47696 699881
rect 59536 699869 59542 699881
rect 47690 699841 59542 699869
rect 47690 699829 47696 699841
rect 59536 699829 59542 699841
rect 59594 699829 59600 699881
rect 673168 699829 673174 699881
rect 673226 699869 673232 699881
rect 679696 699869 679702 699881
rect 673226 699841 679702 699869
rect 673226 699829 673232 699841
rect 679696 699829 679702 699841
rect 679754 699829 679760 699881
rect 42160 699385 42166 699437
rect 42218 699425 42224 699437
rect 42448 699425 42454 699437
rect 42218 699397 42454 699425
rect 42218 699385 42224 699397
rect 42448 699385 42454 699397
rect 42506 699385 42512 699437
rect 654448 696943 654454 696995
rect 654506 696983 654512 696995
rect 670096 696983 670102 696995
rect 654506 696955 670102 696983
rect 654506 696943 654512 696955
rect 670096 696943 670102 696955
rect 670154 696943 670160 696995
rect 41872 694649 41878 694701
rect 41930 694689 41936 694701
rect 46000 694689 46006 694701
rect 41930 694661 46006 694689
rect 41930 694649 41936 694661
rect 46000 694649 46006 694661
rect 46058 694649 46064 694701
rect 673648 693465 673654 693517
rect 673706 693505 673712 693517
rect 675472 693505 675478 693517
rect 673706 693477 675478 693505
rect 673706 693465 673712 693477
rect 675472 693465 675478 693477
rect 675530 693465 675536 693517
rect 673552 692873 673558 692925
rect 673610 692913 673616 692925
rect 675472 692913 675478 692925
rect 673610 692885 675478 692913
rect 673610 692873 673616 692885
rect 675472 692873 675478 692885
rect 675530 692873 675536 692925
rect 655216 692577 655222 692629
rect 655274 692617 655280 692629
rect 674704 692617 674710 692629
rect 655274 692589 674710 692617
rect 655274 692577 655280 692589
rect 674704 692577 674710 692589
rect 674762 692577 674768 692629
rect 672880 689765 672886 689817
rect 672938 689805 672944 689817
rect 675376 689805 675382 689817
rect 672938 689777 675382 689805
rect 672938 689765 672944 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 41776 689469 41782 689521
rect 41834 689509 41840 689521
rect 47920 689509 47926 689521
rect 41834 689481 47926 689509
rect 41834 689469 41840 689481
rect 47920 689469 47926 689481
rect 47978 689469 47984 689521
rect 673264 689099 673270 689151
rect 673322 689139 673328 689151
rect 675376 689139 675382 689151
rect 673322 689111 675382 689139
rect 673322 689099 673328 689111
rect 675376 689099 675382 689111
rect 675434 689099 675440 689151
rect 41776 688877 41782 688929
rect 41834 688917 41840 688929
rect 50512 688917 50518 688929
rect 41834 688889 50518 688917
rect 41834 688877 41840 688889
rect 50512 688877 50518 688889
rect 50570 688877 50576 688929
rect 41584 688581 41590 688633
rect 41642 688621 41648 688633
rect 47728 688621 47734 688633
rect 41642 688593 47734 688621
rect 41642 688581 41648 688593
rect 47728 688581 47734 688593
rect 47786 688581 47792 688633
rect 672976 688581 672982 688633
rect 673034 688621 673040 688633
rect 675472 688621 675478 688633
rect 673034 688593 675478 688621
rect 673034 688581 673040 688593
rect 675472 688581 675478 688593
rect 675530 688581 675536 688633
rect 50416 688359 50422 688411
rect 50474 688399 50480 688411
rect 59536 688399 59542 688411
rect 50474 688371 59542 688399
rect 50474 688359 50480 688371
rect 59536 688359 59542 688371
rect 59594 688359 59600 688411
rect 41584 688137 41590 688189
rect 41642 688177 41648 688189
rect 43216 688177 43222 688189
rect 41642 688149 43222 688177
rect 41642 688137 41648 688149
rect 43216 688137 43222 688149
rect 43274 688137 43280 688189
rect 41584 687175 41590 687227
rect 41642 687215 41648 687227
rect 43216 687215 43222 687227
rect 41642 687187 43222 687215
rect 41642 687175 41648 687187
rect 43216 687175 43222 687187
rect 43274 687175 43280 687227
rect 674704 687027 674710 687079
rect 674762 687067 674768 687079
rect 675472 687067 675478 687079
rect 674762 687039 675478 687067
rect 674762 687027 674768 687039
rect 675472 687027 675478 687039
rect 675530 687027 675536 687079
rect 41776 685917 41782 685969
rect 41834 685957 41840 685969
rect 45904 685957 45910 685969
rect 41834 685929 45910 685957
rect 41834 685917 41840 685929
rect 45904 685917 45910 685929
rect 45962 685917 45968 685969
rect 674224 685473 674230 685525
rect 674282 685513 674288 685525
rect 675472 685513 675478 685525
rect 674282 685485 675478 685513
rect 674282 685473 674288 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 674416 683623 674422 683675
rect 674474 683663 674480 683675
rect 675472 683663 675478 683675
rect 674474 683635 675478 683663
rect 674474 683623 674480 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 41584 682809 41590 682861
rect 41642 682849 41648 682861
rect 42736 682849 42742 682861
rect 41642 682821 42742 682849
rect 41642 682809 41648 682821
rect 42736 682809 42742 682821
rect 42794 682809 42800 682861
rect 654448 682587 654454 682639
rect 654506 682627 654512 682639
rect 666736 682627 666742 682639
rect 654506 682599 666742 682627
rect 654506 682587 654512 682599
rect 666736 682587 666742 682599
rect 666794 682587 666800 682639
rect 41584 680219 41590 680271
rect 41642 680259 41648 680271
rect 42928 680259 42934 680271
rect 41642 680231 42934 680259
rect 41642 680219 41648 680231
rect 42928 680219 42934 680231
rect 42986 680219 42992 680271
rect 41584 679183 41590 679235
rect 41642 679223 41648 679235
rect 42736 679223 42742 679235
rect 41642 679195 42742 679223
rect 41642 679183 41648 679195
rect 42736 679183 42742 679195
rect 42794 679183 42800 679235
rect 41680 678887 41686 678939
rect 41738 678927 41744 678939
rect 42448 678927 42454 678939
rect 41738 678899 42454 678927
rect 41738 678887 41744 678899
rect 42448 678887 42454 678899
rect 42506 678887 42512 678939
rect 42448 678739 42454 678791
rect 42506 678779 42512 678791
rect 42928 678779 42934 678791
rect 42506 678751 42934 678779
rect 42506 678739 42512 678751
rect 42928 678739 42934 678751
rect 42986 678739 42992 678791
rect 41776 678443 41782 678495
rect 41834 678483 41840 678495
rect 42832 678483 42838 678495
rect 41834 678455 42838 678483
rect 41834 678443 41840 678455
rect 42832 678443 42838 678455
rect 42890 678443 42896 678495
rect 41584 676963 41590 677015
rect 41642 677003 41648 677015
rect 43120 677003 43126 677015
rect 41642 676975 43126 677003
rect 41642 676963 41648 676975
rect 43120 676963 43126 676975
rect 43178 676963 43184 677015
rect 41776 676889 41782 676941
rect 41834 676929 41840 676941
rect 45904 676929 45910 676941
rect 41834 676901 45910 676929
rect 41834 676889 41840 676901
rect 45904 676889 45910 676901
rect 45962 676889 45968 676941
rect 53296 673929 53302 673981
rect 53354 673969 53360 673981
rect 59056 673969 59062 673981
rect 53354 673941 59062 673969
rect 53354 673929 53360 673941
rect 59056 673929 59062 673941
rect 59114 673929 59120 673981
rect 670000 672671 670006 672723
rect 670058 672711 670064 672723
rect 676048 672711 676054 672723
rect 670058 672683 676054 672711
rect 670058 672671 670064 672683
rect 676048 672671 676054 672683
rect 676106 672671 676112 672723
rect 661168 672301 661174 672353
rect 661226 672341 661232 672353
rect 676240 672341 676246 672353
rect 661226 672313 676246 672341
rect 661226 672301 661232 672313
rect 676240 672301 676246 672313
rect 676298 672301 676304 672353
rect 41968 671931 41974 671983
rect 42026 671971 42032 671983
rect 42928 671971 42934 671983
rect 42026 671943 42934 671971
rect 42026 671931 42032 671943
rect 42928 671931 42934 671943
rect 42986 671931 42992 671983
rect 663856 671561 663862 671613
rect 663914 671601 663920 671613
rect 676048 671601 676054 671613
rect 663914 671573 676054 671601
rect 663914 671561 663920 671573
rect 676048 671561 676054 671573
rect 676106 671561 676112 671613
rect 673168 671191 673174 671243
rect 673226 671231 673232 671243
rect 676048 671231 676054 671243
rect 673226 671203 676054 671231
rect 673226 671191 673232 671203
rect 676048 671191 676054 671203
rect 676106 671191 676112 671243
rect 43600 671043 43606 671095
rect 43658 671083 43664 671095
rect 53200 671083 53206 671095
rect 43658 671055 53206 671083
rect 43658 671043 43664 671055
rect 53200 671043 53206 671055
rect 53258 671043 53264 671095
rect 41392 670925 41398 670977
rect 41450 670965 41456 670977
rect 43504 670965 43510 670977
rect 41450 670937 43510 670965
rect 41450 670925 41456 670937
rect 43504 670925 43510 670937
rect 43562 670925 43568 670977
rect 41488 670851 41494 670903
rect 41546 670891 41552 670903
rect 43408 670891 43414 670903
rect 41546 670863 43414 670891
rect 41546 670851 41552 670863
rect 43408 670851 43414 670863
rect 43466 670851 43472 670903
rect 42736 670777 42742 670829
rect 42794 670817 42800 670829
rect 43312 670817 43318 670829
rect 42794 670789 43318 670817
rect 42794 670777 42800 670789
rect 43312 670777 43318 670789
rect 43370 670777 43376 670829
rect 41872 670599 41878 670651
rect 41930 670599 41936 670651
rect 42160 670599 42166 670651
rect 42218 670639 42224 670651
rect 42736 670639 42742 670651
rect 42218 670611 42742 670639
rect 42218 670599 42224 670611
rect 42736 670599 42742 670611
rect 42794 670599 42800 670651
rect 672304 670599 672310 670651
rect 672362 670639 672368 670651
rect 676048 670639 676054 670651
rect 672362 670611 676054 670639
rect 672362 670599 672368 670611
rect 676048 670599 676054 670611
rect 676106 670599 676112 670651
rect 41890 670355 41918 670599
rect 41872 670303 41878 670355
rect 41930 670303 41936 670355
rect 670960 670081 670966 670133
rect 671018 670121 671024 670133
rect 676048 670121 676054 670133
rect 671018 670093 676054 670121
rect 671018 670081 671024 670093
rect 676048 670081 676054 670093
rect 676106 670081 676112 670133
rect 667984 669563 667990 669615
rect 668042 669603 668048 669615
rect 676048 669603 676054 669615
rect 668042 669575 676054 669603
rect 668042 669563 668048 669575
rect 676048 669563 676054 669575
rect 676106 669563 676112 669615
rect 670864 669341 670870 669393
rect 670922 669381 670928 669393
rect 676240 669381 676246 669393
rect 670922 669353 676246 669381
rect 670922 669341 670928 669353
rect 676240 669341 676246 669353
rect 676298 669341 676304 669393
rect 42160 668379 42166 668431
rect 42218 668419 42224 668431
rect 43024 668419 43030 668431
rect 42218 668391 43030 668419
rect 42218 668379 42224 668391
rect 43024 668379 43030 668391
rect 43082 668379 43088 668431
rect 43024 668231 43030 668283
rect 43082 668271 43088 668283
rect 43312 668271 43318 668283
rect 43082 668243 43318 668271
rect 43082 668231 43088 668243
rect 43312 668231 43318 668243
rect 43370 668231 43376 668283
rect 674320 668083 674326 668135
rect 674378 668123 674384 668135
rect 676048 668123 676054 668135
rect 674378 668095 676054 668123
rect 674378 668083 674384 668095
rect 676048 668083 676054 668095
rect 676106 668083 676112 668135
rect 674512 668009 674518 668061
rect 674570 668049 674576 668061
rect 676240 668049 676246 668061
rect 674570 668021 676246 668049
rect 674570 668009 674576 668021
rect 676240 668009 676246 668021
rect 676298 668009 676304 668061
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 43600 667901 43606 667913
rect 42218 667873 43606 667901
rect 42218 667861 42224 667873
rect 43600 667861 43606 667873
rect 43658 667861 43664 667913
rect 42160 665345 42166 665397
rect 42218 665385 42224 665397
rect 42832 665385 42838 665397
rect 42218 665357 42838 665385
rect 42218 665345 42224 665357
rect 42832 665345 42838 665357
rect 42890 665345 42896 665397
rect 42160 664827 42166 664879
rect 42218 664867 42224 664879
rect 42928 664867 42934 664879
rect 42218 664839 42934 664867
rect 42218 664827 42224 664839
rect 42928 664827 42934 664839
rect 42986 664827 42992 664879
rect 42928 664679 42934 664731
rect 42986 664719 42992 664731
rect 43408 664719 43414 664731
rect 42986 664691 43414 664719
rect 42986 664679 42992 664691
rect 43408 664679 43414 664691
rect 43466 664679 43472 664731
rect 673840 664605 673846 664657
rect 673898 664645 673904 664657
rect 676048 664645 676054 664657
rect 673898 664617 676054 664645
rect 673898 664605 673904 664617
rect 676048 664605 676054 664617
rect 676106 664605 676112 664657
rect 673456 664309 673462 664361
rect 673514 664349 673520 664361
rect 676240 664349 676246 664361
rect 673514 664321 676246 664349
rect 673514 664309 673520 664321
rect 676240 664309 676246 664321
rect 676298 664309 676304 664361
rect 42064 663939 42070 663991
rect 42122 663979 42128 663991
rect 43120 663979 43126 663991
rect 42122 663951 43126 663979
rect 42122 663939 42128 663951
rect 43120 663939 43126 663951
rect 43178 663939 43184 663991
rect 672688 663865 672694 663917
rect 672746 663905 672752 663917
rect 676240 663905 676246 663917
rect 672746 663877 676246 663905
rect 672746 663865 672752 663877
rect 676240 663865 676246 663877
rect 676298 663865 676304 663917
rect 43120 663791 43126 663843
rect 43178 663831 43184 663843
rect 43504 663831 43510 663843
rect 43178 663803 43510 663831
rect 43178 663791 43184 663803
rect 43504 663791 43510 663803
rect 43562 663791 43568 663843
rect 673360 662607 673366 662659
rect 673418 662647 673424 662659
rect 676048 662647 676054 662659
rect 673418 662619 676054 662647
rect 673418 662607 673424 662619
rect 676048 662607 676054 662619
rect 676106 662607 676112 662659
rect 50320 662385 50326 662437
rect 50378 662425 50384 662437
rect 58096 662425 58102 662437
rect 50378 662397 58102 662425
rect 50378 662385 50384 662397
rect 58096 662385 58102 662397
rect 58154 662385 58160 662437
rect 655408 662311 655414 662363
rect 655466 662351 655472 662363
rect 659056 662351 659062 662363
rect 655466 662323 659062 662351
rect 655466 662311 655472 662323
rect 659056 662311 659062 662323
rect 659114 662311 659120 662363
rect 673744 662237 673750 662289
rect 673802 662277 673808 662289
rect 676048 662277 676054 662289
rect 673802 662249 676054 662277
rect 673802 662237 673808 662249
rect 676048 662237 676054 662249
rect 676106 662237 676112 662289
rect 672784 661645 672790 661697
rect 672842 661685 672848 661697
rect 676048 661685 676054 661697
rect 672842 661657 676054 661685
rect 672842 661645 672848 661657
rect 676048 661645 676054 661657
rect 676106 661645 676112 661697
rect 42064 661053 42070 661105
rect 42122 661093 42128 661105
rect 43024 661093 43030 661105
rect 42122 661065 43030 661093
rect 42122 661053 42128 661065
rect 43024 661053 43030 661065
rect 43082 661053 43088 661105
rect 42064 660387 42070 660439
rect 42122 660427 42128 660439
rect 42832 660427 42838 660439
rect 42122 660399 42838 660427
rect 42122 660387 42128 660399
rect 42832 660387 42838 660399
rect 42890 660387 42896 660439
rect 42160 659869 42166 659921
rect 42218 659909 42224 659921
rect 42736 659909 42742 659921
rect 42218 659881 42742 659909
rect 42218 659869 42224 659881
rect 42736 659869 42742 659881
rect 42794 659869 42800 659921
rect 42736 659721 42742 659773
rect 42794 659761 42800 659773
rect 42928 659761 42934 659773
rect 42794 659733 42934 659761
rect 42794 659721 42800 659733
rect 42928 659721 42934 659733
rect 42986 659721 42992 659773
rect 42928 659573 42934 659625
rect 42986 659613 42992 659625
rect 43120 659613 43126 659625
rect 42986 659585 43126 659613
rect 42986 659573 42992 659585
rect 43120 659573 43126 659585
rect 43178 659573 43184 659625
rect 655216 659499 655222 659551
rect 655274 659539 655280 659551
rect 679792 659539 679798 659551
rect 655274 659511 679798 659539
rect 655274 659499 655280 659511
rect 679792 659499 679798 659511
rect 679850 659499 679856 659551
rect 42064 659055 42070 659107
rect 42122 659095 42128 659107
rect 42928 659095 42934 659107
rect 42122 659067 42934 659095
rect 42122 659055 42128 659067
rect 42928 659055 42934 659067
rect 42986 659055 42992 659107
rect 42064 657205 42070 657257
rect 42122 657245 42128 657257
rect 42832 657245 42838 657257
rect 42122 657217 42838 657245
rect 42122 657205 42128 657217
rect 42832 657205 42838 657217
rect 42890 657205 42896 657257
rect 42160 656687 42166 656739
rect 42218 656727 42224 656739
rect 42928 656727 42934 656739
rect 42218 656699 42934 656727
rect 42218 656687 42224 656699
rect 42928 656687 42934 656699
rect 42986 656687 42992 656739
rect 654448 656687 654454 656739
rect 654506 656727 654512 656739
rect 661072 656727 661078 656739
rect 654506 656699 661078 656727
rect 654506 656687 654512 656699
rect 661072 656687 661078 656699
rect 661130 656687 661136 656739
rect 672496 656687 672502 656739
rect 672554 656727 672560 656739
rect 679888 656727 679894 656739
rect 672554 656699 679894 656727
rect 672554 656687 672560 656699
rect 679888 656687 679894 656699
rect 679946 656687 679952 656739
rect 42160 656169 42166 656221
rect 42218 656209 42224 656221
rect 43024 656209 43030 656221
rect 42218 656181 43030 656209
rect 42218 656169 42224 656181
rect 43024 656169 43030 656181
rect 43082 656169 43088 656221
rect 659056 653801 659062 653853
rect 659114 653841 659120 653853
rect 659114 653813 659534 653841
rect 659114 653801 659120 653813
rect 659506 653767 659534 653813
rect 665008 653767 665014 653779
rect 659506 653739 665014 653767
rect 665008 653727 665014 653739
rect 665066 653727 665072 653779
rect 673744 652099 673750 652151
rect 673802 652139 673808 652151
rect 675472 652139 675478 652151
rect 673802 652111 675478 652139
rect 673802 652099 673808 652111
rect 675472 652099 675478 652111
rect 675530 652099 675536 652151
rect 673072 649065 673078 649117
rect 673130 649105 673136 649117
rect 675472 649105 675478 649117
rect 673130 649077 675478 649105
rect 673130 649065 673136 649077
rect 675472 649065 675478 649077
rect 675530 649065 675536 649117
rect 673168 648251 673174 648303
rect 673226 648291 673232 648303
rect 675376 648291 675382 648303
rect 673226 648263 675382 648291
rect 673226 648251 673232 648263
rect 675376 648251 675382 648263
rect 675434 648251 675440 648303
rect 53200 648029 53206 648081
rect 53258 648069 53264 648081
rect 59536 648069 59542 648081
rect 53258 648041 59542 648069
rect 53258 648029 53264 648041
rect 59536 648029 59542 648041
rect 59594 648029 59600 648081
rect 673840 647881 673846 647933
rect 673898 647921 673904 647933
rect 675472 647921 675478 647933
rect 673898 647893 675478 647921
rect 673898 647881 673904 647893
rect 675472 647881 675478 647893
rect 675530 647881 675536 647933
rect 655504 646549 655510 646601
rect 655562 646589 655568 646601
rect 674704 646589 674710 646601
rect 655562 646561 674710 646589
rect 655562 646549 655568 646561
rect 674704 646549 674710 646561
rect 674762 646549 674768 646601
rect 41776 646253 41782 646305
rect 41834 646293 41840 646305
rect 50416 646293 50422 646305
rect 41834 646265 50422 646293
rect 41834 646253 41840 646265
rect 50416 646253 50422 646265
rect 50474 646253 50480 646305
rect 41776 645735 41782 645787
rect 41834 645775 41840 645787
rect 53296 645775 53302 645787
rect 41834 645747 53302 645775
rect 41834 645735 41840 645747
rect 53296 645735 53302 645747
rect 53354 645735 53360 645787
rect 41584 645365 41590 645417
rect 41642 645405 41648 645417
rect 47632 645405 47638 645417
rect 41642 645377 47638 645405
rect 41642 645365 41648 645377
rect 47632 645365 47638 645377
rect 47690 645365 47696 645417
rect 41776 644773 41782 644825
rect 41834 644813 41840 644825
rect 43216 644813 43222 644825
rect 41834 644785 43222 644813
rect 41834 644773 41840 644785
rect 43216 644773 43222 644785
rect 43274 644773 43280 644825
rect 672784 644773 672790 644825
rect 672842 644813 672848 644825
rect 675376 644813 675382 644825
rect 672842 644785 675382 644813
rect 672842 644773 672848 644785
rect 675376 644773 675382 644785
rect 675434 644773 675440 644825
rect 673456 643959 673462 644011
rect 673514 643999 673520 644011
rect 675472 643999 675478 644011
rect 673514 643971 675478 643999
rect 673514 643959 673520 643971
rect 675472 643959 675478 643971
rect 675530 643959 675536 644011
rect 672688 643367 672694 643419
rect 672746 643407 672752 643419
rect 675376 643407 675382 643419
rect 672746 643379 675382 643407
rect 672746 643367 672752 643379
rect 675376 643367 675382 643379
rect 675434 643367 675440 643419
rect 654448 642257 654454 642309
rect 654506 642297 654512 642309
rect 672592 642297 672598 642309
rect 654506 642269 672598 642297
rect 654506 642257 654512 642269
rect 672592 642257 672598 642269
rect 672650 642257 672656 642309
rect 673360 642257 673366 642309
rect 673418 642297 673424 642309
rect 675472 642297 675478 642309
rect 673418 642269 675478 642297
rect 673418 642257 673424 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 674704 641813 674710 641865
rect 674762 641853 674768 641865
rect 675376 641853 675382 641865
rect 674762 641825 675382 641853
rect 674762 641813 674768 641825
rect 675376 641813 675382 641825
rect 675434 641813 675440 641865
rect 665008 640407 665014 640459
rect 665066 640447 665072 640459
rect 668080 640447 668086 640459
rect 665066 640419 668086 640447
rect 665066 640407 665072 640419
rect 668080 640407 668086 640419
rect 668138 640407 668144 640459
rect 41776 639519 41782 639571
rect 41834 639559 41840 639571
rect 43120 639559 43126 639571
rect 41834 639531 43126 639559
rect 41834 639519 41840 639531
rect 43120 639519 43126 639531
rect 43178 639519 43184 639571
rect 41680 637003 41686 637055
rect 41738 637043 41744 637055
rect 43024 637043 43030 637055
rect 41738 637015 43030 637043
rect 41738 637003 41744 637015
rect 43024 637003 43030 637015
rect 43082 637003 43088 637055
rect 47728 636485 47734 636537
rect 47786 636525 47792 636537
rect 59536 636525 59542 636537
rect 47786 636497 59542 636525
rect 47786 636485 47792 636497
rect 59536 636485 59542 636497
rect 59594 636485 59600 636537
rect 672304 635597 672310 635649
rect 672362 635637 672368 635649
rect 679696 635637 679702 635649
rect 672362 635609 679702 635637
rect 672362 635597 672368 635609
rect 679696 635597 679702 635609
rect 679754 635597 679760 635649
rect 41680 634931 41686 634983
rect 41738 634971 41744 634983
rect 42832 634971 42838 634983
rect 41738 634943 42838 634971
rect 41738 634931 41744 634943
rect 42832 634931 42838 634943
rect 42890 634931 42896 634983
rect 41680 633895 41686 633947
rect 41738 633935 41744 633947
rect 46000 633935 46006 633947
rect 41738 633907 46006 633935
rect 41738 633895 41744 633907
rect 46000 633895 46006 633907
rect 46058 633895 46064 633947
rect 42928 629677 42934 629729
rect 42986 629717 42992 629729
rect 43408 629717 43414 629729
rect 42986 629689 43414 629717
rect 42986 629677 42992 629689
rect 43408 629677 43414 629689
rect 43466 629677 43472 629729
rect 25840 629233 25846 629285
rect 25898 629273 25904 629285
rect 43696 629273 43702 629285
rect 25898 629245 43702 629273
rect 25898 629233 25904 629245
rect 43696 629233 43702 629245
rect 43754 629233 43760 629285
rect 42832 627827 42838 627879
rect 42890 627867 42896 627879
rect 47536 627867 47542 627879
rect 42890 627839 47542 627867
rect 42890 627827 42896 627839
rect 47536 627827 47542 627839
rect 47594 627827 47600 627879
rect 654448 627827 654454 627879
rect 654506 627867 654512 627879
rect 663952 627867 663958 627879
rect 654506 627839 663958 627867
rect 654506 627827 654512 627839
rect 663952 627827 663958 627839
rect 664010 627827 664016 627879
rect 655312 627753 655318 627805
rect 655370 627793 655376 627805
rect 665200 627793 665206 627805
rect 655370 627765 665206 627793
rect 655370 627753 655376 627765
rect 665200 627753 665206 627765
rect 665258 627753 665264 627805
rect 668080 627753 668086 627805
rect 668138 627793 668144 627805
rect 670864 627793 670870 627805
rect 668138 627765 670870 627793
rect 668138 627753 668144 627765
rect 670864 627753 670870 627765
rect 670922 627753 670928 627805
rect 43024 627679 43030 627731
rect 43082 627719 43088 627731
rect 43504 627719 43510 627731
rect 43082 627691 43510 627719
rect 43082 627679 43088 627691
rect 43504 627679 43510 627691
rect 43562 627679 43568 627731
rect 666640 627679 666646 627731
rect 666698 627719 666704 627731
rect 676048 627719 676054 627731
rect 666698 627691 676054 627719
rect 666698 627679 666704 627691
rect 676048 627679 676054 627691
rect 676106 627679 676112 627731
rect 42064 627531 42070 627583
rect 42122 627571 42128 627583
rect 43120 627571 43126 627583
rect 42122 627543 43126 627571
rect 42122 627531 42128 627543
rect 43120 627531 43126 627543
rect 43178 627531 43184 627583
rect 41968 627457 41974 627509
rect 42026 627497 42032 627509
rect 43024 627497 43030 627509
rect 42026 627469 43030 627497
rect 42026 627457 42032 627469
rect 43024 627457 43030 627469
rect 43082 627457 43088 627509
rect 41776 627383 41782 627435
rect 41834 627383 41840 627435
rect 41872 627383 41878 627435
rect 41930 627423 41936 627435
rect 42928 627423 42934 627435
rect 41930 627395 42934 627423
rect 41930 627383 41936 627395
rect 42928 627383 42934 627395
rect 42986 627383 42992 627435
rect 41794 627065 41822 627383
rect 672400 627309 672406 627361
rect 672458 627349 672464 627361
rect 676240 627349 676246 627361
rect 672458 627321 676246 627349
rect 672458 627309 672464 627321
rect 676240 627309 676246 627321
rect 676298 627309 676304 627361
rect 41776 627013 41782 627065
rect 41834 627013 41840 627065
rect 661264 626569 661270 626621
rect 661322 626609 661328 626621
rect 676048 626609 676054 626621
rect 661322 626581 676054 626609
rect 661322 626569 661328 626581
rect 676048 626569 676054 626581
rect 676106 626569 676112 626621
rect 672016 625607 672022 625659
rect 672074 625647 672080 625659
rect 676048 625647 676054 625659
rect 672074 625619 676054 625647
rect 672074 625607 672080 625619
rect 676048 625607 676054 625619
rect 676106 625607 676112 625659
rect 42160 625311 42166 625363
rect 42218 625351 42224 625363
rect 43216 625351 43222 625363
rect 42218 625323 43222 625351
rect 42218 625311 42224 625323
rect 43216 625311 43222 625323
rect 43274 625311 43280 625363
rect 674224 624867 674230 624919
rect 674282 624907 674288 624919
rect 676048 624907 676054 624919
rect 674282 624879 676054 624907
rect 674282 624867 674288 624879
rect 676048 624867 676054 624879
rect 676106 624867 676112 624919
rect 42160 624645 42166 624697
rect 42218 624685 42224 624697
rect 42832 624685 42838 624697
rect 42218 624657 42838 624685
rect 42218 624645 42224 624657
rect 42832 624645 42838 624657
rect 42890 624645 42896 624697
rect 670864 624645 670870 624697
rect 670922 624685 670928 624697
rect 675952 624685 675958 624697
rect 670922 624657 675958 624685
rect 670922 624645 670928 624657
rect 675952 624645 675958 624657
rect 676010 624645 676016 624697
rect 42832 624497 42838 624549
rect 42890 624537 42896 624549
rect 43408 624537 43414 624549
rect 42890 624509 43414 624537
rect 42890 624497 42896 624509
rect 43408 624497 43414 624509
rect 43466 624497 43472 624549
rect 665200 623535 665206 623587
rect 665258 623575 665264 623587
rect 670960 623575 670966 623587
rect 665258 623547 670966 623575
rect 665258 623535 665264 623547
rect 670960 623535 670966 623547
rect 671018 623575 671024 623587
rect 675952 623575 675958 623587
rect 671018 623547 675958 623575
rect 671018 623535 671024 623547
rect 675952 623535 675958 623547
rect 676010 623535 676016 623587
rect 42160 623461 42166 623513
rect 42218 623501 42224 623513
rect 43504 623501 43510 623513
rect 42218 623473 43510 623501
rect 42218 623461 42224 623473
rect 43504 623461 43510 623473
rect 43562 623461 43568 623513
rect 47536 622055 47542 622107
rect 47594 622095 47600 622107
rect 59536 622095 59542 622107
rect 47594 622067 59542 622095
rect 47594 622055 47600 622067
rect 59536 622055 59542 622067
rect 59594 622055 59600 622107
rect 674416 621981 674422 622033
rect 674474 622021 674480 622033
rect 676240 622021 676246 622033
rect 674474 621993 676246 622021
rect 674474 621981 674480 621993
rect 676240 621981 676246 621993
rect 676298 621981 676304 622033
rect 42160 621611 42166 621663
rect 42218 621651 42224 621663
rect 42832 621651 42838 621663
rect 42218 621623 42838 621651
rect 42218 621611 42224 621623
rect 42832 621611 42838 621623
rect 42890 621611 42896 621663
rect 42160 620353 42166 620405
rect 42218 620393 42224 620405
rect 42928 620393 42934 620405
rect 42218 620365 42934 620393
rect 42218 620353 42224 620365
rect 42928 620353 42934 620365
rect 42986 620353 42992 620405
rect 673648 619169 673654 619221
rect 673706 619209 673712 619221
rect 676048 619209 676054 619221
rect 673706 619181 676054 619209
rect 673706 619169 673712 619181
rect 676048 619169 676054 619181
rect 676106 619169 676112 619221
rect 42256 619021 42262 619073
rect 42314 619061 42320 619073
rect 43024 619061 43030 619073
rect 42314 619033 43030 619061
rect 42314 619021 42320 619033
rect 43024 619021 43030 619033
rect 43082 619021 43088 619073
rect 673264 618133 673270 618185
rect 673322 618173 673328 618185
rect 676048 618173 676054 618185
rect 673322 618145 676054 618173
rect 673322 618133 673328 618145
rect 676048 618133 676054 618145
rect 676106 618133 676112 618185
rect 42064 617837 42070 617889
rect 42122 617877 42128 617889
rect 43120 617877 43126 617889
rect 42122 617849 43126 617877
rect 42122 617837 42128 617849
rect 43120 617837 43126 617849
rect 43178 617837 43184 617889
rect 673552 617615 673558 617667
rect 673610 617655 673616 617667
rect 676048 617655 676054 617667
rect 673610 617627 676054 617655
rect 673610 617615 673616 617627
rect 676048 617615 676054 617627
rect 676106 617615 676112 617667
rect 672880 617393 672886 617445
rect 672938 617433 672944 617445
rect 676240 617433 676246 617445
rect 672938 617405 676246 617433
rect 672938 617393 672944 617405
rect 676240 617393 676246 617405
rect 676298 617393 676304 617445
rect 42256 616653 42262 616705
rect 42314 616693 42320 616705
rect 42928 616693 42934 616705
rect 42314 616665 42934 616693
rect 42314 616653 42320 616665
rect 42928 616653 42934 616665
rect 42986 616653 42992 616705
rect 672976 616653 672982 616705
rect 673034 616693 673040 616705
rect 676048 616693 676054 616705
rect 673034 616665 676054 616693
rect 673034 616653 673040 616665
rect 676048 616653 676054 616665
rect 676106 616653 676112 616705
rect 652336 616357 652342 616409
rect 652394 616397 652400 616409
rect 655312 616397 655318 616409
rect 652394 616369 655318 616397
rect 652394 616357 652400 616369
rect 655312 616357 655318 616369
rect 655370 616357 655376 616409
rect 653872 614507 653878 614559
rect 653930 614547 653936 614559
rect 661168 614547 661174 614559
rect 653930 614519 661174 614547
rect 653930 614507 653936 614519
rect 661168 614507 661174 614519
rect 661226 614507 661232 614559
rect 42160 614137 42166 614189
rect 42218 614177 42224 614189
rect 42832 614177 42838 614189
rect 42218 614149 42838 614177
rect 42218 614137 42224 614149
rect 42832 614137 42838 614149
rect 42890 614137 42896 614189
rect 42160 613619 42166 613671
rect 42218 613659 42224 613671
rect 42928 613659 42934 613671
rect 42218 613631 42934 613659
rect 42218 613619 42224 613631
rect 42928 613619 42934 613631
rect 42986 613619 42992 613671
rect 652336 613471 652342 613523
rect 652394 613511 652400 613523
rect 679792 613511 679798 613523
rect 652394 613483 679798 613511
rect 652394 613471 652400 613483
rect 679792 613471 679798 613483
rect 679850 613471 679856 613523
rect 42064 612805 42070 612857
rect 42122 612845 42128 612857
rect 43024 612845 43030 612857
rect 42122 612817 43030 612845
rect 42122 612805 42128 612817
rect 43024 612805 43030 612817
rect 43082 612805 43088 612857
rect 47632 610585 47638 610637
rect 47690 610625 47696 610637
rect 59248 610625 59254 610637
rect 47690 610597 59254 610625
rect 47690 610585 47696 610597
rect 59248 610585 59254 610597
rect 59306 610585 59312 610637
rect 660592 607921 660598 607973
rect 660650 607961 660656 607973
rect 666832 607961 666838 607973
rect 660650 607933 666838 607961
rect 660650 607921 660656 607933
rect 666832 607921 666838 607933
rect 666890 607921 666896 607973
rect 652912 607699 652918 607751
rect 652970 607739 652976 607751
rect 653872 607739 653878 607751
rect 652970 607711 653878 607739
rect 652970 607699 652976 607711
rect 653872 607699 653878 607711
rect 653930 607699 653936 607751
rect 672208 607033 672214 607085
rect 672266 607073 672272 607085
rect 675472 607073 675478 607085
rect 672266 607045 675478 607073
rect 672266 607033 672272 607045
rect 675472 607033 675478 607045
rect 675530 607033 675536 607085
rect 673552 603925 673558 603977
rect 673610 603965 673616 603977
rect 675472 603965 675478 603977
rect 673610 603937 675478 603965
rect 673610 603925 673616 603937
rect 675472 603925 675478 603937
rect 675530 603925 675536 603977
rect 654544 603333 654550 603385
rect 654602 603373 654608 603385
rect 674608 603373 674614 603385
rect 654602 603345 674614 603373
rect 654602 603333 654608 603345
rect 674608 603333 674614 603345
rect 674666 603333 674672 603385
rect 673264 603259 673270 603311
rect 673322 603299 673328 603311
rect 675376 603299 675382 603311
rect 673322 603271 675382 603299
rect 673322 603259 673328 603271
rect 675376 603259 675382 603271
rect 675434 603259 675440 603311
rect 41776 603037 41782 603089
rect 41834 603077 41840 603089
rect 47728 603077 47734 603089
rect 41834 603049 47734 603077
rect 41834 603037 41840 603049
rect 47728 603037 47734 603049
rect 47786 603037 47792 603089
rect 41584 602741 41590 602793
rect 41642 602781 41648 602793
rect 47536 602781 47542 602793
rect 41642 602753 47542 602781
rect 41642 602741 41648 602753
rect 47536 602741 47542 602753
rect 47594 602741 47600 602793
rect 672304 602667 672310 602719
rect 672362 602707 672368 602719
rect 675376 602707 675382 602719
rect 672362 602679 675382 602707
rect 672362 602667 672368 602679
rect 675376 602667 675382 602679
rect 675434 602667 675440 602719
rect 41584 602149 41590 602201
rect 41642 602189 41648 602201
rect 53200 602189 53206 602201
rect 41642 602161 53206 602189
rect 41642 602149 41648 602161
rect 53200 602149 53206 602161
rect 53258 602149 53264 602201
rect 653008 602001 653014 602053
rect 653066 602041 653072 602053
rect 660592 602041 660598 602053
rect 653066 602013 660598 602041
rect 653066 602001 653072 602013
rect 660592 602001 660598 602013
rect 660650 602001 660656 602053
rect 654448 601927 654454 601979
rect 654506 601967 654512 601979
rect 672496 601967 672502 601979
rect 654506 601939 672502 601967
rect 654506 601927 654512 601939
rect 672496 601927 672502 601939
rect 672554 601927 672560 601979
rect 41776 601557 41782 601609
rect 41834 601597 41840 601609
rect 43504 601597 43510 601609
rect 41834 601569 43510 601597
rect 41834 601557 41840 601569
rect 43504 601557 43510 601569
rect 43562 601557 43568 601609
rect 41776 600965 41782 601017
rect 41834 601005 41840 601017
rect 43216 601005 43222 601017
rect 41834 600977 43222 601005
rect 41834 600965 41840 600977
rect 43216 600965 43222 600977
rect 43274 600965 43280 601017
rect 41584 599855 41590 599907
rect 41642 599895 41648 599907
rect 43312 599895 43318 599907
rect 41642 599867 43318 599895
rect 41642 599855 41648 599867
rect 43312 599855 43318 599867
rect 43370 599895 43376 599907
rect 44368 599895 44374 599907
rect 43370 599867 44374 599895
rect 43370 599855 43376 599867
rect 44368 599855 44374 599867
rect 44426 599855 44432 599907
rect 672112 599781 672118 599833
rect 672170 599821 672176 599833
rect 675376 599821 675382 599833
rect 672170 599793 675382 599821
rect 672170 599781 672176 599793
rect 675376 599781 675382 599793
rect 675434 599781 675440 599833
rect 672880 599263 672886 599315
rect 672938 599303 672944 599315
rect 675376 599303 675382 599315
rect 672938 599275 675382 599303
rect 672938 599263 672944 599275
rect 675376 599263 675382 599275
rect 675434 599263 675440 599315
rect 41776 598967 41782 599019
rect 41834 599007 41840 599019
rect 43504 599007 43510 599019
rect 41834 598979 43510 599007
rect 41834 598967 41840 598979
rect 43504 598967 43510 598979
rect 43562 598967 43568 599019
rect 672976 598375 672982 598427
rect 673034 598415 673040 598427
rect 675472 598415 675478 598427
rect 673034 598387 675478 598415
rect 673034 598375 673040 598387
rect 675472 598375 675478 598387
rect 675530 598375 675536 598427
rect 41584 597709 41590 597761
rect 41642 597749 41648 597761
rect 42928 597749 42934 597761
rect 41642 597721 42934 597749
rect 41642 597709 41648 597721
rect 42928 597709 42934 597721
rect 42986 597709 42992 597761
rect 672400 597117 672406 597169
rect 672458 597157 672464 597169
rect 675472 597157 675478 597169
rect 672458 597129 675478 597157
rect 672458 597117 672464 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 674608 596821 674614 596873
rect 674666 596861 674672 596873
rect 675376 596861 675382 596873
rect 674666 596833 675382 596861
rect 674666 596821 674672 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 43504 596155 43510 596207
rect 43562 596195 43568 596207
rect 47536 596195 47542 596207
rect 43562 596167 47542 596195
rect 43562 596155 43568 596167
rect 47536 596155 47542 596167
rect 47594 596155 47600 596207
rect 53200 596155 53206 596207
rect 53258 596195 53264 596207
rect 59344 596195 59350 596207
rect 53258 596167 59350 596195
rect 53258 596155 53264 596167
rect 59344 596155 59350 596167
rect 59402 596155 59408 596207
rect 41776 593935 41782 593987
rect 41834 593975 41840 593987
rect 42736 593975 42742 593987
rect 41834 593947 42742 593975
rect 41834 593935 41840 593947
rect 42736 593935 42742 593947
rect 42794 593935 42800 593987
rect 41776 593491 41782 593543
rect 41834 593531 41840 593543
rect 43120 593531 43126 593543
rect 41834 593503 43126 593531
rect 41834 593491 41840 593503
rect 43120 593491 43126 593503
rect 43178 593491 43184 593543
rect 41776 592529 41782 592581
rect 41834 592569 41840 592581
rect 43024 592569 43030 592581
rect 41834 592541 43030 592569
rect 41834 592529 41840 592541
rect 43024 592529 43030 592541
rect 43082 592529 43088 592581
rect 41776 591197 41782 591249
rect 41834 591237 41840 591249
rect 42832 591237 42838 591249
rect 41834 591209 42838 591237
rect 41834 591197 41840 591209
rect 42832 591197 42838 591209
rect 42890 591197 42896 591249
rect 41584 590679 41590 590731
rect 41642 590719 41648 590731
rect 47440 590719 47446 590731
rect 41642 590691 47446 590719
rect 41642 590679 41648 590691
rect 47440 590679 47446 590691
rect 47498 590679 47504 590731
rect 654448 590383 654454 590435
rect 654506 590423 654512 590435
rect 666832 590423 666838 590435
rect 654506 590395 666838 590423
rect 654506 590383 654512 590395
rect 666832 590383 666838 590395
rect 666890 590383 666896 590435
rect 655312 588607 655318 588659
rect 655370 588647 655376 588659
rect 658864 588647 658870 588659
rect 655370 588619 658870 588647
rect 655370 588607 655376 588619
rect 658864 588607 658870 588619
rect 658922 588607 658928 588659
rect 658864 586017 658870 586069
rect 658922 586057 658928 586069
rect 668080 586057 668086 586069
rect 658922 586029 668086 586057
rect 658922 586017 658928 586029
rect 668080 586017 668086 586029
rect 668138 586017 668144 586069
rect 43504 584685 43510 584737
rect 43562 584725 43568 584737
rect 50320 584725 50326 584737
rect 43562 584697 50326 584725
rect 43562 584685 43568 584697
rect 50320 584685 50326 584697
rect 50378 584685 50384 584737
rect 50416 584685 50422 584737
rect 50474 584725 50480 584737
rect 59536 584725 59542 584737
rect 50474 584697 59542 584725
rect 50474 584685 50480 584697
rect 59536 584685 59542 584697
rect 59594 584685 59600 584737
rect 41776 584315 41782 584367
rect 41834 584355 41840 584367
rect 43696 584355 43702 584367
rect 41834 584327 43702 584355
rect 41834 584315 41840 584327
rect 43696 584315 43702 584327
rect 43754 584315 43760 584367
rect 41968 584241 41974 584293
rect 42026 584281 42032 584293
rect 43792 584281 43798 584293
rect 42026 584253 43798 584281
rect 42026 584241 42032 584253
rect 43792 584241 43798 584253
rect 43850 584241 43856 584293
rect 41872 584167 41878 584219
rect 41930 584167 41936 584219
rect 42160 584167 42166 584219
rect 42218 584207 42224 584219
rect 43408 584207 43414 584219
rect 42218 584179 43414 584207
rect 42218 584167 42224 584179
rect 43408 584167 43414 584179
rect 43466 584167 43472 584219
rect 41890 583997 41918 584167
rect 41872 583945 41878 583997
rect 41930 583945 41936 583997
rect 42448 583649 42454 583701
rect 42506 583689 42512 583701
rect 43312 583689 43318 583701
rect 42506 583661 43318 583689
rect 42506 583649 42512 583661
rect 43312 583649 43318 583661
rect 43370 583649 43376 583701
rect 670096 582465 670102 582517
rect 670154 582505 670160 582517
rect 676048 582505 676054 582517
rect 670154 582477 676054 582505
rect 670154 582465 670160 582477
rect 676048 582465 676054 582477
rect 676106 582465 676112 582517
rect 42160 582095 42166 582147
rect 42218 582135 42224 582147
rect 42928 582135 42934 582147
rect 42218 582107 42934 582135
rect 42218 582095 42224 582107
rect 42928 582095 42934 582107
rect 42986 582095 42992 582147
rect 652816 581947 652822 581999
rect 652874 581987 652880 581999
rect 652874 581959 659534 581987
rect 652874 581947 652880 581959
rect 43024 581873 43030 581925
rect 43082 581913 43088 581925
rect 43312 581913 43318 581925
rect 43082 581885 43318 581913
rect 43082 581873 43088 581885
rect 43312 581873 43318 581885
rect 43370 581873 43376 581925
rect 659506 581765 659534 581959
rect 663760 581947 663766 581999
rect 663818 581987 663824 581999
rect 676048 581987 676054 581999
rect 663818 581959 676054 581987
rect 663818 581947 663824 581959
rect 676048 581947 676054 581959
rect 676106 581947 676112 581999
rect 668080 581799 668086 581851
rect 668138 581839 668144 581851
rect 670768 581839 670774 581851
rect 668138 581811 670774 581839
rect 668138 581799 668144 581811
rect 670768 581799 670774 581811
rect 670826 581799 670832 581851
rect 665872 581765 665878 581777
rect 659506 581737 665878 581765
rect 665872 581725 665878 581737
rect 665930 581725 665936 581777
rect 666736 581577 666742 581629
rect 666794 581617 666800 581629
rect 676240 581617 676246 581629
rect 666794 581589 676246 581617
rect 666794 581577 666800 581589
rect 676240 581577 676246 581589
rect 676298 581577 676304 581629
rect 42064 581355 42070 581407
rect 42122 581395 42128 581407
rect 43504 581395 43510 581407
rect 42122 581367 43510 581395
rect 42122 581355 42128 581367
rect 43504 581355 43510 581367
rect 43562 581355 43568 581407
rect 672016 580985 672022 581037
rect 672074 581025 672080 581037
rect 676048 581025 676054 581037
rect 672074 580997 676054 581025
rect 672074 580985 672080 580997
rect 676048 580985 676054 580997
rect 676106 580985 676112 581037
rect 42064 580245 42070 580297
rect 42122 580285 42128 580297
rect 42736 580285 42742 580297
rect 42122 580257 42742 580285
rect 42122 580245 42128 580257
rect 42736 580245 42742 580257
rect 42794 580245 42800 580297
rect 670576 580171 670582 580223
rect 670634 580211 670640 580223
rect 676240 580211 676246 580223
rect 670634 580183 676246 580211
rect 670634 580171 670640 580183
rect 676240 580171 676246 580183
rect 676298 580171 676304 580223
rect 42736 580097 42742 580149
rect 42794 580137 42800 580149
rect 43120 580137 43126 580149
rect 42794 580109 43126 580137
rect 42794 580097 42800 580109
rect 43120 580097 43126 580109
rect 43178 580097 43184 580149
rect 670864 579949 670870 580001
rect 670922 579989 670928 580001
rect 676048 579989 676054 580001
rect 670922 579961 676054 579989
rect 670922 579949 670928 579961
rect 676048 579949 676054 579961
rect 676106 579949 676112 580001
rect 43024 579801 43030 579853
rect 43082 579841 43088 579853
rect 43408 579841 43414 579853
rect 43082 579813 43414 579841
rect 43082 579801 43088 579813
rect 43408 579801 43414 579813
rect 43466 579801 43472 579853
rect 670768 579431 670774 579483
rect 670826 579471 670832 579483
rect 676048 579471 676054 579483
rect 670826 579443 676054 579471
rect 670826 579431 670832 579443
rect 676048 579431 676054 579443
rect 676106 579431 676112 579483
rect 42160 578987 42166 579039
rect 42218 579027 42224 579039
rect 42832 579027 42838 579039
rect 42218 578999 42838 579027
rect 42218 578987 42224 578999
rect 42832 578987 42838 578999
rect 42890 578987 42896 579039
rect 670960 578913 670966 578965
rect 671018 578953 671024 578965
rect 676048 578953 676054 578965
rect 671018 578925 676054 578953
rect 671018 578913 671024 578925
rect 676048 578913 676054 578925
rect 676106 578913 676112 578965
rect 665872 578395 665878 578447
rect 665930 578435 665936 578447
rect 670672 578435 670678 578447
rect 665930 578407 670678 578435
rect 665930 578395 665936 578407
rect 670672 578395 670678 578407
rect 670730 578435 670736 578447
rect 676048 578435 676054 578447
rect 670730 578407 676054 578435
rect 670730 578395 670736 578407
rect 676048 578395 676054 578407
rect 676106 578395 676112 578447
rect 42064 578247 42070 578299
rect 42122 578287 42128 578299
rect 42736 578287 42742 578299
rect 42122 578259 42742 578287
rect 42122 578247 42128 578259
rect 42736 578247 42742 578259
rect 42794 578247 42800 578299
rect 42160 577655 42166 577707
rect 42218 577695 42224 577707
rect 42928 577695 42934 577707
rect 42218 577667 42934 577695
rect 42218 577655 42224 577667
rect 42928 577655 42934 577667
rect 42986 577655 42992 577707
rect 654448 577285 654454 577337
rect 654506 577325 654512 577337
rect 661168 577325 661174 577337
rect 654506 577297 661174 577325
rect 654506 577285 654512 577297
rect 661168 577285 661174 577297
rect 661226 577285 661232 577337
rect 42160 577137 42166 577189
rect 42218 577177 42224 577189
rect 43504 577177 43510 577189
rect 42218 577149 43510 577177
rect 42218 577137 42224 577149
rect 43504 577137 43510 577149
rect 43562 577137 43568 577189
rect 673744 574991 673750 575043
rect 673802 575031 673808 575043
rect 676048 575031 676054 575043
rect 673802 575003 676054 575031
rect 673802 574991 673808 575003
rect 676048 574991 676054 575003
rect 676106 574991 676112 575043
rect 42160 574621 42166 574673
rect 42218 574661 42224 574673
rect 43120 574661 43126 574673
rect 42218 574633 43126 574661
rect 42218 574621 42224 574633
rect 43120 574621 43126 574633
rect 43178 574621 43184 574673
rect 673072 574621 673078 574673
rect 673130 574661 673136 574673
rect 676240 574661 676246 574673
rect 673130 574633 676246 574661
rect 673130 574621 673136 574633
rect 676240 574621 676246 574633
rect 676298 574621 676304 574673
rect 42160 574103 42166 574155
rect 42218 574143 42224 574155
rect 43024 574143 43030 574155
rect 42218 574115 43030 574143
rect 42218 574103 42224 574115
rect 43024 574103 43030 574115
rect 43082 574103 43088 574155
rect 673168 573881 673174 573933
rect 673226 573921 673232 573933
rect 676048 573921 676054 573933
rect 673226 573893 676054 573921
rect 673226 573881 673232 573893
rect 676048 573881 676054 573893
rect 676106 573881 676112 573933
rect 673360 573511 673366 573563
rect 673418 573551 673424 573563
rect 676048 573551 676054 573563
rect 673418 573523 676054 573551
rect 673418 573511 673424 573523
rect 676048 573511 676054 573523
rect 676106 573511 676112 573563
rect 42160 573437 42166 573489
rect 42218 573477 42224 573489
rect 43600 573477 43606 573489
rect 42218 573449 43606 573477
rect 42218 573437 42224 573449
rect 43600 573437 43606 573449
rect 43658 573437 43664 573489
rect 673456 572993 673462 573045
rect 673514 573033 673520 573045
rect 676048 573033 676054 573045
rect 673514 573005 676054 573033
rect 673514 572993 673520 573005
rect 676048 572993 676054 573005
rect 676106 572993 676112 573045
rect 42160 572771 42166 572823
rect 42218 572811 42224 572823
rect 42832 572811 42838 572823
rect 42218 572783 42838 572811
rect 42218 572771 42224 572783
rect 42832 572771 42838 572783
rect 42890 572771 42896 572823
rect 673840 572401 673846 572453
rect 673898 572441 673904 572453
rect 676048 572441 676054 572453
rect 673898 572413 676054 572441
rect 673898 572401 673904 572413
rect 676048 572401 676054 572413
rect 676106 572401 676112 572453
rect 672784 571957 672790 572009
rect 672842 571997 672848 572009
rect 676048 571997 676054 572009
rect 672842 571969 676054 571997
rect 672842 571957 672848 571969
rect 676048 571957 676054 571969
rect 676106 571957 676112 572009
rect 672688 571661 672694 571713
rect 672746 571701 672752 571713
rect 676240 571701 676246 571713
rect 672746 571673 676246 571701
rect 672746 571661 672752 571673
rect 676240 571661 676246 571673
rect 676298 571661 676304 571713
rect 42160 570847 42166 570899
rect 42218 570887 42224 570899
rect 42928 570887 42934 570899
rect 42218 570859 42934 570887
rect 42218 570847 42224 570859
rect 42928 570847 42934 570859
rect 42986 570847 42992 570899
rect 42160 570403 42166 570455
rect 42218 570443 42224 570455
rect 42352 570443 42358 570455
rect 42218 570415 42358 570443
rect 42218 570403 42224 570415
rect 42352 570403 42358 570415
rect 42410 570403 42416 570455
rect 42352 570255 42358 570307
rect 42410 570295 42416 570307
rect 59536 570295 59542 570307
rect 42410 570267 59542 570295
rect 42410 570255 42416 570267
rect 59536 570255 59542 570267
rect 59594 570255 59600 570307
rect 42064 569663 42070 569715
rect 42122 569703 42128 569715
rect 42736 569703 42742 569715
rect 42122 569675 42742 569703
rect 42122 569663 42128 569675
rect 42736 569663 42742 569675
rect 42794 569663 42800 569715
rect 652816 567369 652822 567421
rect 652874 567409 652880 567421
rect 679984 567409 679990 567421
rect 652874 567381 679990 567409
rect 652874 567369 652880 567381
rect 679984 567369 679990 567381
rect 680042 567369 680048 567421
rect 41776 559821 41782 559873
rect 41834 559861 41840 559873
rect 50416 559861 50422 559873
rect 41834 559833 50422 559861
rect 41834 559821 41840 559833
rect 50416 559821 50422 559833
rect 50474 559821 50480 559873
rect 652720 559821 652726 559873
rect 652778 559861 652784 559873
rect 663760 559861 663766 559873
rect 652778 559833 663766 559861
rect 652778 559821 652784 559833
rect 663760 559821 663766 559833
rect 663818 559821 663824 559873
rect 674608 559377 674614 559429
rect 674666 559417 674672 559429
rect 675376 559417 675382 559429
rect 674666 559389 675382 559417
rect 674666 559377 674672 559389
rect 675376 559377 675382 559389
rect 675434 559377 675440 559429
rect 674512 558933 674518 558985
rect 674570 558973 674576 558985
rect 675472 558973 675478 558985
rect 674570 558945 675478 558973
rect 674570 558933 674576 558945
rect 675472 558933 675478 558945
rect 675530 558933 675536 558985
rect 41776 558785 41782 558837
rect 41834 558825 41840 558837
rect 53200 558825 53206 558837
rect 41834 558797 53206 558825
rect 41834 558785 41840 558797
rect 53200 558785 53206 558797
rect 53258 558785 53264 558837
rect 50320 558711 50326 558763
rect 50378 558751 50384 558763
rect 59536 558751 59542 558763
rect 50378 558723 59542 558751
rect 50378 558711 50384 558723
rect 59536 558711 59542 558723
rect 59594 558711 59600 558763
rect 41776 558341 41782 558393
rect 41834 558381 41840 558393
rect 43216 558381 43222 558393
rect 41834 558353 43222 558381
rect 41834 558341 41840 558353
rect 43216 558341 43222 558353
rect 43274 558341 43280 558393
rect 673840 558045 673846 558097
rect 673898 558085 673904 558097
rect 675376 558085 675382 558097
rect 673898 558057 675382 558085
rect 673898 558045 673904 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 41776 557823 41782 557875
rect 41834 557863 41840 557875
rect 43600 557863 43606 557875
rect 41834 557835 43606 557863
rect 41834 557823 41840 557835
rect 43600 557823 43606 557835
rect 43658 557823 43664 557875
rect 656560 557231 656566 557283
rect 656618 557271 656624 557283
rect 675280 557271 675286 557283
rect 656618 557243 675286 557271
rect 656618 557231 656624 557243
rect 675280 557231 675286 557243
rect 675338 557231 675344 557283
rect 674704 555233 674710 555285
rect 674762 555273 674768 555285
rect 675472 555273 675478 555285
rect 674762 555245 675478 555273
rect 674762 555233 674768 555245
rect 675472 555233 675478 555245
rect 675530 555233 675536 555285
rect 673744 554345 673750 554397
rect 673802 554385 673808 554397
rect 675376 554385 675382 554397
rect 673802 554357 675382 554385
rect 673802 554345 673808 554357
rect 675376 554345 675382 554357
rect 675434 554345 675440 554397
rect 673072 553901 673078 553953
rect 673130 553941 673136 553953
rect 675472 553941 675478 553953
rect 673130 553913 675478 553941
rect 673130 553901 673136 553913
rect 675472 553901 675478 553913
rect 675530 553901 675536 553953
rect 41584 553161 41590 553213
rect 41642 553201 41648 553213
rect 42832 553201 42838 553213
rect 41642 553173 42838 553201
rect 41642 553161 41648 553173
rect 42832 553161 42838 553173
rect 42890 553161 42896 553213
rect 673168 553161 673174 553213
rect 673226 553201 673232 553213
rect 675376 553201 675382 553213
rect 673226 553173 675382 553201
rect 673226 553161 673232 553173
rect 675376 553161 675382 553173
rect 675434 553161 675440 553213
rect 673648 551903 673654 551955
rect 673706 551943 673712 551955
rect 675472 551943 675478 551955
rect 673706 551915 675478 551943
rect 673706 551903 673712 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 41872 550423 41878 550475
rect 41930 550463 41936 550475
rect 43120 550463 43126 550475
rect 41930 550435 43126 550463
rect 41930 550423 41936 550435
rect 43120 550423 43126 550435
rect 43178 550423 43184 550475
rect 652624 550201 652630 550253
rect 652682 550241 652688 550253
rect 656560 550241 656566 550253
rect 652682 550213 656566 550241
rect 652682 550201 652688 550213
rect 656560 550201 656566 550213
rect 656618 550201 656624 550253
rect 41584 550127 41590 550179
rect 41642 550167 41648 550179
rect 42736 550167 42742 550179
rect 41642 550139 42742 550167
rect 41642 550127 41648 550139
rect 42736 550127 42742 550139
rect 42794 550127 42800 550179
rect 654832 550127 654838 550179
rect 654890 550167 654896 550179
rect 666640 550167 666646 550179
rect 654890 550139 666646 550167
rect 654890 550127 654896 550139
rect 666640 550127 666646 550139
rect 666698 550127 666704 550179
rect 674416 548869 674422 548921
rect 674474 548909 674480 548921
rect 675280 548909 675286 548921
rect 674474 548881 675286 548909
rect 674474 548869 674480 548881
rect 675280 548869 675286 548881
rect 675338 548869 675344 548921
rect 41872 548795 41878 548847
rect 41930 548835 41936 548847
rect 42832 548835 42838 548847
rect 41930 548807 42838 548835
rect 41930 548795 41936 548807
rect 42832 548795 42838 548807
rect 42890 548795 42896 548847
rect 674320 548203 674326 548255
rect 674378 548243 674384 548255
rect 675280 548243 675286 548255
rect 674378 548215 675286 548243
rect 674378 548203 674384 548215
rect 675280 548203 675286 548215
rect 675338 548203 675344 548255
rect 41872 547315 41878 547367
rect 41930 547355 41936 547367
rect 44464 547355 44470 547367
rect 41930 547327 44470 547355
rect 41930 547315 41936 547327
rect 44464 547315 44470 547327
rect 44522 547315 44528 547367
rect 670768 547167 670774 547219
rect 670826 547207 670832 547219
rect 679696 547207 679702 547219
rect 670826 547179 679702 547207
rect 670826 547167 670832 547179
rect 679696 547167 679702 547179
rect 679754 547167 679760 547219
rect 53296 544355 53302 544407
rect 53354 544395 53360 544407
rect 59536 544395 59542 544407
rect 53354 544367 59542 544395
rect 53354 544355 53360 544367
rect 59536 544355 59542 544367
rect 59594 544355 59600 544407
rect 42256 542801 42262 542853
rect 42314 542841 42320 542853
rect 43024 542841 43030 542853
rect 42314 542813 43030 542841
rect 42314 542801 42320 542813
rect 43024 542801 43030 542813
rect 43082 542801 43088 542853
rect 42064 541765 42070 541817
rect 42122 541805 42128 541817
rect 43120 541805 43126 541817
rect 42122 541777 43126 541805
rect 42122 541765 42128 541777
rect 43120 541765 43126 541777
rect 43178 541765 43184 541817
rect 656656 541543 656662 541595
rect 656714 541583 656720 541595
rect 656714 541555 659534 541583
rect 656714 541543 656720 541555
rect 42736 541469 42742 541521
rect 42794 541509 42800 541521
rect 47632 541509 47638 541521
rect 42794 541481 47638 541509
rect 42794 541469 42800 541481
rect 47632 541469 47638 541481
rect 47690 541469 47696 541521
rect 659506 541435 659534 541555
rect 670768 541435 670774 541447
rect 659506 541407 670774 541435
rect 670768 541395 670774 541407
rect 670826 541395 670832 541447
rect 41392 541321 41398 541373
rect 41450 541361 41456 541373
rect 43216 541361 43222 541373
rect 41450 541333 43222 541361
rect 41450 541321 41456 541333
rect 43216 541321 43222 541333
rect 43274 541321 43280 541373
rect 663760 541321 663766 541373
rect 663818 541361 663824 541373
rect 676720 541361 676726 541373
rect 663818 541333 676726 541361
rect 663818 541321 663824 541333
rect 676720 541321 676726 541333
rect 676778 541321 676784 541373
rect 41488 541247 41494 541299
rect 41546 541287 41552 541299
rect 43408 541287 43414 541299
rect 41546 541259 43414 541287
rect 41546 541247 41552 541259
rect 43408 541247 43414 541259
rect 43466 541247 43472 541299
rect 41776 540951 41782 541003
rect 41834 540951 41840 541003
rect 41794 540781 41822 540951
rect 41776 540729 41782 540781
rect 41834 540729 41840 540781
rect 42064 538879 42070 538931
rect 42122 538919 42128 538931
rect 42928 538919 42934 538931
rect 42122 538891 42934 538919
rect 42122 538879 42128 538891
rect 42928 538879 42934 538891
rect 42986 538879 42992 538931
rect 42928 538731 42934 538783
rect 42986 538771 42992 538783
rect 43216 538771 43222 538783
rect 42986 538743 43222 538771
rect 42986 538731 42992 538743
rect 43216 538731 43222 538743
rect 43274 538731 43280 538783
rect 42160 538287 42166 538339
rect 42218 538327 42224 538339
rect 42736 538327 42742 538339
rect 42218 538299 42742 538327
rect 42218 538287 42224 538299
rect 42736 538287 42742 538299
rect 42794 538287 42800 538339
rect 654448 537473 654454 537525
rect 654506 537513 654512 537525
rect 663856 537513 663862 537525
rect 654506 537485 663862 537513
rect 654506 537473 654512 537485
rect 663856 537473 663862 537485
rect 663914 537473 663920 537525
rect 672592 537473 672598 537525
rect 672650 537513 672656 537525
rect 676048 537513 676054 537525
rect 672650 537485 676054 537513
rect 672650 537473 672656 537485
rect 676048 537473 676054 537485
rect 676106 537473 676112 537525
rect 670768 537325 670774 537377
rect 670826 537365 670832 537377
rect 676624 537365 676630 537377
rect 670826 537337 676630 537365
rect 670826 537325 670832 537337
rect 676624 537325 676630 537337
rect 676682 537325 676688 537377
rect 42064 537029 42070 537081
rect 42122 537069 42128 537081
rect 43312 537069 43318 537081
rect 42122 537041 43318 537069
rect 42122 537029 42128 537041
rect 43312 537029 43318 537041
rect 43370 537029 43376 537081
rect 661072 536881 661078 536933
rect 661130 536921 661136 536933
rect 676048 536921 676054 536933
rect 661130 536893 676054 536921
rect 661130 536881 661136 536893
rect 676048 536881 676054 536893
rect 676106 536881 676112 536933
rect 663952 536585 663958 536637
rect 664010 536625 664016 536637
rect 676240 536625 676246 536637
rect 664010 536597 676246 536625
rect 664010 536585 664016 536597
rect 676240 536585 676246 536597
rect 676298 536585 676304 536637
rect 42064 535771 42070 535823
rect 42122 535811 42128 535823
rect 42832 535811 42838 535823
rect 42122 535783 42838 535811
rect 42122 535771 42128 535783
rect 42832 535771 42838 535783
rect 42890 535771 42896 535823
rect 670960 534883 670966 534935
rect 671018 534923 671024 534935
rect 676048 534923 676054 534935
rect 671018 534895 676054 534923
rect 671018 534883 671024 534895
rect 676048 534883 676054 534895
rect 676106 534883 676112 534935
rect 42160 534439 42166 534491
rect 42218 534479 42224 534491
rect 42928 534479 42934 534491
rect 42218 534451 42934 534479
rect 42218 534439 42224 534451
rect 42928 534439 42934 534451
rect 42986 534439 42992 534491
rect 42160 533921 42166 533973
rect 42218 533961 42224 533973
rect 43120 533961 43126 533973
rect 42218 533933 43126 533961
rect 42218 533921 42224 533933
rect 43120 533921 43126 533933
rect 43178 533921 43184 533973
rect 670864 533921 670870 533973
rect 670922 533961 670928 533973
rect 676048 533961 676054 533973
rect 670922 533933 676054 533961
rect 670922 533921 670928 533933
rect 676048 533921 676054 533933
rect 676106 533921 676112 533973
rect 47632 532811 47638 532863
rect 47690 532851 47696 532863
rect 59536 532851 59542 532863
rect 47690 532823 59542 532851
rect 47690 532811 47696 532823
rect 59536 532811 59542 532823
rect 59594 532811 59600 532863
rect 42160 531479 42166 531531
rect 42218 531519 42224 531531
rect 42832 531519 42838 531531
rect 42218 531491 42838 531519
rect 42218 531479 42224 531491
rect 42832 531479 42838 531491
rect 42890 531479 42896 531531
rect 42064 530147 42070 530199
rect 42122 530187 42128 530199
rect 43120 530187 43126 530199
rect 42122 530159 43126 530187
rect 42122 530147 42128 530159
rect 43120 530147 43126 530159
rect 43178 530147 43184 530199
rect 672208 529999 672214 530051
rect 672266 530039 672272 530051
rect 676048 530039 676054 530051
rect 672266 530011 676054 530039
rect 672266 529999 672272 530011
rect 676048 529999 676054 530011
rect 676106 529999 676112 530051
rect 673552 529629 673558 529681
rect 673610 529669 673616 529681
rect 676240 529669 676246 529681
rect 673610 529641 676246 529669
rect 673610 529629 673616 529641
rect 676240 529629 676246 529641
rect 676298 529629 676304 529681
rect 673264 528889 673270 528941
rect 673322 528929 673328 528941
rect 676048 528929 676054 528941
rect 673322 528901 676054 528929
rect 673322 528889 673328 528901
rect 676048 528889 676054 528901
rect 676106 528889 676112 528941
rect 674704 528519 674710 528571
rect 674762 528559 674768 528571
rect 674992 528559 674998 528571
rect 674762 528531 674998 528559
rect 674762 528519 674768 528531
rect 674992 528519 674998 528531
rect 675050 528519 675056 528571
rect 672400 528445 672406 528497
rect 672458 528485 672464 528497
rect 676048 528485 676054 528497
rect 672458 528457 676054 528485
rect 672458 528445 672464 528457
rect 676048 528445 676054 528457
rect 676106 528445 676112 528497
rect 672880 528149 672886 528201
rect 672938 528189 672944 528201
rect 676240 528189 676246 528201
rect 672938 528161 676246 528189
rect 672938 528149 672944 528161
rect 676240 528149 676246 528161
rect 676298 528149 676304 528201
rect 672304 527409 672310 527461
rect 672362 527449 672368 527461
rect 676048 527449 676054 527461
rect 672362 527421 676054 527449
rect 672362 527409 672368 527421
rect 676048 527409 676054 527421
rect 676106 527409 676112 527461
rect 42160 527187 42166 527239
rect 42218 527227 42224 527239
rect 43024 527227 43030 527239
rect 42218 527199 43030 527227
rect 42218 527187 42224 527199
rect 43024 527187 43030 527199
rect 43082 527187 43088 527239
rect 42064 527039 42070 527091
rect 42122 527079 42128 527091
rect 42832 527079 42838 527091
rect 42122 527051 42838 527079
rect 42122 527039 42128 527051
rect 42832 527039 42838 527051
rect 42890 527039 42896 527091
rect 672112 526965 672118 527017
rect 672170 527005 672176 527017
rect 676048 527005 676054 527017
rect 672170 526977 676054 527005
rect 672170 526965 672176 526977
rect 676048 526965 676054 526977
rect 676106 526965 676112 527017
rect 672976 526669 672982 526721
rect 673034 526709 673040 526721
rect 676240 526709 676246 526721
rect 673034 526681 676246 526709
rect 673034 526669 673040 526681
rect 676240 526669 676246 526681
rect 676298 526669 676304 526721
rect 654448 524227 654454 524279
rect 654506 524267 654512 524279
rect 663952 524267 663958 524279
rect 654506 524239 663958 524267
rect 654506 524227 654512 524239
rect 663952 524227 663958 524239
rect 664010 524227 664016 524279
rect 661072 524153 661078 524205
rect 661130 524193 661136 524205
rect 679792 524193 679798 524205
rect 661130 524165 679798 524193
rect 661130 524153 661136 524165
rect 679792 524153 679798 524165
rect 679850 524153 679856 524205
rect 47824 518381 47830 518433
rect 47882 518421 47888 518433
rect 59536 518421 59542 518433
rect 47882 518393 59542 518421
rect 47882 518381 47888 518393
rect 59536 518381 59542 518393
rect 59594 518381 59600 518433
rect 654448 509797 654454 509849
rect 654506 509837 654512 509849
rect 672400 509837 672406 509849
rect 654506 509809 672406 509837
rect 654506 509797 654512 509809
rect 672400 509797 672406 509809
rect 672458 509797 672464 509849
rect 47728 504025 47734 504077
rect 47786 504065 47792 504077
rect 59536 504065 59542 504077
rect 47786 504037 59542 504065
rect 47786 504025 47792 504037
rect 59536 504025 59542 504037
rect 59594 504025 59600 504077
rect 676528 498253 676534 498305
rect 676586 498293 676592 498305
rect 679696 498293 679702 498305
rect 676586 498265 679702 498293
rect 676586 498253 676592 498265
rect 679696 498253 679702 498265
rect 679754 498253 679760 498305
rect 654448 495367 654454 495419
rect 654506 495407 654512 495419
rect 670096 495407 670102 495419
rect 654506 495379 670102 495407
rect 654506 495367 654512 495379
rect 670096 495367 670102 495379
rect 670154 495367 670160 495419
rect 666832 493665 666838 493717
rect 666890 493705 666896 493717
rect 676240 493705 676246 493717
rect 666890 493677 676246 493705
rect 666890 493665 666896 493677
rect 676240 493665 676246 493677
rect 676298 493665 676304 493717
rect 672496 492925 672502 492977
rect 672554 492965 672560 492977
rect 676048 492965 676054 492977
rect 672554 492937 676054 492965
rect 672554 492925 672560 492937
rect 676048 492925 676054 492937
rect 676106 492925 676112 492977
rect 50416 492481 50422 492533
rect 50474 492521 50480 492533
rect 59536 492521 59542 492533
rect 50474 492493 59542 492521
rect 50474 492481 50480 492493
rect 59536 492481 59542 492493
rect 59594 492481 59600 492533
rect 661168 492333 661174 492385
rect 661226 492373 661232 492385
rect 676048 492373 676054 492385
rect 661226 492345 676054 492373
rect 661226 492333 661232 492345
rect 676048 492333 676054 492345
rect 676106 492333 676112 492385
rect 674992 489521 674998 489573
rect 675050 489561 675056 489573
rect 676240 489561 676246 489573
rect 675050 489533 676246 489561
rect 675050 489521 675056 489533
rect 676240 489521 676246 489533
rect 676298 489521 676304 489573
rect 674608 489447 674614 489499
rect 674666 489487 674672 489499
rect 676048 489487 676054 489499
rect 674666 489459 676054 489487
rect 674666 489447 674672 489459
rect 676048 489447 676054 489459
rect 676106 489447 676112 489499
rect 674416 489373 674422 489425
rect 674474 489413 674480 489425
rect 676144 489413 676150 489425
rect 674474 489385 676150 489413
rect 674474 489373 674480 489385
rect 676144 489373 676150 489385
rect 676202 489373 676208 489425
rect 674512 486635 674518 486687
rect 674570 486675 674576 486687
rect 676048 486675 676054 486687
rect 674570 486647 676054 486675
rect 674570 486635 674576 486647
rect 676048 486635 676054 486647
rect 676106 486635 676112 486687
rect 674320 486561 674326 486613
rect 674378 486601 674384 486613
rect 676240 486601 676246 486613
rect 674378 486573 676246 486601
rect 674378 486561 674384 486573
rect 676240 486561 676246 486573
rect 676298 486561 676304 486613
rect 673840 485081 673846 485133
rect 673898 485121 673904 485133
rect 676240 485121 676246 485133
rect 673898 485093 676246 485121
rect 673898 485081 673904 485093
rect 676240 485081 676246 485093
rect 676298 485081 676304 485133
rect 673648 484489 673654 484541
rect 673706 484529 673712 484541
rect 676048 484529 676054 484541
rect 673706 484501 676054 484529
rect 673706 484489 673712 484501
rect 676048 484489 676054 484501
rect 676106 484489 676112 484541
rect 654448 484045 654454 484097
rect 654506 484085 654512 484097
rect 661456 484085 661462 484097
rect 654506 484057 661462 484085
rect 654506 484045 654512 484057
rect 661456 484045 661462 484057
rect 661514 484045 661520 484097
rect 673072 483971 673078 484023
rect 673130 484011 673136 484023
rect 676048 484011 676054 484023
rect 673130 483983 676054 484011
rect 673130 483971 673136 483983
rect 676048 483971 676054 483983
rect 676106 483971 676112 484023
rect 673744 483009 673750 483061
rect 673802 483049 673808 483061
rect 676048 483049 676054 483061
rect 673802 483021 676054 483049
rect 673802 483009 673808 483021
rect 676048 483009 676054 483021
rect 676106 483009 676112 483061
rect 673168 482417 673174 482469
rect 673226 482457 673232 482469
rect 676048 482457 676054 482469
rect 673226 482429 676054 482457
rect 673226 482417 673232 482429
rect 676048 482417 676054 482429
rect 676106 482417 676112 482469
rect 661168 479457 661174 479509
rect 661226 479497 661232 479509
rect 679984 479497 679990 479509
rect 661226 479469 679990 479497
rect 661226 479457 661232 479469
rect 679984 479457 679990 479469
rect 680042 479457 680048 479509
rect 48016 478125 48022 478177
rect 48074 478165 48080 478177
rect 59536 478165 59542 478177
rect 48074 478137 59542 478165
rect 48074 478125 48080 478137
rect 59536 478125 59542 478137
rect 59594 478125 59600 478177
rect 654448 469467 654454 469519
rect 654506 469507 654512 469519
rect 666736 469507 666742 469519
rect 654506 469479 666742 469507
rect 654506 469467 654512 469479
rect 666736 469467 666742 469479
rect 666794 469467 666800 469519
rect 53488 466581 53494 466633
rect 53546 466621 53552 466633
rect 57808 466621 57814 466633
rect 53546 466593 57814 466621
rect 53546 466581 53552 466593
rect 57808 466581 57814 466593
rect 57866 466581 57872 466633
rect 654448 455037 654454 455089
rect 654506 455077 654512 455089
rect 661552 455077 661558 455089
rect 654506 455049 661558 455077
rect 654506 455037 654512 455049
rect 661552 455037 661558 455049
rect 661610 455037 661616 455089
rect 53200 452151 53206 452203
rect 53258 452191 53264 452203
rect 59536 452191 59542 452203
rect 53258 452163 59542 452191
rect 53258 452151 53264 452163
rect 59536 452151 59542 452163
rect 59594 452151 59600 452203
rect 654448 443567 654454 443619
rect 654506 443607 654512 443619
rect 672592 443607 672598 443619
rect 654506 443579 672598 443607
rect 654506 443567 654512 443579
rect 672592 443567 672598 443579
rect 672650 443567 672656 443619
rect 47920 440681 47926 440733
rect 47978 440721 47984 440733
rect 57808 440721 57814 440733
rect 47978 440693 57814 440721
rect 47978 440681 47984 440693
rect 57808 440681 57814 440693
rect 57866 440681 57872 440733
rect 41776 432245 41782 432297
rect 41834 432285 41840 432297
rect 47632 432285 47638 432297
rect 41834 432257 47638 432285
rect 41834 432245 41840 432257
rect 47632 432245 47638 432257
rect 47690 432245 47696 432297
rect 41776 431727 41782 431779
rect 41834 431767 41840 431779
rect 47824 431767 47830 431779
rect 41834 431739 47830 431767
rect 41834 431727 41840 431739
rect 47824 431727 47830 431739
rect 47882 431727 47888 431779
rect 41584 431357 41590 431409
rect 41642 431397 41648 431409
rect 53296 431397 53302 431409
rect 41642 431369 53302 431397
rect 41642 431357 41648 431369
rect 53296 431357 53302 431369
rect 53354 431357 53360 431409
rect 41776 430765 41782 430817
rect 41834 430805 41840 430817
rect 43216 430805 43222 430817
rect 41834 430777 43222 430805
rect 41834 430765 41840 430777
rect 43216 430765 43222 430777
rect 43274 430765 43280 430817
rect 41776 430173 41782 430225
rect 41834 430213 41840 430225
rect 43312 430213 43318 430225
rect 41834 430185 43318 430213
rect 41834 430173 41840 430185
rect 43312 430173 43318 430185
rect 43370 430173 43376 430225
rect 654448 429137 654454 429189
rect 654506 429177 654512 429189
rect 663760 429177 663766 429189
rect 654506 429149 663766 429177
rect 654506 429137 654512 429149
rect 663760 429137 663766 429149
rect 663818 429137 663824 429189
rect 41584 428471 41590 428523
rect 41642 428511 41648 428523
rect 43216 428511 43222 428523
rect 41642 428483 43222 428511
rect 41642 428471 41648 428483
rect 43216 428471 43222 428483
rect 43274 428471 43280 428523
rect 53392 426251 53398 426303
rect 53450 426291 53456 426303
rect 59536 426291 59542 426303
rect 53450 426263 59542 426291
rect 53450 426251 53456 426263
rect 59536 426251 59542 426263
rect 59594 426251 59600 426303
rect 41584 421071 41590 421123
rect 41642 421111 41648 421123
rect 43024 421111 43030 421123
rect 41642 421083 43030 421111
rect 41642 421071 41648 421083
rect 43024 421071 43030 421083
rect 43082 421071 43088 421123
rect 41584 420923 41590 420975
rect 41642 420963 41648 420975
rect 42928 420963 42934 420975
rect 41642 420935 42934 420963
rect 41642 420923 41648 420935
rect 42928 420923 42934 420935
rect 42986 420923 42992 420975
rect 41968 420701 41974 420753
rect 42026 420741 42032 420753
rect 43120 420741 43126 420753
rect 42026 420713 43126 420741
rect 42026 420701 42032 420713
rect 43120 420701 43126 420713
rect 43178 420701 43184 420753
rect 41776 420479 41782 420531
rect 41834 420519 41840 420531
rect 42832 420519 42838 420531
rect 41834 420491 42838 420519
rect 41834 420479 41840 420491
rect 42832 420479 42838 420491
rect 42890 420479 42896 420531
rect 41776 419739 41782 419791
rect 41834 419779 41840 419791
rect 47632 419779 47638 419791
rect 41834 419751 47638 419779
rect 41834 419739 41840 419751
rect 47632 419739 47638 419751
rect 47690 419739 47696 419791
rect 654448 417593 654454 417645
rect 654506 417633 654512 417645
rect 672496 417633 672502 417645
rect 654506 417605 672502 417633
rect 654506 417593 654512 417605
rect 672496 417593 672502 417605
rect 672554 417593 672560 417645
rect 40720 417519 40726 417571
rect 40778 417559 40784 417571
rect 44272 417559 44278 417571
rect 40778 417531 44278 417559
rect 40778 417519 40784 417531
rect 44272 417519 44278 417531
rect 44330 417519 44336 417571
rect 50608 414707 50614 414759
rect 50666 414747 50672 414759
rect 59536 414747 59542 414759
rect 50666 414719 59542 414747
rect 50666 414707 50672 414719
rect 59536 414707 59542 414719
rect 59594 414707 59600 414759
rect 41872 413375 41878 413427
rect 41930 413375 41936 413427
rect 41890 413205 41918 413375
rect 41872 413153 41878 413205
rect 41930 413153 41936 413205
rect 42064 410489 42070 410541
rect 42122 410529 42128 410541
rect 50320 410529 50326 410541
rect 42122 410501 50326 410529
rect 42122 410489 42128 410501
rect 50320 410489 50326 410501
rect 50378 410489 50384 410541
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42832 409493 42838 409505
rect 42218 409465 42838 409493
rect 42218 409453 42224 409465
rect 42832 409453 42838 409465
rect 42890 409453 42896 409505
rect 42160 408195 42166 408247
rect 42218 408235 42224 408247
rect 42928 408235 42934 408247
rect 42218 408207 42934 408235
rect 42218 408195 42224 408207
rect 42928 408195 42934 408207
rect 42986 408195 42992 408247
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 43120 407495 43126 407507
rect 42122 407467 43126 407495
rect 42122 407455 42128 407467
rect 43120 407455 43126 407467
rect 43178 407455 43184 407507
rect 42160 406863 42166 406915
rect 42218 406903 42224 406915
rect 43024 406903 43030 406915
rect 42218 406875 43030 406903
rect 42218 406863 42224 406875
rect 43024 406863 43030 406875
rect 43082 406863 43088 406915
rect 663856 405457 663862 405509
rect 663914 405497 663920 405509
rect 676240 405497 676246 405509
rect 663914 405469 676246 405497
rect 663914 405457 663920 405469
rect 676240 405457 676246 405469
rect 676298 405457 676304 405509
rect 666640 404717 666646 404769
rect 666698 404757 666704 404769
rect 676048 404757 676054 404769
rect 666698 404729 676054 404757
rect 666698 404717 666704 404729
rect 676048 404717 676054 404729
rect 676106 404717 676112 404769
rect 663952 404199 663958 404251
rect 664010 404239 664016 404251
rect 676048 404239 676054 404251
rect 664010 404211 676054 404239
rect 664010 404199 664016 404211
rect 676048 404199 676054 404211
rect 676106 404199 676112 404251
rect 654448 403237 654454 403289
rect 654506 403277 654512 403289
rect 666832 403277 666838 403289
rect 654506 403249 666838 403277
rect 654506 403237 654512 403249
rect 666832 403237 666838 403249
rect 666890 403237 666896 403289
rect 673840 403237 673846 403289
rect 673898 403277 673904 403289
rect 676048 403277 676054 403289
rect 673898 403249 676054 403277
rect 673898 403237 673904 403249
rect 676048 403237 676054 403249
rect 676106 403237 676112 403289
rect 670864 402201 670870 402253
rect 670922 402241 670928 402253
rect 676048 402241 676054 402253
rect 670922 402213 676054 402241
rect 670922 402201 670928 402213
rect 676048 402201 676054 402213
rect 676106 402201 676112 402253
rect 676048 402053 676054 402105
rect 676106 402093 676112 402105
rect 676624 402093 676630 402105
rect 676106 402065 676630 402093
rect 676106 402053 676112 402065
rect 676624 402053 676630 402065
rect 676682 402053 676688 402105
rect 666640 401239 666646 401291
rect 666698 401279 666704 401291
rect 676048 401279 676054 401291
rect 666698 401251 676054 401279
rect 666698 401239 666704 401251
rect 676048 401239 676054 401251
rect 676106 401239 676112 401291
rect 670960 400943 670966 400995
rect 671018 400983 671024 400995
rect 676240 400983 676246 400995
rect 671018 400955 676246 400983
rect 671018 400943 671024 400955
rect 676240 400943 676246 400955
rect 676298 400943 676304 400995
rect 50320 400351 50326 400403
rect 50378 400391 50384 400403
rect 59536 400391 59542 400403
rect 50378 400363 59542 400391
rect 50378 400351 50384 400363
rect 59536 400351 59542 400363
rect 59594 400351 59600 400403
rect 674320 400351 674326 400403
rect 674378 400391 674384 400403
rect 676720 400391 676726 400403
rect 674378 400363 676726 400391
rect 674378 400351 674384 400363
rect 676720 400351 676726 400363
rect 676778 400351 676784 400403
rect 673744 395689 673750 395741
rect 673802 395729 673808 395741
rect 676048 395729 676054 395741
rect 673802 395701 676054 395729
rect 673802 395689 673808 395701
rect 676048 395689 676054 395701
rect 676106 395689 676112 395741
rect 673648 393987 673654 394039
rect 673706 394027 673712 394039
rect 676240 394027 676246 394039
rect 673706 393999 676246 394027
rect 673706 393987 673712 393999
rect 676240 393987 676246 393999
rect 676298 393987 676304 394039
rect 661264 391693 661270 391745
rect 661322 391733 661328 391745
rect 679792 391733 679798 391745
rect 661322 391705 679798 391733
rect 661322 391693 661328 391705
rect 679792 391693 679798 391705
rect 679850 391693 679856 391745
rect 654832 390731 654838 390783
rect 654890 390771 654896 390783
rect 661360 390771 661366 390783
rect 654890 390743 661366 390771
rect 654890 390731 654896 390743
rect 661360 390731 661366 390743
rect 661418 390731 661424 390783
rect 41776 389029 41782 389081
rect 41834 389069 41840 389081
rect 48016 389069 48022 389081
rect 41834 389041 48022 389069
rect 41834 389029 41840 389041
rect 48016 389029 48022 389041
rect 48074 389029 48080 389081
rect 53296 388807 53302 388859
rect 53354 388847 53360 388859
rect 59536 388847 59542 388859
rect 53354 388819 59542 388847
rect 53354 388807 53360 388819
rect 59536 388807 59542 388819
rect 59594 388807 59600 388859
rect 41584 388733 41590 388785
rect 41642 388773 41648 388785
rect 53488 388773 53494 388785
rect 41642 388745 53494 388773
rect 41642 388733 41648 388745
rect 53488 388733 53494 388745
rect 53546 388733 53552 388785
rect 41776 387993 41782 388045
rect 41834 388033 41840 388045
rect 50416 388033 50422 388045
rect 41834 388005 50422 388033
rect 41834 387993 41840 388005
rect 50416 387993 50422 388005
rect 50474 387993 50480 388045
rect 41776 387549 41782 387601
rect 41834 387589 41840 387601
rect 43312 387589 43318 387601
rect 41834 387561 43318 387589
rect 41834 387549 41840 387561
rect 43312 387549 43318 387561
rect 43370 387549 43376 387601
rect 41776 386957 41782 387009
rect 41834 386997 41840 387009
rect 43504 386997 43510 387009
rect 41834 386969 43510 386997
rect 41834 386957 41840 386969
rect 43504 386957 43510 386969
rect 43562 386957 43568 387009
rect 670192 385847 670198 385899
rect 670250 385887 670256 385899
rect 674320 385887 674326 385899
rect 670250 385859 674326 385887
rect 670250 385847 670256 385859
rect 674320 385847 674326 385859
rect 674378 385847 674384 385899
rect 41584 385181 41590 385233
rect 41642 385221 41648 385233
rect 43216 385221 43222 385233
rect 41642 385193 43222 385221
rect 41642 385181 41648 385193
rect 43216 385181 43222 385193
rect 43274 385221 43280 385233
rect 44176 385221 44182 385233
rect 43274 385193 44182 385221
rect 43274 385181 43280 385193
rect 44176 385181 44182 385193
rect 44234 385181 44240 385233
rect 34480 381555 34486 381607
rect 34538 381595 34544 381607
rect 43312 381595 43318 381607
rect 34538 381567 43318 381595
rect 34538 381555 34544 381567
rect 43312 381555 43318 381567
rect 43370 381595 43376 381607
rect 61840 381595 61846 381607
rect 43370 381567 61846 381595
rect 43370 381555 43376 381567
rect 61840 381555 61846 381567
rect 61898 381555 61904 381607
rect 41776 380075 41782 380127
rect 41834 380115 41840 380127
rect 42832 380115 42838 380127
rect 41834 380087 42838 380115
rect 41834 380075 41840 380087
rect 42832 380075 42838 380087
rect 42890 380075 42896 380127
rect 655312 378669 655318 378721
rect 655370 378709 655376 378721
rect 666640 378709 666646 378721
rect 655370 378681 666646 378709
rect 655370 378669 655376 378681
rect 666640 378669 666646 378681
rect 666698 378669 666704 378721
rect 41584 378447 41590 378499
rect 41642 378487 41648 378499
rect 43120 378487 43126 378499
rect 41642 378459 43126 378487
rect 41642 378447 41648 378459
rect 43120 378447 43126 378459
rect 43178 378447 43184 378499
rect 41776 378299 41782 378351
rect 41834 378339 41840 378351
rect 42736 378339 42742 378351
rect 41834 378311 42742 378339
rect 41834 378299 41840 378311
rect 42736 378299 42742 378311
rect 42794 378299 42800 378351
rect 41584 378225 41590 378277
rect 41642 378265 41648 378277
rect 43024 378265 43030 378277
rect 41642 378237 43030 378265
rect 41642 378225 41648 378237
rect 43024 378225 43030 378237
rect 43082 378225 43088 378277
rect 41776 377559 41782 377611
rect 41834 377599 41840 377611
rect 42928 377599 42934 377611
rect 41834 377571 42934 377599
rect 41834 377559 41840 377571
rect 42928 377559 42934 377571
rect 42986 377559 42992 377611
rect 654448 377263 654454 377315
rect 654506 377303 654512 377315
rect 670000 377303 670006 377315
rect 654506 377275 670006 377303
rect 654506 377263 654512 377275
rect 670000 377263 670006 377275
rect 670058 377263 670064 377315
rect 673744 377189 673750 377241
rect 673802 377229 673808 377241
rect 675376 377229 675382 377241
rect 673802 377201 675382 377229
rect 673802 377189 673808 377201
rect 675376 377189 675382 377201
rect 675434 377189 675440 377241
rect 673648 376819 673654 376871
rect 673706 376859 673712 376871
rect 675280 376859 675286 376871
rect 673706 376831 675286 376859
rect 673706 376819 673712 376831
rect 675280 376819 675286 376831
rect 675338 376819 675344 376871
rect 40240 376523 40246 376575
rect 40298 376563 40304 376575
rect 41776 376563 41782 376575
rect 40298 376535 41782 376563
rect 40298 376523 40304 376535
rect 41776 376523 41782 376535
rect 41834 376563 41840 376575
rect 47824 376563 47830 376575
rect 41834 376535 47830 376563
rect 41834 376523 41840 376535
rect 47824 376523 47830 376535
rect 47882 376523 47888 376575
rect 50512 374377 50518 374429
rect 50570 374417 50576 374429
rect 59440 374417 59446 374429
rect 50570 374389 59446 374417
rect 50570 374377 50576 374389
rect 59440 374377 59446 374389
rect 59498 374377 59504 374429
rect 41872 370159 41878 370211
rect 41930 370159 41936 370211
rect 41890 369989 41918 370159
rect 652624 370085 652630 370137
rect 652682 370125 652688 370137
rect 670192 370125 670198 370137
rect 652682 370097 670198 370125
rect 652682 370085 652688 370097
rect 670192 370085 670198 370097
rect 670250 370085 670256 370137
rect 41872 369937 41878 369989
rect 41930 369937 41936 369989
rect 42064 367347 42070 367399
rect 42122 367387 42128 367399
rect 47728 367387 47734 367399
rect 42122 367359 47734 367387
rect 42122 367347 42128 367359
rect 47728 367347 47734 367359
rect 47786 367347 47792 367399
rect 42064 366237 42070 366289
rect 42122 366277 42128 366289
rect 42832 366277 42838 366289
rect 42122 366249 42838 366277
rect 42122 366237 42128 366249
rect 42832 366237 42838 366249
rect 42890 366237 42896 366289
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 42928 365019 42934 365031
rect 42218 364991 42934 365019
rect 42218 364979 42224 364991
rect 42928 364979 42934 364991
rect 42986 364979 42992 365031
rect 654448 364831 654454 364883
rect 654506 364871 654512 364883
rect 663856 364871 663862 364883
rect 654506 364843 663862 364871
rect 654506 364831 654512 364843
rect 663856 364831 663862 364843
rect 663914 364831 663920 364883
rect 42064 364387 42070 364439
rect 42122 364427 42128 364439
rect 42736 364427 42742 364439
rect 42122 364399 42742 364427
rect 42122 364387 42128 364399
rect 42736 364387 42742 364399
rect 42794 364387 42800 364439
rect 42160 363647 42166 363699
rect 42218 363687 42224 363699
rect 43024 363687 43030 363699
rect 42218 363659 43030 363687
rect 42218 363647 42224 363659
rect 43024 363647 43030 363659
rect 43082 363647 43088 363699
rect 48016 362907 48022 362959
rect 48074 362947 48080 362959
rect 58384 362947 58390 362959
rect 48074 362919 58390 362947
rect 48074 362907 48080 362919
rect 58384 362907 58390 362919
rect 58442 362907 58448 362959
rect 652720 362833 652726 362885
rect 652778 362873 652784 362885
rect 655312 362873 655318 362885
rect 652778 362845 655318 362873
rect 652778 362833 652784 362845
rect 655312 362833 655318 362845
rect 655370 362833 655376 362885
rect 42160 360613 42166 360665
rect 42218 360653 42224 360665
rect 43120 360653 43126 360665
rect 42218 360625 43126 360653
rect 42218 360613 42224 360625
rect 43120 360613 43126 360625
rect 43178 360613 43184 360665
rect 670096 360021 670102 360073
rect 670154 360061 670160 360073
rect 676048 360061 676054 360073
rect 670154 360033 676054 360061
rect 670154 360021 670160 360033
rect 676048 360021 676054 360033
rect 676106 360021 676112 360073
rect 672400 359725 672406 359777
rect 672458 359765 672464 359777
rect 676240 359765 676246 359777
rect 672458 359737 676246 359765
rect 672458 359725 672464 359737
rect 676240 359725 676246 359737
rect 676298 359725 676304 359777
rect 661456 358985 661462 359037
rect 661514 359025 661520 359037
rect 676048 359025 676054 359037
rect 661514 358997 676054 359025
rect 661514 358985 661520 358997
rect 676048 358985 676054 358997
rect 676106 358985 676112 359037
rect 673840 358541 673846 358593
rect 673898 358581 673904 358593
rect 676048 358581 676054 358593
rect 673898 358553 676054 358581
rect 673898 358541 673904 358553
rect 676048 358541 676054 358553
rect 676106 358541 676112 358593
rect 670096 357727 670102 357779
rect 670154 357767 670160 357779
rect 670864 357767 670870 357779
rect 670154 357739 670870 357767
rect 670154 357727 670160 357739
rect 670864 357727 670870 357739
rect 670922 357767 670928 357779
rect 676240 357767 676246 357779
rect 670922 357739 676246 357767
rect 670922 357727 670928 357739
rect 676240 357727 676246 357739
rect 676298 357727 676304 357779
rect 670960 356543 670966 356595
rect 671018 356583 671024 356595
rect 676048 356583 676054 356595
rect 671018 356555 676054 356583
rect 671018 356543 671024 356555
rect 676048 356543 676054 356555
rect 676106 356543 676112 356595
rect 670288 354249 670294 354301
rect 670346 354289 670352 354301
rect 670960 354289 670966 354301
rect 670346 354261 670966 354289
rect 670346 354249 670352 354261
rect 670960 354249 670966 354261
rect 671018 354249 671024 354301
rect 654448 351363 654454 351415
rect 654506 351403 654512 351415
rect 666640 351403 666646 351415
rect 654506 351375 666646 351403
rect 654506 351363 654512 351375
rect 666640 351363 666646 351375
rect 666698 351363 666704 351415
rect 674800 351363 674806 351415
rect 674858 351403 674864 351415
rect 676048 351403 676054 351415
rect 674858 351375 676054 351403
rect 674858 351363 674864 351375
rect 676048 351363 676054 351375
rect 676106 351363 676112 351415
rect 673936 349883 673942 349935
rect 673994 349923 674000 349935
rect 676240 349923 676246 349935
rect 673994 349895 676246 349923
rect 673994 349883 674000 349895
rect 676240 349883 676246 349895
rect 676298 349883 676304 349935
rect 674032 349143 674038 349195
rect 674090 349183 674096 349195
rect 676048 349183 676054 349195
rect 674090 349155 676054 349183
rect 674090 349143 674096 349155
rect 676048 349143 676054 349155
rect 676106 349143 676112 349195
rect 674224 348551 674230 348603
rect 674282 348591 674288 348603
rect 676240 348591 676246 348603
rect 674282 348563 676246 348591
rect 674282 348551 674288 348563
rect 676240 348551 676246 348563
rect 676298 348551 676304 348603
rect 47728 348477 47734 348529
rect 47786 348517 47792 348529
rect 59536 348517 59542 348529
rect 47786 348489 59542 348517
rect 47786 348477 47792 348489
rect 59536 348477 59542 348489
rect 59594 348477 59600 348529
rect 674704 348477 674710 348529
rect 674762 348517 674768 348529
rect 676048 348517 676054 348529
rect 674762 348489 676054 348517
rect 674762 348477 674768 348489
rect 676048 348477 676054 348489
rect 676106 348477 676112 348529
rect 41776 345887 41782 345939
rect 41834 345927 41840 345939
rect 53392 345927 53398 345939
rect 41834 345899 53398 345927
rect 41834 345887 41840 345899
rect 53392 345887 53398 345899
rect 53450 345887 53456 345939
rect 658576 345591 658582 345643
rect 658634 345631 658640 345643
rect 679792 345631 679798 345643
rect 658634 345603 679798 345631
rect 658634 345591 658640 345603
rect 679792 345591 679798 345603
rect 679850 345591 679856 345643
rect 41584 345517 41590 345569
rect 41642 345557 41648 345569
rect 50608 345557 50614 345569
rect 41642 345529 50614 345557
rect 41642 345517 41648 345529
rect 50608 345517 50614 345529
rect 50666 345517 50672 345569
rect 41776 344777 41782 344829
rect 41834 344817 41840 344829
rect 47920 344817 47926 344829
rect 41834 344789 47926 344817
rect 41834 344777 41840 344789
rect 47920 344777 47926 344789
rect 47978 344777 47984 344829
rect 41776 344333 41782 344385
rect 41834 344373 41840 344385
rect 43504 344373 43510 344385
rect 41834 344345 43510 344373
rect 41834 344333 41840 344345
rect 43504 344333 43510 344345
rect 43562 344333 43568 344385
rect 41776 343815 41782 343867
rect 41834 343855 41840 343867
rect 43216 343855 43222 343867
rect 41834 343827 43222 343855
rect 41834 343815 41840 343827
rect 43216 343815 43222 343827
rect 43274 343815 43280 343867
rect 41776 343297 41782 343349
rect 41834 343337 41840 343349
rect 43408 343337 43414 343349
rect 41834 343309 43414 343337
rect 41834 343297 41840 343309
rect 43408 343297 43414 343309
rect 43466 343337 43472 343349
rect 45328 343337 45334 343349
rect 43466 343309 45334 343337
rect 43466 343297 43472 343309
rect 45328 343297 45334 343309
rect 45386 343297 45392 343349
rect 41776 342335 41782 342387
rect 41834 342375 41840 342387
rect 43504 342375 43510 342387
rect 41834 342347 43510 342375
rect 41834 342335 41840 342347
rect 43504 342335 43510 342347
rect 43562 342375 43568 342387
rect 45232 342375 45238 342387
rect 43562 342347 45238 342375
rect 43562 342335 43568 342347
rect 45232 342335 45238 342347
rect 45290 342335 45296 342387
rect 41584 341965 41590 342017
rect 41642 342005 41648 342017
rect 43312 342005 43318 342017
rect 41642 341977 43318 342005
rect 41642 341965 41648 341977
rect 43312 341965 43318 341977
rect 43370 341965 43376 342017
rect 675760 341151 675766 341203
rect 675818 341151 675824 341203
rect 675778 340981 675806 341151
rect 675760 340929 675766 340981
rect 675818 340929 675824 340981
rect 674800 337895 674806 337947
rect 674858 337935 674864 337947
rect 675472 337935 675478 337947
rect 674858 337907 675478 337935
rect 674858 337895 674864 337907
rect 675472 337895 675478 337907
rect 675530 337895 675536 337947
rect 50416 337007 50422 337059
rect 50474 337047 50480 337059
rect 59536 337047 59542 337059
rect 50474 337019 59542 337047
rect 50474 337007 50480 337019
rect 59536 337007 59542 337019
rect 59594 337007 59600 337059
rect 674224 336045 674230 336097
rect 674282 336085 674288 336097
rect 675376 336085 675382 336097
rect 674282 336057 675382 336085
rect 674282 336045 674288 336057
rect 675376 336045 675382 336057
rect 675434 336045 675440 336097
rect 41584 335231 41590 335283
rect 41642 335271 41648 335283
rect 43120 335271 43126 335283
rect 41642 335243 43126 335271
rect 41642 335231 41648 335243
rect 43120 335231 43126 335243
rect 43178 335231 43184 335283
rect 41776 334935 41782 334987
rect 41834 334975 41840 334987
rect 42928 334975 42934 334987
rect 41834 334947 42934 334975
rect 41834 334935 41840 334947
rect 42928 334935 42934 334947
rect 42986 334935 42992 334987
rect 41584 334639 41590 334691
rect 41642 334679 41648 334691
rect 43024 334679 43030 334691
rect 41642 334651 43030 334679
rect 41642 334639 41648 334651
rect 43024 334639 43030 334651
rect 43082 334639 43088 334691
rect 41776 334491 41782 334543
rect 41834 334531 41840 334543
rect 42832 334531 42838 334543
rect 41834 334503 42838 334531
rect 41834 334491 41840 334503
rect 42832 334491 42838 334503
rect 42890 334491 42896 334543
rect 41776 333307 41782 333359
rect 41834 333347 41840 333359
rect 47920 333347 47926 333359
rect 41834 333319 47926 333347
rect 41834 333307 41840 333319
rect 47920 333307 47926 333319
rect 47978 333307 47984 333359
rect 674032 332715 674038 332767
rect 674090 332755 674096 332767
rect 675376 332755 675382 332767
rect 674090 332727 675382 332755
rect 674090 332715 674096 332727
rect 675376 332715 675382 332727
rect 675434 332715 675440 332767
rect 673936 332197 673942 332249
rect 673994 332237 674000 332249
rect 675472 332237 675478 332249
rect 673994 332209 675478 332237
rect 673994 332197 674000 332209
rect 675472 332197 675478 332209
rect 675530 332197 675536 332249
rect 674704 331753 674710 331805
rect 674762 331793 674768 331805
rect 675376 331793 675382 331805
rect 674762 331765 675382 331793
rect 674762 331753 674768 331765
rect 675376 331753 675382 331765
rect 675434 331753 675440 331805
rect 41872 327017 41878 327069
rect 41930 327017 41936 327069
rect 41890 326773 41918 327017
rect 41872 326721 41878 326773
rect 41930 326721 41936 326773
rect 43024 326647 43030 326699
rect 43082 326687 43088 326699
rect 43312 326687 43318 326699
rect 43082 326659 43318 326687
rect 43082 326647 43088 326659
rect 43312 326647 43318 326659
rect 43370 326647 43376 326699
rect 42448 326499 42454 326551
rect 42506 326539 42512 326551
rect 43024 326539 43030 326551
rect 42506 326511 43030 326539
rect 42506 326499 42512 326511
rect 43024 326499 43030 326511
rect 43082 326499 43088 326551
rect 42160 324131 42166 324183
rect 42218 324171 42224 324183
rect 53200 324171 53206 324183
rect 42218 324143 53206 324171
rect 42218 324131 42224 324143
rect 53200 324131 53206 324143
rect 53258 324131 53264 324183
rect 654832 323243 654838 323295
rect 654890 323283 654896 323295
rect 661456 323283 661462 323295
rect 654890 323255 661462 323283
rect 654890 323243 654896 323255
rect 661456 323243 661462 323255
rect 661514 323243 661520 323295
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 42928 323135 42934 323147
rect 42218 323107 42934 323135
rect 42218 323095 42224 323107
rect 42928 323095 42934 323107
rect 42986 323095 42992 323147
rect 42928 322947 42934 322999
rect 42986 322987 42992 322999
rect 43312 322987 43318 322999
rect 42986 322959 43318 322987
rect 42986 322947 42992 322959
rect 43312 322947 43318 322959
rect 43370 322947 43376 322999
rect 53392 322577 53398 322629
rect 53450 322617 53456 322629
rect 59536 322617 59542 322629
rect 53450 322589 59542 322617
rect 53450 322577 53456 322589
rect 59536 322577 59542 322589
rect 59594 322577 59600 322629
rect 42064 321763 42070 321815
rect 42122 321803 42128 321815
rect 42832 321803 42838 321815
rect 42122 321775 42838 321803
rect 42122 321763 42128 321775
rect 42832 321763 42838 321775
rect 42890 321763 42896 321815
rect 42160 321023 42166 321075
rect 42218 321063 42224 321075
rect 43120 321063 43126 321075
rect 42218 321035 43126 321063
rect 42218 321023 42224 321035
rect 43120 321023 43126 321035
rect 43178 321023 43184 321075
rect 42160 320579 42166 320631
rect 42218 320619 42224 320631
rect 42928 320619 42934 320631
rect 42218 320591 42934 320619
rect 42218 320579 42224 320591
rect 42928 320579 42934 320591
rect 42986 320579 42992 320631
rect 43408 318359 43414 318411
rect 43466 318359 43472 318411
rect 43426 318189 43454 318359
rect 43408 318137 43414 318189
rect 43466 318137 43472 318189
rect 42160 317471 42166 317523
rect 42218 317511 42224 317523
rect 43024 317511 43030 317523
rect 42218 317483 43030 317511
rect 42218 317471 42224 317483
rect 43024 317471 43030 317483
rect 43082 317471 43088 317523
rect 45712 316065 45718 316117
rect 45770 316105 45776 316117
rect 49264 316105 49270 316117
rect 45770 316077 49270 316105
rect 45770 316065 45776 316077
rect 49264 316065 49270 316077
rect 49322 316065 49328 316117
rect 661552 315029 661558 315081
rect 661610 315069 661616 315081
rect 676048 315069 676054 315081
rect 661610 315041 676054 315069
rect 661610 315029 661616 315041
rect 676048 315029 676054 315041
rect 676106 315029 676112 315081
rect 666736 314733 666742 314785
rect 666794 314773 666800 314785
rect 676240 314773 676246 314785
rect 666794 314745 676246 314773
rect 666794 314733 666800 314745
rect 676240 314733 676246 314745
rect 676298 314733 676304 314785
rect 672592 313993 672598 314045
rect 672650 314033 672656 314045
rect 676048 314033 676054 314045
rect 672650 314005 676054 314033
rect 672650 313993 672656 314005
rect 676048 313993 676054 314005
rect 676106 313993 676112 314045
rect 45232 311033 45238 311085
rect 45290 311073 45296 311085
rect 58576 311073 58582 311085
rect 45290 311045 58582 311073
rect 45290 311033 45296 311045
rect 58576 311033 58582 311045
rect 58634 311033 58640 311085
rect 654448 311033 654454 311085
rect 654506 311073 654512 311085
rect 672400 311073 672406 311085
rect 654506 311045 672406 311073
rect 654506 311033 654512 311045
rect 672400 311033 672406 311045
rect 672458 311033 672464 311085
rect 674320 309627 674326 309679
rect 674378 309667 674384 309679
rect 676048 309667 676054 309679
rect 674378 309639 676054 309667
rect 674378 309627 674384 309639
rect 676048 309627 676054 309639
rect 676106 309627 676112 309679
rect 674224 308147 674230 308199
rect 674282 308187 674288 308199
rect 676048 308187 676054 308199
rect 674282 308159 676054 308187
rect 674282 308147 674288 308159
rect 676048 308147 676054 308159
rect 676106 308147 676112 308199
rect 674128 306371 674134 306423
rect 674186 306411 674192 306423
rect 676240 306411 676246 306423
rect 674186 306383 676246 306411
rect 674186 306371 674192 306383
rect 676240 306371 676246 306383
rect 676298 306371 676304 306423
rect 674032 305335 674038 305387
rect 674090 305375 674096 305387
rect 676240 305375 676246 305387
rect 674090 305347 676246 305375
rect 674090 305335 674096 305347
rect 676240 305335 676246 305347
rect 676298 305335 676304 305387
rect 45808 305261 45814 305313
rect 45866 305301 45872 305313
rect 45866 305273 54734 305301
rect 45866 305261 45872 305273
rect 49264 305187 49270 305239
rect 49322 305227 49328 305239
rect 53200 305227 53206 305239
rect 49322 305199 53206 305227
rect 49322 305187 49328 305199
rect 53200 305187 53206 305199
rect 53258 305187 53264 305239
rect 54706 305227 54734 305273
rect 674512 305261 674518 305313
rect 674570 305301 674576 305313
rect 676048 305301 676054 305313
rect 674570 305273 676054 305301
rect 674570 305261 674576 305273
rect 676048 305261 676054 305273
rect 676106 305261 676112 305313
rect 58960 305227 58966 305239
rect 54706 305199 58966 305227
rect 58960 305187 58966 305199
rect 59018 305187 59024 305239
rect 41776 302671 41782 302723
rect 41834 302711 41840 302723
rect 50512 302711 50518 302723
rect 41834 302683 50518 302711
rect 41834 302671 41840 302683
rect 50512 302671 50518 302683
rect 50570 302671 50576 302723
rect 44368 302523 44374 302575
rect 44426 302563 44432 302575
rect 53680 302563 53686 302575
rect 44426 302535 53686 302563
rect 44426 302523 44432 302535
rect 53680 302523 53686 302535
rect 53738 302523 53744 302575
rect 658672 302523 658678 302575
rect 658730 302563 658736 302575
rect 679888 302563 679894 302575
rect 658730 302535 679894 302563
rect 658730 302523 658736 302535
rect 679888 302523 679894 302535
rect 679946 302523 679952 302575
rect 673936 302449 673942 302501
rect 673994 302489 674000 302501
rect 676048 302489 676054 302501
rect 673994 302461 676054 302489
rect 673994 302449 674000 302461
rect 676048 302449 676054 302461
rect 676106 302449 676112 302501
rect 674416 302375 674422 302427
rect 674474 302415 674480 302427
rect 676240 302415 676246 302427
rect 674474 302387 676246 302415
rect 674474 302375 674480 302387
rect 676240 302375 676246 302387
rect 676298 302375 676304 302427
rect 41584 302301 41590 302353
rect 41642 302341 41648 302353
rect 48016 302341 48022 302353
rect 41642 302313 48022 302341
rect 41642 302301 41648 302313
rect 48016 302301 48022 302313
rect 48074 302301 48080 302353
rect 41776 301561 41782 301613
rect 41834 301601 41840 301613
rect 53296 301601 53302 301613
rect 41834 301573 53302 301601
rect 41834 301561 41840 301573
rect 53296 301561 53302 301573
rect 53354 301561 53360 301613
rect 41776 301191 41782 301243
rect 41834 301231 41840 301243
rect 43216 301231 43222 301243
rect 41834 301203 43222 301231
rect 41834 301191 41840 301203
rect 43216 301191 43222 301203
rect 43274 301191 43280 301243
rect 53680 301117 53686 301169
rect 53738 301157 53744 301169
rect 55312 301157 55318 301169
rect 53738 301129 55318 301157
rect 53738 301117 53744 301129
rect 55312 301117 55318 301129
rect 55370 301117 55376 301169
rect 41776 300599 41782 300651
rect 41834 300639 41840 300651
rect 43600 300639 43606 300651
rect 41834 300611 43606 300639
rect 41834 300599 41840 300611
rect 43600 300599 43606 300611
rect 43658 300599 43664 300651
rect 41776 300081 41782 300133
rect 41834 300121 41840 300133
rect 43504 300121 43510 300133
rect 41834 300093 43510 300121
rect 41834 300081 41840 300093
rect 43504 300081 43510 300093
rect 43562 300121 43568 300133
rect 45136 300121 45142 300133
rect 43562 300093 45142 300121
rect 43562 300081 43568 300093
rect 45136 300081 45142 300093
rect 45194 300081 45200 300133
rect 41776 299637 41782 299689
rect 41834 299677 41840 299689
rect 43408 299677 43414 299689
rect 41834 299649 43414 299677
rect 41834 299637 41840 299649
rect 43408 299637 43414 299649
rect 43466 299637 43472 299689
rect 41584 299341 41590 299393
rect 41642 299381 41648 299393
rect 43216 299381 43222 299393
rect 41642 299353 43222 299381
rect 41642 299341 41648 299353
rect 43216 299341 43222 299353
rect 43274 299381 43280 299393
rect 44944 299381 44950 299393
rect 43274 299353 44950 299381
rect 43274 299341 43280 299353
rect 44944 299341 44950 299353
rect 45002 299341 45008 299393
rect 41776 298601 41782 298653
rect 41834 298641 41840 298653
rect 43312 298641 43318 298653
rect 41834 298613 43318 298641
rect 41834 298601 41840 298613
rect 43312 298601 43318 298613
rect 43370 298601 43376 298653
rect 45136 296677 45142 296729
rect 45194 296717 45200 296729
rect 59536 296717 59542 296729
rect 45194 296689 59542 296717
rect 45194 296677 45200 296689
rect 59536 296677 59542 296689
rect 59594 296677 59600 296729
rect 674224 295937 674230 295989
rect 674282 295977 674288 295989
rect 675376 295977 675382 295989
rect 674282 295949 675382 295977
rect 674282 295937 674288 295949
rect 675376 295937 675382 295949
rect 675434 295937 675440 295989
rect 674512 295345 674518 295397
rect 674570 295385 674576 295397
rect 675472 295385 675478 295397
rect 674570 295357 675478 295385
rect 674570 295345 674576 295357
rect 675472 295345 675478 295357
rect 675530 295345 675536 295397
rect 674320 294531 674326 294583
rect 674378 294571 674384 294583
rect 675376 294571 675382 294583
rect 674378 294543 675382 294571
rect 674378 294531 674384 294543
rect 675376 294531 675382 294543
rect 675434 294531 675440 294583
rect 44272 293791 44278 293843
rect 44330 293831 44336 293843
rect 44330 293803 54734 293831
rect 44330 293791 44336 293803
rect 54706 293757 54734 293803
rect 55312 293791 55318 293843
rect 55370 293831 55376 293843
rect 60304 293831 60310 293843
rect 55370 293803 60310 293831
rect 55370 293791 55376 293803
rect 60304 293791 60310 293803
rect 60362 293791 60368 293843
rect 60400 293757 60406 293769
rect 54706 293729 60406 293757
rect 60400 293717 60406 293729
rect 60458 293717 60464 293769
rect 41872 292311 41878 292363
rect 41930 292351 41936 292363
rect 43120 292351 43126 292363
rect 41930 292323 43126 292351
rect 41930 292311 41936 292323
rect 43120 292311 43126 292323
rect 43178 292311 43184 292363
rect 674128 292015 674134 292067
rect 674186 292055 674192 292067
rect 675472 292055 675478 292067
rect 674186 292027 675478 292055
rect 674186 292015 674192 292027
rect 675472 292015 675478 292027
rect 675530 292015 675536 292067
rect 41584 291571 41590 291623
rect 41642 291611 41648 291623
rect 43024 291611 43030 291623
rect 41642 291583 43030 291611
rect 41642 291571 41648 291583
rect 43024 291571 43030 291583
rect 43082 291571 43088 291623
rect 674032 291571 674038 291623
rect 674090 291611 674096 291623
rect 675376 291611 675382 291623
rect 674090 291583 675382 291611
rect 674090 291571 674096 291583
rect 675376 291571 675382 291583
rect 675434 291571 675440 291623
rect 41584 291127 41590 291179
rect 41642 291167 41648 291179
rect 42736 291167 42742 291179
rect 41642 291139 42742 291167
rect 41642 291127 41648 291139
rect 42736 291127 42742 291139
rect 42794 291127 42800 291179
rect 41872 291053 41878 291105
rect 41930 291093 41936 291105
rect 42928 291093 42934 291105
rect 41930 291065 42934 291093
rect 41930 291053 41936 291065
rect 42928 291053 42934 291065
rect 42986 291053 42992 291105
rect 674416 291053 674422 291105
rect 674474 291093 674480 291105
rect 675376 291093 675382 291105
rect 674474 291065 675382 291093
rect 674474 291053 674480 291065
rect 675376 291053 675382 291065
rect 675434 291053 675440 291105
rect 41776 290905 41782 290957
rect 41834 290945 41840 290957
rect 42832 290945 42838 290957
rect 41834 290917 42838 290945
rect 41834 290905 41840 290917
rect 42832 290905 42838 290917
rect 42890 290905 42896 290957
rect 53200 290905 53206 290957
rect 53258 290945 53264 290957
rect 57520 290945 57526 290957
rect 53258 290917 57526 290945
rect 53258 290905 53264 290917
rect 57520 290905 57526 290917
rect 57578 290905 57584 290957
rect 41776 290091 41782 290143
rect 41834 290131 41840 290143
rect 48016 290131 48022 290143
rect 41834 290103 48022 290131
rect 41834 290091 41840 290103
rect 48016 290091 48022 290103
rect 48074 290091 48080 290143
rect 673936 286539 673942 286591
rect 673994 286579 674000 286591
rect 675376 286579 675382 286591
rect 673994 286551 675382 286579
rect 673994 286539 674000 286551
rect 675376 286539 675382 286551
rect 675434 286539 675440 286591
rect 57520 285207 57526 285259
rect 57578 285247 57584 285259
rect 63280 285247 63286 285259
rect 57578 285219 63286 285247
rect 57578 285207 57584 285219
rect 63280 285207 63286 285219
rect 63338 285207 63344 285259
rect 44944 285133 44950 285185
rect 45002 285173 45008 285185
rect 59536 285173 59542 285185
rect 45002 285145 59542 285173
rect 45002 285133 45008 285145
rect 59536 285133 59542 285145
rect 59594 285133 59600 285185
rect 47536 285059 47542 285111
rect 47594 285099 47600 285111
rect 60400 285099 60406 285111
rect 47594 285071 60406 285099
rect 47594 285059 47600 285071
rect 60400 285059 60406 285071
rect 60458 285059 60464 285111
rect 41968 283801 41974 283853
rect 42026 283801 42032 283853
rect 41986 283557 42014 283801
rect 41968 283505 41974 283557
rect 42026 283505 42032 283557
rect 42160 281063 42166 281115
rect 42218 281103 42224 281115
rect 50320 281103 50326 281115
rect 42218 281075 50326 281103
rect 42218 281063 42224 281075
rect 50320 281063 50326 281075
rect 50378 281063 50384 281115
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 42832 279919 42838 279931
rect 42218 279891 42838 279919
rect 42218 279879 42224 279891
rect 42832 279879 42838 279891
rect 42890 279879 42896 279931
rect 60304 278621 60310 278673
rect 60362 278661 60368 278673
rect 652912 278661 652918 278673
rect 60362 278633 652918 278661
rect 60362 278621 60368 278633
rect 652912 278621 652918 278633
rect 652970 278621 652976 278673
rect 42160 278547 42166 278599
rect 42218 278587 42224 278599
rect 42736 278587 42742 278599
rect 42218 278559 42742 278587
rect 42218 278547 42224 278559
rect 42736 278547 42742 278559
rect 42794 278547 42800 278599
rect 58960 278547 58966 278599
rect 59018 278587 59024 278599
rect 652720 278587 652726 278599
rect 59018 278559 652726 278587
rect 59018 278547 59024 278559
rect 652720 278547 652726 278559
rect 652778 278547 652784 278599
rect 60496 278473 60502 278525
rect 60554 278513 60560 278525
rect 653008 278513 653014 278525
rect 60554 278485 653014 278513
rect 60554 278473 60560 278485
rect 653008 278473 653014 278485
rect 653066 278473 653072 278525
rect 60592 278399 60598 278451
rect 60650 278439 60656 278451
rect 652528 278439 652534 278451
rect 60650 278411 652534 278439
rect 60650 278399 60656 278411
rect 652528 278399 652534 278411
rect 652586 278399 652592 278451
rect 320944 278029 320950 278081
rect 321002 278069 321008 278081
rect 422512 278069 422518 278081
rect 321002 278041 422518 278069
rect 321002 278029 321008 278041
rect 422512 278029 422518 278041
rect 422570 278029 422576 278081
rect 317872 277955 317878 278007
rect 317930 277995 317936 278007
rect 415408 277995 415414 278007
rect 317930 277967 415414 277995
rect 317930 277955 317936 277967
rect 415408 277955 415414 277967
rect 415466 277955 415472 278007
rect 319504 277881 319510 277933
rect 319562 277921 319568 277933
rect 419056 277921 419062 277933
rect 319562 277893 419062 277921
rect 319562 277881 319568 277893
rect 419056 277881 419062 277893
rect 419114 277881 419120 277933
rect 42160 277807 42166 277859
rect 42218 277847 42224 277859
rect 43024 277847 43030 277859
rect 42218 277819 43030 277847
rect 42218 277807 42224 277819
rect 43024 277807 43030 277819
rect 43082 277807 43088 277859
rect 322096 277807 322102 277859
rect 322154 277847 322160 277859
rect 426256 277847 426262 277859
rect 322154 277819 426262 277847
rect 322154 277807 322160 277819
rect 426256 277807 426262 277819
rect 426314 277807 426320 277859
rect 323824 277733 323830 277785
rect 323882 277773 323888 277785
rect 429616 277773 429622 277785
rect 323882 277745 429622 277773
rect 323882 277733 323888 277745
rect 429616 277733 429622 277745
rect 429674 277733 429680 277785
rect 324976 277659 324982 277711
rect 325034 277699 325040 277711
rect 433456 277699 433462 277711
rect 325034 277671 433462 277699
rect 325034 277659 325040 277671
rect 433456 277659 433462 277671
rect 433514 277659 433520 277711
rect 328048 277585 328054 277637
rect 328106 277625 328112 277637
rect 440560 277625 440566 277637
rect 328106 277597 440566 277625
rect 328106 277585 328112 277597
rect 440560 277585 440566 277597
rect 440618 277585 440624 277637
rect 408016 277511 408022 277563
rect 408074 277551 408080 277563
rect 546640 277551 546646 277563
rect 408074 277523 546646 277551
rect 408074 277511 408080 277523
rect 546640 277511 546646 277523
rect 546698 277511 546704 277563
rect 316624 277437 316630 277489
rect 316682 277477 316688 277489
rect 412240 277477 412246 277489
rect 316682 277449 412246 277477
rect 316682 277437 316688 277449
rect 412240 277437 412246 277449
rect 412298 277437 412304 277489
rect 42064 277363 42070 277415
rect 42122 277403 42128 277415
rect 42928 277403 42934 277415
rect 42122 277375 42934 277403
rect 42122 277363 42128 277375
rect 42928 277363 42934 277375
rect 42986 277363 42992 277415
rect 326416 277363 326422 277415
rect 326474 277403 326480 277415
rect 437008 277403 437014 277415
rect 326474 277375 437014 277403
rect 326474 277363 326480 277375
rect 437008 277363 437014 277375
rect 437066 277363 437072 277415
rect 329296 277289 329302 277341
rect 329354 277329 329360 277341
rect 444208 277329 444214 277341
rect 329354 277301 444214 277329
rect 329354 277289 329360 277301
rect 444208 277289 444214 277301
rect 444266 277289 444272 277341
rect 332368 277215 332374 277267
rect 332426 277255 332432 277267
rect 451216 277255 451222 277267
rect 332426 277227 451222 277255
rect 332426 277215 332432 277227
rect 451216 277215 451222 277227
rect 451274 277215 451280 277267
rect 330736 277141 330742 277193
rect 330794 277181 330800 277193
rect 447664 277181 447670 277193
rect 330794 277153 447670 277181
rect 330794 277141 330800 277153
rect 447664 277141 447670 277153
rect 447722 277141 447728 277193
rect 333616 277067 333622 277119
rect 333674 277107 333680 277119
rect 454768 277107 454774 277119
rect 333674 277079 454774 277107
rect 333674 277067 333680 277079
rect 454768 277067 454774 277079
rect 454826 277067 454832 277119
rect 336688 276993 336694 277045
rect 336746 277033 336752 277045
rect 461872 277033 461878 277045
rect 336746 277005 461878 277033
rect 336746 276993 336752 277005
rect 461872 276993 461878 277005
rect 461930 276993 461936 277045
rect 405424 276919 405430 276971
rect 405482 276959 405488 276971
rect 612976 276959 612982 276971
rect 405482 276931 612982 276959
rect 405482 276919 405488 276931
rect 612976 276919 612982 276931
rect 613034 276919 613040 276971
rect 393904 276845 393910 276897
rect 393962 276885 393968 276897
rect 603664 276885 603670 276897
rect 393962 276857 603670 276885
rect 393962 276845 393968 276857
rect 603664 276845 603670 276857
rect 603722 276845 603728 276897
rect 396784 276771 396790 276823
rect 396842 276811 396848 276823
rect 610768 276811 610774 276823
rect 396842 276783 610774 276811
rect 396842 276771 396848 276783
rect 610768 276771 610774 276783
rect 610826 276771 610832 276823
rect 398224 276697 398230 276749
rect 398282 276737 398288 276749
rect 614416 276737 614422 276749
rect 398282 276709 614422 276737
rect 398282 276697 398288 276709
rect 614416 276697 614422 276709
rect 614474 276697 614480 276749
rect 401104 276623 401110 276675
rect 401162 276663 401168 276675
rect 621424 276663 621430 276675
rect 401162 276635 621430 276663
rect 401162 276623 401168 276635
rect 621424 276623 621430 276635
rect 621482 276623 621488 276675
rect 399376 276549 399382 276601
rect 399434 276589 399440 276601
rect 617968 276589 617974 276601
rect 399434 276561 617974 276589
rect 399434 276549 399440 276561
rect 617968 276549 617974 276561
rect 618026 276549 618032 276601
rect 402544 276475 402550 276527
rect 402602 276515 402608 276527
rect 625072 276515 625078 276527
rect 402602 276487 625078 276515
rect 402602 276475 402608 276487
rect 625072 276475 625078 276487
rect 625130 276475 625136 276527
rect 350224 276401 350230 276453
rect 350282 276441 350288 276453
rect 496144 276441 496150 276453
rect 350282 276413 496150 276441
rect 350282 276401 350288 276413
rect 496144 276401 496150 276413
rect 496202 276401 496208 276453
rect 353392 276327 353398 276379
rect 353450 276367 353456 276379
rect 503248 276367 503254 276379
rect 353450 276339 503254 276367
rect 353450 276327 353456 276339
rect 503248 276327 503254 276339
rect 503306 276327 503312 276379
rect 357424 276253 357430 276305
rect 357482 276293 357488 276305
rect 513904 276293 513910 276305
rect 357482 276265 513910 276293
rect 357482 276253 357488 276265
rect 513904 276253 513910 276265
rect 513962 276253 513968 276305
rect 293008 276179 293014 276231
rect 293066 276219 293072 276231
rect 354256 276219 354262 276231
rect 293066 276191 354262 276219
rect 293066 276179 293072 276191
rect 354256 276179 354262 276191
rect 354314 276179 354320 276231
rect 356176 276179 356182 276231
rect 356234 276219 356240 276231
rect 510352 276219 510358 276231
rect 356234 276191 510358 276219
rect 356234 276179 356240 276191
rect 510352 276179 510358 276191
rect 510410 276179 510416 276231
rect 294640 276105 294646 276157
rect 294698 276145 294704 276157
rect 357904 276145 357910 276157
rect 294698 276117 357910 276145
rect 294698 276105 294704 276117
rect 357904 276105 357910 276117
rect 357962 276105 357968 276157
rect 360304 276105 360310 276157
rect 360362 276145 360368 276157
rect 521008 276145 521014 276157
rect 360362 276117 521014 276145
rect 360362 276105 360368 276117
rect 521008 276105 521014 276117
rect 521066 276105 521072 276157
rect 295888 276031 295894 276083
rect 295946 276071 295952 276083
rect 361360 276071 361366 276083
rect 295946 276043 361366 276071
rect 295946 276031 295952 276043
rect 361360 276031 361366 276043
rect 361418 276031 361424 276083
rect 363376 276031 363382 276083
rect 363434 276071 363440 276083
rect 528112 276071 528118 276083
rect 363434 276043 528118 276071
rect 363434 276031 363440 276043
rect 528112 276031 528118 276043
rect 528170 276031 528176 276083
rect 297328 275957 297334 276009
rect 297386 275997 297392 276009
rect 364912 275997 364918 276009
rect 297386 275969 364918 275997
rect 297386 275957 297392 275969
rect 364912 275957 364918 275969
rect 364970 275957 364976 276009
rect 365968 275957 365974 276009
rect 366026 275997 366032 276009
rect 535120 275997 535126 276009
rect 366026 275969 535126 275997
rect 366026 275957 366032 275969
rect 535120 275957 535126 275969
rect 535178 275957 535184 276009
rect 298960 275883 298966 275935
rect 299018 275923 299024 275935
rect 368464 275923 368470 275935
rect 299018 275895 368470 275923
rect 299018 275883 299024 275895
rect 368464 275883 368470 275895
rect 368522 275883 368528 275935
rect 372496 275883 372502 275935
rect 372554 275923 372560 275935
rect 550480 275923 550486 275935
rect 372554 275895 550486 275923
rect 372554 275883 372560 275895
rect 550480 275883 550486 275895
rect 550538 275883 550544 275935
rect 300208 275809 300214 275861
rect 300266 275849 300272 275861
rect 372016 275849 372022 275861
rect 300266 275821 372022 275849
rect 300266 275809 300272 275821
rect 372016 275809 372022 275821
rect 372074 275809 372080 275861
rect 375088 275809 375094 275861
rect 375146 275849 375152 275861
rect 557584 275849 557590 275861
rect 375146 275821 557590 275849
rect 375146 275809 375152 275821
rect 557584 275809 557590 275821
rect 557642 275809 557648 275861
rect 301744 275735 301750 275787
rect 301802 275775 301808 275787
rect 375568 275775 375574 275787
rect 301802 275747 375574 275775
rect 301802 275735 301808 275747
rect 375568 275735 375574 275747
rect 375626 275735 375632 275787
rect 380560 275735 380566 275787
rect 380618 275775 380624 275787
rect 380618 275747 399038 275775
rect 380618 275735 380624 275747
rect 303280 275661 303286 275713
rect 303338 275701 303344 275713
rect 379120 275701 379126 275713
rect 303338 275673 379126 275701
rect 303338 275661 303344 275673
rect 379120 275661 379126 275673
rect 379178 275661 379184 275713
rect 381040 275661 381046 275713
rect 381098 275701 381104 275713
rect 399010 275701 399038 275747
rect 399088 275735 399094 275787
rect 399146 275775 399152 275787
rect 564688 275775 564694 275787
rect 399146 275747 564694 275775
rect 399146 275735 399152 275747
rect 564688 275735 564694 275747
rect 564746 275735 564752 275787
rect 570640 275701 570646 275713
rect 381098 275673 398942 275701
rect 399010 275673 570646 275701
rect 381098 275661 381104 275673
rect 303760 275587 303766 275639
rect 303818 275627 303824 275639
rect 380368 275627 380374 275639
rect 303818 275599 380374 275627
rect 303818 275587 303824 275599
rect 380368 275587 380374 275599
rect 380426 275587 380432 275639
rect 383440 275587 383446 275639
rect 383498 275627 383504 275639
rect 398914 275627 398942 275673
rect 570640 275661 570646 275673
rect 570698 275661 570704 275713
rect 571792 275627 571798 275639
rect 383498 275599 398846 275627
rect 398914 275599 571798 275627
rect 383498 275587 383504 275599
rect 304432 275513 304438 275565
rect 304490 275553 304496 275565
rect 382576 275553 382582 275565
rect 304490 275525 382582 275553
rect 304490 275513 304496 275525
rect 382576 275513 382582 275525
rect 382634 275513 382640 275565
rect 386512 275513 386518 275565
rect 386570 275553 386576 275565
rect 398818 275553 398846 275599
rect 571792 275587 571798 275599
rect 571850 275587 571856 275639
rect 577744 275553 577750 275565
rect 386570 275525 398750 275553
rect 398818 275525 577750 275553
rect 386570 275513 386576 275525
rect 305008 275439 305014 275491
rect 305066 275479 305072 275491
rect 383824 275479 383830 275491
rect 305066 275451 383830 275479
rect 305066 275439 305072 275451
rect 383824 275439 383830 275451
rect 383882 275439 383888 275491
rect 398722 275479 398750 275525
rect 577744 275513 577750 275525
rect 577802 275513 577808 275565
rect 586000 275479 586006 275491
rect 398722 275451 586006 275479
rect 586000 275439 586006 275451
rect 586058 275439 586064 275491
rect 306352 275365 306358 275417
rect 306410 275405 306416 275417
rect 387376 275405 387382 275417
rect 306410 275377 387382 275405
rect 306410 275365 306416 275377
rect 387376 275365 387382 275377
rect 387434 275365 387440 275417
rect 584848 275405 584854 275417
rect 387490 275377 584854 275405
rect 306160 275291 306166 275343
rect 306218 275331 306224 275343
rect 386224 275331 386230 275343
rect 306218 275303 386230 275331
rect 306218 275291 306224 275303
rect 386224 275291 386230 275303
rect 386282 275291 386288 275343
rect 386320 275291 386326 275343
rect 386378 275331 386384 275343
rect 387490 275331 387518 275377
rect 584848 275365 584854 275377
rect 584906 275365 584912 275417
rect 386378 275303 387518 275331
rect 386378 275291 386384 275303
rect 390352 275291 390358 275343
rect 390410 275331 390416 275343
rect 390410 275303 407870 275331
rect 390410 275291 390416 275303
rect 308080 275217 308086 275269
rect 308138 275257 308144 275269
rect 390928 275257 390934 275269
rect 308138 275229 390934 275257
rect 308138 275217 308144 275229
rect 390928 275217 390934 275229
rect 390986 275217 390992 275269
rect 395152 275217 395158 275269
rect 395210 275257 395216 275269
rect 407842 275257 407870 275303
rect 407920 275291 407926 275343
rect 407978 275331 407984 275343
rect 591952 275331 591958 275343
rect 407978 275303 591958 275331
rect 407978 275291 407984 275303
rect 591952 275291 591958 275303
rect 592010 275291 592016 275343
rect 595408 275257 595414 275269
rect 395210 275229 407774 275257
rect 407842 275229 595414 275257
rect 395210 275217 395216 275229
rect 310384 275143 310390 275195
rect 310442 275183 310448 275195
rect 396880 275183 396886 275195
rect 310442 275155 396886 275183
rect 310442 275143 310448 275155
rect 396880 275143 396886 275155
rect 396938 275143 396944 275195
rect 404944 275143 404950 275195
rect 405002 275183 405008 275195
rect 407746 275183 407774 275229
rect 595408 275217 595414 275229
rect 595466 275217 595472 275269
rect 607312 275183 607318 275195
rect 405002 275155 407678 275183
rect 407746 275155 607318 275183
rect 405002 275143 405008 275155
rect 314704 275069 314710 275121
rect 314762 275109 314768 275121
rect 407440 275109 407446 275121
rect 314762 275081 407446 275109
rect 314762 275069 314768 275081
rect 407440 275069 407446 275081
rect 407498 275069 407504 275121
rect 313552 274995 313558 275047
rect 313610 275035 313616 275047
rect 405136 275035 405142 275047
rect 313610 275007 405142 275035
rect 313610 274995 313616 275007
rect 405136 274995 405142 275007
rect 405194 274995 405200 275047
rect 407650 275035 407678 275155
rect 607312 275143 607318 275155
rect 607370 275143 607376 275195
rect 407728 275069 407734 275121
rect 407786 275109 407792 275121
rect 634384 275109 634390 275121
rect 407786 275081 634390 275109
rect 407786 275069 407792 275081
rect 634384 275069 634390 275081
rect 634442 275069 634448 275121
rect 630928 275035 630934 275047
rect 407650 275007 630934 275035
rect 630928 274995 630934 275007
rect 630986 274995 630992 275047
rect 347632 274921 347638 274973
rect 347690 274961 347696 274973
rect 489040 274961 489046 274973
rect 347690 274933 489046 274961
rect 347690 274921 347696 274933
rect 489040 274921 489046 274933
rect 489098 274921 489104 274973
rect 344560 274847 344566 274899
rect 344618 274887 344624 274899
rect 481936 274887 481942 274899
rect 344618 274859 481942 274887
rect 344618 274847 344624 274859
rect 481936 274847 481942 274859
rect 481994 274847 482000 274899
rect 341680 274773 341686 274825
rect 341738 274813 341744 274825
rect 474928 274813 474934 274825
rect 341738 274785 474934 274813
rect 341738 274773 341744 274785
rect 474928 274773 474934 274785
rect 474986 274773 474992 274825
rect 339088 274699 339094 274751
rect 339146 274739 339152 274751
rect 467824 274739 467830 274751
rect 339146 274711 467830 274739
rect 339146 274699 339152 274711
rect 467824 274699 467830 274711
rect 467882 274699 467888 274751
rect 336016 274625 336022 274677
rect 336074 274665 336080 274677
rect 460624 274665 460630 274677
rect 336074 274637 460630 274665
rect 336074 274625 336080 274637
rect 460624 274625 460630 274637
rect 460682 274625 460688 274677
rect 333136 274551 333142 274603
rect 333194 274591 333200 274603
rect 453520 274591 453526 274603
rect 333194 274563 453526 274591
rect 333194 274551 333200 274563
rect 453520 274551 453526 274563
rect 453578 274551 453584 274603
rect 330448 274477 330454 274529
rect 330506 274517 330512 274529
rect 446512 274517 446518 274529
rect 330506 274489 446518 274517
rect 330506 274477 330512 274489
rect 446512 274477 446518 274489
rect 446570 274477 446576 274529
rect 327568 274403 327574 274455
rect 327626 274443 327632 274455
rect 439408 274443 439414 274455
rect 327626 274415 439414 274443
rect 327626 274403 327632 274415
rect 439408 274403 439414 274415
rect 439466 274403 439472 274455
rect 325936 274329 325942 274381
rect 325994 274369 326000 274381
rect 435856 274369 435862 274381
rect 325994 274341 435862 274369
rect 325994 274329 326000 274341
rect 435856 274329 435862 274341
rect 435914 274329 435920 274381
rect 42160 274255 42166 274307
rect 42218 274295 42224 274307
rect 43120 274295 43126 274307
rect 42218 274267 43126 274295
rect 42218 274255 42224 274267
rect 43120 274255 43126 274267
rect 43178 274255 43184 274307
rect 321616 274255 321622 274307
rect 321674 274295 321680 274307
rect 425200 274295 425206 274307
rect 321674 274267 425206 274295
rect 321674 274255 321680 274267
rect 425200 274255 425206 274267
rect 425258 274255 425264 274307
rect 320176 274181 320182 274233
rect 320234 274221 320240 274233
rect 421648 274221 421654 274233
rect 320234 274193 421654 274221
rect 320234 274181 320240 274193
rect 421648 274181 421654 274193
rect 421706 274181 421712 274233
rect 317296 274107 317302 274159
rect 317354 274147 317360 274159
rect 414544 274147 414550 274159
rect 317354 274119 414550 274147
rect 317354 274107 317360 274119
rect 414544 274107 414550 274119
rect 414602 274107 414608 274159
rect 315952 274033 315958 274085
rect 316010 274073 316016 274085
rect 411088 274073 411094 274085
rect 316010 274045 411094 274073
rect 316010 274033 316016 274045
rect 411088 274033 411094 274045
rect 411146 274033 411152 274085
rect 311632 273959 311638 274011
rect 311690 273999 311696 274011
rect 400336 273999 400342 274011
rect 311690 273971 400342 273999
rect 311690 273959 311696 273971
rect 400336 273959 400342 273971
rect 400394 273959 400400 274011
rect 307312 273885 307318 273937
rect 307370 273925 307376 273937
rect 389680 273925 389686 273937
rect 307370 273897 389686 273925
rect 307370 273885 307376 273897
rect 389680 273885 389686 273897
rect 389738 273885 389744 273937
rect 378256 273811 378262 273863
rect 378314 273851 378320 273863
rect 399088 273851 399094 273863
rect 378314 273823 399094 273851
rect 378314 273811 378320 273823
rect 399088 273811 399094 273823
rect 399146 273811 399152 273863
rect 388912 273737 388918 273789
rect 388970 273777 388976 273789
rect 407920 273777 407926 273789
rect 388970 273749 407926 273777
rect 388970 273737 388976 273749
rect 407920 273737 407926 273749
rect 407978 273737 407984 273789
rect 406096 273663 406102 273715
rect 406154 273703 406160 273715
rect 407728 273703 407734 273715
rect 406154 273675 407734 273703
rect 406154 273663 406160 273675
rect 407728 273663 407734 273675
rect 407786 273663 407792 273715
rect 409648 273663 409654 273715
rect 409706 273703 409712 273715
rect 480880 273703 480886 273715
rect 409706 273675 480886 273703
rect 409706 273663 409712 273675
rect 480880 273663 480886 273675
rect 480938 273663 480944 273715
rect 403696 273589 403702 273641
rect 403754 273629 403760 273641
rect 506800 273629 506806 273641
rect 403754 273601 506806 273629
rect 403754 273589 403760 273601
rect 506800 273589 506806 273601
rect 506858 273589 506864 273641
rect 84784 273515 84790 273567
rect 84842 273555 84848 273567
rect 142384 273555 142390 273567
rect 84842 273527 142390 273555
rect 84842 273515 84848 273527
rect 142384 273515 142390 273527
rect 142442 273515 142448 273567
rect 149776 273515 149782 273567
rect 149834 273555 149840 273567
rect 207664 273555 207670 273567
rect 149834 273527 207670 273555
rect 149834 273515 149840 273527
rect 207664 273515 207670 273527
rect 207722 273515 207728 273567
rect 277744 273515 277750 273567
rect 277802 273555 277808 273567
rect 316432 273555 316438 273567
rect 277802 273527 316438 273555
rect 277802 273515 277808 273527
rect 316432 273515 316438 273527
rect 316490 273515 316496 273567
rect 342160 273515 342166 273567
rect 342218 273555 342224 273567
rect 476080 273555 476086 273567
rect 342218 273527 476086 273555
rect 342218 273515 342224 273527
rect 476080 273515 476086 273527
rect 476138 273515 476144 273567
rect 480880 273515 480886 273567
rect 480938 273555 480944 273567
rect 642736 273555 642742 273567
rect 480938 273527 642742 273555
rect 480938 273515 480944 273527
rect 642736 273515 642742 273527
rect 642794 273515 642800 273567
rect 80080 273441 80086 273493
rect 80138 273481 80144 273493
rect 142480 273481 142486 273493
rect 80138 273453 142486 273481
rect 80138 273441 80144 273453
rect 142480 273441 142486 273453
rect 142538 273441 142544 273493
rect 146224 273441 146230 273493
rect 146282 273481 146288 273493
rect 210160 273481 210166 273493
rect 146282 273453 210166 273481
rect 146282 273441 146288 273453
rect 210160 273441 210166 273453
rect 210218 273441 210224 273493
rect 275344 273441 275350 273493
rect 275402 273481 275408 273493
rect 310480 273481 310486 273493
rect 275402 273453 310486 273481
rect 275402 273441 275408 273453
rect 310480 273441 310486 273453
rect 310538 273441 310544 273493
rect 312784 273441 312790 273493
rect 312842 273481 312848 273493
rect 402736 273481 402742 273493
rect 312842 273453 402742 273481
rect 312842 273441 312848 273453
rect 402736 273441 402742 273453
rect 402794 273441 402800 273493
rect 402832 273441 402838 273493
rect 402890 273481 402896 273493
rect 545872 273481 545878 273493
rect 402890 273453 545878 273481
rect 402890 273441 402896 273453
rect 545872 273441 545878 273453
rect 545930 273441 545936 273493
rect 546640 273441 546646 273493
rect 546698 273481 546704 273493
rect 639184 273481 639190 273493
rect 546698 273453 639190 273481
rect 546698 273441 546704 273453
rect 639184 273441 639190 273453
rect 639242 273441 639248 273493
rect 139120 273367 139126 273419
rect 139178 273407 139184 273419
rect 207280 273407 207286 273419
rect 139178 273379 207286 273407
rect 139178 273367 139184 273379
rect 207280 273367 207286 273379
rect 207338 273367 207344 273419
rect 276304 273367 276310 273419
rect 276362 273407 276368 273419
rect 312880 273407 312886 273419
rect 276362 273379 312886 273407
rect 276362 273367 276368 273379
rect 312880 273367 312886 273379
rect 312938 273367 312944 273419
rect 313936 273367 313942 273419
rect 313994 273407 314000 273419
rect 329488 273407 329494 273419
rect 313994 273379 329494 273407
rect 313994 273367 314000 273379
rect 329488 273367 329494 273379
rect 329546 273367 329552 273419
rect 350992 273367 350998 273419
rect 351050 273407 351056 273419
rect 497392 273407 497398 273419
rect 351050 273379 497398 273407
rect 351050 273367 351056 273379
rect 497392 273367 497398 273379
rect 497450 273367 497456 273419
rect 506800 273367 506806 273419
rect 506858 273407 506864 273419
rect 628528 273407 628534 273419
rect 506858 273379 628534 273407
rect 506858 273367 506864 273379
rect 628528 273367 628534 273379
rect 628586 273367 628592 273419
rect 119056 273293 119062 273345
rect 119114 273333 119120 273345
rect 120880 273333 120886 273345
rect 119114 273305 120886 273333
rect 119114 273293 119120 273305
rect 120880 273293 120886 273305
rect 120938 273293 120944 273345
rect 132016 273293 132022 273345
rect 132074 273333 132080 273345
rect 206992 273333 206998 273345
rect 132074 273305 206998 273333
rect 132074 273293 132080 273305
rect 206992 273293 206998 273305
rect 207050 273293 207056 273345
rect 278224 273293 278230 273345
rect 278282 273333 278288 273345
rect 317680 273333 317686 273345
rect 278282 273305 317686 273333
rect 278282 273293 278288 273305
rect 317680 273293 317686 273305
rect 317738 273293 317744 273345
rect 352624 273293 352630 273345
rect 352682 273333 352688 273345
rect 502000 273333 502006 273345
rect 352682 273305 502006 273333
rect 352682 273293 352688 273305
rect 502000 273293 502006 273305
rect 502058 273293 502064 273345
rect 612976 273293 612982 273345
rect 613034 273333 613040 273345
rect 632080 273333 632086 273345
rect 613034 273305 632086 273333
rect 613034 273293 613040 273305
rect 632080 273293 632086 273305
rect 632138 273293 632144 273345
rect 127312 273219 127318 273271
rect 127370 273259 127376 273271
rect 209968 273259 209974 273271
rect 127370 273231 209974 273259
rect 127370 273219 127376 273231
rect 209968 273219 209974 273231
rect 210026 273219 210032 273271
rect 219568 273219 219574 273271
rect 219626 273259 219632 273271
rect 238672 273259 238678 273271
rect 219626 273231 238678 273259
rect 219626 273219 219632 273231
rect 238672 273219 238678 273231
rect 238730 273219 238736 273271
rect 281296 273219 281302 273271
rect 281354 273259 281360 273271
rect 324784 273259 324790 273271
rect 281354 273231 324790 273259
rect 281354 273219 281360 273231
rect 324784 273219 324790 273231
rect 324842 273219 324848 273271
rect 353680 273219 353686 273271
rect 353738 273259 353744 273271
rect 504400 273259 504406 273271
rect 353738 273231 504406 273259
rect 353738 273219 353744 273231
rect 504400 273219 504406 273231
rect 504458 273219 504464 273271
rect 123760 273145 123766 273197
rect 123818 273185 123824 273197
rect 209008 273185 209014 273197
rect 123818 273157 209014 273185
rect 123818 273145 123824 273157
rect 209008 273145 209014 273157
rect 209066 273145 209072 273197
rect 279664 273145 279670 273197
rect 279722 273185 279728 273197
rect 321136 273185 321142 273197
rect 279722 273157 321142 273185
rect 279722 273145 279728 273157
rect 321136 273145 321142 273157
rect 321194 273145 321200 273197
rect 355792 273145 355798 273197
rect 355850 273185 355856 273197
rect 509104 273185 509110 273197
rect 355850 273157 509110 273185
rect 355850 273145 355856 273157
rect 509104 273145 509110 273157
rect 509162 273145 509168 273197
rect 509200 273145 509206 273197
rect 509258 273185 509264 273197
rect 635632 273185 635638 273197
rect 509258 273157 635638 273185
rect 509258 273145 509264 273157
rect 635632 273145 635638 273157
rect 635690 273145 635696 273197
rect 116656 273071 116662 273123
rect 116714 273111 116720 273123
rect 207088 273111 207094 273123
rect 116714 273083 207094 273111
rect 116714 273071 116720 273083
rect 207088 273071 207094 273083
rect 207146 273071 207152 273123
rect 217168 273071 217174 273123
rect 217226 273111 217232 273123
rect 237616 273111 237622 273123
rect 217226 273083 237622 273111
rect 217226 273071 217232 273083
rect 237616 273071 237622 273083
rect 237674 273071 237680 273123
rect 280624 273071 280630 273123
rect 280682 273111 280688 273123
rect 323536 273111 323542 273123
rect 280682 273083 323542 273111
rect 280682 273071 280688 273083
rect 323536 273071 323542 273083
rect 323594 273071 323600 273123
rect 356752 273071 356758 273123
rect 356810 273111 356816 273123
rect 511504 273111 511510 273123
rect 356810 273083 511510 273111
rect 356810 273071 356816 273083
rect 511504 273071 511510 273083
rect 511562 273071 511568 273123
rect 113200 272997 113206 273049
rect 113258 273037 113264 273049
rect 205936 273037 205942 273049
rect 113258 273009 205942 273037
rect 113258 272997 113264 273009
rect 205936 272997 205942 273009
rect 205994 272997 206000 273049
rect 218320 272997 218326 273049
rect 218378 273037 218384 273049
rect 238096 273037 238102 273049
rect 218378 273009 238102 273037
rect 218378 272997 218384 273009
rect 238096 272997 238102 273009
rect 238154 272997 238160 273049
rect 279280 272997 279286 273049
rect 279338 273037 279344 273049
rect 319984 273037 319990 273049
rect 279338 273009 319990 273037
rect 279338 272997 279344 273009
rect 319984 272997 319990 273009
rect 320042 272997 320048 273049
rect 359344 272997 359350 273049
rect 359402 273037 359408 273049
rect 359402 273009 375998 273037
rect 359402 272997 359408 273009
rect 120208 272923 120214 272975
rect 120266 272963 120272 272975
rect 207952 272963 207958 272975
rect 120266 272935 207958 272963
rect 120266 272923 120272 272935
rect 207952 272923 207958 272935
rect 208010 272923 208016 272975
rect 220720 272923 220726 272975
rect 220778 272963 220784 272975
rect 239152 272963 239158 272975
rect 220778 272935 239158 272963
rect 220778 272923 220784 272935
rect 239152 272923 239158 272935
rect 239210 272923 239216 272975
rect 288496 272923 288502 272975
rect 288554 272963 288560 272975
rect 342448 272963 342454 272975
rect 288554 272935 342454 272963
rect 288554 272923 288560 272935
rect 342448 272923 342454 272935
rect 342506 272923 342512 272975
rect 361264 272923 361270 272975
rect 361322 272963 361328 272975
rect 375970 272963 375998 273009
rect 376048 272997 376054 273049
rect 376106 273037 376112 273049
rect 516208 273037 516214 273049
rect 376106 273009 516214 273037
rect 376106 272997 376112 273009
rect 516208 272997 516214 273009
rect 516266 272997 516272 273049
rect 518608 272963 518614 272975
rect 361322 272935 375902 272963
rect 375970 272935 518614 272963
rect 361322 272923 361328 272935
rect 109552 272849 109558 272901
rect 109610 272889 109616 272901
rect 205264 272889 205270 272901
rect 109610 272861 205270 272889
rect 109610 272849 109616 272861
rect 205264 272849 205270 272861
rect 205322 272849 205328 272901
rect 214864 272849 214870 272901
rect 214922 272889 214928 272901
rect 236464 272889 236470 272901
rect 214922 272861 236470 272889
rect 214922 272849 214928 272861
rect 236464 272849 236470 272861
rect 236522 272849 236528 272901
rect 284944 272849 284950 272901
rect 285002 272889 285008 272901
rect 334096 272889 334102 272901
rect 285002 272861 334102 272889
rect 285002 272849 285008 272861
rect 334096 272849 334102 272861
rect 334154 272849 334160 272901
rect 362224 272849 362230 272901
rect 362282 272889 362288 272901
rect 375874 272889 375902 272935
rect 518608 272923 518614 272935
rect 518666 272923 518672 272975
rect 523408 272889 523414 272901
rect 362282 272861 375806 272889
rect 375874 272861 523414 272889
rect 362282 272849 362288 272861
rect 107152 272775 107158 272827
rect 107210 272815 107216 272827
rect 204688 272815 204694 272827
rect 107210 272787 204694 272815
rect 107210 272775 107216 272787
rect 204688 272775 204694 272787
rect 204746 272775 204752 272827
rect 213616 272775 213622 272827
rect 213674 272815 213680 272827
rect 236272 272815 236278 272827
rect 213674 272787 236278 272815
rect 213674 272775 213680 272787
rect 236272 272775 236278 272787
rect 236330 272775 236336 272827
rect 287920 272775 287926 272827
rect 287978 272815 287984 272827
rect 341296 272815 341302 272827
rect 287978 272787 341302 272815
rect 287978 272775 287984 272787
rect 341296 272775 341302 272787
rect 341354 272775 341360 272827
rect 364144 272775 364150 272827
rect 364202 272815 364208 272827
rect 375778 272815 375806 272861
rect 523408 272849 523414 272861
rect 523466 272849 523472 272901
rect 525712 272815 525718 272827
rect 364202 272787 375710 272815
rect 375778 272787 525718 272815
rect 364202 272775 364208 272787
rect 102544 272701 102550 272753
rect 102602 272741 102608 272753
rect 203344 272741 203350 272753
rect 102602 272713 203350 272741
rect 102602 272701 102608 272713
rect 203344 272701 203350 272713
rect 203402 272701 203408 272753
rect 215920 272701 215926 272753
rect 215978 272741 215984 272753
rect 236944 272741 236950 272753
rect 215978 272713 236950 272741
rect 215978 272701 215984 272713
rect 236944 272701 236950 272713
rect 237002 272701 237008 272753
rect 271024 272701 271030 272753
rect 271082 272741 271088 272753
rect 299920 272741 299926 272753
rect 271082 272713 299926 272741
rect 271082 272701 271088 272713
rect 299920 272701 299926 272713
rect 299978 272701 299984 272753
rect 301840 272701 301846 272753
rect 301898 272741 301904 272753
rect 358960 272741 358966 272753
rect 301898 272713 358966 272741
rect 301898 272701 301904 272713
rect 358960 272701 358966 272713
rect 359018 272701 359024 272753
rect 365296 272701 365302 272753
rect 365354 272741 365360 272753
rect 375568 272741 375574 272753
rect 365354 272713 375574 272741
rect 365354 272701 365360 272713
rect 375568 272701 375574 272713
rect 375626 272701 375632 272753
rect 375682 272741 375710 272787
rect 525712 272775 525718 272787
rect 525770 272775 525776 272827
rect 530512 272741 530518 272753
rect 375682 272713 530518 272741
rect 530512 272701 530518 272713
rect 530570 272701 530576 272753
rect 95440 272627 95446 272679
rect 95498 272667 95504 272679
rect 201136 272667 201142 272679
rect 95498 272639 201142 272667
rect 95498 272627 95504 272639
rect 201136 272627 201142 272639
rect 201194 272627 201200 272679
rect 233680 272627 233686 272679
rect 233738 272667 233744 272679
rect 244048 272667 244054 272679
rect 233738 272639 244054 272667
rect 233738 272627 233744 272639
rect 244048 272627 244054 272639
rect 244106 272627 244112 272679
rect 292720 272627 292726 272679
rect 292778 272667 292784 272679
rect 353104 272667 353110 272679
rect 292778 272639 353110 272667
rect 292778 272627 292784 272639
rect 353104 272627 353110 272639
rect 353162 272627 353168 272679
rect 367024 272627 367030 272679
rect 367082 272667 367088 272679
rect 537520 272667 537526 272679
rect 367082 272639 537526 272667
rect 367082 272627 367088 272639
rect 537520 272627 537526 272639
rect 537578 272627 537584 272679
rect 100144 272553 100150 272605
rect 100202 272593 100208 272605
rect 202864 272593 202870 272605
rect 100202 272565 202870 272593
rect 100202 272553 100208 272565
rect 202864 272553 202870 272565
rect 202922 272553 202928 272605
rect 212464 272553 212470 272605
rect 212522 272593 212528 272605
rect 235696 272593 235702 272605
rect 212522 272565 235702 272593
rect 212522 272553 212528 272565
rect 235696 272553 235702 272565
rect 235754 272553 235760 272605
rect 295408 272553 295414 272605
rect 295466 272593 295472 272605
rect 360208 272593 360214 272605
rect 295466 272565 360214 272593
rect 295466 272553 295472 272565
rect 360208 272553 360214 272565
rect 360266 272553 360272 272605
rect 367888 272553 367894 272605
rect 367946 272593 367952 272605
rect 367946 272565 375518 272593
rect 367946 272553 367952 272565
rect 93040 272479 93046 272531
rect 93098 272519 93104 272531
rect 200944 272519 200950 272531
rect 93098 272491 200950 272519
rect 93098 272479 93104 272491
rect 200944 272479 200950 272491
rect 201002 272479 201008 272531
rect 208816 272479 208822 272531
rect 208874 272519 208880 272531
rect 234352 272519 234358 272531
rect 208874 272491 234358 272519
rect 208874 272479 208880 272491
rect 234352 272479 234358 272491
rect 234410 272479 234416 272531
rect 270256 272479 270262 272531
rect 270314 272519 270320 272531
rect 297520 272519 297526 272531
rect 270314 272491 297526 272519
rect 270314 272479 270320 272491
rect 297520 272479 297526 272491
rect 297578 272479 297584 272531
rect 298288 272479 298294 272531
rect 298346 272519 298352 272531
rect 367216 272519 367222 272531
rect 298346 272491 367222 272519
rect 298346 272479 298352 272491
rect 367216 272479 367222 272491
rect 367274 272479 367280 272531
rect 374128 272479 374134 272531
rect 374186 272519 374192 272531
rect 375490 272519 375518 272565
rect 375568 272553 375574 272605
rect 375626 272593 375632 272605
rect 532816 272593 532822 272605
rect 375626 272565 532822 272593
rect 375626 272553 375632 272565
rect 532816 272553 532822 272565
rect 532874 272553 532880 272605
rect 539824 272519 539830 272531
rect 374186 272491 374462 272519
rect 375490 272491 539830 272519
rect 374186 272479 374192 272491
rect 90640 272405 90646 272457
rect 90698 272445 90704 272457
rect 199696 272445 199702 272457
rect 90698 272417 199702 272445
rect 90698 272405 90704 272417
rect 199696 272405 199702 272417
rect 199754 272405 199760 272457
rect 232528 272405 232534 272457
rect 232586 272445 232592 272457
rect 243664 272445 243670 272457
rect 232586 272417 243670 272445
rect 232586 272405 232592 272417
rect 243664 272405 243670 272417
rect 243722 272405 243728 272457
rect 271792 272405 271798 272457
rect 271850 272445 271856 272457
rect 301072 272445 301078 272457
rect 271850 272417 301078 272445
rect 271850 272405 271856 272417
rect 301072 272405 301078 272417
rect 301130 272405 301136 272457
rect 301360 272405 301366 272457
rect 301418 272445 301424 272457
rect 374320 272445 374326 272457
rect 301418 272417 374326 272445
rect 301418 272405 301424 272417
rect 374320 272405 374326 272417
rect 374378 272405 374384 272457
rect 374434 272445 374462 272491
rect 539824 272479 539830 272491
rect 539882 272479 539888 272531
rect 555184 272445 555190 272457
rect 374434 272417 555190 272445
rect 555184 272405 555190 272417
rect 555242 272405 555248 272457
rect 87088 272331 87094 272383
rect 87146 272371 87152 272383
rect 199024 272371 199030 272383
rect 87146 272343 199030 272371
rect 87146 272331 87152 272343
rect 199024 272331 199030 272343
rect 199082 272331 199088 272383
rect 207760 272331 207766 272383
rect 207818 272371 207824 272383
rect 233872 272371 233878 272383
rect 207818 272343 233878 272371
rect 207818 272331 207824 272343
rect 233872 272331 233878 272343
rect 233930 272331 233936 272383
rect 236080 272331 236086 272383
rect 236138 272371 236144 272383
rect 245296 272371 245302 272383
rect 236138 272343 245302 272371
rect 236138 272331 236144 272343
rect 245296 272331 245302 272343
rect 245354 272331 245360 272383
rect 272752 272331 272758 272383
rect 272810 272371 272816 272383
rect 303376 272371 303382 272383
rect 272810 272343 303382 272371
rect 272810 272331 272816 272343
rect 303376 272331 303382 272343
rect 303434 272331 303440 272383
rect 303952 272331 303958 272383
rect 304010 272371 304016 272383
rect 381520 272371 381526 272383
rect 304010 272343 381526 272371
rect 304010 272331 304016 272343
rect 381520 272331 381526 272343
rect 381578 272331 381584 272383
rect 382960 272331 382966 272383
rect 383018 272371 383024 272383
rect 576592 272371 576598 272383
rect 383018 272343 576598 272371
rect 383018 272331 383024 272343
rect 576592 272331 576598 272343
rect 576650 272331 576656 272383
rect 81232 272257 81238 272309
rect 81290 272297 81296 272309
rect 196816 272297 196822 272309
rect 81290 272269 196822 272297
rect 81290 272257 81296 272269
rect 196816 272257 196822 272269
rect 196874 272257 196880 272309
rect 210064 272257 210070 272309
rect 210122 272297 210128 272309
rect 234544 272297 234550 272309
rect 210122 272269 234550 272297
rect 210122 272257 210128 272269
rect 234544 272257 234550 272269
rect 234602 272257 234608 272309
rect 234928 272257 234934 272309
rect 234986 272297 234992 272309
rect 244816 272297 244822 272309
rect 234986 272269 244822 272297
rect 234986 272257 234992 272269
rect 244816 272257 244822 272269
rect 244874 272257 244880 272309
rect 273424 272257 273430 272309
rect 273482 272297 273488 272309
rect 305776 272297 305782 272309
rect 273482 272269 305782 272297
rect 273482 272257 273488 272269
rect 305776 272257 305782 272269
rect 305834 272257 305840 272309
rect 306832 272257 306838 272309
rect 306890 272297 306896 272309
rect 388624 272297 388630 272309
rect 306890 272269 388630 272297
rect 306890 272257 306896 272269
rect 388624 272257 388630 272269
rect 388682 272257 388688 272309
rect 388720 272257 388726 272309
rect 388778 272297 388784 272309
rect 590704 272297 590710 272309
rect 388778 272269 590710 272297
rect 388778 272257 388784 272269
rect 590704 272257 590710 272269
rect 590762 272257 590768 272309
rect 82384 272183 82390 272235
rect 82442 272223 82448 272235
rect 197392 272223 197398 272235
rect 82442 272195 197398 272223
rect 82442 272183 82448 272195
rect 197392 272183 197398 272195
rect 197450 272183 197456 272235
rect 228976 272183 228982 272235
rect 229034 272223 229040 272235
rect 242416 272223 242422 272235
rect 229034 272195 242422 272223
rect 229034 272183 229040 272195
rect 242416 272183 242422 272195
rect 242474 272183 242480 272235
rect 275152 272183 275158 272235
rect 275210 272223 275216 272235
rect 309424 272223 309430 272235
rect 275210 272195 309430 272223
rect 275210 272183 275216 272195
rect 309424 272183 309430 272195
rect 309482 272183 309488 272235
rect 309904 272183 309910 272235
rect 309962 272223 309968 272235
rect 395728 272223 395734 272235
rect 309962 272195 395734 272223
rect 309962 272183 309968 272195
rect 395728 272183 395734 272195
rect 395786 272183 395792 272235
rect 397072 272183 397078 272235
rect 397130 272223 397136 272235
rect 612016 272223 612022 272235
rect 397130 272195 612022 272223
rect 397130 272183 397136 272195
rect 612016 272183 612022 272195
rect 612074 272183 612080 272235
rect 72976 272109 72982 272161
rect 73034 272149 73040 272161
rect 194416 272149 194422 272161
rect 73034 272121 194422 272149
rect 73034 272109 73040 272121
rect 194416 272109 194422 272121
rect 194474 272109 194480 272161
rect 194704 272109 194710 272161
rect 194762 272149 194768 272161
rect 224560 272149 224566 272161
rect 194762 272121 224566 272149
rect 194762 272109 194768 272121
rect 224560 272109 224566 272121
rect 224618 272109 224624 272161
rect 227824 272109 227830 272161
rect 227882 272149 227888 272161
rect 242128 272149 242134 272161
rect 227882 272121 242134 272149
rect 227882 272109 227888 272121
rect 242128 272109 242134 272121
rect 242186 272109 242192 272161
rect 277072 272109 277078 272161
rect 277130 272149 277136 272161
rect 314128 272149 314134 272161
rect 277130 272121 314134 272149
rect 277130 272109 277136 272121
rect 314128 272109 314134 272121
rect 314186 272109 314192 272161
rect 315472 272109 315478 272161
rect 315530 272149 315536 272161
rect 409840 272149 409846 272161
rect 315530 272121 409846 272149
rect 315530 272109 315536 272121
rect 409840 272109 409846 272121
rect 409898 272109 409904 272161
rect 410896 272109 410902 272161
rect 410954 272149 410960 272161
rect 646288 272149 646294 272161
rect 410954 272121 646294 272149
rect 410954 272109 410960 272121
rect 646288 272109 646294 272121
rect 646346 272109 646352 272161
rect 101296 272035 101302 272087
rect 101354 272075 101360 272087
rect 159760 272075 159766 272087
rect 101354 272047 159766 272075
rect 101354 272035 101360 272047
rect 159760 272035 159766 272047
rect 159818 272035 159824 272087
rect 163984 272035 163990 272087
rect 164042 272075 164048 272087
rect 207856 272075 207862 272087
rect 164042 272047 207862 272075
rect 164042 272035 164048 272047
rect 207856 272035 207862 272047
rect 207914 272035 207920 272087
rect 230224 272035 230230 272087
rect 230282 272075 230288 272087
rect 242896 272075 242902 272087
rect 230282 272047 242902 272075
rect 230282 272035 230288 272047
rect 242896 272035 242902 272047
rect 242954 272035 242960 272087
rect 273904 272035 273910 272087
rect 273962 272075 273968 272087
rect 307024 272075 307030 272087
rect 273962 272047 307030 272075
rect 273962 272035 273968 272047
rect 307024 272035 307030 272047
rect 307082 272035 307088 272087
rect 348112 272035 348118 272087
rect 348170 272075 348176 272087
rect 490288 272075 490294 272087
rect 348170 272047 490294 272075
rect 348170 272035 348176 272047
rect 490288 272035 490294 272047
rect 490346 272035 490352 272087
rect 97744 271961 97750 272013
rect 97802 272001 97808 272013
rect 151120 272001 151126 272013
rect 97802 271973 151126 272001
rect 97802 271961 97808 271973
rect 151120 271961 151126 271973
rect 151178 271961 151184 272013
rect 156880 271961 156886 272013
rect 156938 272001 156944 272013
rect 207760 272001 207766 272013
rect 156938 271973 207766 272001
rect 156938 271961 156944 271973
rect 207760 271961 207766 271973
rect 207818 271961 207824 272013
rect 231376 271961 231382 272013
rect 231434 272001 231440 272013
rect 243088 272001 243094 272013
rect 231434 271973 243094 272001
rect 231434 271961 231440 271973
rect 243088 271961 243094 271973
rect 243146 271961 243152 272013
rect 272944 271961 272950 272013
rect 273002 272001 273008 272013
rect 304624 272001 304630 272013
rect 273002 271973 304630 272001
rect 273002 271961 273008 271973
rect 304624 271961 304630 271973
rect 304682 271961 304688 272013
rect 350032 271961 350038 272013
rect 350090 272001 350096 272013
rect 494992 272001 494998 272013
rect 350090 271973 494998 272001
rect 350090 271961 350096 271973
rect 494992 271961 494998 271973
rect 495050 271961 495056 272013
rect 89488 271887 89494 271939
rect 89546 271927 89552 271939
rect 142576 271927 142582 271939
rect 89546 271899 142582 271927
rect 89546 271887 89552 271899
rect 142576 271887 142582 271899
rect 142634 271887 142640 271939
rect 168688 271887 168694 271939
rect 168746 271927 168752 271939
rect 169840 271927 169846 271939
rect 168746 271899 169846 271927
rect 168746 271887 168752 271899
rect 169840 271887 169846 271899
rect 169898 271887 169904 271939
rect 179344 271887 179350 271939
rect 179402 271927 179408 271939
rect 181360 271927 181366 271939
rect 179402 271899 181366 271927
rect 179402 271887 179408 271899
rect 181360 271887 181366 271899
rect 181418 271887 181424 271939
rect 182896 271887 182902 271939
rect 182954 271927 182960 271939
rect 184240 271927 184246 271939
rect 182954 271899 184246 271927
rect 182954 271887 182960 271899
rect 184240 271887 184246 271899
rect 184298 271887 184304 271939
rect 207472 271927 207478 271939
rect 187186 271899 207478 271927
rect 111952 271813 111958 271865
rect 112010 271853 112016 271865
rect 162640 271853 162646 271865
rect 112010 271825 162646 271853
rect 112010 271813 112016 271825
rect 162640 271813 162646 271825
rect 162698 271813 162704 271865
rect 170992 271813 170998 271865
rect 171050 271853 171056 271865
rect 187186 271853 187214 271899
rect 207472 271887 207478 271899
rect 207530 271887 207536 271939
rect 211216 271887 211222 271939
rect 211274 271927 211280 271939
rect 235024 271927 235030 271939
rect 211274 271899 235030 271927
rect 211274 271887 211280 271899
rect 235024 271887 235030 271899
rect 235082 271887 235088 271939
rect 270544 271887 270550 271939
rect 270602 271927 270608 271939
rect 298672 271927 298678 271939
rect 270602 271899 298678 271927
rect 270602 271887 270608 271899
rect 298672 271887 298678 271899
rect 298730 271887 298736 271939
rect 299440 271887 299446 271939
rect 299498 271927 299504 271939
rect 327088 271927 327094 271939
rect 299498 271899 327094 271927
rect 299498 271887 299504 271899
rect 327088 271887 327094 271899
rect 327146 271887 327152 271939
rect 346960 271887 346966 271939
rect 347018 271927 347024 271939
rect 487888 271927 487894 271939
rect 347018 271899 487894 271927
rect 347018 271887 347024 271899
rect 487888 271887 487894 271899
rect 487946 271887 487952 271939
rect 171050 271825 187214 271853
rect 171050 271813 171056 271825
rect 191152 271813 191158 271865
rect 191210 271853 191216 271865
rect 227152 271853 227158 271865
rect 191210 271825 227158 271853
rect 191210 271813 191216 271825
rect 227152 271813 227158 271825
rect 227210 271813 227216 271865
rect 272272 271813 272278 271865
rect 272330 271853 272336 271865
rect 302320 271853 302326 271865
rect 272330 271825 302326 271853
rect 272330 271813 272336 271825
rect 302320 271813 302326 271825
rect 302378 271813 302384 271865
rect 345232 271813 345238 271865
rect 345290 271853 345296 271865
rect 483184 271853 483190 271865
rect 345290 271825 483190 271853
rect 345290 271813 345296 271825
rect 483184 271813 483190 271825
rect 483242 271813 483248 271865
rect 94192 271739 94198 271791
rect 94250 271779 94256 271791
rect 142768 271779 142774 271791
rect 94250 271751 142774 271779
rect 94250 271739 94256 271751
rect 142768 271739 142774 271751
rect 142826 271739 142832 271791
rect 155632 271739 155638 271791
rect 155690 271779 155696 271791
rect 155690 271751 161294 271779
rect 155690 271739 155696 271751
rect 104848 271665 104854 271717
rect 104906 271705 104912 271717
rect 154000 271705 154006 271717
rect 104906 271677 154006 271705
rect 104906 271665 104912 271677
rect 154000 271665 154006 271677
rect 154058 271665 154064 271717
rect 108400 271591 108406 271643
rect 108458 271631 108464 271643
rect 156880 271631 156886 271643
rect 108458 271603 156886 271631
rect 108458 271591 108464 271603
rect 156880 271591 156886 271603
rect 156938 271591 156944 271643
rect 126160 271517 126166 271569
rect 126218 271557 126224 271569
rect 143056 271557 143062 271569
rect 126218 271529 143062 271557
rect 126218 271517 126224 271529
rect 143056 271517 143062 271529
rect 143114 271517 143120 271569
rect 161266 271557 161294 271751
rect 162736 271739 162742 271791
rect 162794 271779 162800 271791
rect 192976 271779 192982 271791
rect 162794 271751 192982 271779
rect 162794 271739 162800 271751
rect 192976 271739 192982 271751
rect 193034 271739 193040 271791
rect 195856 271739 195862 271791
rect 195914 271779 195920 271791
rect 221584 271779 221590 271791
rect 195914 271751 221590 271779
rect 195914 271739 195920 271751
rect 221584 271739 221590 271751
rect 221642 271739 221648 271791
rect 344080 271739 344086 271791
rect 344138 271779 344144 271791
rect 480784 271779 480790 271791
rect 344138 271751 480790 271779
rect 344138 271739 344144 271751
rect 480784 271739 480790 271751
rect 480842 271739 480848 271791
rect 178096 271665 178102 271717
rect 178154 271705 178160 271717
rect 207376 271705 207382 271717
rect 178154 271677 207382 271705
rect 178154 271665 178160 271677
rect 207376 271665 207382 271677
rect 207434 271665 207440 271717
rect 341488 271665 341494 271717
rect 341546 271705 341552 271717
rect 473680 271705 473686 271717
rect 341546 271677 473686 271705
rect 341546 271665 341552 271677
rect 473680 271665 473686 271677
rect 473738 271665 473744 271717
rect 161584 271591 161590 271643
rect 161642 271631 161648 271643
rect 164080 271631 164086 271643
rect 161642 271603 164086 271631
rect 161642 271591 161648 271603
rect 164080 271591 164086 271603
rect 164138 271591 164144 271643
rect 185392 271591 185398 271643
rect 185450 271631 185456 271643
rect 186352 271631 186358 271643
rect 185450 271603 186358 271631
rect 185450 271591 185456 271603
rect 186352 271591 186358 271603
rect 186410 271591 186416 271643
rect 193168 271631 193174 271643
rect 187186 271603 193174 271631
rect 187186 271557 187214 271603
rect 193168 271591 193174 271603
rect 193226 271591 193232 271643
rect 201808 271591 201814 271643
rect 201866 271631 201872 271643
rect 224272 271631 224278 271643
rect 201866 271603 224278 271631
rect 201866 271591 201872 271603
rect 224272 271591 224278 271603
rect 224330 271591 224336 271643
rect 338608 271591 338614 271643
rect 338666 271631 338672 271643
rect 466576 271631 466582 271643
rect 338666 271603 466582 271631
rect 338666 271591 338672 271603
rect 466576 271591 466582 271603
rect 466634 271591 466640 271643
rect 161266 271529 187214 271557
rect 192304 271517 192310 271569
rect 192362 271557 192368 271569
rect 221968 271557 221974 271569
rect 192362 271529 221974 271557
rect 192362 271517 192368 271529
rect 221968 271517 221974 271529
rect 222026 271517 222032 271569
rect 335440 271517 335446 271569
rect 335498 271557 335504 271569
rect 459568 271557 459574 271569
rect 335498 271529 459574 271557
rect 335498 271517 335504 271529
rect 459568 271517 459574 271529
rect 459626 271517 459632 271569
rect 129616 271443 129622 271495
rect 129674 271483 129680 271495
rect 142960 271483 142966 271495
rect 129674 271455 142966 271483
rect 129674 271443 129680 271455
rect 142960 271443 142966 271455
rect 143018 271443 143024 271495
rect 181744 271443 181750 271495
rect 181802 271483 181808 271495
rect 210448 271483 210454 271495
rect 181802 271455 210454 271483
rect 181802 271443 181808 271455
rect 210448 271443 210454 271455
rect 210506 271443 210512 271495
rect 332560 271443 332566 271495
rect 332618 271483 332624 271495
rect 452464 271483 452470 271495
rect 332618 271455 452470 271483
rect 332618 271443 332624 271455
rect 452464 271443 452470 271455
rect 452522 271443 452528 271495
rect 133264 271369 133270 271421
rect 133322 271409 133328 271421
rect 142864 271409 142870 271421
rect 133322 271381 142870 271409
rect 133322 271369 133328 271381
rect 142864 271369 142870 271381
rect 142922 271369 142928 271421
rect 169744 271369 169750 271421
rect 169802 271409 169808 271421
rect 198640 271409 198646 271421
rect 169802 271381 198646 271409
rect 169802 271369 169808 271381
rect 198640 271369 198646 271381
rect 198698 271369 198704 271421
rect 199504 271369 199510 271421
rect 199562 271409 199568 271421
rect 221488 271409 221494 271421
rect 199562 271381 221494 271409
rect 199562 271369 199568 271381
rect 221488 271369 221494 271381
rect 221546 271369 221552 271421
rect 329968 271369 329974 271421
rect 330026 271409 330032 271421
rect 445264 271409 445270 271421
rect 330026 271381 445270 271409
rect 330026 271369 330032 271381
rect 445264 271369 445270 271381
rect 445322 271369 445328 271421
rect 185200 271295 185206 271347
rect 185258 271335 185264 271347
rect 210352 271335 210358 271347
rect 185258 271307 210358 271335
rect 185258 271295 185264 271307
rect 210352 271295 210358 271307
rect 210410 271295 210416 271347
rect 237232 271295 237238 271347
rect 237290 271335 237296 271347
rect 245488 271335 245494 271347
rect 237290 271307 245494 271335
rect 237290 271295 237296 271307
rect 245488 271295 245494 271307
rect 245546 271295 245552 271347
rect 326896 271295 326902 271347
rect 326954 271335 326960 271347
rect 438160 271335 438166 271347
rect 326954 271307 438166 271335
rect 326954 271295 326960 271307
rect 438160 271295 438166 271307
rect 438218 271295 438224 271347
rect 136816 271221 136822 271273
rect 136874 271261 136880 271273
rect 143152 271261 143158 271273
rect 136874 271233 143158 271261
rect 136874 271221 136880 271233
rect 143152 271221 143158 271233
rect 143210 271221 143216 271273
rect 193456 271221 193462 271273
rect 193514 271261 193520 271273
rect 221680 271261 221686 271273
rect 193514 271233 221686 271261
rect 193514 271221 193520 271233
rect 221680 271221 221686 271233
rect 221738 271221 221744 271273
rect 238480 271221 238486 271273
rect 238538 271261 238544 271273
rect 246064 271261 246070 271273
rect 238538 271233 246070 271261
rect 238538 271221 238544 271233
rect 246064 271221 246070 271233
rect 246122 271221 246128 271273
rect 324016 271221 324022 271273
rect 324074 271261 324080 271273
rect 431152 271261 431158 271273
rect 324074 271233 431158 271261
rect 324074 271221 324080 271233
rect 431152 271221 431158 271233
rect 431210 271221 431216 271273
rect 75280 271147 75286 271199
rect 75338 271187 75344 271199
rect 77488 271187 77494 271199
rect 75338 271159 77494 271187
rect 75338 271147 75344 271159
rect 77488 271147 77494 271159
rect 77546 271147 77552 271199
rect 176944 271147 176950 271199
rect 177002 271187 177008 271199
rect 204016 271187 204022 271199
rect 177002 271159 204022 271187
rect 177002 271147 177008 271159
rect 204016 271147 204022 271159
rect 204074 271147 204080 271199
rect 205360 271147 205366 271199
rect 205418 271187 205424 271199
rect 232624 271187 232630 271199
rect 205418 271159 232630 271187
rect 205418 271147 205424 271159
rect 232624 271147 232630 271159
rect 232682 271147 232688 271199
rect 239536 271147 239542 271199
rect 239594 271187 239600 271199
rect 246448 271187 246454 271199
rect 239594 271159 246454 271187
rect 239594 271147 239600 271159
rect 246448 271147 246454 271159
rect 246506 271147 246512 271199
rect 321424 271147 321430 271199
rect 321482 271187 321488 271199
rect 424048 271187 424054 271199
rect 321482 271159 424054 271187
rect 321482 271147 321488 271159
rect 424048 271147 424054 271159
rect 424106 271147 424112 271199
rect 140272 271073 140278 271125
rect 140330 271113 140336 271125
rect 143248 271113 143254 271125
rect 140330 271085 143254 271113
rect 140330 271073 140336 271085
rect 143248 271073 143254 271085
rect 143306 271073 143312 271125
rect 175792 271073 175798 271125
rect 175850 271113 175856 271125
rect 178480 271113 178486 271125
rect 175850 271085 178486 271113
rect 175850 271073 175856 271085
rect 178480 271073 178486 271085
rect 178538 271073 178544 271125
rect 188752 271073 188758 271125
rect 188810 271113 188816 271125
rect 210256 271113 210262 271125
rect 188810 271085 210262 271113
rect 188810 271073 188816 271085
rect 210256 271073 210262 271085
rect 210314 271073 210320 271125
rect 240784 271073 240790 271125
rect 240842 271113 240848 271125
rect 247216 271113 247222 271125
rect 240842 271085 247222 271113
rect 240842 271073 240848 271085
rect 247216 271073 247222 271085
rect 247274 271073 247280 271125
rect 318352 271073 318358 271125
rect 318410 271113 318416 271125
rect 416944 271113 416950 271125
rect 318410 271085 416950 271113
rect 318410 271073 318416 271085
rect 416944 271073 416950 271085
rect 417002 271073 417008 271125
rect 187600 270999 187606 271051
rect 187658 271039 187664 271051
rect 205840 271039 205846 271051
rect 187658 271011 205846 271039
rect 187658 270999 187664 271011
rect 205840 270999 205846 271011
rect 205898 270999 205904 271051
rect 221872 270999 221878 271051
rect 221930 271039 221936 271051
rect 239344 271039 239350 271051
rect 221930 271011 239350 271039
rect 221930 270999 221936 271011
rect 239344 270999 239350 271011
rect 239402 270999 239408 271051
rect 241936 270999 241942 271051
rect 241994 271039 242000 271051
rect 247696 271039 247702 271051
rect 241994 271011 247702 271039
rect 241994 270999 242000 271011
rect 247696 270999 247702 271011
rect 247754 270999 247760 271051
rect 358576 270999 358582 271051
rect 358634 271039 358640 271051
rect 376048 271039 376054 271051
rect 358634 271011 376054 271039
rect 358634 270999 358640 271011
rect 376048 270999 376054 271011
rect 376106 270999 376112 271051
rect 198256 270925 198262 270977
rect 198314 270965 198320 270977
rect 198314 270937 216014 270965
rect 198314 270925 198320 270937
rect 68176 270703 68182 270755
rect 68234 270743 68240 270755
rect 69040 270743 69046 270755
rect 68234 270715 69046 270743
rect 68234 270703 68240 270715
rect 69040 270703 69046 270715
rect 69098 270703 69104 270755
rect 115504 270703 115510 270755
rect 115562 270743 115568 270755
rect 118000 270743 118006 270755
rect 115562 270715 118006 270743
rect 115562 270703 115568 270715
rect 118000 270703 118006 270715
rect 118058 270703 118064 270755
rect 122512 270703 122518 270755
rect 122570 270743 122576 270755
rect 123760 270743 123766 270755
rect 122570 270715 123766 270743
rect 122570 270703 122576 270715
rect 123760 270703 123766 270715
rect 123818 270703 123824 270755
rect 143920 270703 143926 270755
rect 143978 270743 143984 270755
rect 145360 270743 145366 270755
rect 143978 270715 145366 270743
rect 143978 270703 143984 270715
rect 145360 270703 145366 270715
rect 145418 270703 145424 270755
rect 147376 270703 147382 270755
rect 147434 270743 147440 270755
rect 149680 270743 149686 270755
rect 147434 270715 149686 270743
rect 147434 270703 147440 270715
rect 149680 270703 149686 270715
rect 149738 270703 149744 270755
rect 151024 270703 151030 270755
rect 151082 270743 151088 270755
rect 152560 270743 152566 270755
rect 151082 270715 152566 270743
rect 151082 270703 151088 270715
rect 152560 270703 152566 270715
rect 152618 270703 152624 270755
rect 154480 270703 154486 270755
rect 154538 270743 154544 270755
rect 155440 270743 155446 270755
rect 154538 270715 155446 270743
rect 154538 270703 154544 270715
rect 155440 270703 155446 270715
rect 155498 270703 155504 270755
rect 165136 270703 165142 270755
rect 165194 270743 165200 270755
rect 166960 270743 166966 270755
rect 165194 270715 166966 270743
rect 165194 270703 165200 270715
rect 166960 270703 166966 270715
rect 167018 270703 167024 270755
rect 215986 270743 216014 270937
rect 223120 270925 223126 270977
rect 223178 270965 223184 270977
rect 240016 270965 240022 270977
rect 223178 270937 240022 270965
rect 223178 270925 223184 270937
rect 240016 270925 240022 270937
rect 240074 270925 240080 270977
rect 243184 270925 243190 270977
rect 243242 270965 243248 270977
rect 247984 270965 247990 270977
rect 243242 270937 247990 270965
rect 243242 270925 243248 270937
rect 247984 270925 247990 270937
rect 248042 270925 248048 270977
rect 224176 270851 224182 270903
rect 224234 270891 224240 270903
rect 240496 270891 240502 270903
rect 224234 270863 240502 270891
rect 224234 270851 224240 270863
rect 240496 270851 240502 270863
rect 240554 270851 240560 270903
rect 244336 270851 244342 270903
rect 244394 270891 244400 270903
rect 248656 270891 248662 270903
rect 244394 270863 248662 270891
rect 244394 270851 244400 270863
rect 248656 270851 248662 270863
rect 248714 270851 248720 270903
rect 225424 270777 225430 270829
rect 225482 270817 225488 270829
rect 241072 270817 241078 270829
rect 225482 270789 241078 270817
rect 225482 270777 225488 270789
rect 241072 270777 241078 270789
rect 241130 270777 241136 270829
rect 245584 270777 245590 270829
rect 245642 270817 245648 270829
rect 249136 270817 249142 270829
rect 245642 270789 249142 270817
rect 245642 270777 245648 270789
rect 249136 270777 249142 270789
rect 249194 270777 249200 270829
rect 340528 270777 340534 270829
rect 340586 270817 340592 270829
rect 348400 270817 348406 270829
rect 340586 270789 348406 270817
rect 340586 270777 340592 270789
rect 348400 270777 348406 270789
rect 348458 270777 348464 270829
rect 215986 270715 224606 270743
rect 142672 270629 142678 270681
rect 142730 270669 142736 270681
rect 214288 270669 214294 270681
rect 142730 270641 214294 270669
rect 142730 270629 142736 270641
rect 214288 270629 214294 270641
rect 214346 270629 214352 270681
rect 224578 270669 224606 270715
rect 226576 270703 226582 270755
rect 226634 270743 226640 270755
rect 241264 270743 241270 270755
rect 226634 270715 241270 270743
rect 226634 270703 226640 270715
rect 241264 270703 241270 270715
rect 241322 270703 241328 270755
rect 246736 270703 246742 270755
rect 246794 270743 246800 270755
rect 249616 270743 249622 270755
rect 246794 270715 249622 270743
rect 246794 270703 246800 270715
rect 249616 270703 249622 270715
rect 249674 270703 249680 270755
rect 337744 270743 337750 270755
rect 336946 270715 337750 270743
rect 230032 270669 230038 270681
rect 224578 270641 230038 270669
rect 230032 270629 230038 270641
rect 230090 270629 230096 270681
rect 262000 270629 262006 270681
rect 262058 270669 262064 270681
rect 262058 270641 276494 270669
rect 262058 270629 262064 270641
rect 137872 270555 137878 270607
rect 137930 270595 137936 270607
rect 212656 270595 212662 270607
rect 137930 270567 212662 270595
rect 137930 270555 137936 270567
rect 212656 270555 212662 270567
rect 212714 270555 212720 270607
rect 262960 270555 262966 270607
rect 263018 270595 263024 270607
rect 263018 270567 270158 270595
rect 263018 270555 263024 270567
rect 134416 270481 134422 270533
rect 134474 270521 134480 270533
rect 211888 270521 211894 270533
rect 134474 270493 211894 270521
rect 134474 270481 134480 270493
rect 211888 270481 211894 270493
rect 211946 270481 211952 270533
rect 124912 270407 124918 270459
rect 124970 270447 124976 270459
rect 209488 270447 209494 270459
rect 124970 270419 209494 270447
rect 124970 270407 124976 270419
rect 209488 270407 209494 270419
rect 209546 270407 209552 270459
rect 262480 270407 262486 270459
rect 262538 270447 262544 270459
rect 262538 270419 270014 270447
rect 262538 270407 262544 270419
rect 121360 270333 121366 270385
rect 121418 270373 121424 270385
rect 208336 270373 208342 270385
rect 121418 270345 208342 270373
rect 121418 270333 121424 270345
rect 208336 270333 208342 270345
rect 208394 270333 208400 270385
rect 117904 270259 117910 270311
rect 117962 270299 117968 270311
rect 207568 270299 207574 270311
rect 117962 270271 207574 270299
rect 117962 270259 117968 270271
rect 207568 270259 207574 270271
rect 207626 270259 207632 270311
rect 207664 270259 207670 270311
rect 207722 270299 207728 270311
rect 216208 270299 216214 270311
rect 207722 270271 216214 270299
rect 207722 270259 207728 270271
rect 216208 270259 216214 270271
rect 216266 270259 216272 270311
rect 253936 270259 253942 270311
rect 253994 270299 254000 270311
rect 257296 270299 257302 270311
rect 253994 270271 257302 270299
rect 253994 270259 254000 270271
rect 257296 270259 257302 270271
rect 257354 270259 257360 270311
rect 264880 270259 264886 270311
rect 264938 270299 264944 270311
rect 269872 270299 269878 270311
rect 264938 270271 269878 270299
rect 264938 270259 264944 270271
rect 269872 270259 269878 270271
rect 269930 270259 269936 270311
rect 269986 270299 270014 270419
rect 270130 270373 270158 270567
rect 276466 270447 276494 270641
rect 283696 270629 283702 270681
rect 283754 270669 283760 270681
rect 330640 270669 330646 270681
rect 283754 270641 330646 270669
rect 283754 270629 283760 270641
rect 330640 270629 330646 270641
rect 330698 270629 330704 270681
rect 284176 270555 284182 270607
rect 284234 270595 284240 270607
rect 331792 270595 331798 270607
rect 284234 270567 331798 270595
rect 284234 270555 284240 270567
rect 331792 270555 331798 270567
rect 331850 270555 331856 270607
rect 285616 270481 285622 270533
rect 285674 270521 285680 270533
rect 335344 270521 335350 270533
rect 285674 270493 335350 270521
rect 285674 270481 285680 270493
rect 335344 270481 335350 270493
rect 335402 270481 335408 270533
rect 277456 270447 277462 270459
rect 276466 270419 277462 270447
rect 277456 270407 277462 270419
rect 277514 270407 277520 270459
rect 286288 270407 286294 270459
rect 286346 270447 286352 270459
rect 336946 270447 336974 270715
rect 337744 270703 337750 270715
rect 337802 270703 337808 270755
rect 348400 270629 348406 270681
rect 348458 270669 348464 270681
rect 491440 270669 491446 270681
rect 348458 270641 491446 270669
rect 348458 270629 348464 270641
rect 491440 270629 491446 270641
rect 491498 270629 491504 270681
rect 349456 270555 349462 270607
rect 349514 270595 349520 270607
rect 493744 270595 493750 270607
rect 349514 270567 493750 270595
rect 349514 270555 349520 270567
rect 493744 270555 493750 270567
rect 493802 270555 493808 270607
rect 352432 270481 352438 270533
rect 352490 270521 352496 270533
rect 500848 270521 500854 270533
rect 352490 270493 500854 270521
rect 352490 270481 352496 270493
rect 500848 270481 500854 270493
rect 500906 270481 500912 270533
rect 286346 270419 336974 270447
rect 286346 270407 286352 270419
rect 351280 270407 351286 270459
rect 351338 270447 351344 270459
rect 498544 270447 498550 270459
rect 351338 270419 498550 270447
rect 351338 270407 351344 270419
rect 498544 270407 498550 270419
rect 498602 270407 498608 270459
rect 279760 270373 279766 270385
rect 270130 270345 279766 270373
rect 279760 270333 279766 270345
rect 279818 270333 279824 270385
rect 286768 270333 286774 270385
rect 286826 270373 286832 270385
rect 338896 270373 338902 270385
rect 286826 270345 338902 270373
rect 286826 270333 286832 270345
rect 338896 270333 338902 270345
rect 338954 270333 338960 270385
rect 355024 270333 355030 270385
rect 355082 270373 355088 270385
rect 507952 270373 507958 270385
rect 355082 270345 507958 270373
rect 355082 270333 355088 270345
rect 507952 270333 507958 270345
rect 508010 270333 508016 270385
rect 278704 270299 278710 270311
rect 269986 270271 278710 270299
rect 278704 270259 278710 270271
rect 278762 270259 278768 270311
rect 290608 270259 290614 270311
rect 290666 270299 290672 270311
rect 340528 270299 340534 270311
rect 290666 270271 340534 270299
rect 290666 270259 290672 270271
rect 340528 270259 340534 270271
rect 340586 270259 340592 270311
rect 354064 270259 354070 270311
rect 354122 270299 354128 270311
rect 505648 270299 505654 270311
rect 354122 270271 505654 270299
rect 354122 270259 354128 270271
rect 505648 270259 505654 270271
rect 505706 270259 505712 270311
rect 114256 270185 114262 270237
rect 114314 270225 114320 270237
rect 206416 270225 206422 270237
rect 114314 270197 206422 270225
rect 114314 270185 114320 270197
rect 206416 270185 206422 270197
rect 206474 270185 206480 270237
rect 210160 270185 210166 270237
rect 210218 270225 210224 270237
rect 214960 270225 214966 270237
rect 210218 270197 214966 270225
rect 210218 270185 210224 270197
rect 214960 270185 214966 270197
rect 215018 270185 215024 270237
rect 255280 270185 255286 270237
rect 255338 270225 255344 270237
rect 260944 270225 260950 270237
rect 255338 270197 260950 270225
rect 255338 270185 255344 270197
rect 260944 270185 260950 270197
rect 261002 270185 261008 270237
rect 266032 270185 266038 270237
rect 266090 270225 266096 270237
rect 286864 270225 286870 270237
rect 266090 270197 286870 270225
rect 266090 270185 266096 270197
rect 286864 270185 286870 270197
rect 286922 270185 286928 270237
rect 289168 270185 289174 270237
rect 289226 270225 289232 270237
rect 344848 270225 344854 270237
rect 289226 270197 344854 270225
rect 289226 270185 289232 270197
rect 344848 270185 344854 270197
rect 344906 270185 344912 270237
rect 357904 270185 357910 270237
rect 357962 270225 357968 270237
rect 515056 270225 515062 270237
rect 357962 270197 515062 270225
rect 357962 270185 357968 270197
rect 515056 270185 515062 270197
rect 515114 270185 515120 270237
rect 110800 270111 110806 270163
rect 110858 270151 110864 270163
rect 205744 270151 205750 270163
rect 110858 270123 205750 270151
rect 110858 270111 110864 270123
rect 205744 270111 205750 270123
rect 205802 270111 205808 270163
rect 207376 270111 207382 270163
rect 207434 270151 207440 270163
rect 223600 270151 223606 270163
rect 207434 270123 223606 270151
rect 207434 270111 207440 270123
rect 223600 270111 223606 270123
rect 223658 270111 223664 270163
rect 264688 270111 264694 270163
rect 264746 270151 264752 270163
rect 264746 270123 269822 270151
rect 264746 270111 264752 270123
rect 103696 270037 103702 270089
rect 103754 270077 103760 270089
rect 203536 270077 203542 270089
rect 103754 270049 203542 270077
rect 103754 270037 103760 270049
rect 203536 270037 203542 270049
rect 203594 270037 203600 270089
rect 210448 270037 210454 270089
rect 210506 270077 210512 270089
rect 224752 270077 224758 270089
rect 210506 270049 224758 270077
rect 210506 270037 210512 270049
rect 224752 270037 224758 270049
rect 224810 270037 224816 270089
rect 265360 270037 265366 270089
rect 265418 270077 265424 270089
rect 269794 270077 269822 270123
rect 269872 270111 269878 270163
rect 269930 270151 269936 270163
rect 284560 270151 284566 270163
rect 269930 270123 284566 270151
rect 269930 270111 269936 270123
rect 284560 270111 284566 270123
rect 284618 270111 284624 270163
rect 289936 270111 289942 270163
rect 289994 270151 290000 270163
rect 346000 270151 346006 270163
rect 289994 270123 346006 270151
rect 289994 270111 290000 270123
rect 346000 270111 346006 270123
rect 346058 270111 346064 270163
rect 356944 270111 356950 270163
rect 357002 270151 357008 270163
rect 512752 270151 512758 270163
rect 357002 270123 512758 270151
rect 357002 270111 357008 270123
rect 512752 270111 512758 270123
rect 512810 270111 512816 270163
rect 283312 270077 283318 270089
rect 265418 270049 269630 270077
rect 269794 270049 283318 270077
rect 265418 270037 265424 270049
rect 106000 269963 106006 270015
rect 106058 270003 106064 270015
rect 204208 270003 204214 270015
rect 106058 269975 204214 270003
rect 106058 269963 106064 269975
rect 204208 269963 204214 269975
rect 204266 269963 204272 270015
rect 210352 269963 210358 270015
rect 210410 270003 210416 270015
rect 225520 270003 225526 270015
rect 210410 269975 225526 270003
rect 210410 269963 210416 269975
rect 225520 269963 225526 269975
rect 225578 269963 225584 270015
rect 266512 269963 266518 270015
rect 266570 270003 266576 270015
rect 269602 270003 269630 270049
rect 283312 270037 283318 270049
rect 283370 270037 283376 270089
rect 291088 270037 291094 270089
rect 291146 270077 291152 270089
rect 349552 270077 349558 270089
rect 291146 270049 349558 270077
rect 291146 270037 291152 270049
rect 349552 270037 349558 270049
rect 349610 270037 349616 270089
rect 359824 270037 359830 270089
rect 359882 270077 359888 270089
rect 519760 270077 519766 270089
rect 359882 270049 519766 270077
rect 359882 270037 359888 270049
rect 519760 270037 519766 270049
rect 519818 270037 519824 270089
rect 672496 270037 672502 270089
rect 672554 270077 672560 270089
rect 676048 270077 676054 270089
rect 672554 270049 676054 270077
rect 672554 270037 672560 270049
rect 676048 270037 676054 270049
rect 676106 270037 676112 270089
rect 285712 270003 285718 270015
rect 266570 269975 269342 270003
rect 269602 269975 285718 270003
rect 266570 269963 266576 269975
rect 98896 269889 98902 269941
rect 98954 269929 98960 269941
rect 202288 269929 202294 269941
rect 98954 269901 202294 269929
rect 98954 269889 98960 269901
rect 202288 269889 202294 269901
rect 202346 269889 202352 269941
rect 207472 269889 207478 269941
rect 207530 269929 207536 269941
rect 221776 269929 221782 269941
rect 207530 269901 221782 269929
rect 207530 269889 207536 269901
rect 221776 269889 221782 269901
rect 221834 269889 221840 269941
rect 96592 269815 96598 269867
rect 96650 269855 96656 269867
rect 201616 269855 201622 269867
rect 96650 269827 201622 269855
rect 96650 269815 96656 269827
rect 201616 269815 201622 269827
rect 201674 269815 201680 269867
rect 210256 269815 210262 269867
rect 210314 269855 210320 269867
rect 226672 269855 226678 269867
rect 210314 269827 226678 269855
rect 210314 269815 210320 269827
rect 226672 269815 226678 269827
rect 226730 269815 226736 269867
rect 258640 269815 258646 269867
rect 258698 269855 258704 269867
rect 269200 269855 269206 269867
rect 258698 269827 269206 269855
rect 258698 269815 258704 269827
rect 269200 269815 269206 269827
rect 269258 269815 269264 269867
rect 269314 269855 269342 269975
rect 285712 269963 285718 269975
rect 285770 269963 285776 270015
rect 293968 269963 293974 270015
rect 294026 270003 294032 270015
rect 356656 270003 356662 270015
rect 294026 269975 356662 270003
rect 294026 269963 294032 269975
rect 356656 269963 356662 269975
rect 356714 269963 356720 270015
rect 360976 269963 360982 270015
rect 361034 270003 361040 270015
rect 522160 270003 522166 270015
rect 361034 269975 522166 270003
rect 361034 269963 361040 269975
rect 522160 269963 522166 269975
rect 522218 269963 522224 270015
rect 269488 269889 269494 269941
rect 269546 269929 269552 269941
rect 289264 269929 289270 269941
rect 269546 269901 289270 269929
rect 269546 269889 269552 269901
rect 289264 269889 289270 269901
rect 289322 269889 289328 269941
rect 292240 269889 292246 269941
rect 292298 269929 292304 269941
rect 351856 269929 351862 269941
rect 292298 269901 351862 269929
rect 292298 269889 292304 269901
rect 351856 269889 351862 269901
rect 351914 269889 351920 269941
rect 363568 269889 363574 269941
rect 363626 269929 363632 269941
rect 529264 269929 529270 269941
rect 363626 269901 529270 269929
rect 363626 269889 363632 269901
rect 529264 269889 529270 269901
rect 529322 269889 529328 269941
rect 288016 269855 288022 269867
rect 269314 269827 288022 269855
rect 288016 269815 288022 269827
rect 288074 269815 288080 269867
rect 293488 269815 293494 269867
rect 293546 269855 293552 269867
rect 355504 269855 355510 269867
rect 293546 269827 355510 269855
rect 293546 269815 293552 269827
rect 355504 269815 355510 269827
rect 355562 269815 355568 269867
rect 362800 269815 362806 269867
rect 362858 269855 362864 269867
rect 526864 269855 526870 269867
rect 362858 269827 526870 269855
rect 362858 269815 362864 269827
rect 526864 269815 526870 269827
rect 526922 269815 526928 269867
rect 91792 269741 91798 269793
rect 91850 269781 91856 269793
rect 177040 269781 177046 269793
rect 91850 269753 177046 269781
rect 91850 269741 91856 269753
rect 177040 269741 177046 269753
rect 177098 269741 177104 269793
rect 204016 269741 204022 269793
rect 204074 269781 204080 269793
rect 223408 269781 223414 269793
rect 204074 269753 223414 269781
rect 204074 269741 204080 269753
rect 223408 269741 223414 269753
rect 223466 269741 223472 269793
rect 268432 269741 268438 269793
rect 268490 269781 268496 269793
rect 292816 269781 292822 269793
rect 268490 269753 292822 269781
rect 268490 269741 268496 269753
rect 292816 269741 292822 269753
rect 292874 269741 292880 269793
rect 296464 269741 296470 269793
rect 296522 269781 296528 269793
rect 362608 269781 362614 269793
rect 296522 269753 362614 269781
rect 296522 269741 296528 269753
rect 362608 269741 362614 269753
rect 362666 269741 362672 269793
rect 365680 269741 365686 269793
rect 365738 269781 365744 269793
rect 533968 269781 533974 269793
rect 365738 269753 533974 269781
rect 365738 269741 365744 269753
rect 533968 269741 533974 269753
rect 534026 269741 534032 269793
rect 663760 269741 663766 269793
rect 663818 269781 663824 269793
rect 676240 269781 676246 269793
rect 663818 269753 676246 269781
rect 663818 269741 663824 269753
rect 676240 269741 676246 269753
rect 676298 269741 676304 269793
rect 88336 269667 88342 269719
rect 88394 269707 88400 269719
rect 199216 269707 199222 269719
rect 88394 269679 199222 269707
rect 88394 269667 88400 269679
rect 199216 269667 199222 269679
rect 199274 269667 199280 269719
rect 205840 269667 205846 269719
rect 205898 269707 205904 269719
rect 226000 269707 226006 269719
rect 205898 269679 226006 269707
rect 205898 269667 205904 269679
rect 226000 269667 226006 269679
rect 226058 269667 226064 269719
rect 255760 269667 255766 269719
rect 255818 269707 255824 269719
rect 262096 269707 262102 269719
rect 255818 269679 262102 269707
rect 255818 269667 255824 269679
rect 262096 269667 262102 269679
rect 262154 269667 262160 269719
rect 267280 269667 267286 269719
rect 267338 269707 267344 269719
rect 290416 269707 290422 269719
rect 267338 269679 290422 269707
rect 267338 269667 267344 269679
rect 290416 269667 290422 269679
rect 290474 269667 290480 269719
rect 297040 269667 297046 269719
rect 297098 269707 297104 269719
rect 363760 269707 363766 269719
rect 297098 269679 363766 269707
rect 297098 269667 297104 269679
rect 363760 269667 363766 269679
rect 363818 269667 363824 269719
rect 366544 269667 366550 269719
rect 366602 269707 366608 269719
rect 536368 269707 536374 269719
rect 366602 269679 536374 269707
rect 366602 269667 366608 269679
rect 536368 269667 536374 269679
rect 536426 269667 536432 269719
rect 85936 269593 85942 269645
rect 85994 269633 86000 269645
rect 198544 269633 198550 269645
rect 85994 269605 198550 269633
rect 85994 269593 86000 269605
rect 198544 269593 198550 269605
rect 198602 269593 198608 269645
rect 198640 269593 198646 269645
rect 198698 269633 198704 269645
rect 221200 269633 221206 269645
rect 198698 269605 221206 269633
rect 198698 269593 198704 269605
rect 221200 269593 221206 269605
rect 221258 269593 221264 269645
rect 249040 269593 249046 269645
rect 249098 269633 249104 269645
rect 250288 269633 250294 269645
rect 249098 269605 250294 269633
rect 249098 269593 249104 269605
rect 250288 269593 250294 269605
rect 250346 269593 250352 269645
rect 269200 269593 269206 269645
rect 269258 269633 269264 269645
rect 295120 269633 295126 269645
rect 269258 269605 295126 269633
rect 269258 269593 269264 269605
rect 295120 269593 295126 269605
rect 295178 269593 295184 269645
rect 299632 269593 299638 269645
rect 299690 269633 299696 269645
rect 299690 269605 367262 269633
rect 299690 269593 299696 269605
rect 83536 269519 83542 269571
rect 83594 269559 83600 269571
rect 198064 269559 198070 269571
rect 83594 269531 198070 269559
rect 83594 269519 83600 269531
rect 198064 269519 198070 269531
rect 198122 269519 198128 269571
rect 206512 269519 206518 269571
rect 206570 269559 206576 269571
rect 233392 269559 233398 269571
rect 206570 269531 233398 269559
rect 206570 269519 206576 269531
rect 233392 269519 233398 269531
rect 233450 269519 233456 269571
rect 253360 269519 253366 269571
rect 253418 269559 253424 269571
rect 256144 269559 256150 269571
rect 253418 269531 256150 269559
rect 253418 269519 253424 269531
rect 256144 269519 256150 269531
rect 256202 269519 256208 269571
rect 267088 269519 267094 269571
rect 267146 269559 267152 269571
rect 269488 269559 269494 269571
rect 267146 269531 269494 269559
rect 267146 269519 267152 269531
rect 269488 269519 269494 269531
rect 269546 269519 269552 269571
rect 269680 269519 269686 269571
rect 269738 269559 269744 269571
rect 296368 269559 296374 269571
rect 269738 269531 296374 269559
rect 269738 269519 269744 269531
rect 296368 269519 296374 269531
rect 296426 269519 296432 269571
rect 302608 269519 302614 269571
rect 302666 269559 302672 269571
rect 367120 269559 367126 269571
rect 302666 269531 367126 269559
rect 302666 269519 302672 269531
rect 367120 269519 367126 269531
rect 367178 269519 367184 269571
rect 367234 269559 367262 269605
rect 369616 269593 369622 269645
rect 369674 269633 369680 269645
rect 543472 269633 543478 269645
rect 369674 269605 543478 269633
rect 369674 269593 369680 269605
rect 543472 269593 543478 269605
rect 543530 269593 543536 269645
rect 370864 269559 370870 269571
rect 367234 269531 370870 269559
rect 370864 269519 370870 269531
rect 370922 269519 370928 269571
rect 384976 269559 384982 269571
rect 377266 269531 384982 269559
rect 76432 269445 76438 269497
rect 76490 269485 76496 269497
rect 195664 269485 195670 269497
rect 76490 269457 195670 269485
rect 76490 269445 76496 269457
rect 195664 269445 195670 269457
rect 195722 269445 195728 269497
rect 204112 269445 204118 269497
rect 204170 269485 204176 269497
rect 232144 269485 232150 269497
rect 204170 269457 232150 269485
rect 204170 269445 204176 269457
rect 232144 269445 232150 269457
rect 232202 269445 232208 269497
rect 256240 269445 256246 269497
rect 256298 269485 256304 269497
rect 263248 269485 263254 269497
rect 256298 269457 263254 269485
rect 256298 269445 256304 269457
rect 263248 269445 263254 269457
rect 263306 269445 263312 269497
rect 267760 269445 267766 269497
rect 267818 269485 267824 269497
rect 291664 269485 291670 269497
rect 267818 269457 291670 269485
rect 267818 269445 267824 269457
rect 291664 269445 291670 269457
rect 291722 269445 291728 269497
rect 305680 269445 305686 269497
rect 305738 269485 305744 269497
rect 377266 269485 377294 269531
rect 384976 269519 384982 269531
rect 385034 269519 385040 269571
rect 567088 269559 567094 269571
rect 385090 269531 567094 269559
rect 305738 269457 377294 269485
rect 305738 269445 305744 269457
rect 78832 269371 78838 269423
rect 78890 269411 78896 269423
rect 196624 269411 196630 269423
rect 78890 269383 196630 269411
rect 78890 269371 78896 269383
rect 196624 269371 196630 269383
rect 196682 269371 196688 269423
rect 202960 269371 202966 269423
rect 203018 269411 203024 269423
rect 231952 269411 231958 269423
rect 203018 269383 231958 269411
rect 203018 269371 203024 269383
rect 231952 269371 231958 269383
rect 232010 269371 232016 269423
rect 268624 269371 268630 269423
rect 268682 269411 268688 269423
rect 294064 269411 294070 269423
rect 268682 269383 294070 269411
rect 268682 269371 268688 269383
rect 294064 269371 294070 269383
rect 294122 269371 294128 269423
rect 308272 269371 308278 269423
rect 308330 269411 308336 269423
rect 308330 269383 379070 269411
rect 308330 269371 308336 269383
rect 74032 269297 74038 269349
rect 74090 269337 74096 269349
rect 194992 269337 194998 269349
rect 74090 269309 194998 269337
rect 74090 269297 74096 269309
rect 194992 269297 194998 269309
rect 195050 269297 195056 269349
rect 200560 269297 200566 269349
rect 200618 269337 200624 269349
rect 230992 269337 230998 269349
rect 200618 269309 230998 269337
rect 200618 269297 200624 269309
rect 230992 269297 230998 269309
rect 231050 269297 231056 269349
rect 258160 269297 258166 269349
rect 258218 269337 258224 269349
rect 267952 269337 267958 269349
rect 258218 269309 267958 269337
rect 258218 269297 258224 269309
rect 267952 269297 267958 269309
rect 268010 269297 268016 269349
rect 274672 269297 274678 269349
rect 274730 269337 274736 269349
rect 308176 269337 308182 269349
rect 274730 269309 308182 269337
rect 274730 269297 274736 269309
rect 308176 269297 308182 269309
rect 308234 269297 308240 269349
rect 367120 269297 367126 269349
rect 367178 269337 367184 269349
rect 377968 269337 377974 269349
rect 367178 269309 377974 269337
rect 367178 269297 367184 269309
rect 377968 269297 377974 269309
rect 378026 269297 378032 269349
rect 379042 269337 379070 269383
rect 379120 269371 379126 269423
rect 379178 269411 379184 269423
rect 385090 269411 385118 269531
rect 567088 269519 567094 269531
rect 567146 269519 567152 269571
rect 580048 269485 580054 269497
rect 379178 269383 385118 269411
rect 392674 269457 580054 269485
rect 379178 269371 379184 269383
rect 392080 269337 392086 269349
rect 379042 269309 392086 269337
rect 392080 269297 392086 269309
rect 392138 269297 392144 269349
rect 77680 269223 77686 269275
rect 77738 269263 77744 269275
rect 196144 269263 196150 269275
rect 77738 269235 196150 269263
rect 77738 269223 77744 269235
rect 196144 269223 196150 269235
rect 196202 269223 196208 269275
rect 197104 269223 197110 269275
rect 197162 269263 197168 269275
rect 229552 269263 229558 269275
rect 197162 269235 229558 269263
rect 197162 269223 197168 269235
rect 229552 269223 229558 269235
rect 229610 269223 229616 269275
rect 260080 269223 260086 269275
rect 260138 269263 260144 269275
rect 272656 269263 272662 269275
rect 260138 269235 272662 269263
rect 260138 269223 260144 269235
rect 272656 269223 272662 269235
rect 272714 269223 272720 269275
rect 384112 269223 384118 269275
rect 384170 269263 384176 269275
rect 392674 269263 392702 269457
rect 580048 269445 580054 269457
rect 580106 269445 580112 269497
rect 392752 269371 392758 269423
rect 392810 269411 392816 269423
rect 601360 269411 601366 269423
rect 392810 269383 601366 269411
rect 392810 269371 392816 269383
rect 601360 269371 601366 269383
rect 601418 269371 601424 269423
rect 398992 269297 398998 269349
rect 399050 269337 399056 269349
rect 615568 269337 615574 269349
rect 399050 269309 615574 269337
rect 399050 269297 399056 269309
rect 615568 269297 615574 269309
rect 615626 269297 615632 269349
rect 384170 269235 392702 269263
rect 384170 269223 384176 269235
rect 407248 269223 407254 269275
rect 407306 269263 407312 269275
rect 636784 269263 636790 269275
rect 407306 269235 636790 269263
rect 407306 269223 407312 269235
rect 636784 269223 636790 269235
rect 636842 269223 636848 269275
rect 135664 269149 135670 269201
rect 135722 269189 135728 269201
rect 212368 269189 212374 269201
rect 135722 269161 212374 269189
rect 135722 269149 135728 269161
rect 212368 269149 212374 269161
rect 212426 269149 212432 269201
rect 260560 269149 260566 269201
rect 260618 269189 260624 269201
rect 273808 269189 273814 269201
rect 260618 269161 273814 269189
rect 260618 269149 260624 269161
rect 273808 269149 273814 269161
rect 273866 269149 273872 269201
rect 281776 269149 281782 269201
rect 281834 269189 281840 269201
rect 325360 269189 325366 269201
rect 281834 269161 325366 269189
rect 281834 269149 281840 269161
rect 325360 269149 325366 269161
rect 325418 269149 325424 269201
rect 345424 269149 345430 269201
rect 345482 269189 345488 269201
rect 484240 269189 484246 269201
rect 345482 269161 484246 269189
rect 345482 269149 345488 269161
rect 484240 269149 484246 269161
rect 484298 269149 484304 269201
rect 666832 269149 666838 269201
rect 666890 269189 666896 269201
rect 676240 269189 676246 269201
rect 666890 269161 676246 269189
rect 666890 269149 666896 269161
rect 676240 269149 676246 269161
rect 676298 269149 676304 269201
rect 141520 269075 141526 269127
rect 141578 269115 141584 269127
rect 213808 269115 213814 269127
rect 141578 269087 213814 269115
rect 141578 269075 141584 269087
rect 213808 269075 213814 269087
rect 213866 269075 213872 269127
rect 259888 269075 259894 269127
rect 259946 269115 259952 269127
rect 271504 269115 271510 269127
rect 259946 269087 271510 269115
rect 259946 269075 259952 269087
rect 271504 269075 271510 269087
rect 271562 269075 271568 269127
rect 282544 269075 282550 269127
rect 282602 269115 282608 269127
rect 328240 269115 328246 269127
rect 282602 269087 328246 269115
rect 282602 269075 282608 269087
rect 328240 269075 328246 269087
rect 328298 269075 328304 269127
rect 346480 269075 346486 269127
rect 346538 269115 346544 269127
rect 486640 269115 486646 269127
rect 346538 269087 486646 269115
rect 346538 269075 346544 269087
rect 486640 269075 486646 269087
rect 486698 269075 486704 269127
rect 144976 269001 144982 269053
rect 145034 269041 145040 269053
rect 214480 269041 214486 269053
rect 145034 269013 214486 269041
rect 145034 269001 145040 269013
rect 214480 269001 214486 269013
rect 214538 269001 214544 269053
rect 261808 269001 261814 269053
rect 261866 269041 261872 269053
rect 276208 269041 276214 269053
rect 261866 269013 276214 269041
rect 261866 269001 261872 269013
rect 276208 269001 276214 269013
rect 276266 269001 276272 269053
rect 280144 269001 280150 269053
rect 280202 269041 280208 269053
rect 322384 269041 322390 269053
rect 280202 269013 322390 269041
rect 280202 269001 280208 269013
rect 322384 269001 322390 269013
rect 322442 269001 322448 269053
rect 343600 269001 343606 269053
rect 343658 269041 343664 269053
rect 479632 269041 479638 269053
rect 343658 269013 479638 269041
rect 343658 269001 343664 269013
rect 479632 269001 479638 269013
rect 479690 269001 479696 269053
rect 148624 268927 148630 268979
rect 148682 268967 148688 268979
rect 215728 268967 215734 268979
rect 148682 268939 215734 268967
rect 148682 268927 148688 268939
rect 215728 268927 215734 268939
rect 215786 268927 215792 268979
rect 278896 268927 278902 268979
rect 278954 268967 278960 268979
rect 318736 268967 318742 268979
rect 278954 268939 318742 268967
rect 278954 268927 278960 268939
rect 318736 268927 318742 268939
rect 318794 268927 318800 268979
rect 342640 268927 342646 268979
rect 342698 268967 342704 268979
rect 477232 268967 477238 268979
rect 342698 268939 477238 268967
rect 342698 268927 342704 268939
rect 477232 268927 477238 268939
rect 477290 268927 477296 268979
rect 152176 268853 152182 268905
rect 152234 268893 152240 268905
rect 216688 268893 216694 268905
rect 152234 268865 216694 268893
rect 152234 268853 152240 268865
rect 216688 268853 216694 268865
rect 216746 268853 216752 268905
rect 264112 268853 264118 268905
rect 264170 268893 264176 268905
rect 264170 268865 276494 268893
rect 264170 268853 264176 268865
rect 153328 268779 153334 268831
rect 153386 268819 153392 268831
rect 216880 268819 216886 268831
rect 153386 268791 216886 268819
rect 153386 268779 153392 268791
rect 216880 268779 216886 268791
rect 216938 268779 216944 268831
rect 257008 268779 257014 268831
rect 257066 268819 257072 268831
rect 264400 268819 264406 268831
rect 257066 268791 264406 268819
rect 257066 268779 257072 268791
rect 264400 268779 264406 268791
rect 264458 268779 264464 268831
rect 276466 268819 276494 268865
rect 277552 268853 277558 268905
rect 277610 268893 277616 268905
rect 315280 268893 315286 268905
rect 277610 268865 315286 268893
rect 277610 268853 277616 268865
rect 315280 268853 315286 268865
rect 315338 268853 315344 268905
rect 339760 268853 339766 268905
rect 339818 268893 339824 268905
rect 470128 268893 470134 268905
rect 339818 268865 470134 268893
rect 339818 268853 339824 268865
rect 470128 268853 470134 268865
rect 470186 268853 470192 268905
rect 282160 268819 282166 268831
rect 276466 268791 282166 268819
rect 282160 268779 282166 268791
rect 282218 268779 282224 268831
rect 283024 268779 283030 268831
rect 283082 268819 283088 268831
rect 313936 268819 313942 268831
rect 283082 268791 313942 268819
rect 283082 268779 283088 268791
rect 313936 268779 313942 268791
rect 313994 268779 314000 268831
rect 341008 268779 341014 268831
rect 341066 268819 341072 268831
rect 472528 268819 472534 268831
rect 341066 268791 472534 268819
rect 341066 268779 341072 268791
rect 472528 268779 472534 268791
rect 472586 268779 472592 268831
rect 160432 268705 160438 268757
rect 160490 268745 160496 268757
rect 218896 268745 218902 268757
rect 160490 268717 218902 268745
rect 160490 268705 160496 268717
rect 218896 268705 218902 268717
rect 218954 268705 218960 268757
rect 257680 268705 257686 268757
rect 257738 268745 257744 268757
rect 266800 268745 266806 268757
rect 257738 268717 266806 268745
rect 257738 268705 257744 268717
rect 266800 268705 266806 268717
rect 266858 268705 266864 268757
rect 282064 268705 282070 268757
rect 282122 268745 282128 268757
rect 299440 268745 299446 268757
rect 282122 268717 299446 268745
rect 282122 268705 282128 268717
rect 299440 268705 299446 268717
rect 299498 268705 299504 268757
rect 336880 268705 336886 268757
rect 336938 268745 336944 268757
rect 463024 268745 463030 268757
rect 336938 268717 463030 268745
rect 336938 268705 336944 268717
rect 463024 268705 463030 268717
rect 463082 268705 463088 268757
rect 159280 268631 159286 268683
rect 159338 268671 159344 268683
rect 218608 268671 218614 268683
rect 159338 268643 218614 268671
rect 159338 268631 159344 268643
rect 218608 268631 218614 268643
rect 218666 268631 218672 268683
rect 275824 268631 275830 268683
rect 275882 268671 275888 268683
rect 311728 268671 311734 268683
rect 275882 268643 311734 268671
rect 275882 268631 275888 268643
rect 311728 268631 311734 268643
rect 311786 268631 311792 268683
rect 334288 268631 334294 268683
rect 334346 268671 334352 268683
rect 455920 268671 455926 268683
rect 334346 268643 455926 268671
rect 334346 268631 334352 268643
rect 455920 268631 455926 268643
rect 455978 268631 455984 268683
rect 166384 268557 166390 268609
rect 166442 268597 166448 268609
rect 220528 268597 220534 268609
rect 166442 268569 220534 268597
rect 166442 268557 166448 268569
rect 220528 268557 220534 268569
rect 220586 268557 220592 268609
rect 331216 268557 331222 268609
rect 331274 268597 331280 268609
rect 448816 268597 448822 268609
rect 331274 268569 448822 268597
rect 331274 268557 331280 268569
rect 448816 268557 448822 268569
rect 448874 268557 448880 268609
rect 167536 268483 167542 268535
rect 167594 268523 167600 268535
rect 221008 268523 221014 268535
rect 167594 268495 221014 268523
rect 167594 268483 167600 268495
rect 221008 268483 221014 268495
rect 221066 268483 221072 268535
rect 253168 268483 253174 268535
rect 253226 268523 253232 268535
rect 254992 268523 254998 268535
rect 253226 268495 254998 268523
rect 253226 268483 253232 268495
rect 254992 268483 254998 268495
rect 255050 268483 255056 268535
rect 259408 268483 259414 268535
rect 259466 268523 259472 268535
rect 270352 268523 270358 268535
rect 259466 268495 270358 268523
rect 259466 268483 259472 268495
rect 270352 268483 270358 268495
rect 270410 268483 270416 268535
rect 328336 268483 328342 268535
rect 328394 268523 328400 268535
rect 441808 268523 441814 268535
rect 328394 268495 441814 268523
rect 328394 268483 328400 268495
rect 441808 268483 441814 268495
rect 441866 268483 441872 268535
rect 173392 268409 173398 268461
rect 173450 268449 173456 268461
rect 222352 268449 222358 268461
rect 173450 268421 222358 268449
rect 173450 268409 173456 268421
rect 222352 268409 222358 268421
rect 222410 268409 222416 268461
rect 325744 268409 325750 268461
rect 325802 268449 325808 268461
rect 434704 268449 434710 268461
rect 325802 268421 434710 268449
rect 325802 268409 325808 268421
rect 434704 268409 434710 268421
rect 434762 268409 434768 268461
rect 174640 268335 174646 268387
rect 174698 268375 174704 268387
rect 222832 268375 222838 268387
rect 174698 268347 222838 268375
rect 174698 268335 174704 268347
rect 222832 268335 222838 268347
rect 222890 268335 222896 268387
rect 247888 268335 247894 268387
rect 247946 268375 247952 268387
rect 249808 268375 249814 268387
rect 247946 268347 249814 268375
rect 247946 268335 247952 268347
rect 249808 268335 249814 268347
rect 249866 268335 249872 268387
rect 252688 268335 252694 268387
rect 252746 268375 252752 268387
rect 253840 268375 253846 268387
rect 252746 268347 253846 268375
rect 252746 268335 252752 268347
rect 253840 268335 253846 268347
rect 253898 268335 253904 268387
rect 261232 268335 261238 268387
rect 261290 268375 261296 268387
rect 275056 268375 275062 268387
rect 261290 268347 275062 268375
rect 261290 268335 261296 268347
rect 275056 268335 275062 268347
rect 275114 268335 275120 268387
rect 322576 268335 322582 268387
rect 322634 268375 322640 268387
rect 427600 268375 427606 268387
rect 322634 268347 427606 268375
rect 322634 268335 322640 268347
rect 427600 268335 427606 268347
rect 427658 268335 427664 268387
rect 177040 268261 177046 268313
rect 177098 268301 177104 268313
rect 200464 268301 200470 268313
rect 177098 268273 200470 268301
rect 177098 268261 177104 268273
rect 200464 268261 200470 268273
rect 200522 268261 200528 268313
rect 205360 268261 205366 268313
rect 205418 268301 205424 268313
rect 225232 268301 225238 268313
rect 205418 268273 225238 268301
rect 205418 268261 205424 268273
rect 225232 268261 225238 268273
rect 225290 268261 225296 268313
rect 257488 268261 257494 268313
rect 257546 268301 257552 268313
rect 265552 268301 265558 268313
rect 257546 268273 265558 268301
rect 257546 268261 257552 268273
rect 265552 268261 265558 268273
rect 265610 268261 265616 268313
rect 319696 268261 319702 268313
rect 319754 268301 319760 268313
rect 420496 268301 420502 268313
rect 319754 268273 420502 268301
rect 319754 268261 319760 268273
rect 420496 268261 420502 268273
rect 420554 268261 420560 268313
rect 180496 268187 180502 268239
rect 180554 268227 180560 268239
rect 205456 268227 205462 268239
rect 180554 268199 205462 268227
rect 180554 268187 180560 268199
rect 205456 268187 205462 268199
rect 205514 268187 205520 268239
rect 205648 268187 205654 268239
rect 205706 268227 205712 268239
rect 224080 268227 224086 268239
rect 205706 268199 224086 268227
rect 205706 268187 205712 268199
rect 224080 268187 224086 268199
rect 224138 268187 224144 268239
rect 224272 268187 224278 268239
rect 224330 268227 224336 268239
rect 231472 268227 231478 268239
rect 224330 268199 231478 268227
rect 224330 268187 224336 268199
rect 231472 268187 231478 268199
rect 231530 268187 231536 268239
rect 254608 268187 254614 268239
rect 254666 268227 254672 268239
rect 258544 268227 258550 268239
rect 254666 268199 258550 268227
rect 254666 268187 254672 268199
rect 258544 268187 258550 268199
rect 258602 268187 258608 268239
rect 263632 268187 263638 268239
rect 263690 268227 263696 268239
rect 281008 268227 281014 268239
rect 263690 268199 281014 268227
rect 263690 268187 263696 268199
rect 281008 268187 281014 268199
rect 281066 268187 281072 268239
rect 317104 268187 317110 268239
rect 317162 268227 317168 268239
rect 413392 268227 413398 268239
rect 317162 268199 413398 268227
rect 317162 268187 317168 268199
rect 413392 268187 413398 268199
rect 413450 268187 413456 268239
rect 184144 268113 184150 268165
rect 184202 268153 184208 268165
rect 205360 268153 205366 268165
rect 184202 268125 205366 268153
rect 184202 268113 184208 268125
rect 205360 268113 205366 268125
rect 205418 268113 205424 268165
rect 219280 268153 219286 268165
rect 205858 268125 219286 268153
rect 192976 268039 192982 268091
rect 193034 268079 193040 268091
rect 205858 268079 205886 268125
rect 219280 268113 219286 268125
rect 219338 268113 219344 268165
rect 224560 268113 224566 268165
rect 224618 268153 224624 268165
rect 228400 268153 228406 268165
rect 224618 268125 228406 268153
rect 224618 268113 224624 268125
rect 228400 268113 228406 268125
rect 228458 268113 228464 268165
rect 311152 268113 311158 268165
rect 311210 268153 311216 268165
rect 399184 268153 399190 268165
rect 311210 268125 399190 268153
rect 311210 268113 311216 268125
rect 399184 268113 399190 268125
rect 399242 268113 399248 268165
rect 193034 268051 205886 268079
rect 193034 268039 193040 268051
rect 207280 268039 207286 268091
rect 207338 268079 207344 268091
rect 213328 268079 213334 268091
rect 207338 268051 213334 268079
rect 207338 268039 207344 268051
rect 213328 268039 213334 268051
rect 213386 268039 213392 268091
rect 221488 268039 221494 268091
rect 221546 268079 221552 268091
rect 230416 268079 230422 268091
rect 221546 268051 230422 268079
rect 221546 268039 221552 268051
rect 230416 268039 230422 268051
rect 230474 268039 230480 268091
rect 314224 268039 314230 268091
rect 314282 268079 314288 268091
rect 406288 268079 406294 268091
rect 314282 268051 406294 268079
rect 314282 268039 314288 268051
rect 406288 268039 406294 268051
rect 406346 268039 406352 268091
rect 193168 267965 193174 268017
rect 193226 268005 193232 268017
rect 217360 268005 217366 268017
rect 193226 267977 217366 268005
rect 193226 267965 193232 267977
rect 217360 267965 217366 267977
rect 217418 267965 217424 268017
rect 221584 267965 221590 268017
rect 221642 268005 221648 268017
rect 229072 268005 229078 268017
rect 221642 267977 229078 268005
rect 221642 267965 221648 267977
rect 229072 267965 229078 267977
rect 229130 267965 229136 268017
rect 334960 267965 334966 268017
rect 335018 268005 335024 268017
rect 346864 268005 346870 268017
rect 335018 267977 346870 268005
rect 335018 267965 335024 267977
rect 346864 267965 346870 267977
rect 346922 267965 346928 268017
rect 207856 267891 207862 267943
rect 207914 267931 207920 267943
rect 219952 267931 219958 267943
rect 207914 267903 219958 267931
rect 207914 267891 207920 267903
rect 219952 267891 219958 267903
rect 220010 267891 220016 267943
rect 221968 267891 221974 267943
rect 222026 267931 222032 267943
rect 227632 267931 227638 267943
rect 222026 267903 227638 267931
rect 222026 267891 222032 267903
rect 227632 267891 227638 267903
rect 227690 267891 227696 267943
rect 255088 267891 255094 267943
rect 255146 267931 255152 267943
rect 259696 267931 259702 267943
rect 255146 267903 259702 267931
rect 255146 267891 255152 267903
rect 259696 267891 259702 267903
rect 259754 267891 259760 267943
rect 337840 267891 337846 267943
rect 337898 267931 337904 267943
rect 337898 267903 357134 267931
rect 337898 267891 337904 267903
rect 207760 267817 207766 267869
rect 207818 267857 207824 267869
rect 218128 267857 218134 267869
rect 207818 267829 218134 267857
rect 207818 267817 207824 267829
rect 218128 267817 218134 267829
rect 218186 267817 218192 267869
rect 221680 267817 221686 267869
rect 221738 267857 221744 267869
rect 227824 267857 227830 267869
rect 221738 267829 227830 267857
rect 221738 267817 221744 267829
rect 227824 267817 227830 267829
rect 227882 267817 227888 267869
rect 295216 267817 295222 267869
rect 295274 267857 295280 267869
rect 301840 267857 301846 267869
rect 295274 267829 301846 267857
rect 295274 267817 295280 267829
rect 301840 267817 301846 267829
rect 301898 267817 301904 267869
rect 339280 267817 339286 267869
rect 339338 267857 339344 267869
rect 354256 267857 354262 267869
rect 339338 267829 354262 267857
rect 339338 267817 339344 267829
rect 354256 267817 354262 267829
rect 354314 267817 354320 267869
rect 357106 267857 357134 267903
rect 359920 267857 359926 267869
rect 357106 267829 359926 267857
rect 359920 267817 359926 267829
rect 359978 267817 359984 267869
rect 359152 267743 359158 267795
rect 359210 267783 359216 267795
rect 517360 267783 517366 267795
rect 359210 267755 517366 267783
rect 359210 267743 359216 267755
rect 517360 267743 517366 267755
rect 517418 267743 517424 267795
rect 361744 267669 361750 267721
rect 361802 267709 361808 267721
rect 524464 267709 524470 267721
rect 361802 267681 524470 267709
rect 361802 267669 361808 267681
rect 524464 267669 524470 267681
rect 524522 267669 524528 267721
rect 364624 267595 364630 267647
rect 364682 267635 364688 267647
rect 531568 267635 531574 267647
rect 364682 267607 531574 267635
rect 364682 267595 364688 267607
rect 531568 267595 531574 267607
rect 531626 267595 531632 267647
rect 367696 267521 367702 267573
rect 367754 267561 367760 267573
rect 538768 267561 538774 267573
rect 367754 267533 538774 267561
rect 367754 267521 367760 267533
rect 538768 267521 538774 267533
rect 538826 267521 538832 267573
rect 370768 267447 370774 267499
rect 370826 267487 370832 267499
rect 547024 267487 547030 267499
rect 370826 267459 547030 267487
rect 370826 267447 370832 267459
rect 547024 267447 547030 267459
rect 547082 267447 547088 267499
rect 286096 267373 286102 267425
rect 286154 267413 286160 267425
rect 336496 267413 336502 267425
rect 286154 267385 336502 267413
rect 286154 267373 286160 267385
rect 336496 267373 336502 267385
rect 336554 267373 336560 267425
rect 372016 267373 372022 267425
rect 372074 267413 372080 267425
rect 549328 267413 549334 267425
rect 372074 267385 549334 267413
rect 372074 267373 372080 267385
rect 549328 267373 549334 267385
rect 549386 267373 549392 267425
rect 284464 267299 284470 267351
rect 284522 267339 284528 267351
rect 333040 267339 333046 267351
rect 284522 267311 333046 267339
rect 284522 267299 284528 267311
rect 333040 267299 333046 267311
rect 333098 267299 333104 267351
rect 373168 267299 373174 267351
rect 373226 267339 373232 267351
rect 552880 267339 552886 267351
rect 373226 267311 552886 267339
rect 373226 267299 373232 267311
rect 552880 267299 552886 267311
rect 552938 267299 552944 267351
rect 288688 267225 288694 267277
rect 288746 267265 288752 267277
rect 343312 267265 343318 267277
rect 288746 267237 343318 267265
rect 288746 267225 288752 267237
rect 343312 267225 343318 267237
rect 343370 267225 343376 267277
rect 373840 267225 373846 267277
rect 373898 267265 373904 267277
rect 554128 267265 554134 267277
rect 373898 267237 554134 267265
rect 373898 267225 373904 267237
rect 554128 267225 554134 267237
rect 554186 267225 554192 267277
rect 287344 267151 287350 267203
rect 287402 267191 287408 267203
rect 340144 267191 340150 267203
rect 287402 267163 340150 267191
rect 287402 267151 287408 267163
rect 340144 267151 340150 267163
rect 340202 267151 340208 267203
rect 374608 267151 374614 267203
rect 374666 267191 374672 267203
rect 556432 267191 556438 267203
rect 374666 267163 556438 267191
rect 374666 267151 374672 267163
rect 556432 267151 556438 267163
rect 556490 267151 556496 267203
rect 291568 267077 291574 267129
rect 291626 267117 291632 267129
rect 350704 267117 350710 267129
rect 291626 267089 350710 267117
rect 291626 267077 291632 267089
rect 350704 267077 350710 267089
rect 350762 267077 350768 267129
rect 377488 267077 377494 267129
rect 377546 267117 377552 267129
rect 563536 267117 563542 267129
rect 377546 267089 563542 267117
rect 377546 267077 377552 267089
rect 563536 267077 563542 267089
rect 563594 267077 563600 267129
rect 290416 267003 290422 267055
rect 290474 267043 290480 267055
rect 347248 267043 347254 267055
rect 290474 267015 347254 267043
rect 290474 267003 290480 267015
rect 347248 267003 347254 267015
rect 347306 267003 347312 267055
rect 376816 267003 376822 267055
rect 376874 267043 376880 267055
rect 561232 267043 561238 267055
rect 376874 267015 561238 267043
rect 376874 267003 376880 267015
rect 561232 267003 561238 267015
rect 561290 267003 561296 267055
rect 297808 266929 297814 266981
rect 297866 266969 297872 266981
rect 366064 266969 366070 266981
rect 297866 266941 366070 266969
rect 297866 266929 297872 266941
rect 366064 266929 366070 266941
rect 366122 266929 366128 266981
rect 376240 266929 376246 266981
rect 376298 266969 376304 266981
rect 559984 266969 559990 266981
rect 376298 266941 559990 266969
rect 376298 266929 376304 266941
rect 559984 266929 559990 266941
rect 560042 266929 560048 266981
rect 300688 266855 300694 266907
rect 300746 266895 300752 266907
rect 373264 266895 373270 266907
rect 300746 266867 373270 266895
rect 300746 266855 300752 266867
rect 373264 266855 373270 266867
rect 373322 266855 373328 266907
rect 379408 266855 379414 266907
rect 379466 266895 379472 266907
rect 568240 266895 568246 266907
rect 379466 266867 568246 266895
rect 379466 266855 379472 266867
rect 568240 266855 568246 266867
rect 568298 266855 568304 266907
rect 299440 266781 299446 266833
rect 299498 266821 299504 266833
rect 369328 266821 369334 266833
rect 299498 266793 369334 266821
rect 299498 266781 299504 266793
rect 369328 266781 369334 266793
rect 369386 266781 369392 266833
rect 382288 266781 382294 266833
rect 382346 266821 382352 266833
rect 575344 266821 575350 266833
rect 382346 266793 575350 266821
rect 382346 266781 382352 266793
rect 575344 266781 575350 266793
rect 575402 266781 575408 266833
rect 302032 266707 302038 266759
rect 302090 266747 302096 266759
rect 376720 266747 376726 266759
rect 302090 266719 376726 266747
rect 302090 266707 302096 266719
rect 376720 266707 376726 266719
rect 376778 266707 376784 266759
rect 385360 266707 385366 266759
rect 385418 266747 385424 266759
rect 582448 266747 582454 266759
rect 385418 266719 582454 266747
rect 385418 266707 385424 266719
rect 582448 266707 582454 266719
rect 582506 266707 582512 266759
rect 308752 266633 308758 266685
rect 308810 266673 308816 266685
rect 308810 266645 379454 266673
rect 308810 266633 308816 266645
rect 309232 266559 309238 266611
rect 309290 266599 309296 266611
rect 379426 266599 379454 266645
rect 392272 266633 392278 266685
rect 392330 266673 392336 266685
rect 600208 266673 600214 266685
rect 392330 266645 600214 266673
rect 392330 266633 392336 266645
rect 600208 266633 600214 266645
rect 600266 266633 600272 266685
rect 393328 266599 393334 266611
rect 309290 266571 379358 266599
rect 379426 266571 393334 266599
rect 309290 266559 309296 266571
rect 310672 266485 310678 266537
rect 310730 266525 310736 266537
rect 379330 266525 379358 266571
rect 393328 266559 393334 266571
rect 393386 266559 393392 266611
rect 394672 266559 394678 266611
rect 394730 266599 394736 266611
rect 606064 266599 606070 266611
rect 394730 266571 606070 266599
rect 394730 266559 394736 266571
rect 606064 266559 606070 266571
rect 606122 266559 606128 266611
rect 394480 266525 394486 266537
rect 310730 266497 377294 266525
rect 379330 266497 394486 266525
rect 310730 266485 310736 266497
rect 377266 266451 377294 266497
rect 394480 266485 394486 266497
rect 394538 266485 394544 266537
rect 398896 266485 398902 266537
rect 398954 266525 398960 266537
rect 616720 266525 616726 266537
rect 398954 266497 616726 266525
rect 398954 266485 398960 266497
rect 616720 266485 616726 266497
rect 616778 266485 616784 266537
rect 398032 266451 398038 266463
rect 377266 266423 398038 266451
rect 398032 266411 398038 266423
rect 398090 266411 398096 266463
rect 400624 266411 400630 266463
rect 400682 266451 400688 266463
rect 620272 266451 620278 266463
rect 400682 266423 620278 266451
rect 400682 266411 400688 266423
rect 620272 266411 620278 266423
rect 620330 266411 620336 266463
rect 187216 266337 187222 266389
rect 187274 266377 187280 266389
rect 189712 266377 189718 266389
rect 187274 266349 189718 266377
rect 187274 266337 187280 266349
rect 189712 266337 189718 266349
rect 189770 266337 189776 266389
rect 312304 266337 312310 266389
rect 312362 266377 312368 266389
rect 401584 266377 401590 266389
rect 312362 266349 401590 266377
rect 312362 266337 312368 266349
rect 401584 266337 401590 266349
rect 401642 266337 401648 266389
rect 403216 266337 403222 266389
rect 403274 266377 403280 266389
rect 627376 266377 627382 266389
rect 403274 266349 627382 266377
rect 403274 266337 403280 266349
rect 627376 266337 627382 266349
rect 627434 266337 627440 266389
rect 354832 266263 354838 266315
rect 354890 266303 354896 266315
rect 506512 266303 506518 266315
rect 354890 266275 506518 266303
rect 354890 266263 354896 266275
rect 506512 266263 506518 266275
rect 506570 266263 506576 266315
rect 351952 266189 351958 266241
rect 352010 266229 352016 266241
rect 499696 266229 499702 266241
rect 352010 266201 499702 266229
rect 352010 266189 352016 266201
rect 499696 266189 499702 266201
rect 499754 266189 499760 266241
rect 348880 266115 348886 266167
rect 348938 266155 348944 266167
rect 492592 266155 492598 266167
rect 348938 266127 492598 266155
rect 348938 266115 348944 266127
rect 492592 266115 492598 266127
rect 492650 266115 492656 266167
rect 346000 266041 346006 266093
rect 346058 266081 346064 266093
rect 485488 266081 485494 266093
rect 346058 266053 485494 266081
rect 346058 266041 346064 266053
rect 485488 266041 485494 266053
rect 485546 266041 485552 266093
rect 343312 265967 343318 266019
rect 343370 266007 343376 266019
rect 478384 266007 478390 266019
rect 343370 265979 478390 266007
rect 343370 265967 343376 265979
rect 478384 265967 478390 265979
rect 478442 265967 478448 266019
rect 340240 265893 340246 265945
rect 340298 265933 340304 265945
rect 471280 265933 471286 265945
rect 340298 265905 471286 265933
rect 340298 265893 340304 265905
rect 471280 265893 471286 265905
rect 471338 265893 471344 265945
rect 337360 265819 337366 265871
rect 337418 265859 337424 265871
rect 464272 265859 464278 265871
rect 337418 265831 464278 265859
rect 337418 265819 337424 265831
rect 464272 265819 464278 265831
rect 464330 265819 464336 265871
rect 334768 265745 334774 265797
rect 334826 265785 334832 265797
rect 457168 265785 457174 265797
rect 334826 265757 457174 265785
rect 334826 265745 334832 265757
rect 457168 265745 457174 265757
rect 457226 265745 457232 265797
rect 331888 265671 331894 265723
rect 331946 265711 331952 265723
rect 450064 265711 450070 265723
rect 331946 265683 450070 265711
rect 331946 265671 331952 265683
rect 450064 265671 450070 265683
rect 450122 265671 450128 265723
rect 328816 265597 328822 265649
rect 328874 265637 328880 265649
rect 442960 265637 442966 265649
rect 328874 265609 442966 265637
rect 328874 265597 328880 265609
rect 442960 265597 442966 265609
rect 443018 265597 443024 265649
rect 324496 265523 324502 265575
rect 324554 265563 324560 265575
rect 432304 265563 432310 265575
rect 324554 265535 432310 265563
rect 324554 265523 324560 265535
rect 432304 265523 432310 265535
rect 432362 265523 432368 265575
rect 323344 265449 323350 265501
rect 323402 265489 323408 265501
rect 428848 265489 428854 265501
rect 323402 265461 428854 265489
rect 323402 265449 323408 265461
rect 428848 265449 428854 265461
rect 428906 265449 428912 265501
rect 313072 265375 313078 265427
rect 313130 265415 313136 265427
rect 403984 265415 403990 265427
rect 313130 265387 403990 265415
rect 313130 265375 313136 265387
rect 403984 265375 403990 265387
rect 404042 265375 404048 265427
rect 406576 265375 406582 265427
rect 406634 265415 406640 265427
rect 509200 265415 509206 265427
rect 406634 265387 509206 265415
rect 406634 265375 406640 265387
rect 509200 265375 509206 265387
rect 509258 265375 509264 265427
rect 319024 265301 319030 265353
rect 319082 265341 319088 265353
rect 418096 265341 418102 265353
rect 319082 265313 418102 265341
rect 319082 265301 319088 265313
rect 418096 265301 418102 265313
rect 418154 265301 418160 265353
rect 314896 265227 314902 265279
rect 314954 265267 314960 265279
rect 408688 265267 408694 265279
rect 314954 265239 408694 265267
rect 314954 265227 314960 265239
rect 408688 265227 408694 265239
rect 408746 265227 408752 265279
rect 354256 264931 354262 264983
rect 354314 264971 354320 264983
rect 468880 264971 468886 264983
rect 354314 264943 468886 264971
rect 354314 264931 354320 264943
rect 468880 264931 468886 264943
rect 468938 264931 468944 264983
rect 346864 264857 346870 264909
rect 346922 264897 346928 264909
rect 458320 264897 458326 264909
rect 346922 264869 458326 264897
rect 346922 264857 346928 264869
rect 458320 264857 458326 264869
rect 458378 264857 458384 264909
rect 359920 264783 359926 264835
rect 359978 264823 359984 264835
rect 465424 264823 465430 264835
rect 359978 264795 465430 264823
rect 359978 264783 359984 264795
rect 465424 264783 465430 264795
rect 465482 264783 465488 264835
rect 142384 262415 142390 262467
rect 142442 262455 142448 262467
rect 142672 262455 142678 262467
rect 142442 262427 142678 262455
rect 142442 262415 142448 262427
rect 142672 262415 142678 262427
rect 142730 262415 142736 262467
rect 420400 262119 420406 262171
rect 420458 262159 420464 262171
rect 606160 262159 606166 262171
rect 420458 262131 606166 262159
rect 420458 262119 420464 262131
rect 606160 262119 606166 262131
rect 606218 262119 606224 262171
rect 674608 261379 674614 261431
rect 674666 261419 674672 261431
rect 676240 261419 676246 261431
rect 674666 261391 676246 261419
rect 674666 261379 674672 261391
rect 676240 261379 676246 261391
rect 676298 261379 676304 261431
rect 41584 259677 41590 259729
rect 41642 259717 41648 259729
rect 50416 259717 50422 259729
rect 41642 259689 50422 259717
rect 41642 259677 41648 259689
rect 50416 259677 50422 259689
rect 50474 259677 50480 259729
rect 674704 259307 674710 259359
rect 674762 259347 674768 259359
rect 676048 259347 676054 259359
rect 674762 259319 676054 259347
rect 674762 259307 674768 259319
rect 676048 259307 676054 259319
rect 676106 259307 676112 259359
rect 420400 259233 420406 259285
rect 420458 259273 420464 259285
rect 603280 259273 603286 259285
rect 420458 259245 603286 259273
rect 420458 259233 420464 259245
rect 603280 259233 603286 259245
rect 603338 259233 603344 259285
rect 43216 259159 43222 259211
rect 43274 259199 43280 259211
rect 44848 259199 44854 259211
rect 43274 259171 44854 259199
rect 43274 259159 43280 259171
rect 44848 259159 44854 259171
rect 44906 259159 44912 259211
rect 41776 258937 41782 258989
rect 41834 258977 41840 258989
rect 53392 258977 53398 258989
rect 41834 258949 53398 258977
rect 41834 258937 41840 258949
rect 53392 258937 53398 258949
rect 53450 258937 53456 258989
rect 41776 258345 41782 258397
rect 41834 258385 41840 258397
rect 47728 258385 47734 258397
rect 41834 258357 47734 258385
rect 41834 258345 41840 258357
rect 47728 258345 47734 258357
rect 47786 258345 47792 258397
rect 41776 257975 41782 258027
rect 41834 258015 41840 258027
rect 43600 258015 43606 258027
rect 41834 257987 43606 258015
rect 41834 257975 41840 257987
rect 43600 257975 43606 257987
rect 43658 257975 43664 258027
rect 41776 257383 41782 257435
rect 41834 257423 41840 257435
rect 43504 257423 43510 257435
rect 41834 257395 43510 257423
rect 41834 257383 41840 257395
rect 43504 257383 43510 257395
rect 43562 257383 43568 257435
rect 41776 256865 41782 256917
rect 41834 256905 41840 256917
rect 43216 256905 43222 256917
rect 41834 256877 43222 256905
rect 41834 256865 41840 256877
rect 43216 256865 43222 256877
rect 43274 256865 43280 256917
rect 41776 256495 41782 256547
rect 41834 256535 41840 256547
rect 43408 256535 43414 256547
rect 41834 256507 43414 256535
rect 41834 256495 41840 256507
rect 43408 256495 43414 256507
rect 43466 256495 43472 256547
rect 674032 256421 674038 256473
rect 674090 256461 674096 256473
rect 676048 256461 676054 256473
rect 674090 256433 676054 256461
rect 674090 256421 674096 256433
rect 676048 256421 676054 256433
rect 676106 256421 676112 256473
rect 420400 256347 420406 256399
rect 420458 256387 420464 256399
rect 603376 256387 603382 256399
rect 420458 256359 603382 256387
rect 420458 256347 420464 256359
rect 603376 256347 603382 256359
rect 603434 256347 603440 256399
rect 646480 256347 646486 256399
rect 646538 256387 646544 256399
rect 679696 256387 679702 256399
rect 646538 256359 679702 256387
rect 646538 256347 646544 256359
rect 679696 256347 679702 256359
rect 679754 256347 679760 256399
rect 41776 255903 41782 255955
rect 41834 255943 41840 255955
rect 43408 255943 43414 255955
rect 41834 255915 43414 255943
rect 41834 255903 41840 255915
rect 43408 255903 43414 255915
rect 43466 255903 43472 255955
rect 41776 255385 41782 255437
rect 41834 255425 41840 255437
rect 43312 255425 43318 255437
rect 41834 255397 43318 255425
rect 41834 255385 41840 255397
rect 43312 255385 43318 255397
rect 43370 255385 43376 255437
rect 43408 255385 43414 255437
rect 43466 255425 43472 255437
rect 44752 255425 44758 255437
rect 43466 255397 44758 255425
rect 43466 255385 43472 255397
rect 44752 255385 44758 255397
rect 44810 255385 44816 255437
rect 420400 253461 420406 253513
rect 420458 253501 420464 253513
rect 603472 253501 603478 253513
rect 420458 253473 603478 253501
rect 420458 253461 420464 253473
rect 603472 253461 603478 253473
rect 603530 253461 603536 253513
rect 675664 251167 675670 251219
rect 675722 251167 675728 251219
rect 675760 251167 675766 251219
rect 675818 251167 675824 251219
rect 675682 250997 675710 251167
rect 675664 250945 675670 250997
rect 675722 250945 675728 250997
rect 420400 250575 420406 250627
rect 420458 250615 420464 250627
rect 603568 250615 603574 250627
rect 420458 250587 603574 250615
rect 420458 250575 420464 250587
rect 603568 250575 603574 250587
rect 603626 250575 603632 250627
rect 675778 250257 675806 251167
rect 675760 250205 675766 250257
rect 675818 250205 675824 250257
rect 120880 249465 120886 249517
rect 120938 249505 120944 249517
rect 145552 249505 145558 249517
rect 120938 249477 145558 249505
rect 120938 249465 120944 249477
rect 145552 249465 145558 249477
rect 145610 249465 145616 249517
rect 48016 249391 48022 249443
rect 48074 249431 48080 249443
rect 186832 249431 186838 249443
rect 48074 249403 186838 249431
rect 48074 249391 48080 249403
rect 186832 249391 186838 249403
rect 186890 249391 186896 249443
rect 47632 249317 47638 249369
rect 47690 249357 47696 249369
rect 186736 249357 186742 249369
rect 47690 249329 186742 249357
rect 47690 249317 47696 249329
rect 186736 249317 186742 249329
rect 186794 249317 186800 249369
rect 41584 249243 41590 249295
rect 41642 249283 41648 249295
rect 43120 249283 43126 249295
rect 41642 249255 43126 249283
rect 41642 249243 41648 249255
rect 43120 249243 43126 249255
rect 43178 249243 43184 249295
rect 47824 249243 47830 249295
rect 47882 249283 47888 249295
rect 186928 249283 186934 249295
rect 47882 249255 186934 249283
rect 47882 249243 47888 249255
rect 186928 249243 186934 249255
rect 186986 249243 186992 249295
rect 47920 249169 47926 249221
rect 47978 249209 47984 249221
rect 187024 249209 187030 249221
rect 47978 249181 187030 249209
rect 47978 249169 47984 249181
rect 187024 249169 187030 249181
rect 187082 249169 187088 249221
rect 44464 249095 44470 249147
rect 44522 249135 44528 249147
rect 186448 249135 186454 249147
rect 44522 249107 186454 249135
rect 44522 249095 44528 249107
rect 186448 249095 186454 249107
rect 186506 249095 186512 249147
rect 41584 248355 41590 248407
rect 41642 248395 41648 248407
rect 42832 248395 42838 248407
rect 41642 248367 42838 248395
rect 41642 248355 41648 248367
rect 42832 248355 42838 248367
rect 42890 248355 42896 248407
rect 41584 248059 41590 248111
rect 41642 248099 41648 248111
rect 42928 248099 42934 248111
rect 41642 248071 42934 248099
rect 41642 248059 41648 248071
rect 42928 248059 42934 248071
rect 42986 248059 42992 248111
rect 41776 247911 41782 247963
rect 41834 247951 41840 247963
rect 42736 247951 42742 247963
rect 41834 247923 42742 247951
rect 41834 247911 41840 247923
rect 42736 247911 42742 247923
rect 42794 247911 42800 247963
rect 41968 247837 41974 247889
rect 42026 247877 42032 247889
rect 43024 247877 43030 247889
rect 42026 247849 43030 247877
rect 42026 247837 42032 247849
rect 43024 247837 43030 247849
rect 43082 247837 43088 247889
rect 420304 247763 420310 247815
rect 420362 247803 420368 247815
rect 600400 247803 600406 247815
rect 420362 247775 600406 247803
rect 420362 247763 420368 247775
rect 600400 247763 600406 247775
rect 600458 247763 600464 247815
rect 41584 247689 41590 247741
rect 41642 247729 41648 247741
rect 157072 247729 157078 247741
rect 41642 247701 157078 247729
rect 41642 247689 41648 247701
rect 157072 247689 157078 247701
rect 157130 247689 157136 247741
rect 420400 247689 420406 247741
rect 420458 247729 420464 247741
rect 626320 247729 626326 247741
rect 420458 247701 626326 247729
rect 420458 247689 420464 247701
rect 626320 247689 626326 247701
rect 626378 247689 626384 247741
rect 674608 247023 674614 247075
rect 674666 247063 674672 247075
rect 675472 247063 675478 247075
rect 674666 247035 675478 247063
rect 674666 247023 674672 247035
rect 675472 247023 675478 247035
rect 675530 247023 675536 247075
rect 118000 246949 118006 247001
rect 118058 246989 118064 247001
rect 145648 246989 145654 247001
rect 118058 246961 145654 246989
rect 118058 246949 118064 246961
rect 145648 246949 145654 246961
rect 145706 246949 145712 247001
rect 123760 246875 123766 246927
rect 123818 246915 123824 246927
rect 168496 246915 168502 246927
rect 123818 246887 168502 246915
rect 123818 246875 123824 246887
rect 168496 246875 168502 246887
rect 168554 246875 168560 246927
rect 77488 246801 77494 246853
rect 77546 246841 77552 246853
rect 145456 246841 145462 246853
rect 77546 246813 145462 246841
rect 77546 246801 77552 246813
rect 145456 246801 145462 246813
rect 145514 246801 145520 246853
rect 69040 246727 69046 246779
rect 69098 246767 69104 246779
rect 145744 246767 145750 246779
rect 69098 246739 145750 246767
rect 69098 246727 69104 246739
rect 145744 246727 145750 246739
rect 145802 246727 145808 246779
rect 47440 246653 47446 246705
rect 47498 246693 47504 246705
rect 186640 246693 186646 246705
rect 47498 246665 186646 246693
rect 47498 246653 47504 246665
rect 186640 246653 186646 246665
rect 186698 246653 186704 246705
rect 45904 246579 45910 246631
rect 45962 246619 45968 246631
rect 186160 246619 186166 246631
rect 45962 246591 186166 246619
rect 45962 246579 45968 246591
rect 186160 246579 186166 246591
rect 186218 246579 186224 246631
rect 46000 246505 46006 246557
rect 46058 246545 46064 246557
rect 186544 246545 186550 246557
rect 46058 246517 186550 246545
rect 46058 246505 46064 246517
rect 186544 246505 186550 246517
rect 186602 246505 186608 246557
rect 45424 246431 45430 246483
rect 45482 246471 45488 246483
rect 186064 246471 186070 246483
rect 45482 246443 186070 246471
rect 45482 246431 45488 246443
rect 186064 246431 186070 246443
rect 186122 246431 186128 246483
rect 45616 246357 45622 246409
rect 45674 246397 45680 246409
rect 186352 246397 186358 246409
rect 45674 246369 186358 246397
rect 45674 246357 45680 246369
rect 186352 246357 186358 246369
rect 186410 246357 186416 246409
rect 45520 246283 45526 246335
rect 45578 246323 45584 246335
rect 186256 246323 186262 246335
rect 45578 246295 186262 246323
rect 45578 246283 45584 246295
rect 186256 246283 186262 246295
rect 186314 246283 186320 246335
rect 45040 246209 45046 246261
rect 45098 246249 45104 246261
rect 185872 246249 185878 246261
rect 45098 246221 185878 246249
rect 45098 246209 45104 246221
rect 185872 246209 185878 246221
rect 185930 246209 185936 246261
rect 41584 244803 41590 244855
rect 41642 244843 41648 244855
rect 156976 244843 156982 244855
rect 41642 244815 156982 244843
rect 41642 244803 41648 244815
rect 156976 244803 156982 244815
rect 157034 244803 157040 244855
rect 420400 244803 420406 244855
rect 420458 244843 420464 244855
rect 629200 244843 629206 244855
rect 420458 244815 629206 244843
rect 420458 244803 420464 244815
rect 629200 244803 629206 244815
rect 629258 244803 629264 244855
rect 41680 243323 41686 243375
rect 41738 243363 41744 243375
rect 185584 243363 185590 243375
rect 41738 243335 185590 243363
rect 41738 243323 41744 243335
rect 185584 243323 185590 243335
rect 185642 243323 185648 243375
rect 674704 242953 674710 243005
rect 674762 242993 674768 243005
rect 675376 242993 675382 243005
rect 674762 242965 675382 242993
rect 674762 242953 674768 242965
rect 675376 242953 675382 242965
rect 675434 242953 675440 243005
rect 45040 242805 45046 242857
rect 45098 242845 45104 242857
rect 185296 242845 185302 242857
rect 45098 242817 185302 242845
rect 45098 242805 45104 242817
rect 185296 242805 185302 242817
rect 185354 242805 185360 242857
rect 45328 242731 45334 242783
rect 45386 242771 45392 242783
rect 185968 242771 185974 242783
rect 45386 242743 185974 242771
rect 45386 242731 45392 242743
rect 185968 242731 185974 242743
rect 186026 242731 186032 242783
rect 44848 242657 44854 242709
rect 44906 242697 44912 242709
rect 185488 242697 185494 242709
rect 44906 242669 185494 242697
rect 44906 242657 44912 242669
rect 185488 242657 185494 242669
rect 185546 242657 185552 242709
rect 44752 242583 44758 242635
rect 44810 242623 44816 242635
rect 185776 242623 185782 242635
rect 44810 242595 185782 242623
rect 44810 242583 44816 242595
rect 185776 242583 185782 242595
rect 185834 242583 185840 242635
rect 149392 241917 149398 241969
rect 149450 241957 149456 241969
rect 168400 241957 168406 241969
rect 149450 241929 168406 241957
rect 149450 241917 149456 241929
rect 168400 241917 168406 241929
rect 168458 241917 168464 241969
rect 420400 241917 420406 241969
rect 420458 241957 420464 241969
rect 600496 241957 600502 241969
rect 420458 241929 600502 241957
rect 420458 241917 420464 241929
rect 600496 241917 600502 241929
rect 600554 241917 600560 241969
rect 674032 241769 674038 241821
rect 674090 241809 674096 241821
rect 675280 241809 675286 241821
rect 674090 241781 675286 241809
rect 674090 241769 674096 241781
rect 675280 241769 675286 241781
rect 675338 241769 675344 241821
rect 41872 240585 41878 240637
rect 41930 240585 41936 240637
rect 41890 240415 41918 240585
rect 41872 240363 41878 240415
rect 41930 240363 41936 240415
rect 383056 239623 383062 239675
rect 383114 239663 383120 239675
rect 464752 239663 464758 239675
rect 383114 239635 464758 239663
rect 383114 239623 383120 239635
rect 464752 239623 464758 239635
rect 464810 239623 464816 239675
rect 352816 239549 352822 239601
rect 352874 239589 352880 239601
rect 439120 239589 439126 239601
rect 352874 239561 439126 239589
rect 352874 239549 352880 239561
rect 439120 239549 439126 239561
rect 439178 239549 439184 239601
rect 363232 239475 363238 239527
rect 363290 239515 363296 239527
rect 378832 239515 378838 239527
rect 363290 239487 378838 239515
rect 363290 239475 363296 239487
rect 378832 239475 378838 239487
rect 378890 239475 378896 239527
rect 383152 239475 383158 239527
rect 383210 239515 383216 239527
rect 473872 239515 473878 239527
rect 383210 239487 473878 239515
rect 383210 239475 383216 239487
rect 473872 239475 473878 239487
rect 473930 239475 473936 239527
rect 369280 239401 369286 239453
rect 369338 239441 369344 239453
rect 376144 239441 376150 239453
rect 369338 239413 376150 239441
rect 369338 239401 369344 239413
rect 376144 239401 376150 239413
rect 376202 239401 376208 239453
rect 394480 239401 394486 239453
rect 394538 239441 394544 239453
rect 496528 239441 496534 239453
rect 394538 239413 496534 239441
rect 394538 239401 394544 239413
rect 496528 239401 496534 239413
rect 496586 239401 496592 239453
rect 365008 239327 365014 239379
rect 365066 239367 365072 239379
rect 505648 239367 505654 239379
rect 365066 239339 505654 239367
rect 365066 239327 365072 239339
rect 505648 239327 505654 239339
rect 505706 239327 505712 239379
rect 372112 239253 372118 239305
rect 372170 239293 372176 239305
rect 523792 239293 523798 239305
rect 372170 239265 523798 239293
rect 372170 239253 372176 239265
rect 523792 239253 523798 239265
rect 523850 239253 523856 239305
rect 388528 239179 388534 239231
rect 388586 239219 388592 239231
rect 413392 239219 413398 239231
rect 388586 239191 413398 239219
rect 388586 239179 388592 239191
rect 413392 239179 413398 239191
rect 413450 239179 413456 239231
rect 420400 239179 420406 239231
rect 420458 239219 420464 239231
rect 596176 239219 596182 239231
rect 420458 239191 596182 239219
rect 420458 239179 420464 239191
rect 596176 239179 596182 239191
rect 596234 239179 596240 239231
rect 367216 239105 367222 239157
rect 367274 239145 367280 239157
rect 542608 239145 542614 239157
rect 367274 239117 542614 239145
rect 367274 239105 367280 239117
rect 542608 239105 542614 239117
rect 542666 239105 542672 239157
rect 149392 239031 149398 239083
rect 149450 239071 149456 239083
rect 174160 239071 174166 239083
rect 149450 239043 174166 239071
rect 149450 239031 149456 239043
rect 174160 239031 174166 239043
rect 174218 239031 174224 239083
rect 377584 239031 377590 239083
rect 377642 239071 377648 239083
rect 561712 239071 561718 239083
rect 377642 239043 561718 239071
rect 377642 239031 377648 239043
rect 561712 239031 561718 239043
rect 561770 239031 561776 239083
rect 323920 238957 323926 239009
rect 323978 238997 323984 239009
rect 455056 238997 455062 239009
rect 323978 238969 455062 238997
rect 323978 238957 323984 238969
rect 455056 238957 455062 238969
rect 455114 238957 455120 239009
rect 327664 238883 327670 238935
rect 327722 238923 327728 238935
rect 461872 238923 461878 238935
rect 327722 238895 461878 238923
rect 327722 238883 327728 238895
rect 461872 238883 461878 238895
rect 461930 238883 461936 238935
rect 326704 238809 326710 238861
rect 326762 238849 326768 238861
rect 462544 238849 462550 238861
rect 326762 238821 462550 238849
rect 326762 238809 326768 238821
rect 462544 238809 462550 238821
rect 462602 238809 462608 238861
rect 329872 238735 329878 238787
rect 329930 238775 329936 238787
rect 468592 238775 468598 238787
rect 329930 238747 468598 238775
rect 329930 238735 329936 238747
rect 468592 238735 468598 238747
rect 468650 238735 468656 238787
rect 332656 238661 332662 238713
rect 332714 238701 332720 238713
rect 474640 238701 474646 238713
rect 332714 238673 474646 238701
rect 332714 238661 332720 238673
rect 474640 238661 474646 238673
rect 474698 238661 474704 238713
rect 335728 238587 335734 238639
rect 335786 238627 335792 238639
rect 480688 238627 480694 238639
rect 335786 238599 480694 238627
rect 335786 238587 335792 238599
rect 480688 238587 480694 238599
rect 480746 238587 480752 238639
rect 338992 238513 338998 238565
rect 339050 238553 339056 238565
rect 486736 238553 486742 238565
rect 339050 238525 486742 238553
rect 339050 238513 339056 238525
rect 486736 238513 486742 238525
rect 486794 238513 486800 238565
rect 341776 238439 341782 238491
rect 341834 238479 341840 238491
rect 492784 238479 492790 238491
rect 341834 238451 492790 238479
rect 341834 238439 341840 238451
rect 492784 238439 492790 238451
rect 492842 238439 492848 238491
rect 345904 238365 345910 238417
rect 345962 238405 345968 238417
rect 498256 238405 498262 238417
rect 345962 238377 498262 238405
rect 345962 238365 345968 238377
rect 498256 238365 498262 238377
rect 498314 238365 498320 238417
rect 345328 238291 345334 238343
rect 345386 238331 345392 238343
rect 500272 238331 500278 238343
rect 345386 238303 500278 238331
rect 345386 238291 345392 238303
rect 500272 238291 500278 238303
rect 500330 238291 500336 238343
rect 348112 238217 348118 238269
rect 348170 238257 348176 238269
rect 504112 238257 504118 238269
rect 348170 238229 504118 238257
rect 348170 238217 348176 238229
rect 504112 238217 504118 238229
rect 504170 238217 504176 238269
rect 351184 238143 351190 238195
rect 351242 238183 351248 238195
rect 512368 238183 512374 238195
rect 351242 238155 512374 238183
rect 351242 238143 351248 238155
rect 512368 238143 512374 238155
rect 512426 238143 512432 238195
rect 354160 238069 354166 238121
rect 354218 238109 354224 238121
rect 518512 238109 518518 238121
rect 354218 238081 518518 238109
rect 354218 238069 354224 238081
rect 518512 238069 518518 238081
rect 518570 238069 518576 238121
rect 361360 237995 361366 238047
rect 361418 238035 361424 238047
rect 532048 238035 532054 238047
rect 361418 238007 532054 238035
rect 361418 237995 361424 238007
rect 532048 237995 532054 238007
rect 532106 237995 532112 238047
rect 363088 237921 363094 237973
rect 363146 237961 363152 237973
rect 535120 237961 535126 237973
rect 363146 237933 535126 237961
rect 363146 237921 363152 237933
rect 535120 237921 535126 237933
rect 535178 237921 535184 237973
rect 360304 237847 360310 237899
rect 360362 237887 360368 237899
rect 530512 237887 530518 237899
rect 360362 237859 530518 237887
rect 360362 237847 360368 237859
rect 530512 237847 530518 237859
rect 530570 237847 530576 237899
rect 364432 237773 364438 237825
rect 364490 237813 364496 237825
rect 538000 237813 538006 237825
rect 364490 237785 538006 237813
rect 364490 237773 364496 237785
rect 538000 237773 538006 237785
rect 538058 237773 538064 237825
rect 365872 237699 365878 237751
rect 365930 237739 365936 237751
rect 538576 237739 538582 237751
rect 365930 237711 538582 237739
rect 365930 237699 365936 237711
rect 538576 237699 538582 237711
rect 538634 237699 538640 237751
rect 367600 237625 367606 237677
rect 367658 237665 367664 237677
rect 541552 237665 541558 237677
rect 367658 237637 541558 237665
rect 367658 237625 367664 237637
rect 541552 237625 541558 237637
rect 541610 237625 541616 237677
rect 370384 237551 370390 237603
rect 370442 237591 370448 237603
rect 550864 237591 550870 237603
rect 370442 237563 550870 237591
rect 370442 237551 370448 237563
rect 550864 237551 550870 237563
rect 550922 237551 550928 237603
rect 323152 237477 323158 237529
rect 323210 237517 323216 237529
rect 452752 237517 452758 237529
rect 323210 237489 452758 237517
rect 323210 237477 323216 237489
rect 452752 237477 452758 237489
rect 452810 237477 452816 237529
rect 320848 237403 320854 237455
rect 320906 237443 320912 237455
rect 450448 237443 450454 237455
rect 320906 237415 450454 237443
rect 320906 237403 320912 237415
rect 450448 237403 450454 237415
rect 450506 237403 450512 237455
rect 317584 237329 317590 237381
rect 317642 237369 317648 237381
rect 444496 237369 444502 237381
rect 317642 237341 444502 237369
rect 317642 237329 317648 237341
rect 444496 237329 444502 237341
rect 444554 237329 444560 237381
rect 314800 237255 314806 237307
rect 314858 237295 314864 237307
rect 438352 237295 438358 237307
rect 314858 237267 438358 237295
rect 314858 237255 314864 237267
rect 438352 237255 438358 237267
rect 438410 237255 438416 237307
rect 313840 237181 313846 237233
rect 313898 237221 313904 237233
rect 434608 237221 434614 237233
rect 313898 237193 434614 237221
rect 313898 237181 313904 237193
rect 434608 237181 434614 237193
rect 434666 237181 434672 237233
rect 310768 237107 310774 237159
rect 310826 237147 310832 237159
rect 428656 237147 428662 237159
rect 310826 237119 428662 237147
rect 310826 237107 310832 237119
rect 428656 237107 428662 237119
rect 428714 237107 428720 237159
rect 307024 237033 307030 237085
rect 307082 237073 307088 237085
rect 423280 237073 423286 237085
rect 307082 237045 423286 237073
rect 307082 237033 307088 237045
rect 423280 237033 423286 237045
rect 423338 237033 423344 237085
rect 304816 236959 304822 237011
rect 304874 236999 304880 237011
rect 304874 236971 410654 236999
rect 304874 236959 304880 236971
rect 301744 236885 301750 236937
rect 301802 236925 301808 236937
rect 409648 236925 409654 236937
rect 301802 236897 409654 236925
rect 301802 236885 301808 236897
rect 409648 236885 409654 236897
rect 409706 236885 409712 236937
rect 286192 236811 286198 236863
rect 286250 236851 286256 236863
rect 381040 236851 381046 236863
rect 286250 236823 381046 236851
rect 286250 236811 286256 236823
rect 381040 236811 381046 236823
rect 381098 236811 381104 236863
rect 410626 236851 410654 236971
rect 411568 236959 411574 237011
rect 411626 236999 411632 237011
rect 413968 236999 413974 237011
rect 411626 236971 413974 236999
rect 411626 236959 411632 236971
rect 413968 236959 413974 236971
rect 414026 236959 414032 237011
rect 410704 236885 410710 236937
rect 410762 236925 410768 236937
rect 413680 236925 413686 236937
rect 410762 236897 413686 236925
rect 410762 236885 410768 236897
rect 413680 236885 413686 236897
rect 413738 236885 413744 236937
rect 416464 236851 416470 236863
rect 410626 236823 416470 236851
rect 416464 236811 416470 236823
rect 416522 236811 416528 236863
rect 281584 236737 281590 236789
rect 281642 236777 281648 236789
rect 372400 236777 372406 236789
rect 281642 236749 372406 236777
rect 281642 236737 281648 236749
rect 372400 236737 372406 236749
rect 372458 236737 372464 236789
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 42736 236703 42742 236715
rect 42218 236675 42742 236703
rect 42218 236663 42224 236675
rect 42736 236663 42742 236675
rect 42794 236663 42800 236715
rect 278416 236663 278422 236715
rect 278474 236703 278480 236715
rect 366736 236703 366742 236715
rect 278474 236675 366742 236703
rect 278474 236663 278480 236675
rect 366736 236663 366742 236675
rect 366794 236663 366800 236715
rect 388816 236663 388822 236715
rect 388874 236703 388880 236715
rect 390352 236703 390358 236715
rect 388874 236675 390358 236703
rect 388874 236663 388880 236675
rect 390352 236663 390358 236675
rect 390410 236663 390416 236715
rect 279856 236589 279862 236641
rect 279914 236629 279920 236641
rect 368944 236629 368950 236641
rect 279914 236601 368950 236629
rect 279914 236589 279920 236601
rect 368944 236589 368950 236601
rect 369002 236589 369008 236641
rect 388624 236589 388630 236641
rect 388682 236629 388688 236641
rect 389008 236629 389014 236641
rect 388682 236601 389014 236629
rect 388682 236589 388688 236601
rect 389008 236589 389014 236601
rect 389066 236589 389072 236641
rect 390352 236515 390358 236567
rect 390410 236555 390416 236567
rect 476944 236555 476950 236567
rect 390410 236527 476950 236555
rect 390410 236515 390416 236527
rect 476944 236515 476950 236527
rect 477002 236515 477008 236567
rect 42832 236441 42838 236493
rect 42890 236481 42896 236493
rect 43120 236481 43126 236493
rect 42890 236453 43126 236481
rect 42890 236441 42896 236453
rect 43120 236441 43126 236453
rect 43178 236441 43184 236493
rect 397360 236441 397366 236493
rect 397418 236481 397424 236493
rect 483856 236481 483862 236493
rect 397418 236453 483862 236481
rect 397418 236441 397424 236453
rect 483856 236441 483862 236453
rect 483914 236441 483920 236493
rect 508624 236407 508630 236419
rect 398914 236379 508630 236407
rect 363568 236293 363574 236345
rect 363626 236333 363632 236345
rect 381424 236333 381430 236345
rect 363626 236305 381430 236333
rect 363626 236293 363632 236305
rect 381424 236293 381430 236305
rect 381482 236293 381488 236345
rect 346288 236145 346294 236197
rect 346346 236185 346352 236197
rect 361648 236185 361654 236197
rect 346346 236157 361654 236185
rect 346346 236145 346352 236157
rect 361648 236145 361654 236157
rect 361706 236145 361712 236197
rect 383824 236145 383830 236197
rect 383882 236185 383888 236197
rect 388720 236185 388726 236197
rect 383882 236157 388726 236185
rect 383882 236145 383888 236157
rect 388720 236145 388726 236157
rect 388778 236145 388784 236197
rect 231184 236071 231190 236123
rect 231242 236111 231248 236123
rect 253552 236111 253558 236123
rect 231242 236083 253558 236111
rect 231242 236071 231248 236083
rect 253552 236071 253558 236083
rect 253610 236071 253616 236123
rect 255280 236071 255286 236123
rect 255338 236111 255344 236123
rect 273712 236111 273718 236123
rect 255338 236083 273718 236111
rect 255338 236071 255344 236083
rect 273712 236071 273718 236083
rect 273770 236071 273776 236123
rect 285136 236071 285142 236123
rect 285194 236111 285200 236123
rect 326800 236111 326806 236123
rect 285194 236083 326806 236111
rect 285194 236071 285200 236083
rect 326800 236071 326806 236083
rect 326858 236071 326864 236123
rect 350416 236071 350422 236123
rect 350474 236111 350480 236123
rect 398914 236111 398942 236379
rect 508624 236367 508630 236379
rect 508682 236367 508688 236419
rect 403312 236293 403318 236345
rect 403370 236333 403376 236345
rect 520720 236333 520726 236345
rect 403370 236305 520726 236333
rect 403370 236293 403376 236305
rect 520720 236293 520726 236305
rect 520778 236293 520784 236345
rect 403216 236219 403222 236271
rect 403274 236259 403280 236271
rect 526672 236259 526678 236271
rect 403274 236231 526678 236259
rect 403274 236219 403280 236231
rect 526672 236219 526678 236231
rect 526730 236219 526736 236271
rect 411664 236145 411670 236197
rect 411722 236185 411728 236197
rect 544336 236185 544342 236197
rect 411722 236157 544342 236185
rect 411722 236145 411728 236157
rect 544336 236145 544342 236157
rect 544394 236145 544400 236197
rect 350474 236083 398942 236111
rect 350474 236071 350480 236083
rect 400240 236071 400246 236123
rect 400298 236111 400304 236123
rect 485584 236111 485590 236123
rect 400298 236083 485590 236111
rect 400298 236071 400304 236083
rect 485584 236071 485590 236083
rect 485642 236071 485648 236123
rect 250480 235997 250486 236049
rect 250538 236037 250544 236049
rect 272368 236037 272374 236049
rect 250538 236009 272374 236037
rect 250538 235997 250544 236009
rect 272368 235997 272374 236009
rect 272426 235997 272432 236049
rect 282160 235997 282166 236049
rect 282218 236037 282224 236049
rect 325360 236037 325366 236049
rect 282218 236009 325366 236037
rect 282218 235997 282224 236009
rect 325360 235997 325366 236009
rect 325418 235997 325424 236049
rect 333808 235997 333814 236049
rect 333866 236037 333872 236049
rect 466480 236037 466486 236049
rect 333866 236009 466486 236037
rect 333866 235997 333872 236009
rect 466480 235997 466486 236009
rect 466538 235997 466544 236049
rect 211216 235923 211222 235975
rect 211274 235963 211280 235975
rect 229264 235963 229270 235975
rect 211274 235935 229270 235963
rect 211274 235923 211280 235935
rect 229264 235923 229270 235935
rect 229322 235923 229328 235975
rect 241648 235923 241654 235975
rect 241706 235963 241712 235975
rect 266320 235963 266326 235975
rect 241706 235935 266326 235963
rect 241706 235923 241712 235935
rect 266320 235923 266326 235935
rect 266378 235923 266384 235975
rect 286672 235923 286678 235975
rect 286730 235963 286736 235975
rect 331120 235963 331126 235975
rect 286730 235935 331126 235963
rect 286730 235923 286736 235935
rect 331120 235923 331126 235935
rect 331178 235923 331184 235975
rect 339856 235923 339862 235975
rect 339914 235963 339920 235975
rect 475216 235963 475222 235975
rect 339914 235935 475222 235963
rect 339914 235923 339920 235935
rect 475216 235923 475222 235935
rect 475274 235923 475280 235975
rect 210640 235849 210646 235901
rect 210698 235889 210704 235901
rect 230032 235889 230038 235901
rect 210698 235861 230038 235889
rect 210698 235849 210704 235861
rect 230032 235849 230038 235861
rect 230090 235849 230096 235901
rect 244336 235849 244342 235901
rect 244394 235889 244400 235901
rect 268144 235889 268150 235901
rect 244394 235861 268150 235889
rect 244394 235849 244400 235861
rect 268144 235849 268150 235861
rect 268202 235849 268208 235901
rect 271984 235849 271990 235901
rect 272042 235889 272048 235901
rect 282352 235889 282358 235901
rect 272042 235861 282358 235889
rect 272042 235849 272048 235861
rect 282352 235849 282358 235861
rect 282410 235849 282416 235901
rect 287440 235849 287446 235901
rect 287498 235889 287504 235901
rect 341968 235889 341974 235901
rect 287498 235861 341974 235889
rect 287498 235849 287504 235861
rect 341968 235849 341974 235861
rect 342026 235849 342032 235901
rect 343120 235849 343126 235901
rect 343178 235889 343184 235901
rect 483760 235889 483766 235901
rect 343178 235861 483766 235889
rect 343178 235849 343184 235861
rect 483760 235849 483766 235861
rect 483818 235849 483824 235901
rect 212944 235775 212950 235827
rect 213002 235815 213008 235827
rect 232336 235815 232342 235827
rect 213002 235787 232342 235815
rect 213002 235775 213008 235787
rect 232336 235775 232342 235787
rect 232394 235775 232400 235827
rect 233488 235775 233494 235827
rect 233546 235815 233552 235827
rect 233546 235787 236174 235815
rect 233546 235775 233552 235787
rect 211984 235701 211990 235753
rect 212042 235741 212048 235753
rect 233008 235741 233014 235753
rect 212042 235713 233014 235741
rect 212042 235701 212048 235713
rect 233008 235701 233014 235713
rect 233066 235701 233072 235753
rect 211600 235627 211606 235679
rect 211658 235667 211664 235679
rect 230704 235667 230710 235679
rect 211658 235639 230710 235667
rect 211658 235627 211664 235639
rect 230704 235627 230710 235639
rect 230762 235627 230768 235679
rect 236146 235667 236174 235787
rect 238000 235775 238006 235827
rect 238058 235815 238064 235827
rect 264688 235815 264694 235827
rect 238058 235787 264694 235815
rect 238058 235775 238064 235787
rect 264688 235775 264694 235787
rect 264746 235775 264752 235827
rect 265744 235775 265750 235827
rect 265802 235815 265808 235827
rect 290992 235815 290998 235827
rect 265802 235787 290998 235815
rect 265802 235775 265808 235787
rect 290992 235775 290998 235787
rect 291050 235775 291056 235827
rect 294448 235775 294454 235827
rect 294506 235815 294512 235827
rect 338512 235815 338518 235827
rect 294506 235787 338518 235815
rect 294506 235775 294512 235787
rect 338512 235775 338518 235787
rect 338570 235775 338576 235827
rect 339472 235775 339478 235827
rect 339530 235815 339536 235827
rect 397360 235815 397366 235827
rect 339530 235787 397366 235815
rect 339530 235775 339536 235787
rect 397360 235775 397366 235787
rect 397418 235775 397424 235827
rect 398224 235775 398230 235827
rect 398282 235815 398288 235827
rect 400240 235815 400246 235827
rect 398282 235787 400246 235815
rect 398282 235775 398288 235787
rect 400240 235775 400246 235787
rect 400298 235775 400304 235827
rect 400336 235775 400342 235827
rect 400394 235815 400400 235827
rect 559216 235815 559222 235827
rect 400394 235787 559222 235815
rect 400394 235775 400400 235787
rect 559216 235775 559222 235787
rect 559274 235775 559280 235827
rect 257968 235701 257974 235753
rect 258026 235741 258032 235753
rect 279184 235741 279190 235753
rect 258026 235713 279190 235741
rect 258026 235701 258032 235713
rect 279184 235701 279190 235713
rect 279242 235701 279248 235753
rect 283888 235701 283894 235753
rect 283946 235741 283952 235753
rect 325840 235741 325846 235753
rect 283946 235713 325846 235741
rect 283946 235701 283952 235713
rect 325840 235701 325846 235713
rect 325898 235701 325904 235753
rect 328912 235701 328918 235753
rect 328970 235741 328976 235753
rect 328970 235713 374462 235741
rect 328970 235701 328976 235713
rect 262000 235667 262006 235679
rect 236146 235639 262006 235667
rect 262000 235627 262006 235639
rect 262058 235627 262064 235679
rect 279280 235627 279286 235679
rect 279338 235667 279344 235679
rect 322480 235667 322486 235679
rect 279338 235639 322486 235667
rect 279338 235627 279344 235639
rect 322480 235627 322486 235639
rect 322538 235627 322544 235679
rect 348880 235627 348886 235679
rect 348938 235667 348944 235679
rect 365008 235667 365014 235679
rect 348938 235639 365014 235667
rect 348938 235627 348944 235639
rect 365008 235627 365014 235639
rect 365066 235627 365072 235679
rect 214192 235553 214198 235605
rect 214250 235593 214256 235605
rect 235312 235593 235318 235605
rect 214250 235565 235318 235593
rect 214250 235553 214256 235565
rect 235312 235553 235318 235565
rect 235370 235553 235376 235605
rect 249712 235553 249718 235605
rect 249770 235593 249776 235605
rect 293776 235593 293782 235605
rect 249770 235565 293782 235593
rect 249770 235553 249776 235565
rect 293776 235553 293782 235565
rect 293834 235553 293840 235605
rect 298000 235553 298006 235605
rect 298058 235593 298064 235605
rect 338320 235593 338326 235605
rect 298058 235565 338326 235593
rect 298058 235553 298064 235565
rect 338320 235553 338326 235565
rect 338378 235553 338384 235605
rect 358000 235553 358006 235605
rect 358058 235593 358064 235605
rect 372112 235593 372118 235605
rect 358058 235565 372118 235593
rect 358058 235553 358064 235565
rect 372112 235553 372118 235565
rect 372170 235553 372176 235605
rect 374434 235593 374462 235713
rect 378640 235701 378646 235753
rect 378698 235741 378704 235753
rect 398512 235741 398518 235753
rect 378698 235713 398518 235741
rect 378698 235701 378704 235713
rect 398512 235701 398518 235713
rect 398570 235701 398576 235753
rect 398608 235701 398614 235753
rect 398666 235741 398672 235753
rect 564304 235741 564310 235753
rect 398666 235713 564310 235741
rect 398666 235701 398672 235713
rect 564304 235701 564310 235713
rect 564362 235701 564368 235753
rect 374512 235627 374518 235679
rect 374570 235667 374576 235679
rect 410704 235667 410710 235679
rect 374570 235639 410710 235667
rect 374570 235627 374576 235639
rect 410704 235627 410710 235639
rect 410762 235627 410768 235679
rect 410800 235627 410806 235679
rect 410858 235667 410864 235679
rect 585232 235667 585238 235679
rect 410858 235639 585238 235667
rect 410858 235627 410864 235639
rect 585232 235627 585238 235639
rect 585290 235627 585296 235679
rect 383056 235593 383062 235605
rect 374434 235565 383062 235593
rect 383056 235553 383062 235565
rect 383114 235553 383120 235605
rect 411568 235593 411574 235605
rect 384322 235565 411574 235593
rect 211024 235479 211030 235531
rect 211082 235519 211088 235531
rect 231568 235519 231574 235531
rect 211082 235491 231574 235519
rect 211082 235479 211088 235491
rect 231568 235479 231574 235491
rect 231626 235479 231632 235531
rect 234256 235479 234262 235531
rect 234314 235519 234320 235531
rect 264880 235519 264886 235531
rect 234314 235491 264886 235519
rect 234314 235479 234320 235491
rect 264880 235479 264886 235491
rect 264938 235479 264944 235531
rect 273424 235479 273430 235531
rect 273482 235519 273488 235531
rect 336496 235519 336502 235531
rect 273482 235491 336502 235519
rect 273482 235479 273488 235491
rect 336496 235479 336502 235491
rect 336554 235479 336560 235531
rect 341200 235479 341206 235531
rect 341258 235519 341264 235531
rect 341258 235491 383102 235519
rect 341258 235479 341264 235491
rect 383074 235457 383102 235491
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 42928 235445 42934 235457
rect 42218 235417 42934 235445
rect 42218 235405 42224 235417
rect 42928 235405 42934 235417
rect 42986 235405 42992 235457
rect 220624 235405 220630 235457
rect 220682 235445 220688 235457
rect 235888 235445 235894 235457
rect 220682 235417 235894 235445
rect 220682 235405 220688 235417
rect 235888 235405 235894 235417
rect 235946 235405 235952 235457
rect 235984 235405 235990 235457
rect 236042 235445 236048 235457
rect 240688 235445 240694 235457
rect 236042 235417 240694 235445
rect 236042 235405 236048 235417
rect 240688 235405 240694 235417
rect 240746 235405 240752 235457
rect 245200 235405 245206 235457
rect 245258 235445 245264 235457
rect 278224 235445 278230 235457
rect 245258 235417 278230 235445
rect 245258 235405 245264 235417
rect 278224 235405 278230 235417
rect 278282 235405 278288 235457
rect 284752 235405 284758 235457
rect 284810 235445 284816 235457
rect 345616 235445 345622 235457
rect 284810 235417 345622 235445
rect 284810 235405 284816 235417
rect 345616 235405 345622 235417
rect 345674 235405 345680 235457
rect 347632 235405 347638 235457
rect 347690 235445 347696 235457
rect 378640 235445 378646 235457
rect 347690 235417 378646 235445
rect 347690 235405 347696 235417
rect 378640 235405 378646 235417
rect 378698 235405 378704 235457
rect 383056 235405 383062 235457
rect 383114 235405 383120 235457
rect 219376 235331 219382 235383
rect 219434 235371 219440 235383
rect 244528 235371 244534 235383
rect 219434 235343 244534 235371
rect 219434 235331 219440 235343
rect 244528 235331 244534 235343
rect 244586 235331 244592 235383
rect 251152 235331 251158 235383
rect 251210 235371 251216 235383
rect 299248 235371 299254 235383
rect 251210 235343 299254 235371
rect 251210 235331 251216 235343
rect 299248 235331 299254 235343
rect 299306 235331 299312 235383
rect 311536 235331 311542 235383
rect 311594 235371 311600 235383
rect 325264 235371 325270 235383
rect 311594 235343 325270 235371
rect 311594 235331 311600 235343
rect 325264 235331 325270 235343
rect 325322 235331 325328 235383
rect 332176 235331 332182 235383
rect 332234 235371 332240 235383
rect 372880 235371 372886 235383
rect 332234 235343 372886 235371
rect 332234 235331 332240 235343
rect 372880 235331 372886 235343
rect 372938 235331 372944 235383
rect 373072 235331 373078 235383
rect 373130 235371 373136 235383
rect 384322 235371 384350 235565
rect 411568 235553 411574 235565
rect 411626 235553 411632 235605
rect 397648 235479 397654 235531
rect 397706 235519 397712 235531
rect 400240 235519 400246 235531
rect 397706 235491 400246 235519
rect 397706 235479 397712 235491
rect 400240 235479 400246 235491
rect 400298 235479 400304 235531
rect 401776 235479 401782 235531
rect 401834 235519 401840 235531
rect 410608 235519 410614 235531
rect 401834 235491 410614 235519
rect 401834 235479 401840 235491
rect 410608 235479 410614 235491
rect 410666 235479 410672 235531
rect 411760 235479 411766 235531
rect 411818 235519 411824 235531
rect 587440 235519 587446 235531
rect 411818 235491 587446 235519
rect 411818 235479 411824 235491
rect 587440 235479 587446 235491
rect 587498 235479 587504 235531
rect 409168 235405 409174 235457
rect 409226 235445 409232 235457
rect 588880 235445 588886 235457
rect 409226 235417 588886 235445
rect 409226 235405 409232 235417
rect 588880 235405 588886 235417
rect 588938 235405 588944 235457
rect 373130 235343 384350 235371
rect 373130 235331 373136 235343
rect 384400 235331 384406 235383
rect 384458 235371 384464 235383
rect 398800 235371 398806 235383
rect 384458 235343 398806 235371
rect 384458 235331 384464 235343
rect 398800 235331 398806 235343
rect 398858 235331 398864 235383
rect 403600 235331 403606 235383
rect 403658 235371 403664 235383
rect 585136 235371 585142 235383
rect 403658 235343 585142 235371
rect 403658 235331 403664 235343
rect 585136 235331 585142 235343
rect 585194 235331 585200 235383
rect 210064 235257 210070 235309
rect 210122 235297 210128 235309
rect 227824 235297 227830 235309
rect 210122 235269 227830 235297
rect 210122 235257 210128 235269
rect 227824 235257 227830 235269
rect 227882 235257 227888 235309
rect 228400 235257 228406 235309
rect 228458 235297 228464 235309
rect 264016 235297 264022 235309
rect 228458 235269 264022 235297
rect 228458 235257 228464 235269
rect 264016 235257 264022 235269
rect 264074 235257 264080 235309
rect 267472 235257 267478 235309
rect 267530 235297 267536 235309
rect 328336 235297 328342 235309
rect 267530 235269 328342 235297
rect 267530 235257 267536 235269
rect 328336 235257 328342 235269
rect 328394 235257 328400 235309
rect 330448 235257 330454 235309
rect 330506 235297 330512 235309
rect 392848 235297 392854 235309
rect 330506 235269 392854 235297
rect 330506 235257 330512 235269
rect 392848 235257 392854 235269
rect 392906 235257 392912 235309
rect 396304 235257 396310 235309
rect 396362 235297 396368 235309
rect 587344 235297 587350 235309
rect 396362 235269 587350 235297
rect 396362 235257 396368 235269
rect 587344 235257 587350 235269
rect 587402 235257 587408 235309
rect 213424 235183 213430 235235
rect 213482 235223 213488 235235
rect 213482 235195 232862 235223
rect 213482 235183 213488 235195
rect 209296 235109 209302 235161
rect 209354 235149 209360 235161
rect 228496 235149 228502 235161
rect 209354 235121 228502 235149
rect 209354 235109 209360 235121
rect 228496 235109 228502 235121
rect 228554 235109 228560 235161
rect 208912 235035 208918 235087
rect 208970 235075 208976 235087
rect 226960 235075 226966 235087
rect 208970 235047 226966 235075
rect 208970 235035 208976 235047
rect 226960 235035 226966 235047
rect 227018 235035 227024 235087
rect 232834 235075 232862 235195
rect 235696 235183 235702 235235
rect 235754 235223 235760 235235
rect 271120 235223 271126 235235
rect 235754 235195 271126 235223
rect 235754 235183 235760 235195
rect 271120 235183 271126 235195
rect 271178 235183 271184 235235
rect 275248 235183 275254 235235
rect 275306 235223 275312 235235
rect 291088 235223 291094 235235
rect 275306 235195 291094 235223
rect 275306 235183 275312 235195
rect 291088 235183 291094 235195
rect 291146 235183 291152 235235
rect 293488 235183 293494 235235
rect 293546 235223 293552 235235
rect 359920 235223 359926 235235
rect 293546 235195 359926 235223
rect 293546 235183 293552 235195
rect 359920 235183 359926 235195
rect 359978 235183 359984 235235
rect 390832 235183 390838 235235
rect 390890 235223 390896 235235
rect 590128 235223 590134 235235
rect 390890 235195 590134 235223
rect 390890 235183 390896 235195
rect 590128 235183 590134 235195
rect 590186 235183 590192 235235
rect 232912 235109 232918 235161
rect 232970 235149 232976 235161
rect 259024 235149 259030 235161
rect 232970 235121 259030 235149
rect 232970 235109 232976 235121
rect 259024 235109 259030 235121
rect 259082 235109 259088 235161
rect 290704 235109 290710 235161
rect 290762 235149 290768 235161
rect 354352 235149 354358 235161
rect 290762 235121 354358 235149
rect 290762 235109 290768 235121
rect 354352 235109 354358 235121
rect 354410 235109 354416 235161
rect 389776 235109 389782 235161
rect 389834 235149 389840 235161
rect 587920 235149 587926 235161
rect 389834 235121 587926 235149
rect 389834 235109 389840 235121
rect 587920 235109 587926 235121
rect 587978 235109 587984 235161
rect 235792 235075 235798 235087
rect 232834 235047 235798 235075
rect 235792 235035 235798 235047
rect 235850 235035 235856 235087
rect 235888 235035 235894 235087
rect 235946 235075 235952 235087
rect 245008 235075 245014 235087
rect 235946 235047 245014 235075
rect 235946 235035 235952 235047
rect 245008 235035 245014 235047
rect 245066 235035 245072 235087
rect 246640 235035 246646 235087
rect 246698 235075 246704 235087
rect 290896 235075 290902 235087
rect 246698 235047 290902 235075
rect 246698 235035 246704 235047
rect 290896 235035 290902 235047
rect 290954 235035 290960 235087
rect 296080 235035 296086 235087
rect 296138 235075 296144 235087
rect 362704 235075 362710 235087
rect 296138 235047 362710 235075
rect 296138 235035 296144 235047
rect 362704 235035 362710 235047
rect 362762 235035 362768 235087
rect 372880 235035 372886 235087
rect 372938 235075 372944 235087
rect 392080 235075 392086 235087
rect 372938 235047 392086 235075
rect 372938 235035 372944 235047
rect 392080 235035 392086 235047
rect 392138 235035 392144 235087
rect 392272 235035 392278 235087
rect 392330 235075 392336 235087
rect 593104 235075 593110 235087
rect 392330 235047 593110 235075
rect 392330 235035 392336 235047
rect 593104 235035 593110 235047
rect 593162 235035 593168 235087
rect 225136 234961 225142 235013
rect 225194 235001 225200 235013
rect 250576 235001 250582 235013
rect 225194 234973 250582 235001
rect 225194 234961 225200 234973
rect 250576 234961 250582 234973
rect 250634 234961 250640 235013
rect 254224 234961 254230 235013
rect 254282 235001 254288 235013
rect 305104 235001 305110 235013
rect 254282 234973 305110 235001
rect 254282 234961 254288 234973
rect 305104 234961 305110 234973
rect 305162 234961 305168 235013
rect 318352 234961 318358 235013
rect 318410 235001 318416 235013
rect 393904 235001 393910 235013
rect 318410 234973 393910 235001
rect 318410 234961 318416 234973
rect 393904 234961 393910 234973
rect 393962 234961 393968 235013
rect 396688 234961 396694 235013
rect 396746 235001 396752 235013
rect 408304 235001 408310 235013
rect 396746 234973 408310 235001
rect 396746 234961 396752 234973
rect 408304 234961 408310 234973
rect 408362 234961 408368 235013
rect 410416 234961 410422 235013
rect 410474 235001 410480 235013
rect 609040 235001 609046 235013
rect 410474 234973 609046 235001
rect 410474 234961 410480 234973
rect 609040 234961 609046 234973
rect 609098 234961 609104 235013
rect 204400 234887 204406 234939
rect 204458 234927 204464 234939
rect 217936 234927 217942 234939
rect 204458 234899 217942 234927
rect 204458 234887 204464 234899
rect 217936 234887 217942 234899
rect 217994 234887 218000 234939
rect 225520 234887 225526 234939
rect 225578 234927 225584 234939
rect 260176 234927 260182 234939
rect 225578 234899 260182 234927
rect 225578 234887 225584 234899
rect 260176 234887 260182 234899
rect 260234 234887 260240 234939
rect 261904 234887 261910 234939
rect 261962 234927 261968 234939
rect 311056 234927 311062 234939
rect 261962 234899 311062 234927
rect 261962 234887 261968 234899
rect 311056 234887 311062 234899
rect 311114 234887 311120 234939
rect 313072 234887 313078 234939
rect 313130 234927 313136 234939
rect 323440 234927 323446 234939
rect 313130 234899 323446 234927
rect 313130 234887 313136 234899
rect 323440 234887 323446 234899
rect 323498 234887 323504 234939
rect 324400 234887 324406 234939
rect 324458 234927 324464 234939
rect 391408 234927 391414 234939
rect 324458 234899 391414 234927
rect 324458 234887 324464 234899
rect 391408 234887 391414 234899
rect 391466 234887 391472 234939
rect 393040 234887 393046 234939
rect 393098 234927 393104 234939
rect 594640 234927 594646 234939
rect 393098 234899 594646 234927
rect 393098 234887 393104 234899
rect 594640 234887 594646 234899
rect 594698 234887 594704 234939
rect 42160 234813 42166 234865
rect 42218 234853 42224 234865
rect 42832 234853 42838 234865
rect 42218 234825 42838 234853
rect 42218 234813 42224 234825
rect 42832 234813 42838 234825
rect 42890 234813 42896 234865
rect 203248 234813 203254 234865
rect 203306 234853 203312 234865
rect 216496 234853 216502 234865
rect 203306 234825 216502 234853
rect 203306 234813 203312 234825
rect 216496 234813 216502 234825
rect 216554 234813 216560 234865
rect 222352 234813 222358 234865
rect 222410 234853 222416 234865
rect 250480 234853 250486 234865
rect 222410 234825 250486 234853
rect 222410 234813 222416 234825
rect 250480 234813 250486 234825
rect 250538 234813 250544 234865
rect 258736 234813 258742 234865
rect 258794 234853 258800 234865
rect 308176 234853 308182 234865
rect 258794 234825 308182 234853
rect 258794 234813 258800 234825
rect 308176 234813 308182 234825
rect 308234 234813 308240 234865
rect 317104 234813 317110 234865
rect 317162 234853 317168 234865
rect 391504 234853 391510 234865
rect 317162 234825 391510 234853
rect 317162 234813 317168 234825
rect 391504 234813 391510 234825
rect 391562 234813 391568 234865
rect 392656 234813 392662 234865
rect 392714 234853 392720 234865
rect 593968 234853 593974 234865
rect 392714 234825 593974 234853
rect 392714 234813 392720 234825
rect 593968 234813 593974 234825
rect 594026 234813 594032 234865
rect 206992 234739 206998 234791
rect 207050 234779 207056 234791
rect 221776 234779 221782 234791
rect 207050 234751 221782 234779
rect 207050 234739 207056 234751
rect 221776 234739 221782 234751
rect 221834 234739 221840 234791
rect 223888 234739 223894 234791
rect 223946 234779 223952 234791
rect 250768 234779 250774 234791
rect 223946 234751 250774 234779
rect 223946 234739 223952 234751
rect 250768 234739 250774 234751
rect 250826 234739 250832 234791
rect 255760 234739 255766 234791
rect 255818 234779 255824 234791
rect 305776 234779 305782 234791
rect 255818 234751 305782 234779
rect 255818 234739 255824 234751
rect 305776 234739 305782 234751
rect 305834 234739 305840 234791
rect 309328 234739 309334 234791
rect 309386 234779 309392 234791
rect 394192 234779 394198 234791
rect 309386 234751 394198 234779
rect 309386 234739 309392 234751
rect 394192 234739 394198 234751
rect 394250 234739 394256 234791
rect 394384 234739 394390 234791
rect 394442 234779 394448 234791
rect 596944 234779 596950 234791
rect 394442 234751 596950 234779
rect 394442 234739 394448 234751
rect 596944 234739 596950 234751
rect 597002 234739 597008 234791
rect 206512 234665 206518 234717
rect 206570 234705 206576 234717
rect 222448 234705 222454 234717
rect 206570 234677 222454 234705
rect 206570 234665 206576 234677
rect 222448 234665 222454 234677
rect 222506 234665 222512 234717
rect 227056 234665 227062 234717
rect 227114 234705 227120 234717
rect 263248 234705 263254 234717
rect 227114 234677 263254 234705
rect 227114 234665 227120 234677
rect 263248 234665 263254 234677
rect 263306 234665 263312 234717
rect 264400 234665 264406 234717
rect 264458 234705 264464 234717
rect 319600 234705 319606 234717
rect 264458 234677 319606 234705
rect 264458 234665 264464 234677
rect 319600 234665 319606 234677
rect 319658 234665 319664 234717
rect 319888 234665 319894 234717
rect 319946 234705 319952 234717
rect 403408 234705 403414 234717
rect 319946 234677 403414 234705
rect 319946 234665 319952 234677
rect 403408 234665 403414 234677
rect 403466 234665 403472 234717
rect 407728 234665 407734 234717
rect 407786 234705 407792 234717
rect 624112 234705 624118 234717
rect 407786 234677 624118 234705
rect 407786 234665 407792 234677
rect 624112 234665 624118 234677
rect 624170 234665 624176 234717
rect 204784 234591 204790 234643
rect 204842 234631 204848 234643
rect 207280 234631 207286 234643
rect 204842 234603 207286 234631
rect 204842 234591 204848 234603
rect 207280 234591 207286 234603
rect 207338 234591 207344 234643
rect 207856 234591 207862 234643
rect 207914 234631 207920 234643
rect 225520 234631 225526 234643
rect 207914 234603 225526 234631
rect 207914 234591 207920 234603
rect 225520 234591 225526 234603
rect 225578 234591 225584 234643
rect 235984 234631 235990 234643
rect 228706 234603 235990 234631
rect 202864 234517 202870 234569
rect 202922 234557 202928 234569
rect 214864 234557 214870 234569
rect 202922 234529 214870 234557
rect 202922 234517 202928 234529
rect 214864 234517 214870 234529
rect 214922 234517 214928 234569
rect 217840 234517 217846 234569
rect 217898 234557 217904 234569
rect 228706 234557 228734 234603
rect 235984 234591 235990 234603
rect 236042 234591 236048 234643
rect 246544 234591 246550 234643
rect 246602 234631 246608 234643
rect 267952 234631 267958 234643
rect 246602 234603 267958 234631
rect 246602 234591 246608 234603
rect 267952 234591 267958 234603
rect 268010 234591 268016 234643
rect 277552 234591 277558 234643
rect 277610 234631 277616 234643
rect 318160 234631 318166 234643
rect 277610 234603 318166 234631
rect 277610 234591 277616 234603
rect 318160 234591 318166 234603
rect 318218 234591 318224 234643
rect 326224 234591 326230 234643
rect 326282 234631 326288 234643
rect 449296 234631 449302 234643
rect 326282 234603 449302 234631
rect 326282 234591 326288 234603
rect 449296 234591 449302 234603
rect 449354 234591 449360 234643
rect 217898 234529 228734 234557
rect 217898 234517 217904 234529
rect 228784 234517 228790 234569
rect 228842 234557 228848 234569
rect 266224 234557 266230 234569
rect 228842 234529 266230 234557
rect 228842 234517 228848 234529
rect 266224 234517 266230 234529
rect 266282 234517 266288 234569
rect 267088 234517 267094 234569
rect 267146 234557 267152 234569
rect 298192 234557 298198 234569
rect 267146 234529 298198 234557
rect 267146 234517 267152 234529
rect 298192 234517 298198 234529
rect 298250 234517 298256 234569
rect 303472 234517 303478 234569
rect 303530 234557 303536 234569
rect 354256 234557 354262 234569
rect 303530 234529 354262 234557
rect 303530 234517 303536 234529
rect 354256 234517 354262 234529
rect 354314 234517 354320 234569
rect 391216 234517 391222 234569
rect 391274 234557 391280 234569
rect 512656 234557 512662 234569
rect 391274 234529 512662 234557
rect 391274 234517 391280 234529
rect 512656 234517 512662 234529
rect 512714 234517 512720 234569
rect 202000 234443 202006 234495
rect 202058 234483 202064 234495
rect 213424 234483 213430 234495
rect 202058 234455 213430 234483
rect 202058 234443 202064 234455
rect 213424 234443 213430 234455
rect 213482 234443 213488 234495
rect 249328 234443 249334 234495
rect 249386 234483 249392 234495
rect 271024 234483 271030 234495
rect 249386 234455 271030 234483
rect 249386 234443 249392 234455
rect 271024 234443 271030 234455
rect 271082 234443 271088 234495
rect 280624 234443 280630 234495
rect 280682 234483 280688 234495
rect 322192 234483 322198 234495
rect 280682 234455 322198 234483
rect 280682 234443 280688 234455
rect 322192 234443 322198 234455
rect 322250 234443 322256 234495
rect 323536 234443 323542 234495
rect 323594 234483 323600 234495
rect 446320 234483 446326 234495
rect 323594 234455 446326 234483
rect 323594 234443 323600 234455
rect 446320 234443 446326 234455
rect 446378 234443 446384 234495
rect 149392 234369 149398 234421
rect 149450 234409 149456 234421
rect 159856 234409 159862 234421
rect 149450 234381 159862 234409
rect 149450 234369 149456 234381
rect 159856 234369 159862 234381
rect 159914 234369 159920 234421
rect 206128 234369 206134 234421
rect 206186 234409 206192 234421
rect 220912 234409 220918 234421
rect 206186 234381 220918 234409
rect 206186 234369 206192 234381
rect 220912 234369 220918 234381
rect 220970 234369 220976 234421
rect 252592 234369 252598 234421
rect 252650 234409 252656 234421
rect 273616 234409 273622 234421
rect 252650 234381 273622 234409
rect 252650 234369 252656 234381
rect 273616 234369 273622 234381
rect 273674 234369 273680 234421
rect 276112 234369 276118 234421
rect 276170 234409 276176 234421
rect 313936 234409 313942 234421
rect 276170 234381 313942 234409
rect 276170 234369 276176 234381
rect 313936 234369 313942 234381
rect 313994 234369 314000 234421
rect 320272 234369 320278 234421
rect 320330 234409 320336 234421
rect 443440 234409 443446 234421
rect 320330 234381 443446 234409
rect 320330 234369 320336 234381
rect 443440 234369 443446 234381
rect 443498 234369 443504 234421
rect 207376 234295 207382 234347
rect 207434 234335 207440 234347
rect 219376 234335 219382 234347
rect 207434 234307 219382 234335
rect 207434 234295 207440 234307
rect 219376 234295 219382 234307
rect 219434 234295 219440 234347
rect 247408 234295 247414 234347
rect 247466 234335 247472 234347
rect 269392 234335 269398 234347
rect 247466 234307 269398 234335
rect 247466 234295 247472 234307
rect 269392 234295 269398 234307
rect 269450 234295 269456 234347
rect 270256 234295 270262 234347
rect 270314 234335 270320 234347
rect 304336 234335 304342 234347
rect 270314 234307 304342 234335
rect 270314 234295 270320 234307
rect 304336 234295 304342 234307
rect 304394 234295 304400 234347
rect 314416 234295 314422 234347
rect 314474 234335 314480 234347
rect 436144 234335 436150 234347
rect 314474 234307 436150 234335
rect 314474 234295 314480 234307
rect 436144 234295 436150 234307
rect 436202 234295 436208 234347
rect 200272 234221 200278 234273
rect 200330 234261 200336 234273
rect 210352 234261 210358 234273
rect 200330 234233 210358 234261
rect 200330 234221 200336 234233
rect 210352 234221 210358 234233
rect 210410 234221 210416 234273
rect 253456 234221 253462 234273
rect 253514 234261 253520 234273
rect 270832 234261 270838 234273
rect 253514 234233 270838 234261
rect 253514 234221 253520 234233
rect 270832 234221 270838 234233
rect 270890 234221 270896 234273
rect 273040 234221 273046 234273
rect 273098 234261 273104 234273
rect 306640 234261 306646 234273
rect 273098 234233 306646 234261
rect 273098 234221 273104 234233
rect 306640 234221 306646 234233
rect 306698 234221 306704 234273
rect 317200 234221 317206 234273
rect 317258 234261 317264 234273
rect 434896 234261 434902 234273
rect 317258 234233 434902 234261
rect 317258 234221 317264 234233
rect 434896 234221 434902 234233
rect 434954 234221 434960 234273
rect 200176 234147 200182 234199
rect 200234 234187 200240 234199
rect 208816 234187 208822 234199
rect 200234 234159 208822 234187
rect 200234 234147 200240 234159
rect 208816 234147 208822 234159
rect 208874 234147 208880 234199
rect 209680 234147 209686 234199
rect 209738 234187 209744 234199
rect 226288 234187 226294 234199
rect 209738 234159 226294 234187
rect 209738 234147 209744 234159
rect 226288 234147 226294 234159
rect 226346 234147 226352 234199
rect 268528 234147 268534 234199
rect 268586 234187 268592 234199
rect 293968 234187 293974 234199
rect 268586 234159 293974 234187
rect 268586 234147 268592 234159
rect 293968 234147 293974 234159
rect 294026 234147 294032 234199
rect 295696 234147 295702 234199
rect 295754 234187 295760 234199
rect 303568 234187 303574 234199
rect 295754 234159 303574 234187
rect 295754 234147 295760 234159
rect 303568 234147 303574 234159
rect 303626 234147 303632 234199
rect 308464 234147 308470 234199
rect 308522 234187 308528 234199
rect 424048 234187 424054 234199
rect 308522 234159 424054 234187
rect 308522 234147 308528 234159
rect 424048 234147 424054 234159
rect 424106 234147 424112 234199
rect 198736 234073 198742 234125
rect 198794 234113 198800 234125
rect 207376 234113 207382 234125
rect 198794 234085 207382 234113
rect 198794 234073 198800 234085
rect 207376 234073 207382 234085
rect 207434 234073 207440 234125
rect 207472 234073 207478 234125
rect 207530 234113 207536 234125
rect 223984 234113 223990 234125
rect 207530 234085 223990 234113
rect 207530 234073 207536 234085
rect 223984 234073 223990 234085
rect 224042 234073 224048 234125
rect 264304 234073 264310 234125
rect 264362 234113 264368 234125
rect 289840 234113 289846 234125
rect 264362 234085 289846 234113
rect 264362 234073 264368 234085
rect 289840 234073 289846 234085
rect 289898 234073 289904 234125
rect 298960 234073 298966 234125
rect 299018 234113 299024 234125
rect 348496 234113 348502 234125
rect 299018 234085 348502 234113
rect 299018 234073 299024 234085
rect 348496 234073 348502 234085
rect 348554 234073 348560 234125
rect 352144 234073 352150 234125
rect 352202 234113 352208 234125
rect 400432 234113 400438 234125
rect 352202 234085 400438 234113
rect 352202 234073 352208 234085
rect 400432 234073 400438 234085
rect 400490 234073 400496 234125
rect 403504 234073 403510 234125
rect 403562 234113 403568 234125
rect 509776 234113 509782 234125
rect 403562 234085 509782 234113
rect 403562 234073 403568 234085
rect 509776 234073 509782 234085
rect 509834 234073 509840 234125
rect 42064 233999 42070 234051
rect 42122 234039 42128 234051
rect 43024 234039 43030 234051
rect 42122 234011 43030 234039
rect 42122 233999 42128 234011
rect 43024 233999 43030 234011
rect 43082 233999 43088 234051
rect 198352 233999 198358 234051
rect 198410 234039 198416 234051
rect 205936 234039 205942 234051
rect 198410 234011 205942 234039
rect 198410 233999 198416 234011
rect 205936 233999 205942 234011
rect 205994 233999 206000 234051
rect 206896 233999 206902 234051
rect 206954 234039 206960 234051
rect 220240 234039 220246 234051
rect 206954 234011 220246 234039
rect 206954 233999 206960 234011
rect 220240 233999 220246 234011
rect 220298 233999 220304 234051
rect 261232 233999 261238 234051
rect 261290 234039 261296 234051
rect 279664 234039 279670 234051
rect 261290 234011 279670 234039
rect 261290 233999 261296 234011
rect 279664 233999 279670 234011
rect 279722 233999 279728 234051
rect 281200 233999 281206 234051
rect 281258 234039 281264 234051
rect 300784 234039 300790 234051
rect 281258 234011 300790 234039
rect 281258 233999 281264 234011
rect 300784 233999 300790 234011
rect 300842 233999 300848 234051
rect 311152 233999 311158 234051
rect 311210 234039 311216 234051
rect 420400 234039 420406 234051
rect 311210 234011 420406 234039
rect 311210 233999 311216 234011
rect 420400 233999 420406 234011
rect 420458 233999 420464 234051
rect 197488 233925 197494 233977
rect 197546 233965 197552 233977
rect 204304 233965 204310 233977
rect 197546 233937 204310 233965
rect 197546 233925 197552 233937
rect 204304 233925 204310 233937
rect 204362 233925 204368 233977
rect 205168 233925 205174 233977
rect 205226 233965 205232 233977
rect 207280 233965 207286 233977
rect 205226 233937 207286 233965
rect 205226 233925 205232 233937
rect 207280 233925 207286 233937
rect 207338 233925 207344 233977
rect 208720 233925 208726 233977
rect 208778 233965 208784 233977
rect 224752 233965 224758 233977
rect 208778 233937 224758 233965
rect 208778 233925 208784 233937
rect 224752 233925 224758 233937
rect 224810 233925 224816 233977
rect 258352 233925 258358 233977
rect 258410 233965 258416 233977
rect 278128 233965 278134 233977
rect 258410 233937 278134 233965
rect 258410 233925 258416 233937
rect 278128 233925 278134 233937
rect 278186 233925 278192 233977
rect 287056 233925 287062 233977
rect 287114 233965 287120 233977
rect 321136 233965 321142 233977
rect 287114 233937 321142 233965
rect 287114 233925 287120 233937
rect 321136 233925 321142 233937
rect 321194 233925 321200 233977
rect 326128 233925 326134 233977
rect 326186 233965 326192 233977
rect 374608 233965 374614 233977
rect 326186 233937 374614 233965
rect 326186 233925 326192 233937
rect 374608 233925 374614 233937
rect 374666 233925 374672 233977
rect 387184 233965 387190 233977
rect 377890 233937 387190 233965
rect 199120 233851 199126 233903
rect 199178 233891 199184 233903
rect 205072 233891 205078 233903
rect 199178 233863 205078 233891
rect 199178 233851 199184 233863
rect 205072 233851 205078 233863
rect 205130 233851 205136 233903
rect 205552 233851 205558 233903
rect 205610 233891 205616 233903
rect 218704 233891 218710 233903
rect 205610 233863 218710 233891
rect 205610 233851 205616 233863
rect 218704 233851 218710 233863
rect 218762 233851 218768 233903
rect 299344 233851 299350 233903
rect 299402 233891 299408 233903
rect 344656 233891 344662 233903
rect 299402 233863 344662 233891
rect 299402 233851 299408 233863
rect 344656 233851 344662 233863
rect 344714 233851 344720 233903
rect 354928 233851 354934 233903
rect 354986 233891 354992 233903
rect 377890 233891 377918 233937
rect 387184 233925 387190 233937
rect 387242 233925 387248 233977
rect 403312 233965 403318 233977
rect 388786 233937 403318 233965
rect 388786 233891 388814 233937
rect 403312 233925 403318 233937
rect 403370 233925 403376 233977
rect 492496 233965 492502 233977
rect 404770 233937 492502 233965
rect 354986 233863 377918 233891
rect 378706 233863 388814 233891
rect 354986 233851 354992 233863
rect 196912 233777 196918 233829
rect 196970 233817 196976 233829
rect 202864 233817 202870 233829
rect 196970 233789 202870 233817
rect 196970 233777 196976 233789
rect 202864 233777 202870 233789
rect 202922 233777 202928 233829
rect 204208 233777 204214 233829
rect 204266 233817 204272 233829
rect 215536 233817 215542 233829
rect 204266 233789 215542 233817
rect 204266 233777 204272 233789
rect 215536 233777 215542 233789
rect 215594 233777 215600 233829
rect 261616 233777 261622 233829
rect 261674 233817 261680 233829
rect 279280 233817 279286 233829
rect 261674 233789 279286 233817
rect 261674 233777 261680 233789
rect 279280 233777 279286 233789
rect 279338 233777 279344 233829
rect 292912 233777 292918 233829
rect 292970 233817 292976 233829
rect 325456 233817 325462 233829
rect 292970 233789 325462 233817
rect 292970 233777 292976 233789
rect 325456 233777 325462 233789
rect 325514 233777 325520 233829
rect 339856 233817 339862 233829
rect 325570 233789 339862 233817
rect 196528 233703 196534 233755
rect 196586 233743 196592 233755
rect 200560 233743 200566 233755
rect 196586 233715 200566 233743
rect 196586 233703 196592 233715
rect 200560 233703 200566 233715
rect 200618 233703 200624 233755
rect 201520 233703 201526 233755
rect 201578 233743 201584 233755
rect 211888 233743 211894 233755
rect 201578 233715 211894 233743
rect 201578 233703 201584 233715
rect 211888 233703 211894 233715
rect 211946 233703 211952 233755
rect 299824 233703 299830 233755
rect 299882 233743 299888 233755
rect 325570 233743 325598 233789
rect 339856 233777 339862 233789
rect 339914 233777 339920 233829
rect 356752 233777 356758 233829
rect 356810 233817 356816 233829
rect 378706 233817 378734 233863
rect 392080 233851 392086 233903
rect 392138 233891 392144 233903
rect 396976 233891 396982 233903
rect 392138 233863 396982 233891
rect 392138 233851 392144 233863
rect 396976 233851 396982 233863
rect 397034 233851 397040 233903
rect 401200 233851 401206 233903
rect 401258 233891 401264 233903
rect 404770 233891 404798 233937
rect 492496 233925 492502 233937
rect 492554 233925 492560 233977
rect 401258 233863 404798 233891
rect 401258 233851 401264 233863
rect 406192 233851 406198 233903
rect 406250 233891 406256 233903
rect 489616 233891 489622 233903
rect 406250 233863 489622 233891
rect 406250 233851 406256 233863
rect 489616 233851 489622 233863
rect 489674 233851 489680 233903
rect 356810 233789 378734 233817
rect 356810 233777 356816 233789
rect 385360 233777 385366 233829
rect 385418 233817 385424 233829
rect 385418 233789 409502 233817
rect 385418 233777 385424 233789
rect 299882 233715 325598 233743
rect 299882 233703 299888 233715
rect 334960 233703 334966 233755
rect 335018 233743 335024 233755
rect 390352 233743 390358 233755
rect 335018 233715 390358 233743
rect 335018 233703 335024 233715
rect 390352 233703 390358 233715
rect 390410 233703 390416 233755
rect 399472 233703 399478 233755
rect 399530 233743 399536 233755
rect 406192 233743 406198 233755
rect 399530 233715 406198 233743
rect 399530 233703 399536 233715
rect 406192 233703 406198 233715
rect 406250 233703 406256 233755
rect 409474 233743 409502 233789
rect 409552 233777 409558 233829
rect 409610 233817 409616 233829
rect 582544 233817 582550 233829
rect 409610 233789 582550 233817
rect 409610 233777 409616 233789
rect 582544 233777 582550 233789
rect 582602 233777 582608 233829
rect 455248 233743 455254 233755
rect 409474 233715 455254 233743
rect 455248 233703 455254 233715
rect 455306 233703 455312 233755
rect 195664 233629 195670 233681
rect 195722 233669 195728 233681
rect 201328 233669 201334 233681
rect 195722 233641 201334 233669
rect 195722 233629 195728 233641
rect 201328 233629 201334 233641
rect 201386 233629 201392 233681
rect 202480 233629 202486 233681
rect 202538 233669 202544 233681
rect 212560 233669 212566 233681
rect 202538 233641 212566 233669
rect 202538 233629 202544 233641
rect 212560 233629 212566 233641
rect 212618 233629 212624 233681
rect 305200 233629 305206 233681
rect 305258 233669 305264 233681
rect 305258 233641 338270 233669
rect 305258 233629 305264 233641
rect 192880 233555 192886 233607
rect 192938 233595 192944 233607
rect 195280 233595 195286 233607
rect 192938 233567 195286 233595
rect 192938 233555 192944 233567
rect 195280 233555 195286 233567
rect 195338 233555 195344 233607
rect 195568 233555 195574 233607
rect 195626 233595 195632 233607
rect 199792 233595 199798 233607
rect 195626 233567 199798 233595
rect 195626 233555 195632 233567
rect 199792 233555 199798 233567
rect 199850 233555 199856 233607
rect 201040 233555 201046 233607
rect 201098 233595 201104 233607
rect 209680 233595 209686 233607
rect 201098 233567 209686 233595
rect 201098 233555 201104 233567
rect 209680 233555 209686 233567
rect 209738 233555 209744 233607
rect 290320 233555 290326 233607
rect 290378 233595 290384 233607
rect 325168 233595 325174 233607
rect 290378 233567 325174 233595
rect 290378 233555 290384 233567
rect 325168 233555 325174 233567
rect 325226 233555 325232 233607
rect 325456 233555 325462 233607
rect 325514 233595 325520 233607
rect 336304 233595 336310 233607
rect 325514 233567 336310 233595
rect 325514 233555 325520 233567
rect 336304 233555 336310 233567
rect 336362 233555 336368 233607
rect 338242 233595 338270 233641
rect 338320 233629 338326 233681
rect 338378 233669 338384 233681
rect 358480 233669 358486 233681
rect 338378 233641 358486 233669
rect 338378 233629 338384 233641
rect 358480 233629 358486 233641
rect 358538 233629 358544 233681
rect 358576 233629 358582 233681
rect 358634 233669 358640 233681
rect 429136 233669 429142 233681
rect 358634 233641 429142 233669
rect 358634 233629 358640 233641
rect 429136 233629 429142 233641
rect 429194 233629 429200 233681
rect 342928 233595 342934 233607
rect 338242 233567 342934 233595
rect 342928 233555 342934 233567
rect 342986 233555 342992 233607
rect 343504 233555 343510 233607
rect 343562 233595 343568 233607
rect 348688 233595 348694 233607
rect 343562 233567 348694 233595
rect 343562 233555 343568 233567
rect 348688 233555 348694 233567
rect 348746 233555 348752 233607
rect 365680 233555 365686 233607
rect 365738 233595 365744 233607
rect 408976 233595 408982 233607
rect 365738 233567 408982 233595
rect 365738 233555 365744 233567
rect 408976 233555 408982 233567
rect 409034 233555 409040 233607
rect 194224 233481 194230 233533
rect 194282 233521 194288 233533
rect 198352 233521 198358 233533
rect 194282 233493 198358 233521
rect 194282 233481 194288 233493
rect 198352 233481 198358 233493
rect 198410 233481 198416 233533
rect 200656 233481 200662 233533
rect 200714 233521 200720 233533
rect 208144 233521 208150 233533
rect 200714 233493 208150 233521
rect 200714 233481 200720 233493
rect 208144 233481 208150 233493
rect 208202 233481 208208 233533
rect 208432 233481 208438 233533
rect 208490 233521 208496 233533
rect 223216 233521 223222 233533
rect 208490 233493 223222 233521
rect 208490 233481 208496 233493
rect 223216 233481 223222 233493
rect 223274 233481 223280 233533
rect 256528 233481 256534 233533
rect 256586 233521 256592 233533
rect 274672 233521 274678 233533
rect 256586 233493 274678 233521
rect 256586 233481 256592 233493
rect 274672 233481 274678 233493
rect 274730 233481 274736 233533
rect 304432 233481 304438 233533
rect 304490 233521 304496 233533
rect 334000 233521 334006 233533
rect 304490 233493 334006 233521
rect 304490 233481 304496 233493
rect 334000 233481 334006 233493
rect 334058 233481 334064 233533
rect 336688 233481 336694 233533
rect 336746 233521 336752 233533
rect 363952 233521 363958 233533
rect 336746 233493 363958 233521
rect 336746 233481 336752 233493
rect 363952 233481 363958 233493
rect 364010 233481 364016 233533
rect 364048 233481 364054 233533
rect 364106 233521 364112 233533
rect 406096 233521 406102 233533
rect 364106 233493 406102 233521
rect 364106 233481 364112 233493
rect 406096 233481 406102 233493
rect 406154 233481 406160 233533
rect 194608 233407 194614 233459
rect 194666 233447 194672 233459
rect 196048 233447 196054 233459
rect 194666 233419 196054 233447
rect 194666 233407 194672 233419
rect 196048 233407 196054 233419
rect 196106 233407 196112 233459
rect 196144 233407 196150 233459
rect 196202 233447 196208 233459
rect 199120 233447 199126 233459
rect 196202 233419 199126 233447
rect 196202 233407 196208 233419
rect 199120 233407 199126 233419
rect 199178 233407 199184 233459
rect 199696 233407 199702 233459
rect 199754 233447 199760 233459
rect 206608 233447 206614 233459
rect 199754 233419 206614 233447
rect 199754 233407 199760 233419
rect 206608 233407 206614 233419
rect 206666 233407 206672 233459
rect 207280 233407 207286 233459
rect 207338 233447 207344 233459
rect 217168 233447 217174 233459
rect 207338 233419 217174 233447
rect 207338 233407 207344 233419
rect 217168 233407 217174 233419
rect 217226 233407 217232 233459
rect 268912 233407 268918 233459
rect 268970 233447 268976 233459
rect 273424 233447 273430 233459
rect 268970 233419 273430 233447
rect 268970 233407 268976 233419
rect 273424 233407 273430 233419
rect 273482 233407 273488 233459
rect 277936 233407 277942 233459
rect 277994 233447 278000 233459
rect 294448 233447 294454 233459
rect 277994 233419 294454 233447
rect 277994 233407 278000 233419
rect 294448 233407 294454 233419
rect 294506 233407 294512 233459
rect 315760 233407 315766 233459
rect 315818 233447 315824 233459
rect 352816 233447 352822 233459
rect 315818 233419 352822 233447
rect 315818 233407 315824 233419
rect 352816 233407 352822 233419
rect 352874 233407 352880 233459
rect 361264 233407 361270 233459
rect 361322 233447 361328 233459
rect 400336 233447 400342 233459
rect 361322 233419 400342 233447
rect 361322 233407 361328 233419
rect 400336 233407 400342 233419
rect 400394 233407 400400 233459
rect 410032 233407 410038 233459
rect 410090 233447 410096 233459
rect 411664 233447 411670 233459
rect 410090 233419 411670 233447
rect 410090 233407 410096 233419
rect 411664 233407 411670 233419
rect 411722 233407 411728 233459
rect 192400 233333 192406 233385
rect 192458 233373 192464 233385
rect 193744 233373 193750 233385
rect 192458 233345 193750 233373
rect 192458 233333 192464 233345
rect 193744 233333 193750 233345
rect 193802 233333 193808 233385
rect 193840 233333 193846 233385
rect 193898 233373 193904 233385
rect 196816 233373 196822 233385
rect 193898 233345 196822 233373
rect 193898 233333 193904 233345
rect 196816 233333 196822 233345
rect 196874 233333 196880 233385
rect 197968 233333 197974 233385
rect 198026 233373 198032 233385
rect 203632 233373 203638 233385
rect 198026 233345 203638 233373
rect 198026 233333 198032 233345
rect 203632 233333 203638 233345
rect 203690 233333 203696 233385
rect 203920 233333 203926 233385
rect 203978 233373 203984 233385
rect 214192 233373 214198 233385
rect 203978 233345 214198 233373
rect 203978 233333 203984 233345
rect 214192 233333 214198 233345
rect 214250 233333 214256 233385
rect 262864 233333 262870 233385
rect 262922 233373 262928 233385
rect 281200 233373 281206 233385
rect 262922 233345 281206 233373
rect 262922 233333 262928 233345
rect 281200 233333 281206 233345
rect 281258 233333 281264 233385
rect 285712 233333 285718 233385
rect 285770 233373 285776 233385
rect 290704 233373 290710 233385
rect 285770 233345 290710 233373
rect 285770 233333 285776 233345
rect 290704 233333 290710 233345
rect 290762 233333 290768 233385
rect 291568 233333 291574 233385
rect 291626 233373 291632 233385
rect 291626 233345 296654 233373
rect 291626 233333 291632 233345
rect 193456 233259 193462 233311
rect 193514 233299 193520 233311
rect 194608 233299 194614 233311
rect 193514 233271 194614 233299
rect 193514 233259 193520 233271
rect 194608 233259 194614 233271
rect 194666 233259 194672 233311
rect 195184 233259 195190 233311
rect 195242 233299 195248 233311
rect 197488 233299 197494 233311
rect 195242 233271 197494 233299
rect 195242 233259 195248 233271
rect 197488 233259 197494 233271
rect 197546 233259 197552 233311
rect 197872 233259 197878 233311
rect 197930 233299 197936 233311
rect 202096 233299 202102 233311
rect 197930 233271 202102 233299
rect 197930 233259 197936 233271
rect 202096 233259 202102 233271
rect 202154 233259 202160 233311
rect 202384 233259 202390 233311
rect 202442 233299 202448 233311
rect 211120 233299 211126 233311
rect 202442 233271 211126 233299
rect 202442 233259 202448 233271
rect 211120 233259 211126 233271
rect 211178 233259 211184 233311
rect 266128 233259 266134 233311
rect 266186 233299 266192 233311
rect 280912 233299 280918 233311
rect 266186 233271 280918 233299
rect 266186 233259 266192 233271
rect 280912 233259 280918 233271
rect 280970 233259 280976 233311
rect 288496 233259 288502 233311
rect 288554 233299 288560 233311
rect 292816 233299 292822 233311
rect 288554 233271 292822 233299
rect 288554 233259 288560 233271
rect 292816 233259 292822 233271
rect 292874 233259 292880 233311
rect 296626 233299 296654 233345
rect 297232 233333 297238 233385
rect 297290 233373 297296 233385
rect 312688 233373 312694 233385
rect 297290 233345 312694 233373
rect 297290 233333 297296 233345
rect 312688 233333 312694 233345
rect 312746 233333 312752 233385
rect 321712 233333 321718 233385
rect 321770 233373 321776 233385
rect 332080 233373 332086 233385
rect 321770 233345 332086 233373
rect 321770 233333 321776 233345
rect 332080 233333 332086 233345
rect 332138 233333 332144 233385
rect 333424 233333 333430 233385
rect 333482 233373 333488 233385
rect 383152 233373 383158 233385
rect 333482 233345 383158 233373
rect 333482 233333 333488 233345
rect 383152 233333 383158 233345
rect 383210 233333 383216 233385
rect 406288 233333 406294 233385
rect 406346 233373 406352 233385
rect 409168 233373 409174 233385
rect 406346 233345 409174 233373
rect 406346 233333 406352 233345
rect 409168 233333 409174 233345
rect 409226 233333 409232 233385
rect 409936 233333 409942 233385
rect 409994 233373 410000 233385
rect 411760 233373 411766 233385
rect 409994 233345 411766 233373
rect 409994 233333 410000 233345
rect 411760 233333 411766 233345
rect 411818 233333 411824 233385
rect 301552 233299 301558 233311
rect 296626 233271 301558 233299
rect 301552 233259 301558 233271
rect 301610 233259 301616 233311
rect 301648 233259 301654 233311
rect 301706 233299 301712 233311
rect 310192 233299 310198 233311
rect 301706 233271 310198 233299
rect 301706 233259 301712 233271
rect 310192 233259 310198 233271
rect 310250 233259 310256 233311
rect 325168 233259 325174 233311
rect 325226 233299 325232 233311
rect 326896 233299 326902 233311
rect 325226 233271 326902 233299
rect 325226 233259 325232 233271
rect 326896 233259 326902 233271
rect 326954 233259 326960 233311
rect 329296 233259 329302 233311
rect 329354 233299 329360 233311
rect 460720 233299 460726 233311
rect 329354 233271 460726 233299
rect 329354 233259 329360 233271
rect 460720 233259 460726 233271
rect 460778 233259 460784 233311
rect 259120 233185 259126 233237
rect 259178 233225 259184 233237
rect 328144 233225 328150 233237
rect 259178 233197 328150 233225
rect 259178 233185 259184 233197
rect 328144 233185 328150 233197
rect 328202 233185 328208 233237
rect 331600 233185 331606 233237
rect 331658 233225 331664 233237
rect 343408 233225 343414 233237
rect 331658 233197 343414 233225
rect 331658 233185 331664 233197
rect 343408 233185 343414 233197
rect 343466 233185 343472 233237
rect 350320 233185 350326 233237
rect 350378 233225 350384 233237
rect 350378 233197 367166 233225
rect 350378 233185 350384 233197
rect 263536 233111 263542 233163
rect 263594 233151 263600 233163
rect 335728 233151 335734 233163
rect 263594 233123 335734 233151
rect 263594 233111 263600 233123
rect 335728 233111 335734 233123
rect 335786 233111 335792 233163
rect 337936 233111 337942 233163
rect 337994 233151 338000 233163
rect 355312 233151 355318 233163
rect 337994 233123 355318 233151
rect 337994 233111 338000 233123
rect 355312 233111 355318 233123
rect 355370 233111 355376 233163
rect 367138 233151 367166 233197
rect 367216 233185 367222 233237
rect 367274 233225 367280 233237
rect 497968 233225 497974 233237
rect 367274 233197 497974 233225
rect 367274 233185 367280 233197
rect 497968 233185 497974 233197
rect 498026 233185 498032 233237
rect 507088 233151 507094 233163
rect 367138 233123 507094 233151
rect 507088 233111 507094 233123
rect 507146 233111 507152 233163
rect 513136 233151 513142 233163
rect 512578 233123 513142 233151
rect 262096 233037 262102 233089
rect 262154 233077 262160 233089
rect 334192 233077 334198 233089
rect 262154 233049 334198 233077
rect 262154 233037 262160 233049
rect 334192 233037 334198 233049
rect 334250 233037 334256 233089
rect 334288 233037 334294 233089
rect 334346 233077 334352 233089
rect 346288 233077 346294 233089
rect 334346 233049 346294 233077
rect 334346 233037 334352 233049
rect 346288 233037 346294 233049
rect 346346 233037 346352 233089
rect 353104 233037 353110 233089
rect 353162 233077 353168 233089
rect 512578 233077 512606 233123
rect 513136 233111 513142 233123
rect 513194 233111 513200 233163
rect 353162 233049 512606 233077
rect 353162 233037 353168 233049
rect 512656 233037 512662 233089
rect 512714 233077 512720 233089
rect 590896 233077 590902 233089
rect 512714 233049 590902 233077
rect 512714 233037 512720 233049
rect 590896 233037 590902 233049
rect 590954 233037 590960 233089
rect 325360 232963 325366 233015
rect 325418 233003 325424 233015
rect 360784 233003 360790 233015
rect 325418 232975 352478 233003
rect 325418 232963 325424 232975
rect 265168 232889 265174 232941
rect 265226 232929 265232 232941
rect 335440 232929 335446 232941
rect 265226 232901 335446 232929
rect 265226 232889 265232 232901
rect 335440 232889 335446 232901
rect 335498 232889 335504 232941
rect 338032 232889 338038 232941
rect 338090 232929 338096 232941
rect 352336 232929 352342 232941
rect 338090 232901 352342 232929
rect 338090 232889 338096 232901
rect 352336 232889 352342 232901
rect 352394 232889 352400 232941
rect 352450 232929 352478 232975
rect 357106 232975 360790 233003
rect 357106 232929 357134 232975
rect 360784 232963 360790 232975
rect 360842 232963 360848 233015
rect 360880 232963 360886 233015
rect 360938 233003 360944 233015
rect 360938 232975 378878 233003
rect 360938 232963 360944 232975
rect 352450 232901 357134 232929
rect 378850 232929 378878 232975
rect 378928 232963 378934 233015
rect 378986 233003 378992 233015
rect 522160 233003 522166 233015
rect 378986 232975 522166 233003
rect 378986 232963 378992 232975
rect 522160 232963 522166 232975
rect 522218 232963 522224 233015
rect 528304 232929 528310 232941
rect 378850 232901 528310 232929
rect 528304 232889 528310 232901
rect 528362 232889 528368 232941
rect 277456 232815 277462 232867
rect 277514 232855 277520 232867
rect 295600 232855 295606 232867
rect 277514 232827 295606 232855
rect 277514 232815 277520 232827
rect 295600 232815 295606 232827
rect 295658 232815 295664 232867
rect 322480 232815 322486 232867
rect 322538 232855 322544 232867
rect 363376 232855 363382 232867
rect 322538 232827 337886 232855
rect 322538 232815 322544 232827
rect 268432 232741 268438 232793
rect 268490 232781 268496 232793
rect 334288 232781 334294 232793
rect 268490 232753 334294 232781
rect 268490 232741 268496 232753
rect 334288 232741 334294 232753
rect 334346 232741 334352 232793
rect 337858 232781 337886 232827
rect 342706 232827 363382 232855
rect 342706 232781 342734 232827
rect 363376 232815 363382 232827
rect 363434 232815 363440 232867
rect 375376 232815 375382 232867
rect 375434 232855 375440 232867
rect 378448 232855 378454 232867
rect 375434 232827 378454 232855
rect 375434 232815 375440 232827
rect 378448 232815 378454 232827
rect 378506 232815 378512 232867
rect 381424 232815 381430 232867
rect 381482 232855 381488 232867
rect 534256 232855 534262 232867
rect 381482 232827 534262 232855
rect 381482 232815 381488 232827
rect 534256 232815 534262 232827
rect 534314 232815 534320 232867
rect 337858 232753 342734 232781
rect 345520 232741 345526 232793
rect 345578 232781 345584 232793
rect 367216 232781 367222 232793
rect 345578 232753 367222 232781
rect 345578 232741 345584 232753
rect 367216 232741 367222 232753
rect 367274 232741 367280 232793
rect 378832 232741 378838 232793
rect 378890 232781 378896 232793
rect 536560 232781 536566 232793
rect 378890 232753 536566 232781
rect 378890 232741 378896 232753
rect 536560 232741 536566 232753
rect 536618 232741 536624 232793
rect 266608 232667 266614 232719
rect 266666 232707 266672 232719
rect 338224 232707 338230 232719
rect 266666 232679 338230 232707
rect 266666 232667 266672 232679
rect 338224 232667 338230 232679
rect 338282 232667 338288 232719
rect 338320 232667 338326 232719
rect 338378 232707 338384 232719
rect 356080 232707 356086 232719
rect 338378 232679 356086 232707
rect 338378 232667 338384 232679
rect 356080 232667 356086 232679
rect 356138 232667 356144 232719
rect 366640 232667 366646 232719
rect 366698 232707 366704 232719
rect 540304 232707 540310 232719
rect 366698 232679 540310 232707
rect 366698 232667 366704 232679
rect 540304 232667 540310 232679
rect 540362 232667 540368 232719
rect 271600 232593 271606 232645
rect 271658 232633 271664 232645
rect 350032 232633 350038 232645
rect 271658 232605 350038 232633
rect 271658 232593 271664 232605
rect 350032 232593 350038 232605
rect 350090 232593 350096 232645
rect 360784 232593 360790 232645
rect 360842 232633 360848 232645
rect 371248 232633 371254 232645
rect 360842 232605 371254 232633
rect 360842 232593 360848 232605
rect 371248 232593 371254 232605
rect 371306 232593 371312 232645
rect 371824 232593 371830 232645
rect 371882 232633 371888 232645
rect 380176 232633 380182 232645
rect 371882 232605 380182 232633
rect 371882 232593 371888 232605
rect 380176 232593 380182 232605
rect 380234 232593 380240 232645
rect 380272 232593 380278 232645
rect 380330 232633 380336 232645
rect 546352 232633 546358 232645
rect 380330 232605 546358 232633
rect 380330 232593 380336 232605
rect 546352 232593 546358 232605
rect 546410 232593 546416 232645
rect 219760 232519 219766 232571
rect 219818 232559 219824 232571
rect 248080 232559 248086 232571
rect 219818 232531 248086 232559
rect 219818 232519 219824 232531
rect 248080 232519 248086 232531
rect 248138 232519 248144 232571
rect 274864 232519 274870 232571
rect 274922 232559 274928 232571
rect 338320 232559 338326 232571
rect 274922 232531 338326 232559
rect 274922 232519 274928 232531
rect 338320 232519 338326 232531
rect 338378 232519 338384 232571
rect 338416 232519 338422 232571
rect 338474 232559 338480 232571
rect 358288 232559 358294 232571
rect 338474 232531 358294 232559
rect 338474 232519 338480 232531
rect 358288 232519 358294 232531
rect 358346 232519 358352 232571
rect 364912 232519 364918 232571
rect 364970 232559 364976 232571
rect 539536 232559 539542 232571
rect 364970 232531 539542 232559
rect 364970 232519 364976 232531
rect 539536 232519 539542 232531
rect 539594 232519 539600 232571
rect 218224 232445 218230 232497
rect 218282 232485 218288 232497
rect 245104 232485 245110 232497
rect 218282 232457 245110 232485
rect 218282 232445 218288 232457
rect 245104 232445 245110 232457
rect 245162 232445 245168 232497
rect 271216 232445 271222 232497
rect 271274 232485 271280 232497
rect 338032 232485 338038 232497
rect 271274 232457 338038 232485
rect 271274 232445 271280 232457
rect 338032 232445 338038 232457
rect 338090 232445 338096 232497
rect 338704 232445 338710 232497
rect 338762 232485 338768 232497
rect 361264 232485 361270 232497
rect 338762 232457 361270 232485
rect 338762 232445 338768 232457
rect 361264 232445 361270 232457
rect 361322 232445 361328 232497
rect 366256 232445 366262 232497
rect 366314 232485 366320 232497
rect 542608 232485 542614 232497
rect 366314 232457 542614 232485
rect 366314 232445 366320 232457
rect 542608 232445 542614 232457
rect 542666 232445 542672 232497
rect 221008 232371 221014 232423
rect 221066 232411 221072 232423
rect 251152 232411 251158 232423
rect 221066 232383 251158 232411
rect 221066 232371 221072 232383
rect 251152 232371 251158 232383
rect 251210 232371 251216 232423
rect 269680 232371 269686 232423
rect 269738 232411 269744 232423
rect 269738 232383 338462 232411
rect 269738 232371 269744 232383
rect 222544 232297 222550 232349
rect 222602 232337 222608 232349
rect 254224 232337 254230 232349
rect 222602 232309 254230 232337
rect 222602 232297 222608 232309
rect 254224 232297 254230 232309
rect 254282 232297 254288 232349
rect 272944 232297 272950 232349
rect 273002 232337 273008 232349
rect 337936 232337 337942 232349
rect 273002 232309 337942 232337
rect 273002 232297 273008 232309
rect 337936 232297 337942 232309
rect 337994 232297 338000 232349
rect 338434 232337 338462 232383
rect 345616 232371 345622 232423
rect 345674 232411 345680 232423
rect 379504 232411 379510 232423
rect 345674 232383 379510 232411
rect 345674 232371 345680 232383
rect 379504 232371 379510 232383
rect 379562 232371 379568 232423
rect 349360 232337 349366 232349
rect 338434 232309 349366 232337
rect 349360 232297 349366 232309
rect 349418 232297 349424 232349
rect 357616 232297 357622 232349
rect 357674 232337 357680 232349
rect 378928 232337 378934 232349
rect 357674 232309 378934 232337
rect 357674 232297 357680 232309
rect 378928 232297 378934 232309
rect 378986 232297 378992 232349
rect 380176 232297 380182 232349
rect 380234 232337 380240 232349
rect 550864 232337 550870 232349
rect 380234 232309 550870 232337
rect 380234 232297 380240 232309
rect 550864 232297 550870 232309
rect 550922 232297 550928 232349
rect 224272 232223 224278 232275
rect 224330 232263 224336 232275
rect 257200 232263 257206 232275
rect 224330 232235 257206 232263
rect 224330 232223 224336 232235
rect 257200 232223 257206 232235
rect 257258 232223 257264 232275
rect 274192 232223 274198 232275
rect 274250 232263 274256 232275
rect 338320 232263 338326 232275
rect 274250 232235 338326 232263
rect 274250 232223 274256 232235
rect 338320 232223 338326 232235
rect 338378 232223 338384 232275
rect 338416 232223 338422 232275
rect 338474 232263 338480 232275
rect 362032 232263 362038 232275
rect 338474 232235 362038 232263
rect 338474 232223 338480 232235
rect 362032 232223 362038 232235
rect 362090 232223 362096 232275
rect 363184 232223 363190 232275
rect 363242 232263 363248 232275
rect 363242 232235 368030 232263
rect 363242 232223 363248 232235
rect 224368 232149 224374 232201
rect 224426 232189 224432 232201
rect 258736 232189 258742 232201
rect 224426 232161 258742 232189
rect 224426 232149 224432 232161
rect 258736 232149 258742 232161
rect 258794 232149 258800 232201
rect 278992 232149 278998 232201
rect 279050 232189 279056 232201
rect 295504 232189 295510 232201
rect 279050 232161 295510 232189
rect 279050 232149 279056 232161
rect 295504 232149 295510 232161
rect 295562 232149 295568 232201
rect 295600 232149 295606 232201
rect 295658 232189 295664 232201
rect 364432 232189 364438 232201
rect 295658 232161 364438 232189
rect 295658 232149 295664 232161
rect 364432 232149 364438 232161
rect 364490 232149 364496 232201
rect 227440 232075 227446 232127
rect 227498 232115 227504 232127
rect 264784 232115 264790 232127
rect 227498 232087 264790 232115
rect 227498 232075 227504 232087
rect 264784 232075 264790 232087
rect 264842 232075 264848 232127
rect 275728 232075 275734 232127
rect 275786 232115 275792 232127
rect 338704 232115 338710 232127
rect 275786 232087 338710 232115
rect 275786 232075 275792 232087
rect 338704 232075 338710 232087
rect 338762 232075 338768 232127
rect 354256 232075 354262 232127
rect 354314 232115 354320 232127
rect 367120 232115 367126 232127
rect 354314 232087 367126 232115
rect 354314 232075 354320 232087
rect 367120 232075 367126 232087
rect 367178 232075 367184 232127
rect 368002 232115 368030 232235
rect 368080 232223 368086 232275
rect 368138 232263 368144 232275
rect 545584 232263 545590 232275
rect 368138 232235 545590 232263
rect 368138 232223 368144 232235
rect 545584 232223 545590 232235
rect 545642 232223 545648 232275
rect 369904 232149 369910 232201
rect 369962 232189 369968 232201
rect 380272 232189 380278 232201
rect 369962 232161 380278 232189
rect 369962 232149 369968 232161
rect 380272 232149 380278 232161
rect 380330 232149 380336 232201
rect 554704 232189 554710 232201
rect 380578 232161 554710 232189
rect 376432 232115 376438 232127
rect 368002 232087 376438 232115
rect 376432 232075 376438 232087
rect 376490 232075 376496 232127
rect 380578 232115 380606 232161
rect 554704 232149 554710 232161
rect 554762 232149 554768 232201
rect 377026 232087 380606 232115
rect 233200 232001 233206 232053
rect 233258 232041 233264 232053
rect 275344 232041 275350 232053
rect 233258 232013 275350 232041
rect 233258 232001 233264 232013
rect 275344 232001 275350 232013
rect 275402 232001 275408 232053
rect 280240 232001 280246 232053
rect 280298 232041 280304 232053
rect 370384 232041 370390 232053
rect 280298 232013 370390 232041
rect 280298 232001 280304 232013
rect 370384 232001 370390 232013
rect 370442 232001 370448 232053
rect 372304 232001 372310 232053
rect 372362 232041 372368 232053
rect 377026 232041 377054 232087
rect 380656 232075 380662 232127
rect 380714 232115 380720 232127
rect 551632 232115 551638 232127
rect 380714 232087 551638 232115
rect 380714 232075 380720 232087
rect 551632 232075 551638 232087
rect 551690 232075 551696 232127
rect 372362 232013 377054 232041
rect 372362 232001 372368 232013
rect 378448 232001 378454 232053
rect 378506 232041 378512 232053
rect 560752 232041 560758 232053
rect 378506 232013 560758 232041
rect 378506 232001 378512 232013
rect 560752 232001 560758 232013
rect 560810 232001 560816 232053
rect 234832 231927 234838 231979
rect 234890 231967 234896 231979
rect 278320 231967 278326 231979
rect 234890 231939 278326 231967
rect 234890 231927 234896 231939
rect 278320 231927 278326 231939
rect 278378 231927 278384 231979
rect 283504 231927 283510 231979
rect 283562 231967 283568 231979
rect 283562 231939 295454 231967
rect 283562 231927 283568 231939
rect 237616 231853 237622 231905
rect 237674 231893 237680 231905
rect 284368 231893 284374 231905
rect 237674 231865 284374 231893
rect 237674 231853 237680 231865
rect 284368 231853 284374 231865
rect 284426 231853 284432 231905
rect 295426 231893 295454 231939
rect 295504 231927 295510 231979
rect 295562 231967 295568 231979
rect 367408 231967 367414 231979
rect 295562 231939 367414 231967
rect 295562 231927 295568 231939
rect 367408 231927 367414 231939
rect 367466 231927 367472 231979
rect 377200 231927 377206 231979
rect 377258 231967 377264 231979
rect 561424 231967 561430 231979
rect 377258 231939 561430 231967
rect 377258 231927 377264 231939
rect 561424 231927 561430 231939
rect 561482 231927 561488 231979
rect 363184 231893 363190 231905
rect 295426 231865 363190 231893
rect 363184 231853 363190 231865
rect 363242 231853 363248 231905
rect 363298 231865 366878 231893
rect 236080 231779 236086 231831
rect 236138 231819 236144 231831
rect 281296 231819 281302 231831
rect 236138 231791 281302 231819
rect 236138 231779 236144 231791
rect 281296 231779 281302 231791
rect 281354 231779 281360 231831
rect 281968 231779 281974 231831
rect 282026 231819 282032 231831
rect 363298 231819 363326 231865
rect 282026 231791 363326 231819
rect 282026 231779 282032 231791
rect 363376 231779 363382 231831
rect 363434 231819 363440 231831
rect 365104 231819 365110 231831
rect 363434 231791 365110 231819
rect 363434 231779 363440 231791
rect 365104 231779 365110 231791
rect 365162 231779 365168 231831
rect 366850 231819 366878 231865
rect 366928 231853 366934 231905
rect 366986 231893 366992 231905
rect 377104 231893 377110 231905
rect 366986 231865 377110 231893
rect 366986 231853 366992 231865
rect 377104 231853 377110 231865
rect 377162 231853 377168 231905
rect 378544 231853 378550 231905
rect 378602 231893 378608 231905
rect 566704 231893 566710 231905
rect 378602 231865 566710 231893
rect 378602 231853 378608 231865
rect 566704 231853 566710 231865
rect 566762 231853 566768 231905
rect 373456 231819 373462 231831
rect 366850 231791 373462 231819
rect 373456 231779 373462 231791
rect 373514 231779 373520 231831
rect 376816 231779 376822 231831
rect 376874 231819 376880 231831
rect 563632 231819 563638 231831
rect 376874 231791 563638 231819
rect 376874 231779 376880 231791
rect 563632 231779 563638 231791
rect 563690 231779 563696 231831
rect 260272 231705 260278 231757
rect 260330 231745 260336 231757
rect 329584 231745 329590 231757
rect 260330 231717 329590 231745
rect 260330 231705 260336 231717
rect 329584 231705 329590 231717
rect 329642 231705 329648 231757
rect 338224 231705 338230 231757
rect 338282 231745 338288 231757
rect 343216 231745 343222 231757
rect 338282 231717 343222 231745
rect 338282 231705 338288 231717
rect 343216 231705 343222 231717
rect 343274 231705 343280 231757
rect 479152 231745 479158 231757
rect 343330 231717 479158 231745
rect 257488 231631 257494 231683
rect 257546 231671 257552 231683
rect 323632 231671 323638 231683
rect 257546 231643 323638 231671
rect 257546 231631 257552 231643
rect 323632 231631 323638 231643
rect 323690 231631 323696 231683
rect 334864 231631 334870 231683
rect 334922 231671 334928 231683
rect 343330 231671 343358 231717
rect 479152 231705 479158 231717
rect 479210 231705 479216 231757
rect 334922 231643 343358 231671
rect 334922 231631 334928 231643
rect 343408 231631 343414 231683
rect 343466 231671 343472 231683
rect 473104 231671 473110 231683
rect 343466 231643 473110 231671
rect 343466 231631 343472 231643
rect 473104 231631 473110 231643
rect 473162 231631 473168 231683
rect 243856 231557 243862 231609
rect 243914 231597 243920 231609
rect 289744 231597 289750 231609
rect 243914 231569 289750 231597
rect 243914 231557 243920 231569
rect 289744 231557 289750 231569
rect 289802 231557 289808 231609
rect 290416 231597 290422 231609
rect 289858 231569 290422 231597
rect 240592 231483 240598 231535
rect 240650 231523 240656 231535
rect 289858 231523 289886 231569
rect 290416 231557 290422 231569
rect 290474 231557 290480 231609
rect 297136 231557 297142 231609
rect 297194 231597 297200 231609
rect 400240 231597 400246 231609
rect 297194 231569 400246 231597
rect 297194 231557 297200 231569
rect 400240 231557 400246 231569
rect 400298 231557 400304 231609
rect 408976 231557 408982 231609
rect 409034 231597 409040 231609
rect 538864 231597 538870 231609
rect 409034 231569 538870 231597
rect 409034 231557 409040 231569
rect 538864 231557 538870 231569
rect 538922 231557 538928 231609
rect 240650 231495 289886 231523
rect 240650 231483 240656 231495
rect 289936 231483 289942 231535
rect 289994 231523 290000 231535
rect 386320 231523 386326 231535
rect 289994 231495 386326 231523
rect 289994 231483 290000 231495
rect 386320 231483 386326 231495
rect 386378 231483 386384 231535
rect 400336 231483 400342 231535
rect 400394 231523 400400 231535
rect 529744 231523 529750 231535
rect 400394 231495 529750 231523
rect 400394 231483 400400 231495
rect 529744 231483 529750 231495
rect 529802 231483 529808 231535
rect 248368 231409 248374 231461
rect 248426 231449 248432 231461
rect 305488 231449 305494 231461
rect 248426 231421 305494 231449
rect 248426 231409 248432 231421
rect 305488 231409 305494 231421
rect 305546 231409 305552 231461
rect 312208 231409 312214 231461
rect 312266 231449 312272 231461
rect 433840 231449 433846 231461
rect 312266 231421 433846 231449
rect 312266 231409 312272 231421
rect 433840 231409 433846 231421
rect 433898 231409 433904 231461
rect 242128 231335 242134 231387
rect 242186 231375 242192 231387
rect 242186 231347 290750 231375
rect 242186 231335 242192 231347
rect 239344 231261 239350 231313
rect 239402 231301 239408 231313
rect 287440 231301 287446 231313
rect 239402 231273 287446 231301
rect 239402 231261 239408 231273
rect 287440 231261 287446 231273
rect 287498 231261 287504 231313
rect 290722 231227 290750 231347
rect 290896 231335 290902 231387
rect 290954 231375 290960 231387
rect 302512 231375 302518 231387
rect 290954 231347 302518 231375
rect 290954 231335 290960 231347
rect 302512 231335 302518 231347
rect 302570 231335 302576 231387
rect 307600 231335 307606 231387
rect 307658 231375 307664 231387
rect 424720 231375 424726 231387
rect 307658 231347 424726 231375
rect 307658 231335 307664 231347
rect 424720 231335 424726 231347
rect 424778 231335 424784 231387
rect 290800 231261 290806 231313
rect 290858 231301 290864 231313
rect 374512 231301 374518 231313
rect 290858 231273 374518 231301
rect 290858 231261 290864 231273
rect 374512 231261 374518 231273
rect 374570 231261 374576 231313
rect 383056 231261 383062 231313
rect 383114 231301 383120 231313
rect 383114 231273 399038 231301
rect 383114 231261 383120 231273
rect 293488 231227 293494 231239
rect 290722 231199 293494 231227
rect 293488 231187 293494 231199
rect 293546 231187 293552 231239
rect 293872 231187 293878 231239
rect 293930 231227 293936 231239
rect 379984 231227 379990 231239
rect 293930 231199 379990 231227
rect 293930 231187 293936 231199
rect 379984 231187 379990 231199
rect 380042 231187 380048 231239
rect 387760 231187 387766 231239
rect 387818 231227 387824 231239
rect 392560 231227 392566 231239
rect 387818 231199 392566 231227
rect 387818 231187 387824 231199
rect 392560 231187 392566 231199
rect 392618 231187 392624 231239
rect 392848 231187 392854 231239
rect 392906 231227 392912 231239
rect 399010 231227 399038 231273
rect 403216 231261 403222 231313
rect 403274 231301 403280 231313
rect 514672 231301 514678 231313
rect 403274 231273 514678 231301
rect 403274 231261 403280 231273
rect 514672 231261 514678 231273
rect 514730 231261 514736 231313
rect 488944 231227 488950 231239
rect 392906 231199 398942 231227
rect 399010 231199 488950 231227
rect 392906 231187 392912 231199
rect 252976 231113 252982 231165
rect 253034 231153 253040 231165
rect 314512 231153 314518 231165
rect 253034 231125 314518 231153
rect 253034 231113 253040 231125
rect 314512 231113 314518 231125
rect 314570 231113 314576 231165
rect 334000 231113 334006 231165
rect 334058 231153 334064 231165
rect 334058 231125 398846 231153
rect 334058 231113 334064 231125
rect 42064 231039 42070 231091
rect 42122 231079 42128 231091
rect 42736 231079 42742 231091
rect 42122 231051 42742 231079
rect 42122 231039 42128 231051
rect 42736 231039 42742 231051
rect 42794 231039 42800 231091
rect 278224 231039 278230 231091
rect 278282 231079 278288 231091
rect 299440 231079 299446 231091
rect 278282 231051 299446 231079
rect 278282 231039 278288 231051
rect 299440 231039 299446 231051
rect 299498 231039 299504 231091
rect 299536 231039 299542 231091
rect 299594 231079 299600 231091
rect 368656 231079 368662 231091
rect 299594 231051 368662 231079
rect 299594 231039 299600 231051
rect 368656 231039 368662 231051
rect 368714 231039 368720 231091
rect 370768 231039 370774 231091
rect 370826 231079 370832 231091
rect 380656 231079 380662 231091
rect 370826 231051 380662 231079
rect 370826 231039 370832 231051
rect 380656 231039 380662 231051
rect 380714 231039 380720 231091
rect 289744 230965 289750 231017
rect 289802 231005 289808 231017
rect 296464 231005 296470 231017
rect 289802 230977 296470 231005
rect 289802 230965 289808 230977
rect 296464 230965 296470 230977
rect 296522 230965 296528 231017
rect 311056 230965 311062 231017
rect 311114 231005 311120 231017
rect 332656 231005 332662 231017
rect 311114 230977 332662 231005
rect 311114 230965 311120 230977
rect 332656 230965 332662 230977
rect 332714 230965 332720 231017
rect 339856 230965 339862 231017
rect 339914 231005 339920 231017
rect 398704 231005 398710 231017
rect 339914 230977 398710 231005
rect 339914 230965 339920 230977
rect 398704 230965 398710 230977
rect 398762 230965 398768 231017
rect 398818 231005 398846 231125
rect 398914 231079 398942 231199
rect 488944 231187 488950 231199
rect 489002 231187 489008 231239
rect 467824 231079 467830 231091
rect 398914 231051 467830 231079
rect 467824 231039 467830 231051
rect 467882 231039 467888 231091
rect 418768 231005 418774 231017
rect 398818 230977 418774 231005
rect 418768 230965 418774 230977
rect 418826 230965 418832 231017
rect 293776 230891 293782 230943
rect 293834 230931 293840 230943
rect 293834 230903 296654 230931
rect 293834 230891 293840 230903
rect 296626 230783 296654 230903
rect 308176 230891 308182 230943
rect 308234 230931 308240 230943
rect 326704 230931 326710 230943
rect 308234 230903 326710 230931
rect 308234 230891 308240 230903
rect 326704 230891 326710 230903
rect 326762 230891 326768 230943
rect 326800 230891 326806 230943
rect 326858 230931 326864 230943
rect 338320 230931 338326 230943
rect 326858 230903 338326 230931
rect 326858 230891 326864 230903
rect 338320 230891 338326 230903
rect 338378 230891 338384 230943
rect 338512 230891 338518 230943
rect 338570 230931 338576 230943
rect 395344 230931 395350 230943
rect 338570 230903 395350 230931
rect 338570 230891 338576 230903
rect 395344 230891 395350 230903
rect 395402 230891 395408 230943
rect 403408 230891 403414 230943
rect 403466 230931 403472 230943
rect 446608 230931 446614 230943
rect 403466 230903 446614 230931
rect 403466 230891 403472 230903
rect 446608 230891 446614 230903
rect 446666 230891 446672 230943
rect 305776 230817 305782 230869
rect 305834 230857 305840 230869
rect 320656 230857 320662 230869
rect 305834 230829 320662 230857
rect 305834 230817 305840 230829
rect 320656 230817 320662 230829
rect 320714 230817 320720 230869
rect 336304 230817 336310 230869
rect 336362 230857 336368 230869
rect 392368 230857 392374 230869
rect 336362 230829 392374 230857
rect 336362 230817 336368 230829
rect 392368 230817 392374 230829
rect 392426 230817 392432 230869
rect 393904 230817 393910 230869
rect 393962 230857 393968 230869
rect 443728 230857 443734 230869
rect 393962 230829 443734 230857
rect 393962 230817 393968 230829
rect 443728 230817 443734 230829
rect 443786 230817 443792 230869
rect 308560 230783 308566 230795
rect 296626 230755 308566 230783
rect 308560 230743 308566 230755
rect 308618 230743 308624 230795
rect 325840 230743 325846 230795
rect 325898 230783 325904 230795
rect 374224 230783 374230 230795
rect 325898 230755 374230 230783
rect 325898 230743 325904 230755
rect 374224 230743 374230 230755
rect 374282 230743 374288 230795
rect 376144 230743 376150 230795
rect 376202 230783 376208 230795
rect 548560 230783 548566 230795
rect 376202 230755 548566 230783
rect 376202 230743 376208 230755
rect 548560 230743 548566 230755
rect 548618 230743 548624 230795
rect 299248 230669 299254 230721
rect 299306 230709 299312 230721
rect 311632 230709 311638 230721
rect 299306 230681 311638 230709
rect 299306 230669 299312 230681
rect 311632 230669 311638 230681
rect 311690 230669 311696 230721
rect 318160 230669 318166 230721
rect 318218 230709 318224 230721
rect 338416 230709 338422 230721
rect 318218 230681 338422 230709
rect 318218 230669 318224 230681
rect 338416 230669 338422 230681
rect 338474 230669 338480 230721
rect 348496 230669 348502 230721
rect 348554 230709 348560 230721
rect 348554 230681 380414 230709
rect 348554 230669 348560 230681
rect 263920 230595 263926 230647
rect 263978 230635 263984 230647
rect 337264 230635 337270 230647
rect 263978 230607 337270 230635
rect 263978 230595 263984 230607
rect 337264 230595 337270 230607
rect 337322 230595 337328 230647
rect 380272 230635 380278 230647
rect 337378 230607 380278 230635
rect 260656 230521 260662 230573
rect 260714 230561 260720 230573
rect 331216 230561 331222 230573
rect 260714 230533 331222 230561
rect 260714 230521 260720 230533
rect 331216 230521 331222 230533
rect 331274 230521 331280 230573
rect 331312 230521 331318 230573
rect 331370 230561 331376 230573
rect 337378 230561 337406 230607
rect 380272 230595 380278 230607
rect 380330 230595 380336 230647
rect 380386 230635 380414 230681
rect 383026 230681 388814 230709
rect 383026 230635 383054 230681
rect 380386 230607 383054 230635
rect 388786 230635 388814 230681
rect 398704 230669 398710 230721
rect 398762 230709 398768 230721
rect 409648 230709 409654 230721
rect 398762 230681 409654 230709
rect 398762 230669 398768 230681
rect 409648 230669 409654 230681
rect 409706 230669 409712 230721
rect 404464 230635 404470 230647
rect 388786 230607 404470 230635
rect 404464 230595 404470 230607
rect 404522 230595 404528 230647
rect 425584 230635 425590 230647
rect 408946 230607 425590 230635
rect 331370 230533 337406 230561
rect 331370 230521 331376 230533
rect 338320 230521 338326 230573
rect 338378 230561 338384 230573
rect 366928 230561 366934 230573
rect 338378 230533 366934 230561
rect 338378 230521 338384 230533
rect 366928 230521 366934 230533
rect 366986 230521 366992 230573
rect 368080 230561 368086 230573
rect 367042 230533 368086 230561
rect 305104 230447 305110 230499
rect 305162 230487 305168 230499
rect 317584 230487 317590 230499
rect 305162 230459 317590 230487
rect 305162 230447 305168 230459
rect 317584 230447 317590 230459
rect 317642 230447 317648 230499
rect 322192 230447 322198 230499
rect 322250 230487 322256 230499
rect 367042 230487 367070 230533
rect 368080 230521 368086 230533
rect 368138 230521 368144 230573
rect 394192 230521 394198 230573
rect 394250 230561 394256 230573
rect 408946 230561 408974 230607
rect 425584 230595 425590 230607
rect 425642 230595 425648 230647
rect 394250 230533 408974 230561
rect 394250 230521 394256 230533
rect 322250 230459 367070 230487
rect 322250 230447 322256 230459
rect 367120 230447 367126 230499
rect 367178 230487 367184 230499
rect 413488 230487 413494 230499
rect 367178 230459 413494 230487
rect 367178 230447 367184 230459
rect 413488 230447 413494 230459
rect 413546 230447 413552 230499
rect 420400 230447 420406 230499
rect 420458 230487 420464 230499
rect 430096 230487 430102 230499
rect 420458 230459 430102 230487
rect 420458 230447 420464 230459
rect 430096 230447 430102 230459
rect 430154 230447 430160 230499
rect 246160 230373 246166 230425
rect 246218 230413 246224 230425
rect 298672 230413 298678 230425
rect 246218 230385 298678 230413
rect 246218 230373 246224 230385
rect 298672 230373 298678 230385
rect 298730 230373 298736 230425
rect 300208 230373 300214 230425
rect 300266 230413 300272 230425
rect 313264 230413 313270 230425
rect 300266 230385 313270 230413
rect 300266 230373 300272 230385
rect 313264 230373 313270 230385
rect 313322 230373 313328 230425
rect 325744 230373 325750 230425
rect 325802 230413 325808 230425
rect 461008 230413 461014 230425
rect 325802 230385 461014 230413
rect 325802 230373 325808 230385
rect 461008 230373 461014 230385
rect 461066 230373 461072 230425
rect 471280 230373 471286 230425
rect 471338 230413 471344 230425
rect 481456 230413 481462 230425
rect 471338 230385 481462 230413
rect 471338 230373 471344 230385
rect 481456 230373 481462 230385
rect 481514 230373 481520 230425
rect 248944 230299 248950 230351
rect 249002 230339 249008 230351
rect 304816 230339 304822 230351
rect 249002 230311 304822 230339
rect 249002 230299 249008 230311
rect 304816 230299 304822 230311
rect 304874 230299 304880 230351
rect 330256 230299 330262 230351
rect 330314 230339 330320 230351
rect 330314 230311 343550 230339
rect 330314 230299 330320 230311
rect 251920 230225 251926 230277
rect 251978 230265 251984 230277
rect 310768 230265 310774 230277
rect 251978 230237 310774 230265
rect 251978 230225 251984 230237
rect 310768 230225 310774 230237
rect 310826 230225 310832 230277
rect 336208 230225 336214 230277
rect 336266 230265 336272 230277
rect 343522 230265 343550 230311
rect 343696 230299 343702 230351
rect 343754 230339 343760 230351
rect 467056 230339 467062 230351
rect 343754 230311 467062 230339
rect 343754 230299 343760 230311
rect 467056 230299 467062 230311
rect 467114 230299 467120 230351
rect 475216 230299 475222 230351
rect 475274 230339 475280 230351
rect 487504 230339 487510 230351
rect 475274 230311 487510 230339
rect 475274 230299 475280 230311
rect 487504 230299 487510 230311
rect 487562 230299 487568 230351
rect 470128 230265 470134 230277
rect 336266 230237 342734 230265
rect 343522 230237 470134 230265
rect 336266 230225 336272 230237
rect 298192 230151 298198 230203
rect 298250 230191 298256 230203
rect 341008 230191 341014 230203
rect 298250 230163 341014 230191
rect 298250 230151 298256 230163
rect 341008 230151 341014 230163
rect 341066 230151 341072 230203
rect 342706 230191 342734 230237
rect 470128 230225 470134 230237
rect 470186 230225 470192 230277
rect 352720 230191 352726 230203
rect 342706 230163 352726 230191
rect 352720 230151 352726 230163
rect 352778 230151 352784 230203
rect 492496 230151 492502 230203
rect 492554 230191 492560 230203
rect 610480 230191 610486 230203
rect 492554 230163 610486 230191
rect 492554 230151 492560 230163
rect 610480 230151 610486 230163
rect 610538 230151 610544 230203
rect 290992 230077 290998 230129
rect 291050 230117 291056 230129
rect 338032 230117 338038 230129
rect 291050 230089 338038 230117
rect 291050 230077 291056 230089
rect 338032 230077 338038 230089
rect 338090 230077 338096 230129
rect 485200 230117 485206 230129
rect 352642 230089 485206 230117
rect 250288 230003 250294 230055
rect 250346 230043 250352 230055
rect 310000 230043 310006 230055
rect 250346 230015 310006 230043
rect 250346 230003 250352 230015
rect 310000 230003 310006 230015
rect 310058 230003 310064 230055
rect 313936 230003 313942 230055
rect 313994 230043 314000 230055
rect 321616 230043 321622 230055
rect 313994 230015 321622 230043
rect 313994 230003 314000 230015
rect 321616 230003 321622 230015
rect 321674 230003 321680 230055
rect 337552 230003 337558 230055
rect 337610 230043 337616 230055
rect 352642 230043 352670 230089
rect 485200 230077 485206 230089
rect 485258 230077 485264 230129
rect 501040 230077 501046 230129
rect 501098 230117 501104 230129
rect 613552 230117 613558 230129
rect 501098 230089 613558 230117
rect 501098 230077 501104 230089
rect 613552 230077 613558 230089
rect 613610 230077 613616 230129
rect 337610 230015 352670 230043
rect 337610 230003 337616 230015
rect 352720 230003 352726 230055
rect 352778 230043 352784 230055
rect 482128 230043 482134 230055
rect 352778 230015 482134 230043
rect 352778 230003 352784 230015
rect 482128 230003 482134 230015
rect 482186 230003 482192 230055
rect 485584 230003 485590 230055
rect 485642 230043 485648 230055
rect 604528 230043 604534 230055
rect 485642 230015 604534 230043
rect 485642 230003 485648 230015
rect 604528 230003 604534 230015
rect 604586 230003 604592 230055
rect 247024 229929 247030 229981
rect 247082 229969 247088 229981
rect 303952 229969 303958 229981
rect 247082 229941 303958 229969
rect 247082 229929 247088 229941
rect 303952 229929 303958 229941
rect 304010 229929 304016 229981
rect 304336 229929 304342 229981
rect 304394 229969 304400 229981
rect 347152 229969 347158 229981
rect 304394 229941 347158 229969
rect 304394 229929 304400 229941
rect 347152 229929 347158 229941
rect 347210 229929 347216 229981
rect 357232 229929 357238 229981
rect 357290 229969 357296 229981
rect 378928 229969 378934 229981
rect 357290 229941 378934 229969
rect 357290 229929 357296 229941
rect 378928 229929 378934 229941
rect 378986 229929 378992 229981
rect 489616 229929 489622 229981
rect 489674 229969 489680 229981
rect 607504 229969 607510 229981
rect 489674 229941 607510 229969
rect 489674 229929 489680 229941
rect 607504 229929 607510 229941
rect 607562 229929 607568 229981
rect 255184 229855 255190 229907
rect 255242 229895 255248 229907
rect 316816 229895 316822 229907
rect 255242 229867 316822 229895
rect 255242 229855 255248 229867
rect 316816 229855 316822 229867
rect 316874 229855 316880 229907
rect 317968 229855 317974 229907
rect 318026 229895 318032 229907
rect 338512 229895 338518 229907
rect 318026 229867 338518 229895
rect 318026 229855 318032 229867
rect 338512 229855 338518 229867
rect 338570 229855 338576 229907
rect 343984 229855 343990 229907
rect 344042 229895 344048 229907
rect 495088 229895 495094 229907
rect 344042 229867 495094 229895
rect 344042 229855 344048 229867
rect 495088 229855 495094 229867
rect 495146 229855 495152 229907
rect 254800 229781 254806 229833
rect 254858 229821 254864 229833
rect 319120 229821 319126 229833
rect 254858 229793 319126 229821
rect 254858 229781 254864 229793
rect 319120 229781 319126 229793
rect 319178 229781 319184 229833
rect 323440 229781 323446 229833
rect 323498 229821 323504 229833
rect 338416 229821 338422 229833
rect 323498 229793 338422 229821
rect 323498 229781 323504 229793
rect 338416 229781 338422 229793
rect 338474 229781 338480 229833
rect 347056 229781 347062 229833
rect 347114 229821 347120 229833
rect 501040 229821 501046 229833
rect 347114 229793 501046 229821
rect 347114 229781 347120 229793
rect 501040 229781 501046 229793
rect 501098 229781 501104 229833
rect 506128 229781 506134 229833
rect 506186 229821 506192 229833
rect 516112 229821 516118 229833
rect 506186 229793 516118 229821
rect 506186 229781 506192 229793
rect 516112 229781 516118 229793
rect 516170 229781 516176 229833
rect 245680 229707 245686 229759
rect 245738 229747 245744 229759
rect 300976 229747 300982 229759
rect 245738 229719 300982 229747
rect 245738 229707 245744 229719
rect 300976 229707 300982 229719
rect 301034 229707 301040 229759
rect 306640 229707 306646 229759
rect 306698 229747 306704 229759
rect 306698 229719 313214 229747
rect 306698 229707 306704 229719
rect 251536 229633 251542 229685
rect 251594 229673 251600 229685
rect 313072 229673 313078 229685
rect 251594 229645 313078 229673
rect 251594 229633 251600 229645
rect 313072 229633 313078 229645
rect 313130 229633 313136 229685
rect 313186 229673 313214 229719
rect 313264 229707 313270 229759
rect 313322 229747 313328 229759
rect 407440 229747 407446 229759
rect 313322 229719 407446 229747
rect 313322 229707 313328 229719
rect 407440 229707 407446 229719
rect 407498 229707 407504 229759
rect 416944 229707 416950 229759
rect 417002 229747 417008 229759
rect 572080 229747 572086 229759
rect 417002 229719 572086 229747
rect 417002 229707 417008 229719
rect 572080 229707 572086 229719
rect 572138 229707 572144 229759
rect 313186 229645 351710 229673
rect 220144 229559 220150 229611
rect 220202 229599 220208 229611
rect 249712 229599 249718 229611
rect 220202 229571 249718 229599
rect 220202 229559 220208 229571
rect 249712 229559 249718 229571
rect 249770 229559 249776 229611
rect 257584 229559 257590 229611
rect 257642 229599 257648 229611
rect 325168 229599 325174 229611
rect 257642 229571 325174 229599
rect 257642 229559 257648 229571
rect 325168 229559 325174 229571
rect 325226 229559 325232 229611
rect 325264 229559 325270 229611
rect 325322 229599 325328 229611
rect 338320 229599 338326 229611
rect 325322 229571 338326 229599
rect 325322 229559 325328 229571
rect 338320 229559 338326 229571
rect 338378 229559 338384 229611
rect 351682 229599 351710 229645
rect 351760 229633 351766 229685
rect 351818 229673 351824 229685
rect 351818 229645 506270 229673
rect 351818 229633 351824 229645
rect 353104 229599 353110 229611
rect 351682 229571 353110 229599
rect 353104 229559 353110 229571
rect 353162 229559 353168 229611
rect 354832 229559 354838 229611
rect 354890 229599 354896 229611
rect 506128 229599 506134 229611
rect 354890 229571 506134 229599
rect 354890 229559 354896 229571
rect 506128 229559 506134 229571
rect 506186 229559 506192 229611
rect 506242 229599 506270 229645
rect 509776 229633 509782 229685
rect 509834 229673 509840 229685
rect 614992 229673 614998 229685
rect 509834 229645 614998 229673
rect 509834 229633 509840 229645
rect 614992 229633 614998 229645
rect 615050 229633 615056 229685
rect 510160 229599 510166 229611
rect 506242 229571 510166 229599
rect 510160 229559 510166 229571
rect 510218 229559 510224 229611
rect 516208 229559 516214 229611
rect 516266 229599 516272 229611
rect 618064 229599 618070 229611
rect 516266 229571 618070 229599
rect 516266 229559 516272 229571
rect 618064 229559 618070 229571
rect 618122 229559 618128 229611
rect 222928 229485 222934 229537
rect 222986 229525 222992 229537
rect 255664 229525 255670 229537
rect 222986 229497 255670 229525
rect 222986 229485 222992 229497
rect 255664 229485 255670 229497
rect 255722 229485 255728 229537
rect 259792 229485 259798 229537
rect 259850 229525 259856 229537
rect 321424 229525 321430 229537
rect 259850 229497 321430 229525
rect 259850 229485 259856 229497
rect 321424 229485 321430 229497
rect 321482 229485 321488 229537
rect 322096 229525 322102 229537
rect 321538 229497 322102 229525
rect 221584 229411 221590 229463
rect 221642 229451 221648 229463
rect 252592 229451 252598 229463
rect 221642 229423 252598 229451
rect 221642 229411 221648 229423
rect 252592 229411 252598 229423
rect 252650 229411 252656 229463
rect 256144 229411 256150 229463
rect 256202 229451 256208 229463
rect 321538 229451 321566 229497
rect 322096 229485 322102 229497
rect 322154 229485 322160 229537
rect 328528 229485 328534 229537
rect 328586 229525 328592 229537
rect 343696 229525 343702 229537
rect 328586 229497 343702 229525
rect 328586 229485 328592 229497
rect 343696 229485 343702 229497
rect 343754 229485 343760 229537
rect 362128 229485 362134 229537
rect 362186 229525 362192 229537
rect 362186 229497 378878 229525
rect 362186 229485 362192 229497
rect 256202 229423 321566 229451
rect 256202 229411 256208 229423
rect 321616 229411 321622 229463
rect 321674 229451 321680 229463
rect 359152 229451 359158 229463
rect 321674 229423 359158 229451
rect 321674 229411 321680 229423
rect 359152 229411 359158 229423
rect 359210 229411 359216 229463
rect 365392 229411 365398 229463
rect 365450 229451 365456 229463
rect 378850 229451 378878 229497
rect 378928 229485 378934 229537
rect 378986 229525 378992 229537
rect 524464 229525 524470 229537
rect 378986 229497 524470 229525
rect 378986 229485 378992 229497
rect 524464 229485 524470 229497
rect 524522 229485 524528 229537
rect 531280 229451 531286 229463
rect 365450 229423 378734 229451
rect 378850 229423 531286 229451
rect 365450 229411 365456 229423
rect 216688 229337 216694 229389
rect 216746 229377 216752 229389
rect 242128 229377 242134 229389
rect 216746 229349 242134 229377
rect 216746 229337 216752 229349
rect 242128 229337 242134 229349
rect 242186 229337 242192 229389
rect 242800 229337 242806 229389
rect 242858 229377 242864 229389
rect 294928 229377 294934 229389
rect 242858 229349 294934 229377
rect 242858 229337 242864 229349
rect 294928 229337 294934 229349
rect 294986 229337 294992 229389
rect 296560 229337 296566 229389
rect 296618 229377 296624 229389
rect 361360 229377 361366 229389
rect 296618 229349 361366 229377
rect 296618 229337 296624 229349
rect 361360 229337 361366 229349
rect 361418 229337 361424 229389
rect 368176 229337 368182 229389
rect 368234 229377 368240 229389
rect 378706 229377 378734 229423
rect 531280 229411 531286 229423
rect 531338 229411 531344 229463
rect 537232 229377 537238 229389
rect 368234 229349 378590 229377
rect 378706 229349 537238 229377
rect 368234 229337 368240 229349
rect 226192 229263 226198 229315
rect 226250 229303 226256 229315
rect 261712 229303 261718 229315
rect 226250 229275 261718 229303
rect 226250 229263 226256 229275
rect 261712 229263 261718 229275
rect 261770 229263 261776 229315
rect 262768 229263 262774 229315
rect 262826 229303 262832 229315
rect 321328 229303 321334 229315
rect 262826 229275 321334 229303
rect 262826 229263 262832 229275
rect 321328 229263 321334 229275
rect 321386 229263 321392 229315
rect 321424 229263 321430 229315
rect 321482 229303 321488 229315
rect 325840 229303 325846 229315
rect 321482 229275 325846 229303
rect 321482 229263 321488 229275
rect 325840 229263 325846 229275
rect 325898 229263 325904 229315
rect 333040 229263 333046 229315
rect 333098 229303 333104 229315
rect 344752 229303 344758 229315
rect 333098 229275 344758 229303
rect 333098 229263 333104 229275
rect 344752 229263 344758 229275
rect 344810 229263 344816 229315
rect 371536 229303 371542 229315
rect 367138 229275 371542 229303
rect 231952 229189 231958 229241
rect 232010 229229 232016 229241
rect 273808 229229 273814 229241
rect 232010 229201 273814 229229
rect 232010 229189 232016 229201
rect 273808 229189 273814 229201
rect 273866 229189 273872 229241
rect 287920 229189 287926 229241
rect 287978 229229 287984 229241
rect 287978 229201 301886 229229
rect 287978 229189 287984 229201
rect 235216 229115 235222 229167
rect 235274 229155 235280 229167
rect 279856 229155 279862 229167
rect 235274 229127 279862 229155
rect 235274 229115 235280 229127
rect 279856 229115 279862 229127
rect 279914 229115 279920 229167
rect 286288 229115 286294 229167
rect 286346 229155 286352 229167
rect 286346 229127 289310 229155
rect 286346 229115 286352 229127
rect 239728 229041 239734 229093
rect 239786 229081 239792 229093
rect 288880 229081 288886 229093
rect 239786 229053 288886 229081
rect 239786 229041 239792 229053
rect 288880 229041 288886 229053
rect 288938 229041 288944 229093
rect 289282 229081 289310 229127
rect 289360 229115 289366 229167
rect 289418 229155 289424 229167
rect 301858 229155 301886 229201
rect 306640 229189 306646 229241
rect 306698 229229 306704 229241
rect 367024 229229 367030 229241
rect 306698 229201 367030 229229
rect 306698 229189 306704 229201
rect 367024 229189 367030 229201
rect 367082 229189 367088 229241
rect 367138 229155 367166 229275
rect 371536 229263 371542 229275
rect 371594 229263 371600 229315
rect 378562 229303 378590 229349
rect 537232 229337 537238 229349
rect 537290 229337 537296 229389
rect 543376 229303 543382 229315
rect 378562 229275 543382 229303
rect 543376 229263 543382 229275
rect 543434 229263 543440 229315
rect 564400 229263 564406 229315
rect 564458 229303 564464 229315
rect 606736 229303 606742 229315
rect 564458 229275 606742 229303
rect 564458 229263 564464 229275
rect 606736 229263 606742 229275
rect 606794 229263 606800 229315
rect 372688 229189 372694 229241
rect 372746 229229 372752 229241
rect 552400 229229 552406 229241
rect 372746 229201 552406 229229
rect 372746 229189 372752 229201
rect 552400 229189 552406 229201
rect 552458 229189 552464 229241
rect 559216 229189 559222 229241
rect 559274 229229 559280 229241
rect 603664 229229 603670 229241
rect 559274 229201 603670 229229
rect 559274 229189 559280 229201
rect 603664 229189 603670 229201
rect 603722 229189 603728 229241
rect 374416 229155 374422 229167
rect 289418 229127 298430 229155
rect 301858 229127 367166 229155
rect 367330 229127 374422 229155
rect 289418 229115 289424 229127
rect 298402 229081 298430 229127
rect 367330 229081 367358 229127
rect 374416 229115 374422 229127
rect 374474 229115 374480 229167
rect 375760 229115 375766 229167
rect 375818 229155 375824 229167
rect 558448 229155 558454 229167
rect 375818 229127 558454 229155
rect 375818 229115 375824 229127
rect 558448 229115 558454 229127
rect 558506 229115 558512 229167
rect 564304 229115 564310 229167
rect 564362 229155 564368 229167
rect 605296 229155 605302 229167
rect 564362 229127 605302 229155
rect 564362 229115 564368 229127
rect 605296 229115 605302 229127
rect 605354 229115 605360 229167
rect 289282 229053 298334 229081
rect 298402 229053 367358 229081
rect 215248 228967 215254 229019
rect 215306 229007 215312 229019
rect 239056 229007 239062 229019
rect 215306 228979 239062 229007
rect 215306 228967 215312 228979
rect 239056 228967 239062 228979
rect 239114 228967 239120 229019
rect 244144 228967 244150 229019
rect 244202 229007 244208 229019
rect 298000 229007 298006 229019
rect 244202 228979 298006 229007
rect 244202 228967 244208 228979
rect 298000 228967 298006 228979
rect 298058 228967 298064 229019
rect 298306 229007 298334 229053
rect 378736 229041 378742 229093
rect 378794 229081 378800 229093
rect 564496 229081 564502 229093
rect 378794 229053 564502 229081
rect 378794 229041 378800 229053
rect 564496 229041 564502 229053
rect 564554 229041 564560 229093
rect 306640 229007 306646 229019
rect 298306 228979 306646 229007
rect 306640 228967 306646 228979
rect 306698 228967 306704 229019
rect 312688 228967 312694 229019
rect 312746 229007 312752 229019
rect 316240 229007 316246 229019
rect 312746 228979 316246 229007
rect 312746 228967 312752 228979
rect 316240 228967 316246 228979
rect 316298 228967 316304 229019
rect 406000 229007 406006 229019
rect 316786 228979 406006 229007
rect 241072 228893 241078 228945
rect 241130 228933 241136 228945
rect 291952 228933 291958 228945
rect 241130 228905 291958 228933
rect 241130 228893 241136 228905
rect 291952 228893 291958 228905
rect 292010 228893 292016 228945
rect 298384 228893 298390 228945
rect 298442 228933 298448 228945
rect 316786 228933 316814 228979
rect 406000 228967 406006 228979
rect 406058 228967 406064 229019
rect 408304 228967 408310 229019
rect 408362 229007 408368 229019
rect 601456 229007 601462 229019
rect 408362 228979 601462 229007
rect 408362 228967 408368 228979
rect 601456 228967 601462 228979
rect 601514 228967 601520 229019
rect 298442 228905 316814 228933
rect 298442 228893 298448 228905
rect 321328 228893 321334 228945
rect 321386 228933 321392 228945
rect 331888 228933 331894 228945
rect 321386 228905 331894 228933
rect 321386 228893 321392 228905
rect 331888 228893 331894 228905
rect 331946 228893 331952 228945
rect 455152 228933 455158 228945
rect 332578 228905 455158 228933
rect 243184 228819 243190 228871
rect 243242 228859 243248 228871
rect 292624 228859 292630 228871
rect 243242 228831 292630 228859
rect 243242 228819 243248 228831
rect 292624 228819 292630 228831
rect 292682 228819 292688 228871
rect 295312 228819 295318 228871
rect 295370 228859 295376 228871
rect 332464 228859 332470 228871
rect 295370 228831 332470 228859
rect 295370 228819 295376 228831
rect 332464 228819 332470 228831
rect 332522 228819 332528 228871
rect 228880 228745 228886 228797
rect 228938 228785 228944 228797
rect 267856 228785 267862 228797
rect 228938 228757 267862 228785
rect 228938 228745 228944 228757
rect 267856 228745 267862 228757
rect 267914 228745 267920 228797
rect 274672 228745 274678 228797
rect 274730 228785 274736 228797
rect 319888 228785 319894 228797
rect 274730 228757 319894 228785
rect 274730 228745 274736 228757
rect 319888 228745 319894 228757
rect 319946 228745 319952 228797
rect 322384 228745 322390 228797
rect 322442 228785 322448 228797
rect 332578 228785 332606 228905
rect 455152 228893 455158 228905
rect 455210 228893 455216 228945
rect 455248 228893 455254 228945
rect 455306 228933 455312 228945
rect 578032 228933 578038 228945
rect 455306 228905 578038 228933
rect 455306 228893 455312 228905
rect 578032 228893 578038 228905
rect 578090 228893 578096 228945
rect 338704 228819 338710 228871
rect 338762 228859 338768 228871
rect 394576 228859 394582 228871
rect 338762 228831 394582 228859
rect 338762 228819 338768 228831
rect 394576 228819 394582 228831
rect 394634 228819 394640 228871
rect 406096 228819 406102 228871
rect 406154 228859 406160 228871
rect 535792 228859 535798 228871
rect 406154 228831 535798 228859
rect 406154 228819 406160 228831
rect 535792 228819 535798 228831
rect 535850 228819 535856 228871
rect 451984 228785 451990 228797
rect 322442 228757 332606 228785
rect 338386 228757 451990 228785
rect 322442 228745 322448 228757
rect 230800 228671 230806 228723
rect 230858 228711 230864 228723
rect 270736 228711 270742 228723
rect 230858 228683 270742 228711
rect 230858 228671 230864 228683
rect 270736 228671 270742 228683
rect 270794 228671 270800 228723
rect 270832 228671 270838 228723
rect 270890 228711 270896 228723
rect 313840 228711 313846 228723
rect 270890 228683 313846 228711
rect 270890 228671 270896 228683
rect 313840 228671 313846 228683
rect 313898 228671 313904 228723
rect 321232 228671 321238 228723
rect 321290 228711 321296 228723
rect 338386 228711 338414 228757
rect 451984 228745 451990 228757
rect 452042 228745 452048 228797
rect 321290 228683 338414 228711
rect 321290 228671 321296 228683
rect 338512 228671 338518 228723
rect 338570 228711 338576 228723
rect 445936 228711 445942 228723
rect 338570 228683 445942 228711
rect 338570 228671 338576 228683
rect 445936 228671 445942 228683
rect 445994 228671 446000 228723
rect 231664 228597 231670 228649
rect 231722 228637 231728 228649
rect 272272 228637 272278 228649
rect 231722 228609 272278 228637
rect 231722 228597 231728 228609
rect 272272 228597 272278 228609
rect 272330 228597 272336 228649
rect 272368 228597 272374 228649
rect 272426 228637 272432 228649
rect 307696 228637 307702 228649
rect 272426 228609 307702 228637
rect 272426 228597 272432 228609
rect 307696 228597 307702 228609
rect 307754 228597 307760 228649
rect 313456 228597 313462 228649
rect 313514 228637 313520 228649
rect 436912 228637 436918 228649
rect 313514 228609 436918 228637
rect 313514 228597 313520 228609
rect 436912 228597 436918 228609
rect 436970 228597 436976 228649
rect 230320 228523 230326 228575
rect 230378 228563 230384 228575
rect 269296 228563 269302 228575
rect 230378 228535 269302 228563
rect 230378 228523 230384 228535
rect 269296 228523 269302 228535
rect 269354 228523 269360 228575
rect 269392 228523 269398 228575
rect 269450 228563 269456 228575
rect 301744 228563 301750 228575
rect 269450 228535 301750 228563
rect 269450 228523 269456 228535
rect 301744 228523 301750 228535
rect 301802 228523 301808 228575
rect 308944 228523 308950 228575
rect 309002 228563 309008 228575
rect 427792 228563 427798 228575
rect 309002 228535 427798 228563
rect 309002 228523 309008 228535
rect 427792 228523 427798 228535
rect 427850 228523 427856 228575
rect 429136 228523 429142 228575
rect 429194 228563 429200 228575
rect 526000 228563 526006 228575
rect 429194 228535 526006 228563
rect 429194 228523 429200 228535
rect 526000 228523 526006 228535
rect 526058 228523 526064 228575
rect 538576 228523 538582 228575
rect 538634 228563 538640 228575
rect 541072 228563 541078 228575
rect 538634 228535 541078 228563
rect 538634 228523 538640 228535
rect 541072 228523 541078 228535
rect 541130 228523 541136 228575
rect 561712 228523 561718 228575
rect 561770 228563 561776 228575
rect 562960 228563 562966 228575
rect 561770 228535 562966 228563
rect 561770 228523 561776 228535
rect 562960 228523 562966 228535
rect 563018 228523 563024 228575
rect 567376 228523 567382 228575
rect 567434 228563 567440 228575
rect 569008 228563 569014 228575
rect 567434 228535 569014 228563
rect 567434 228523 567440 228535
rect 569008 228523 569014 228535
rect 569066 228523 569072 228575
rect 268144 228449 268150 228501
rect 268202 228489 268208 228501
rect 295696 228489 295702 228501
rect 268202 228461 295702 228489
rect 268202 228449 268208 228461
rect 295696 228449 295702 228461
rect 295754 228449 295760 228501
rect 306160 228449 306166 228501
rect 306218 228489 306224 228501
rect 421840 228489 421846 228501
rect 306218 228461 421846 228489
rect 306218 228449 306224 228461
rect 421840 228449 421846 228461
rect 421898 228449 421904 228501
rect 455056 228449 455062 228501
rect 455114 228489 455120 228501
rect 456496 228489 456502 228501
rect 455114 228461 456502 228489
rect 455114 228449 455120 228461
rect 456496 228449 456502 228461
rect 456554 228449 456560 228501
rect 466480 228449 466486 228501
rect 466538 228489 466544 228501
rect 475312 228489 475318 228501
rect 466538 228461 475318 228489
rect 466538 228449 466544 228461
rect 475312 228449 475318 228461
rect 475370 228449 475376 228501
rect 483856 228449 483862 228501
rect 483914 228489 483920 228501
rect 485968 228489 485974 228501
rect 483914 228461 485974 228489
rect 483914 228449 483920 228461
rect 485968 228449 485974 228461
rect 486026 228449 486032 228501
rect 266320 228375 266326 228427
rect 266378 228415 266384 228427
rect 289744 228415 289750 228427
rect 266378 228387 289750 228415
rect 266378 228375 266384 228387
rect 289744 228375 289750 228387
rect 289802 228375 289808 228427
rect 289840 228375 289846 228427
rect 289898 228415 289904 228427
rect 334960 228415 334966 228427
rect 289898 228387 334966 228415
rect 289898 228375 289904 228387
rect 334960 228375 334966 228387
rect 335018 228375 335024 228427
rect 340816 228375 340822 228427
rect 340874 228415 340880 228427
rect 344560 228415 344566 228427
rect 340874 228387 344566 228415
rect 340874 228375 340880 228387
rect 344560 228375 344566 228387
rect 344618 228375 344624 228427
rect 344752 228375 344758 228427
rect 344810 228415 344816 228427
rect 476176 228415 476182 228427
rect 344810 228387 476182 228415
rect 344810 228375 344816 228387
rect 476176 228375 476182 228387
rect 476234 228375 476240 228427
rect 483760 228375 483766 228427
rect 483818 228415 483824 228427
rect 493456 228415 493462 228427
rect 483818 228387 493462 228415
rect 483818 228375 483824 228387
rect 493456 228375 493462 228387
rect 493514 228375 493520 228427
rect 262000 228301 262006 228353
rect 262058 228341 262064 228353
rect 276784 228341 276790 228353
rect 262058 228313 276790 228341
rect 262058 228301 262064 228313
rect 276784 228301 276790 228313
rect 276842 228301 276848 228353
rect 279184 228301 279190 228353
rect 279242 228341 279248 228353
rect 322960 228341 322966 228353
rect 279242 228313 322966 228341
rect 279242 228301 279248 228313
rect 322960 228301 322966 228313
rect 323018 228301 323024 228353
rect 338320 228301 338326 228353
rect 338378 228341 338384 228353
rect 432400 228341 432406 228353
rect 338378 228313 432406 228341
rect 338378 228301 338384 228313
rect 432400 228301 432406 228313
rect 432458 228301 432464 228353
rect 449296 228301 449302 228353
rect 449354 228341 449360 228353
rect 460240 228341 460246 228353
rect 449354 228313 460246 228341
rect 449354 228301 449360 228313
rect 460240 228301 460246 228313
rect 460298 228301 460304 228353
rect 264688 228227 264694 228279
rect 264746 228267 264752 228279
rect 285904 228267 285910 228279
rect 264746 228239 285910 228267
rect 264746 228227 264752 228239
rect 285904 228227 285910 228239
rect 285962 228227 285968 228279
rect 291472 228227 291478 228279
rect 291530 228267 291536 228279
rect 389296 228267 389302 228279
rect 291530 228239 389302 228267
rect 291530 228227 291536 228239
rect 389296 228227 389302 228239
rect 389354 228227 389360 228279
rect 400432 228227 400438 228279
rect 400490 228267 400496 228279
rect 511600 228267 511606 228279
rect 400490 228239 511606 228267
rect 400490 228227 400496 228239
rect 511600 228227 511606 228239
rect 511658 228227 511664 228279
rect 248752 228153 248758 228205
rect 248810 228193 248816 228205
rect 307024 228193 307030 228205
rect 248810 228165 307030 228193
rect 248810 228153 248816 228165
rect 307024 228153 307030 228165
rect 307082 228153 307088 228205
rect 310192 228153 310198 228205
rect 310250 228193 310256 228205
rect 412720 228193 412726 228205
rect 310250 228165 412726 228193
rect 310250 228153 310256 228165
rect 412720 228153 412726 228165
rect 412778 228153 412784 228205
rect 303568 228079 303574 228131
rect 303626 228119 303632 228131
rect 398320 228119 398326 228131
rect 303626 228091 398326 228119
rect 303626 228079 303632 228091
rect 398320 228079 398326 228091
rect 398378 228079 398384 228131
rect 400624 228079 400630 228131
rect 400682 228119 400688 228131
rect 492016 228119 492022 228131
rect 400682 228091 492022 228119
rect 400682 228079 400688 228091
rect 492016 228079 492022 228091
rect 492074 228079 492080 228131
rect 288400 228005 288406 228057
rect 288458 228045 288464 228057
rect 383248 228045 383254 228057
rect 288458 228017 383254 228045
rect 288458 228005 288464 228017
rect 383248 228005 383254 228017
rect 383306 228005 383312 228057
rect 396976 228005 396982 228057
rect 397034 228045 397040 228057
rect 470896 228045 470902 228057
rect 397034 228017 470902 228045
rect 397034 228005 397040 228017
rect 470896 228005 470902 228017
rect 470954 228005 470960 228057
rect 253072 227931 253078 227983
rect 253130 227971 253136 227983
rect 316144 227971 316150 227983
rect 253130 227943 316150 227971
rect 253130 227931 253136 227943
rect 316144 227931 316150 227943
rect 316202 227931 316208 227983
rect 316240 227931 316246 227983
rect 316298 227971 316304 227983
rect 401392 227971 401398 227983
rect 316298 227943 401398 227971
rect 316298 227931 316304 227943
rect 401392 227931 401398 227943
rect 401450 227931 401456 227983
rect 434896 227931 434902 227983
rect 434954 227971 434960 227983
rect 442192 227971 442198 227983
rect 434954 227943 442198 227971
rect 434954 227931 434960 227943
rect 442192 227931 442198 227943
rect 442250 227931 442256 227983
rect 292528 227857 292534 227909
rect 292586 227897 292592 227909
rect 380080 227897 380086 227909
rect 292586 227869 380086 227897
rect 292586 227857 292592 227869
rect 380080 227857 380086 227869
rect 380138 227857 380144 227909
rect 391408 227857 391414 227909
rect 391466 227897 391472 227909
rect 455728 227897 455734 227909
rect 391466 227869 455734 227897
rect 391466 227857 391472 227869
rect 455728 227857 455734 227869
rect 455786 227857 455792 227909
rect 301168 227783 301174 227835
rect 301226 227823 301232 227835
rect 363280 227823 363286 227835
rect 301226 227795 363286 227823
rect 301226 227783 301232 227795
rect 363280 227783 363286 227795
rect 363338 227783 363344 227835
rect 391504 227783 391510 227835
rect 391562 227823 391568 227835
rect 440656 227823 440662 227835
rect 391562 227795 440662 227823
rect 391562 227783 391568 227795
rect 440656 227783 440662 227795
rect 440714 227783 440720 227835
rect 292144 227709 292150 227761
rect 292202 227749 292208 227761
rect 354256 227749 354262 227761
rect 292202 227721 354262 227749
rect 292202 227709 292208 227721
rect 354256 227709 354262 227721
rect 354314 227709 354320 227761
rect 385840 227709 385846 227761
rect 385898 227749 385904 227761
rect 401968 227749 401974 227761
rect 385898 227721 401974 227749
rect 385898 227709 385904 227721
rect 401968 227709 401974 227721
rect 402026 227709 402032 227761
rect 407152 227709 407158 227761
rect 407210 227749 407216 227761
rect 413200 227749 413206 227761
rect 407210 227721 413206 227749
rect 407210 227709 407216 227721
rect 413200 227709 413206 227721
rect 413258 227709 413264 227761
rect 446320 227709 446326 227761
rect 446378 227749 446384 227761
rect 454288 227749 454294 227761
rect 446378 227721 454294 227749
rect 446378 227709 446384 227721
rect 454288 227709 454294 227721
rect 454346 227709 454352 227761
rect 293968 227635 293974 227687
rect 294026 227675 294032 227687
rect 343984 227675 343990 227687
rect 294026 227647 343990 227675
rect 294026 227635 294032 227647
rect 343984 227635 343990 227647
rect 344042 227635 344048 227687
rect 344560 227635 344566 227687
rect 344618 227675 344624 227687
rect 491248 227675 491254 227687
rect 344618 227647 491254 227675
rect 344618 227635 344624 227647
rect 491248 227635 491254 227647
rect 491306 227635 491312 227687
rect 279664 227561 279670 227613
rect 279722 227601 279728 227613
rect 328912 227601 328918 227613
rect 279722 227573 328918 227601
rect 279722 227561 279728 227573
rect 328912 227561 328918 227573
rect 328970 227561 328976 227613
rect 338416 227561 338422 227613
rect 338474 227601 338480 227613
rect 435376 227601 435382 227613
rect 338474 227573 435382 227601
rect 338474 227561 338480 227573
rect 435376 227561 435382 227573
rect 435434 227561 435440 227613
rect 443440 227561 443446 227613
rect 443498 227601 443504 227613
rect 448240 227601 448246 227613
rect 443498 227573 448246 227601
rect 443498 227561 443504 227573
rect 448240 227561 448246 227573
rect 448298 227561 448304 227613
rect 460720 227561 460726 227613
rect 460778 227601 460784 227613
rect 466384 227601 466390 227613
rect 460778 227573 466390 227601
rect 460778 227561 460784 227573
rect 466384 227561 466390 227573
rect 466442 227561 466448 227613
rect 190000 227487 190006 227539
rect 190058 227527 190064 227539
rect 191536 227527 191542 227539
rect 190058 227499 191542 227527
rect 190058 227487 190064 227499
rect 191536 227487 191542 227499
rect 191594 227487 191600 227539
rect 228016 227487 228022 227539
rect 228074 227527 228080 227539
rect 262480 227527 262486 227539
rect 228074 227499 262486 227527
rect 228074 227487 228080 227499
rect 262480 227487 262486 227499
rect 262538 227487 262544 227539
rect 291088 227487 291094 227539
rect 291146 227527 291152 227539
rect 357616 227527 357622 227539
rect 291146 227499 357622 227527
rect 291146 227487 291152 227499
rect 357616 227487 357622 227499
rect 357674 227487 357680 227539
rect 392176 227487 392182 227539
rect 392234 227527 392240 227539
rect 392234 227499 394814 227527
rect 392234 227487 392240 227499
rect 226576 227413 226582 227465
rect 226634 227453 226640 227465
rect 259408 227453 259414 227465
rect 226634 227425 259414 227453
rect 226634 227413 226640 227425
rect 259408 227413 259414 227425
rect 259466 227413 259472 227465
rect 282352 227413 282358 227465
rect 282410 227453 282416 227465
rect 351568 227453 351574 227465
rect 282410 227425 351574 227453
rect 282410 227413 282416 227425
rect 351568 227413 351574 227425
rect 351626 227413 351632 227465
rect 354256 227413 354262 227465
rect 354314 227453 354320 227465
rect 393136 227453 393142 227465
rect 354314 227425 393142 227453
rect 354314 227413 354320 227425
rect 393136 227413 393142 227425
rect 393194 227413 393200 227465
rect 394786 227453 394814 227499
rect 395056 227487 395062 227539
rect 395114 227527 395120 227539
rect 584848 227527 584854 227539
rect 395114 227499 584854 227527
rect 395114 227487 395120 227499
rect 584848 227487 584854 227499
rect 584906 227487 584912 227539
rect 585232 227487 585238 227539
rect 585290 227527 585296 227539
rect 630160 227527 630166 227539
rect 585290 227499 630166 227527
rect 585290 227487 585296 227499
rect 630160 227487 630166 227499
rect 630218 227487 630224 227539
rect 592336 227453 592342 227465
rect 394786 227425 592342 227453
rect 592336 227413 592342 227425
rect 592394 227413 592400 227465
rect 606160 227413 606166 227465
rect 606218 227453 606224 227465
rect 606218 227425 619214 227453
rect 606218 227413 606224 227425
rect 232912 227339 232918 227391
rect 232970 227379 232976 227391
rect 261040 227379 261046 227391
rect 232970 227351 261046 227379
rect 232970 227339 232976 227351
rect 261040 227339 261046 227351
rect 261098 227339 261104 227391
rect 294448 227339 294454 227391
rect 294506 227379 294512 227391
rect 363664 227379 363670 227391
rect 294506 227351 363670 227379
rect 294506 227339 294512 227351
rect 363664 227339 363670 227351
rect 363722 227339 363728 227391
rect 390064 227339 390070 227391
rect 390122 227339 390128 227391
rect 390448 227339 390454 227391
rect 390506 227379 390512 227391
rect 407632 227379 407638 227391
rect 390506 227351 407638 227379
rect 390506 227339 390512 227351
rect 407632 227339 407638 227351
rect 407690 227339 407696 227391
rect 407824 227339 407830 227391
rect 407882 227379 407888 227391
rect 585616 227379 585622 227391
rect 407882 227351 585622 227379
rect 407882 227339 407888 227351
rect 585616 227339 585622 227351
rect 585674 227339 585680 227391
rect 588976 227339 588982 227391
rect 589034 227379 589040 227391
rect 599152 227379 599158 227391
rect 589034 227351 599158 227379
rect 589034 227339 589040 227351
rect 599152 227339 599158 227351
rect 599210 227339 599216 227391
rect 619186 227379 619214 227425
rect 639952 227379 639958 227391
rect 619186 227351 639958 227379
rect 639952 227339 639958 227351
rect 640010 227339 640016 227391
rect 229552 227265 229558 227317
rect 229610 227305 229616 227317
rect 265552 227305 265558 227317
rect 229610 227277 265558 227305
rect 229610 227265 229616 227277
rect 265552 227265 265558 227277
rect 265610 227265 265616 227317
rect 267952 227265 267958 227317
rect 268010 227305 268016 227317
rect 300208 227305 300214 227317
rect 268010 227277 300214 227305
rect 268010 227265 268016 227277
rect 300208 227265 300214 227277
rect 300266 227265 300272 227317
rect 300784 227265 300790 227317
rect 300842 227305 300848 227317
rect 369616 227305 369622 227317
rect 300842 227277 369622 227305
rect 300842 227265 300848 227277
rect 369616 227265 369622 227277
rect 369674 227265 369680 227317
rect 371536 227265 371542 227317
rect 371594 227305 371600 227317
rect 385552 227305 385558 227317
rect 371594 227277 385558 227305
rect 371594 227265 371600 227277
rect 385552 227265 385558 227277
rect 385610 227265 385616 227317
rect 390082 227305 390110 227339
rect 407152 227305 407158 227317
rect 390082 227277 407158 227305
rect 407152 227265 407158 227277
rect 407210 227265 407216 227317
rect 413200 227265 413206 227317
rect 413258 227305 413264 227317
rect 588592 227305 588598 227317
rect 413258 227277 588598 227305
rect 413258 227265 413264 227277
rect 588592 227265 588598 227277
rect 588650 227265 588656 227317
rect 600496 227265 600502 227317
rect 600554 227305 600560 227317
rect 634672 227305 634678 227317
rect 600554 227277 634678 227305
rect 600554 227265 600560 227277
rect 634672 227265 634678 227277
rect 634730 227265 634736 227317
rect 229744 227191 229750 227243
rect 229802 227231 229808 227243
rect 266992 227231 266998 227243
rect 229802 227203 266998 227231
rect 229802 227191 229808 227203
rect 266992 227191 266998 227203
rect 267050 227191 267056 227243
rect 273424 227191 273430 227243
rect 273482 227231 273488 227243
rect 345520 227231 345526 227243
rect 273482 227203 345526 227231
rect 273482 227191 273488 227203
rect 345520 227191 345526 227203
rect 345578 227191 345584 227243
rect 354352 227191 354358 227243
rect 354410 227231 354416 227243
rect 390064 227231 390070 227243
rect 354410 227203 390070 227231
rect 354410 227191 354416 227203
rect 390064 227191 390070 227203
rect 390122 227191 390128 227243
rect 394960 227191 394966 227243
rect 395018 227231 395024 227243
rect 395018 227203 397454 227231
rect 395018 227191 395024 227203
rect 231088 227117 231094 227169
rect 231146 227157 231152 227169
rect 268528 227157 268534 227169
rect 231146 227129 268534 227157
rect 231146 227117 231152 227129
rect 268528 227117 268534 227129
rect 268586 227117 268592 227169
rect 270640 227117 270646 227169
rect 270698 227157 270704 227169
rect 348592 227157 348598 227169
rect 270698 227129 348598 227157
rect 270698 227117 270704 227129
rect 348592 227117 348598 227129
rect 348650 227117 348656 227169
rect 359920 227117 359926 227169
rect 359978 227157 359984 227169
rect 396112 227157 396118 227169
rect 359978 227129 396118 227157
rect 359978 227117 359984 227129
rect 396112 227117 396118 227129
rect 396170 227117 396176 227169
rect 397426 227157 397454 227203
rect 399952 227191 399958 227243
rect 400010 227231 400016 227243
rect 407344 227231 407350 227243
rect 400010 227203 407350 227231
rect 400010 227191 400016 227203
rect 407344 227191 407350 227203
rect 407402 227191 407408 227243
rect 407632 227191 407638 227243
rect 407690 227231 407696 227243
rect 589360 227231 589366 227243
rect 407690 227203 589366 227231
rect 407690 227191 407696 227203
rect 589360 227191 589366 227203
rect 589418 227191 589424 227243
rect 596176 227191 596182 227243
rect 596234 227231 596240 227243
rect 633136 227231 633142 227243
rect 596234 227203 633142 227231
rect 596234 227191 596240 227203
rect 633136 227191 633142 227203
rect 633194 227191 633200 227243
rect 598480 227157 598486 227169
rect 397426 227129 598486 227157
rect 598480 227117 598486 227129
rect 598538 227117 598544 227169
rect 603376 227117 603382 227169
rect 603434 227157 603440 227169
rect 638512 227157 638518 227169
rect 603434 227129 638518 227157
rect 603434 227117 603440 227129
rect 638512 227117 638518 227129
rect 638570 227117 638576 227169
rect 233872 227043 233878 227095
rect 233930 227083 233936 227095
rect 274480 227083 274486 227095
rect 233930 227055 274486 227083
rect 233930 227043 233936 227055
rect 274480 227043 274486 227055
rect 274538 227043 274544 227095
rect 276688 227043 276694 227095
rect 276746 227083 276752 227095
rect 360592 227083 360598 227095
rect 276746 227055 360598 227083
rect 276746 227043 276752 227055
rect 360592 227043 360598 227055
rect 360650 227043 360656 227095
rect 394864 227043 394870 227095
rect 394922 227083 394928 227095
rect 597712 227083 597718 227095
rect 394922 227055 597718 227083
rect 394922 227043 394928 227055
rect 597712 227043 597718 227055
rect 597770 227043 597776 227095
rect 232528 226969 232534 227021
rect 232586 227009 232592 227021
rect 271600 227009 271606 227021
rect 232586 226981 271606 227009
rect 232586 226969 232592 226981
rect 271600 226969 271606 226981
rect 271658 226969 271664 227021
rect 279760 226969 279766 227021
rect 279818 227009 279824 227021
rect 366736 227009 366742 227021
rect 279818 226981 366742 227009
rect 279818 226969 279824 226981
rect 366736 226969 366742 226981
rect 366794 226969 366800 227021
rect 368656 226969 368662 227021
rect 368714 227009 368720 227021
rect 408208 227009 408214 227021
rect 368714 226981 408214 227009
rect 368714 226969 368720 226981
rect 408208 226969 408214 226981
rect 408266 226969 408272 227021
rect 410608 226969 410614 227021
rect 410666 227009 410672 227021
rect 612112 227009 612118 227021
rect 410666 226981 612118 227009
rect 410666 226969 410672 226981
rect 612112 226969 612118 226981
rect 612170 226969 612176 227021
rect 235600 226895 235606 226947
rect 235658 226935 235664 226947
rect 277552 226935 277558 226947
rect 235658 226907 277558 226935
rect 235658 226895 235664 226907
rect 277552 226895 277558 226907
rect 277610 226895 277616 226947
rect 282544 226895 282550 226947
rect 282602 226935 282608 226947
rect 372688 226935 372694 226947
rect 282602 226907 372694 226935
rect 282602 226895 282608 226907
rect 372688 226895 372694 226907
rect 372746 226895 372752 226947
rect 374512 226895 374518 226947
rect 374570 226935 374576 226947
rect 390736 226935 390742 226947
rect 374570 226907 390742 226935
rect 374570 226895 374576 226907
rect 390736 226895 390742 226907
rect 390794 226895 390800 226947
rect 401968 226895 401974 226947
rect 402026 226935 402032 226947
rect 406480 226935 406486 226947
rect 402026 226907 406486 226935
rect 402026 226895 402032 226907
rect 406480 226895 406486 226907
rect 406538 226895 406544 226947
rect 407344 226895 407350 226947
rect 407402 226935 407408 226947
rect 418960 226935 418966 226947
rect 407402 226907 418966 226935
rect 407402 226895 407408 226907
rect 418960 226895 418966 226907
rect 419018 226895 419024 226947
rect 419248 226895 419254 226947
rect 419306 226935 419312 226947
rect 609808 226935 609814 226947
rect 419306 226907 609814 226935
rect 419306 226895 419312 226907
rect 609808 226895 609814 226907
rect 609866 226895 609872 226947
rect 213040 226821 213046 226873
rect 213098 226861 213104 226873
rect 233776 226861 233782 226873
rect 213098 226833 233782 226861
rect 213098 226821 213104 226833
rect 233776 226821 233782 226833
rect 233834 226821 233840 226873
rect 237424 226821 237430 226873
rect 237482 226861 237488 226873
rect 282064 226861 282070 226873
rect 237482 226833 282070 226861
rect 237482 226821 237488 226833
rect 282064 226821 282070 226833
rect 282122 226821 282128 226873
rect 301552 226821 301558 226873
rect 301610 226861 301616 226873
rect 390832 226861 390838 226873
rect 301610 226833 390838 226861
rect 301610 226821 301616 226833
rect 390832 226821 390838 226833
rect 390890 226821 390896 226873
rect 401680 226821 401686 226873
rect 401738 226861 401744 226873
rect 611248 226861 611254 226873
rect 401738 226833 418910 226861
rect 401738 226821 401744 226833
rect 213808 226747 213814 226799
rect 213866 226787 213872 226799
rect 237520 226787 237526 226799
rect 213866 226759 237526 226787
rect 213866 226747 213872 226759
rect 237520 226747 237526 226759
rect 237578 226747 237584 226799
rect 238384 226747 238390 226799
rect 238442 226787 238448 226799
rect 252208 226787 252214 226799
rect 238442 226759 252214 226787
rect 238442 226747 238448 226759
rect 252208 226747 252214 226759
rect 252266 226747 252272 226799
rect 280624 226787 280630 226799
rect 252322 226759 280630 226787
rect 214576 226673 214582 226725
rect 214634 226713 214640 226725
rect 236848 226713 236854 226725
rect 214634 226685 236854 226713
rect 214634 226673 214640 226685
rect 236848 226673 236854 226685
rect 236906 226673 236912 226725
rect 252322 226713 252350 226759
rect 280624 226747 280630 226759
rect 280682 226747 280688 226799
rect 290704 226747 290710 226799
rect 290762 226787 290768 226799
rect 290762 226759 368654 226787
rect 290762 226747 290768 226759
rect 247810 226685 252350 226713
rect 216112 226599 216118 226651
rect 216170 226639 216176 226651
rect 239824 226639 239830 226651
rect 216170 226611 239830 226639
rect 216170 226599 216176 226611
rect 239824 226599 239830 226611
rect 239882 226599 239888 226651
rect 240112 226599 240118 226651
rect 240170 226639 240176 226651
rect 247696 226639 247702 226651
rect 240170 226611 247702 226639
rect 240170 226599 240176 226611
rect 247696 226599 247702 226611
rect 247754 226599 247760 226651
rect 212368 226525 212374 226577
rect 212426 226565 212432 226577
rect 234544 226565 234550 226577
rect 212426 226537 234550 226565
rect 212426 226525 212432 226537
rect 234544 226525 234550 226537
rect 234602 226525 234608 226577
rect 237040 226525 237046 226577
rect 237098 226565 237104 226577
rect 247810 226565 247838 226685
rect 252400 226673 252406 226725
rect 252458 226713 252464 226725
rect 282928 226713 282934 226725
rect 252458 226685 282934 226713
rect 252458 226673 252464 226685
rect 282928 226673 282934 226685
rect 282986 226673 282992 226725
rect 283984 226673 283990 226725
rect 284042 226713 284048 226725
rect 358480 226713 358486 226725
rect 284042 226685 358486 226713
rect 284042 226673 284048 226685
rect 358480 226673 358486 226685
rect 358538 226673 358544 226725
rect 368626 226713 368654 226759
rect 388144 226747 388150 226799
rect 388202 226787 388208 226799
rect 395056 226787 395062 226799
rect 388202 226759 395062 226787
rect 388202 226747 388208 226759
rect 395056 226747 395062 226759
rect 395114 226747 395120 226799
rect 400816 226747 400822 226799
rect 400874 226787 400880 226799
rect 413200 226787 413206 226799
rect 400874 226759 413206 226787
rect 400874 226747 400880 226759
rect 413200 226747 413206 226759
rect 413258 226747 413264 226799
rect 418882 226787 418910 226833
rect 419074 226833 611254 226861
rect 419074 226787 419102 226833
rect 611248 226821 611254 226833
rect 611306 226821 611312 226873
rect 418882 226759 419102 226787
rect 419152 226747 419158 226799
rect 419210 226787 419216 226799
rect 608944 226787 608950 226799
rect 419210 226759 608950 226787
rect 419210 226747 419216 226759
rect 608944 226747 608950 226759
rect 609002 226747 609008 226799
rect 609040 226747 609046 226799
rect 609098 226787 609104 226799
rect 629392 226787 629398 226799
rect 609098 226759 629398 226787
rect 609098 226747 609104 226759
rect 629392 226747 629398 226759
rect 629450 226747 629456 226799
rect 378736 226713 378742 226725
rect 368626 226685 378742 226713
rect 378736 226673 378742 226685
rect 378794 226673 378800 226725
rect 379984 226673 379990 226725
rect 380042 226713 380048 226725
rect 397648 226713 397654 226725
rect 380042 226685 397654 226713
rect 380042 226673 380048 226685
rect 397648 226673 397654 226685
rect 397706 226673 397712 226725
rect 402832 226673 402838 226725
rect 402890 226713 402896 226725
rect 402890 226685 419006 226713
rect 402890 226673 402896 226685
rect 247888 226599 247894 226651
rect 247946 226639 247952 226651
rect 286672 226639 286678 226651
rect 247946 226611 286678 226639
rect 247946 226599 247952 226611
rect 286672 226599 286678 226611
rect 286730 226599 286736 226651
rect 292816 226599 292822 226651
rect 292874 226639 292880 226651
rect 384784 226639 384790 226651
rect 292874 226611 384790 226639
rect 292874 226599 292880 226611
rect 384784 226599 384790 226611
rect 384842 226599 384848 226651
rect 388528 226599 388534 226651
rect 388586 226639 388592 226651
rect 407632 226639 407638 226651
rect 388586 226611 407638 226639
rect 388586 226599 388592 226611
rect 407632 226599 407638 226611
rect 407690 226599 407696 226651
rect 407728 226599 407734 226651
rect 407786 226639 407792 226651
rect 418864 226639 418870 226651
rect 407786 226611 418870 226639
rect 407786 226599 407792 226611
rect 418864 226599 418870 226611
rect 418922 226599 418928 226651
rect 418978 226639 419006 226685
rect 419056 226673 419062 226725
rect 419114 226713 419120 226725
rect 608272 226713 608278 226725
rect 419114 226685 608278 226713
rect 419114 226673 419120 226685
rect 608272 226673 608278 226685
rect 608330 226673 608336 226725
rect 609136 226673 609142 226725
rect 609194 226713 609200 226725
rect 630928 226713 630934 226725
rect 609194 226685 630934 226713
rect 609194 226673 609200 226685
rect 630928 226673 630934 226685
rect 630986 226673 630992 226725
rect 614320 226639 614326 226651
rect 418978 226611 614326 226639
rect 614320 226599 614326 226611
rect 614378 226599 614384 226651
rect 237098 226537 247838 226565
rect 237098 226525 237104 226537
rect 247984 226525 247990 226577
rect 248042 226565 248048 226577
rect 248042 226537 252158 226565
rect 248042 226525 248048 226537
rect 221680 226451 221686 226503
rect 221738 226491 221744 226503
rect 250384 226491 250390 226503
rect 221738 226463 250390 226491
rect 221738 226451 221744 226463
rect 250384 226451 250390 226463
rect 250442 226451 250448 226503
rect 252130 226491 252158 226537
rect 252208 226525 252214 226577
rect 252266 226565 252272 226577
rect 283600 226565 283606 226577
rect 252266 226537 283606 226565
rect 252266 226525 252272 226537
rect 283600 226525 283606 226537
rect 283658 226525 283664 226577
rect 293104 226525 293110 226577
rect 293162 226565 293168 226577
rect 393808 226565 393814 226577
rect 293162 226537 393814 226565
rect 293162 226525 293168 226537
rect 393808 226525 393814 226537
rect 393866 226525 393872 226577
rect 406672 226525 406678 226577
rect 406730 226565 406736 226577
rect 621808 226565 621814 226577
rect 406730 226537 621814 226565
rect 406730 226525 406736 226537
rect 621808 226525 621814 226537
rect 621866 226525 621872 226577
rect 303184 226491 303190 226503
rect 252130 226463 303190 226491
rect 303184 226451 303190 226463
rect 303242 226451 303248 226503
rect 304240 226451 304246 226503
rect 304298 226491 304304 226503
rect 409552 226491 409558 226503
rect 304298 226463 409558 226491
rect 304298 226451 304304 226463
rect 409552 226451 409558 226463
rect 409610 226451 409616 226503
rect 411952 226491 411958 226503
rect 409666 226463 411958 226491
rect 217456 226377 217462 226429
rect 217514 226417 217520 226429
rect 217514 226389 240158 226417
rect 217514 226377 217520 226389
rect 215728 226303 215734 226355
rect 215786 226343 215792 226355
rect 238384 226343 238390 226355
rect 215786 226315 238390 226343
rect 215786 226303 215792 226315
rect 238384 226303 238390 226315
rect 238442 226303 238448 226355
rect 240130 226343 240158 226389
rect 240208 226377 240214 226429
rect 240266 226417 240272 226429
rect 288112 226417 288118 226429
rect 240266 226389 288118 226417
rect 240266 226377 240272 226389
rect 288112 226377 288118 226389
rect 288170 226377 288176 226429
rect 294832 226377 294838 226429
rect 294890 226417 294896 226429
rect 396880 226417 396886 226429
rect 294890 226389 396886 226417
rect 294890 226377 294896 226389
rect 396880 226377 396886 226389
rect 396938 226377 396944 226429
rect 397552 226377 397558 226429
rect 397610 226417 397616 226429
rect 409666 226417 409694 226463
rect 411952 226451 411958 226463
rect 412010 226451 412016 226503
rect 413200 226451 413206 226503
rect 413258 226491 413264 226503
rect 419248 226491 419254 226503
rect 413258 226463 419254 226491
rect 413258 226451 413264 226463
rect 419248 226451 419254 226463
rect 419306 226451 419312 226503
rect 588880 226451 588886 226503
rect 588938 226491 588944 226503
rect 626416 226491 626422 226503
rect 588938 226463 626422 226491
rect 588938 226451 588944 226463
rect 626416 226451 626422 226463
rect 626474 226451 626480 226503
rect 629200 226451 629206 226503
rect 629258 226491 629264 226503
rect 634000 226491 634006 226503
rect 629258 226463 634006 226491
rect 629258 226451 629264 226463
rect 634000 226451 634006 226463
rect 634058 226451 634064 226503
rect 397610 226389 409694 226417
rect 397610 226377 397616 226389
rect 409744 226377 409750 226429
rect 409802 226417 409808 226429
rect 619600 226417 619606 226429
rect 409802 226389 619606 226417
rect 409802 226377 409808 226389
rect 619600 226377 619606 226389
rect 619658 226377 619664 226429
rect 241264 226343 241270 226355
rect 240130 226315 241270 226343
rect 241264 226303 241270 226315
rect 241322 226303 241328 226355
rect 243280 226303 243286 226355
rect 243338 226343 243344 226355
rect 243338 226315 250814 226343
rect 243338 226303 243344 226315
rect 217072 226229 217078 226281
rect 217130 226269 217136 226281
rect 243568 226269 243574 226281
rect 217130 226241 243574 226269
rect 217130 226229 217136 226241
rect 243568 226229 243574 226241
rect 243626 226229 243632 226281
rect 244912 226229 244918 226281
rect 244970 226269 244976 226281
rect 250786 226269 250814 226315
rect 250864 226303 250870 226355
rect 250922 226343 250928 226355
rect 285136 226343 285142 226355
rect 250922 226315 285142 226343
rect 250922 226303 250928 226315
rect 285136 226303 285142 226315
rect 285194 226303 285200 226355
rect 297616 226303 297622 226355
rect 297674 226343 297680 226355
rect 402832 226343 402838 226355
rect 297674 226315 402838 226343
rect 297674 226303 297680 226315
rect 402832 226303 402838 226315
rect 402890 226303 402896 226355
rect 407248 226303 407254 226355
rect 407306 226343 407312 226355
rect 622672 226343 622678 226355
rect 407306 226315 622678 226343
rect 407306 226303 407312 226315
rect 622672 226303 622678 226315
rect 622730 226303 622736 226355
rect 294256 226269 294262 226281
rect 244970 226241 250718 226269
rect 250786 226241 294262 226269
rect 244970 226229 244976 226241
rect 218320 226155 218326 226207
rect 218378 226195 218384 226207
rect 246640 226195 246646 226207
rect 218378 226167 246646 226195
rect 218378 226155 218384 226167
rect 246640 226155 246646 226167
rect 246698 226155 246704 226207
rect 250690 226195 250718 226241
rect 294256 226229 294262 226241
rect 294314 226229 294320 226281
rect 295216 226229 295222 226281
rect 295274 226269 295280 226281
rect 399088 226269 399094 226281
rect 295274 226241 399094 226269
rect 295274 226229 295280 226241
rect 399088 226229 399094 226241
rect 399146 226229 399152 226281
rect 400240 226229 400246 226281
rect 400298 226269 400304 226281
rect 403696 226269 403702 226281
rect 400298 226241 403702 226269
rect 400298 226229 400304 226241
rect 403696 226229 403702 226241
rect 403754 226229 403760 226281
rect 415024 226269 415030 226281
rect 411682 226241 415030 226269
rect 297232 226195 297238 226207
rect 250690 226167 297238 226195
rect 297232 226155 297238 226167
rect 297290 226155 297296 226207
rect 302128 226155 302134 226207
rect 302186 226195 302192 226207
rect 397552 226195 397558 226207
rect 302186 226167 397558 226195
rect 302186 226155 302192 226167
rect 397552 226155 397558 226167
rect 397610 226155 397616 226207
rect 408976 226195 408982 226207
rect 397666 226167 408982 226195
rect 215632 226081 215638 226133
rect 215690 226121 215696 226133
rect 240592 226121 240598 226133
rect 215690 226093 240598 226121
rect 215690 226081 215696 226093
rect 240592 226081 240598 226093
rect 240650 226081 240656 226133
rect 241840 226081 241846 226133
rect 241898 226121 241904 226133
rect 291184 226121 291190 226133
rect 241898 226093 291190 226121
rect 241898 226081 241904 226093
rect 291184 226081 291190 226093
rect 291242 226081 291248 226133
rect 300880 226081 300886 226133
rect 300938 226121 300944 226133
rect 397666 226121 397694 226167
rect 408976 226155 408982 226167
rect 409034 226155 409040 226207
rect 300938 226093 397694 226121
rect 300938 226081 300944 226093
rect 397744 226081 397750 226133
rect 397802 226121 397808 226133
rect 411682 226121 411710 226241
rect 415024 226229 415030 226241
rect 415082 226229 415088 226281
rect 418864 226229 418870 226281
rect 418922 226269 418928 226281
rect 623344 226269 623350 226281
rect 418922 226241 623350 226269
rect 418922 226229 418928 226241
rect 623344 226229 623350 226241
rect 623402 226229 623408 226281
rect 412144 226155 412150 226207
rect 412202 226195 412208 226207
rect 632368 226195 632374 226207
rect 412202 226167 632374 226195
rect 412202 226155 412208 226167
rect 632368 226155 632374 226167
rect 632426 226155 632432 226207
rect 397802 226093 411710 226121
rect 397802 226081 397808 226093
rect 411760 226081 411766 226133
rect 411818 226121 411824 226133
rect 627856 226121 627862 226133
rect 411818 226093 627862 226121
rect 411818 226081 411824 226093
rect 627856 226081 627862 226093
rect 627914 226081 627920 226133
rect 226672 226007 226678 226059
rect 226730 226047 226736 226059
rect 232912 226047 232918 226059
rect 226730 226019 232918 226047
rect 226730 226007 226736 226019
rect 232912 226007 232918 226019
rect 232970 226007 232976 226059
rect 250768 226007 250774 226059
rect 250826 226047 250832 226059
rect 254896 226047 254902 226059
rect 250826 226019 254902 226047
rect 250826 226007 250832 226019
rect 254896 226007 254902 226019
rect 254954 226007 254960 226059
rect 264880 226007 264886 226059
rect 264938 226047 264944 226059
rect 276112 226047 276118 226059
rect 264938 226019 276118 226047
rect 264938 226007 264944 226019
rect 276112 226007 276118 226019
rect 276170 226007 276176 226059
rect 321328 226047 321334 226059
rect 276466 226019 321334 226047
rect 224944 225933 224950 225985
rect 225002 225973 225008 225985
rect 256432 225973 256438 225985
rect 225002 225945 256438 225973
rect 225002 225933 225008 225945
rect 256432 225933 256438 225945
rect 256490 225933 256496 225985
rect 257104 225933 257110 225985
rect 257162 225973 257168 225985
rect 276466 225973 276494 226019
rect 321328 226007 321334 226019
rect 321386 226007 321392 226059
rect 326896 226007 326902 226059
rect 326954 226047 326960 226059
rect 387760 226047 387766 226059
rect 326954 226019 387766 226047
rect 326954 226007 326960 226019
rect 387760 226007 387766 226019
rect 387818 226007 387824 226059
rect 583408 226047 583414 226059
rect 389410 226019 583414 226047
rect 257162 225945 276494 225973
rect 257162 225933 257168 225945
rect 321136 225933 321142 225985
rect 321194 225973 321200 225985
rect 381808 225973 381814 225985
rect 321194 225945 381814 225973
rect 321194 225933 321200 225945
rect 381808 225933 381814 225945
rect 381866 225933 381872 225985
rect 387664 225933 387670 225985
rect 387722 225973 387728 225985
rect 389410 225973 389438 226019
rect 583408 226007 583414 226019
rect 583466 226007 583472 226059
rect 587440 226007 587446 226059
rect 587498 226047 587504 226059
rect 631696 226047 631702 226059
rect 587498 226019 631702 226047
rect 587498 226007 587504 226019
rect 631696 226007 631702 226019
rect 631754 226007 631760 226059
rect 387722 225945 389438 225973
rect 387722 225933 387728 225945
rect 389488 225933 389494 225985
rect 389546 225973 389552 225985
rect 587152 225973 587158 225985
rect 389546 225945 587158 225973
rect 389546 225933 389552 225945
rect 587152 225933 587158 225945
rect 587210 225933 587216 225985
rect 600400 225933 600406 225985
rect 600458 225973 600464 225985
rect 636208 225973 636214 225985
rect 600458 225945 636214 225973
rect 600458 225933 600464 225945
rect 636208 225933 636214 225945
rect 636266 225933 636272 225985
rect 218800 225859 218806 225911
rect 218858 225899 218864 225911
rect 244336 225899 244342 225911
rect 218858 225871 244342 225899
rect 218858 225859 218864 225871
rect 244336 225859 244342 225871
rect 244394 225859 244400 225911
rect 253840 225859 253846 225911
rect 253898 225899 253904 225911
rect 315376 225899 315382 225911
rect 253898 225871 315382 225899
rect 253898 225859 253904 225871
rect 315376 225859 315382 225871
rect 315434 225859 315440 225911
rect 335440 225859 335446 225911
rect 335498 225899 335504 225911
rect 340240 225899 340246 225911
rect 335498 225871 340246 225899
rect 335498 225859 335504 225871
rect 340240 225859 340246 225871
rect 340298 225859 340304 225911
rect 341968 225859 341974 225911
rect 342026 225899 342032 225911
rect 384016 225899 384022 225911
rect 342026 225871 384022 225899
rect 342026 225859 342032 225871
rect 384016 225859 384022 225871
rect 384074 225859 384080 225911
rect 387376 225859 387382 225911
rect 387434 225899 387440 225911
rect 387434 225871 388862 225899
rect 387434 225859 387440 225871
rect 220336 225785 220342 225837
rect 220394 225825 220400 225837
rect 247408 225825 247414 225837
rect 220394 225797 247414 225825
rect 220394 225785 220400 225797
rect 247408 225785 247414 225797
rect 247466 225785 247472 225837
rect 250864 225825 250870 225837
rect 250498 225797 250870 225825
rect 238768 225711 238774 225763
rect 238826 225751 238832 225763
rect 250498 225751 250526 225797
rect 250864 225785 250870 225797
rect 250922 225785 250928 225837
rect 251056 225785 251062 225837
rect 251114 225825 251120 225837
rect 251114 225797 261758 225825
rect 251114 225785 251120 225797
rect 238826 225723 250526 225751
rect 238826 225711 238832 225723
rect 250576 225711 250582 225763
rect 250634 225751 250640 225763
rect 257968 225751 257974 225763
rect 250634 225723 257974 225751
rect 250634 225711 250640 225723
rect 257968 225711 257974 225723
rect 258026 225711 258032 225763
rect 261730 225751 261758 225797
rect 271120 225785 271126 225837
rect 271178 225825 271184 225837
rect 279088 225825 279094 225837
rect 271178 225797 279094 225825
rect 271178 225785 271184 225797
rect 279088 225785 279094 225797
rect 279146 225785 279152 225837
rect 280912 225785 280918 225837
rect 280970 225825 280976 225837
rect 339472 225825 339478 225837
rect 280970 225797 339478 225825
rect 280970 225785 280976 225797
rect 339472 225785 339478 225797
rect 339530 225785 339536 225837
rect 374416 225785 374422 225837
rect 374474 225825 374480 225837
rect 388624 225825 388630 225837
rect 374474 225797 388630 225825
rect 374474 225785 374480 225797
rect 388624 225785 388630 225797
rect 388682 225785 388688 225837
rect 388834 225825 388862 225871
rect 388912 225859 388918 225911
rect 388970 225899 388976 225911
rect 586384 225899 586390 225911
rect 388970 225871 586390 225899
rect 388970 225859 388976 225871
rect 586384 225859 586390 225871
rect 586442 225859 586448 225911
rect 603280 225859 603286 225911
rect 603338 225899 603344 225911
rect 639184 225899 639190 225911
rect 603338 225871 639190 225899
rect 603338 225859 603344 225871
rect 639184 225859 639190 225871
rect 639242 225859 639248 225911
rect 582640 225825 582646 225837
rect 388834 225797 582646 225825
rect 582640 225785 582646 225797
rect 582698 225785 582704 225837
rect 603568 225785 603574 225837
rect 603626 225825 603632 225837
rect 636880 225825 636886 225837
rect 603626 225797 636886 225825
rect 603626 225785 603632 225797
rect 636880 225785 636886 225797
rect 636938 225785 636944 225837
rect 309328 225751 309334 225763
rect 261730 225723 309334 225751
rect 309328 225711 309334 225723
rect 309386 225711 309392 225763
rect 319600 225711 319606 225763
rect 319658 225751 319664 225763
rect 336400 225751 336406 225763
rect 319658 225723 336406 225751
rect 319658 225711 319664 225723
rect 336400 225711 336406 225723
rect 336458 225711 336464 225763
rect 336496 225711 336502 225763
rect 336554 225751 336560 225763
rect 354544 225751 354550 225763
rect 336554 225723 354550 225751
rect 336554 225711 336560 225723
rect 354544 225711 354550 225723
rect 354602 225711 354608 225763
rect 358480 225711 358486 225763
rect 358538 225751 358544 225763
rect 375760 225751 375766 225763
rect 358538 225723 375766 225751
rect 358538 225711 358544 225723
rect 375760 225711 375766 225723
rect 375818 225711 375824 225763
rect 390736 225711 390742 225763
rect 390794 225751 390800 225763
rect 391504 225751 391510 225763
rect 390794 225723 391510 225751
rect 390794 225711 390800 225723
rect 391504 225711 391510 225723
rect 391562 225711 391568 225763
rect 392560 225711 392566 225763
rect 392618 225751 392624 225763
rect 392618 225723 394814 225751
rect 392618 225711 392624 225723
rect 223312 225637 223318 225689
rect 223370 225677 223376 225689
rect 253456 225677 253462 225689
rect 223370 225649 253462 225677
rect 223370 225637 223376 225649
rect 253456 225637 253462 225649
rect 253514 225637 253520 225689
rect 253552 225637 253558 225689
rect 253610 225677 253616 225689
rect 269968 225677 269974 225689
rect 253610 225649 269974 225677
rect 253610 225637 253616 225649
rect 269968 225637 269974 225649
rect 270026 225637 270032 225689
rect 281200 225637 281206 225689
rect 281258 225677 281264 225689
rect 333520 225677 333526 225689
rect 281258 225649 333526 225677
rect 281258 225637 281264 225649
rect 333520 225637 333526 225649
rect 333578 225637 333584 225689
rect 380080 225637 380086 225689
rect 380138 225677 380144 225689
rect 394384 225677 394390 225689
rect 380138 225649 394390 225677
rect 380138 225637 380144 225649
rect 394384 225637 394390 225649
rect 394442 225637 394448 225689
rect 394786 225677 394814 225723
rect 394864 225711 394870 225763
rect 394922 225751 394928 225763
rect 394922 225723 398078 225751
rect 394922 225711 394928 225723
rect 398050 225677 398078 225723
rect 406480 225711 406486 225763
rect 406538 225751 406544 225763
rect 580336 225751 580342 225763
rect 406538 225723 580342 225751
rect 406538 225711 406544 225723
rect 580336 225711 580342 225723
rect 580394 225711 580400 225763
rect 603472 225711 603478 225763
rect 603530 225751 603536 225763
rect 603530 225723 619214 225751
rect 603530 225711 603536 225723
rect 581104 225677 581110 225689
rect 394786 225649 397982 225677
rect 398050 225649 581110 225677
rect 236464 225563 236470 225615
rect 236522 225603 236528 225615
rect 252400 225603 252406 225615
rect 236522 225575 252406 225603
rect 236522 225563 236528 225575
rect 252400 225563 252406 225575
rect 252458 225563 252464 225615
rect 259024 225563 259030 225615
rect 259082 225603 259088 225615
rect 273040 225603 273046 225615
rect 259082 225575 273046 225603
rect 259082 225563 259088 225575
rect 273040 225563 273046 225575
rect 273098 225563 273104 225615
rect 279280 225563 279286 225615
rect 279338 225603 279344 225615
rect 330448 225603 330454 225615
rect 279338 225575 330454 225603
rect 279338 225563 279344 225575
rect 330448 225563 330454 225575
rect 330506 225563 330512 225615
rect 367024 225563 367030 225615
rect 367082 225603 367088 225615
rect 382576 225603 382582 225615
rect 367082 225575 382582 225603
rect 367082 225563 367088 225575
rect 382576 225563 382582 225575
rect 382634 225563 382640 225615
rect 386608 225563 386614 225615
rect 386666 225603 386672 225615
rect 394480 225603 394486 225615
rect 386666 225575 394486 225603
rect 386666 225563 386672 225575
rect 394480 225563 394486 225575
rect 394538 225563 394544 225615
rect 394576 225563 394582 225615
rect 394634 225603 394640 225615
rect 397840 225603 397846 225615
rect 394634 225575 397846 225603
rect 394634 225563 394640 225575
rect 397840 225563 397846 225575
rect 397898 225563 397904 225615
rect 397954 225603 397982 225649
rect 581104 225637 581110 225649
rect 581162 225637 581168 225689
rect 585136 225637 585142 225689
rect 585194 225677 585200 225689
rect 615856 225677 615862 225689
rect 585194 225649 615862 225677
rect 585194 225637 585200 225649
rect 615856 225637 615862 225649
rect 615914 225637 615920 225689
rect 619186 225677 619214 225723
rect 626320 225711 626326 225763
rect 626378 225751 626384 225763
rect 635440 225751 635446 225763
rect 626378 225723 635446 225751
rect 626378 225711 626384 225723
rect 635440 225711 635446 225723
rect 635498 225711 635504 225763
rect 637744 225677 637750 225689
rect 619186 225649 637750 225677
rect 637744 225637 637750 225649
rect 637802 225637 637808 225689
rect 584080 225603 584086 225615
rect 397954 225575 584086 225603
rect 584080 225563 584086 225575
rect 584138 225563 584144 225615
rect 587344 225563 587350 225615
rect 587402 225603 587408 225615
rect 600784 225603 600790 225615
rect 587402 225575 600790 225603
rect 587402 225563 587408 225575
rect 600784 225563 600790 225575
rect 600842 225563 600848 225615
rect 273712 225489 273718 225541
rect 273770 225529 273776 225541
rect 318352 225529 318358 225541
rect 273770 225501 318358 225529
rect 273770 225489 273776 225501
rect 318352 225489 318358 225501
rect 318410 225489 318416 225541
rect 318928 225489 318934 225541
rect 318986 225529 318992 225541
rect 445168 225529 445174 225541
rect 318986 225501 445174 225529
rect 318986 225489 318992 225501
rect 445168 225489 445174 225501
rect 445226 225489 445232 225541
rect 582544 225489 582550 225541
rect 582602 225529 582608 225541
rect 627184 225529 627190 225541
rect 582602 225501 627190 225529
rect 582602 225489 582608 225501
rect 627184 225489 627190 225501
rect 627242 225489 627248 225541
rect 273616 225415 273622 225467
rect 273674 225455 273680 225467
rect 312304 225455 312310 225467
rect 273674 225427 312310 225455
rect 273674 225415 273680 225427
rect 312304 225415 312310 225427
rect 312362 225415 312368 225467
rect 312976 225415 312982 225467
rect 313034 225455 313040 225467
rect 433168 225455 433174 225467
rect 313034 225427 433174 225455
rect 313034 225415 313040 225427
rect 433168 225415 433174 225427
rect 433226 225415 433232 225467
rect 278128 225341 278134 225393
rect 278186 225381 278192 225393
rect 324400 225381 324406 225393
rect 278186 225353 324406 225381
rect 278186 225341 278192 225353
rect 324400 225341 324406 225353
rect 324458 225341 324464 225393
rect 332080 225341 332086 225393
rect 332138 225381 332144 225393
rect 451216 225381 451222 225393
rect 332138 225353 451222 225381
rect 332138 225341 332144 225353
rect 451216 225341 451222 225353
rect 451274 225341 451280 225393
rect 271024 225267 271030 225319
rect 271082 225307 271088 225319
rect 306256 225307 306262 225319
rect 271082 225279 306262 225307
rect 271082 225267 271088 225279
rect 306256 225267 306262 225279
rect 306314 225267 306320 225319
rect 309904 225267 309910 225319
rect 309962 225307 309968 225319
rect 427024 225307 427030 225319
rect 309962 225279 427030 225307
rect 309962 225267 309968 225279
rect 427024 225267 427030 225279
rect 427082 225267 427088 225319
rect 306736 225193 306742 225245
rect 306794 225233 306800 225245
rect 420976 225233 420982 225245
rect 306794 225205 420982 225233
rect 306794 225193 306800 225205
rect 420976 225193 420982 225205
rect 421034 225193 421040 225245
rect 303856 225119 303862 225171
rect 303914 225159 303920 225171
rect 397744 225159 397750 225171
rect 303914 225131 397750 225159
rect 303914 225119 303920 225131
rect 397744 225119 397750 225131
rect 397802 225119 397808 225171
rect 397840 225119 397846 225171
rect 397898 225159 397904 225171
rect 400624 225159 400630 225171
rect 397898 225131 400630 225159
rect 397898 225119 397904 225131
rect 400624 225119 400630 225131
rect 400682 225119 400688 225171
rect 415408 225119 415414 225171
rect 415466 225159 415472 225171
rect 628624 225159 628630 225171
rect 415466 225131 628630 225159
rect 415466 225119 415472 225131
rect 628624 225119 628630 225131
rect 628682 225119 628688 225171
rect 259888 225045 259894 225097
rect 259946 225085 259952 225097
rect 327376 225085 327382 225097
rect 259946 225057 327382 225085
rect 259946 225045 259952 225057
rect 327376 225045 327382 225057
rect 327434 225045 327440 225097
rect 328336 225045 328342 225097
rect 328394 225085 328400 225097
rect 342544 225085 342550 225097
rect 328394 225057 342550 225085
rect 328394 225045 328400 225057
rect 342544 225045 342550 225057
rect 342602 225045 342608 225097
rect 342928 225045 342934 225097
rect 342986 225085 342992 225097
rect 418000 225085 418006 225097
rect 342986 225057 418006 225085
rect 342986 225045 342992 225057
rect 418000 225045 418006 225057
rect 418058 225045 418064 225097
rect 670000 225045 670006 225097
rect 670058 225085 670064 225097
rect 676240 225085 676246 225097
rect 670058 225057 676246 225085
rect 670058 225045 670064 225057
rect 676240 225045 676246 225057
rect 676298 225045 676304 225097
rect 344656 224971 344662 225023
rect 344714 225011 344720 225023
rect 405904 225011 405910 225023
rect 344714 224983 405910 225011
rect 344714 224971 344720 224983
rect 405904 224971 405910 224983
rect 405962 224971 405968 225023
rect 406000 224971 406006 225023
rect 406058 225011 406064 225023
rect 406768 225011 406774 225023
rect 406058 224983 406774 225011
rect 406058 224971 406064 224983
rect 406768 224971 406774 224983
rect 406826 224971 406832 225023
rect 409552 224971 409558 225023
rect 409610 225011 409616 225023
rect 417232 225011 417238 225023
rect 409610 224983 417238 225011
rect 409610 224971 409616 224983
rect 417232 224971 417238 224983
rect 417290 224971 417296 225023
rect 189904 224897 189910 224949
rect 189962 224937 189968 224949
rect 192304 224937 192310 224949
rect 189962 224909 192310 224937
rect 189962 224897 189968 224909
rect 192304 224897 192310 224909
rect 192362 224897 192368 224949
rect 363280 224897 363286 224949
rect 363338 224937 363344 224949
rect 411280 224937 411286 224949
rect 363338 224909 411286 224937
rect 363338 224897 363344 224909
rect 411280 224897 411286 224909
rect 411338 224897 411344 224949
rect 250480 224823 250486 224875
rect 250538 224863 250544 224875
rect 251920 224863 251926 224875
rect 250538 224835 251926 224863
rect 250538 224823 250544 224835
rect 251920 224823 251926 224835
rect 251978 224823 251984 224875
rect 358576 224823 358582 224875
rect 358634 224863 358640 224875
rect 405136 224863 405142 224875
rect 358634 224835 405142 224863
rect 358634 224823 358640 224835
rect 405136 224823 405142 224835
rect 405194 224823 405200 224875
rect 405520 224823 405526 224875
rect 405578 224863 405584 224875
rect 409744 224863 409750 224875
rect 405578 224835 409750 224863
rect 405578 224823 405584 224835
rect 409744 224823 409750 224835
rect 409802 224823 409808 224875
rect 245008 224749 245014 224801
rect 245066 224789 245072 224801
rect 248848 224789 248854 224801
rect 245066 224761 248854 224789
rect 245066 224749 245072 224761
rect 248848 224749 248854 224761
rect 248906 224749 248912 224801
rect 361360 224749 361366 224801
rect 361418 224789 361424 224801
rect 402160 224789 402166 224801
rect 361418 224761 402166 224789
rect 361418 224749 361424 224761
rect 402160 224749 402166 224761
rect 402218 224749 402224 224801
rect 185680 224675 185686 224727
rect 185738 224715 185744 224727
rect 187120 224715 187126 224727
rect 185738 224687 187126 224715
rect 185738 224675 185744 224687
rect 187120 224675 187126 224687
rect 187178 224715 187184 224727
rect 190768 224715 190774 224727
rect 187178 224687 190774 224715
rect 187178 224675 187184 224687
rect 190768 224675 190774 224687
rect 190826 224675 190832 224727
rect 240688 224675 240694 224727
rect 240746 224715 240752 224727
rect 242896 224715 242902 224727
rect 240746 224687 242902 224715
rect 240746 224675 240752 224687
rect 242896 224675 242902 224687
rect 242954 224675 242960 224727
rect 244528 224675 244534 224727
rect 244586 224715 244592 224727
rect 245872 224715 245878 224727
rect 244586 224687 245878 224715
rect 244586 224675 244592 224687
rect 245872 224675 245878 224687
rect 245930 224675 245936 224727
rect 362704 224675 362710 224727
rect 362762 224715 362768 224727
rect 399952 224715 399958 224727
rect 362762 224687 399958 224715
rect 362762 224675 362768 224687
rect 399952 224675 399958 224687
rect 400010 224675 400016 224727
rect 400048 224675 400054 224727
rect 400106 224715 400112 224727
rect 419056 224715 419062 224727
rect 400106 224687 419062 224715
rect 400106 224675 400112 224687
rect 419056 224675 419062 224687
rect 419114 224675 419120 224727
rect 289072 224601 289078 224653
rect 289130 224641 289136 224653
rect 386992 224641 386998 224653
rect 289130 224613 386998 224641
rect 289130 224601 289136 224613
rect 386992 224601 386998 224613
rect 387050 224601 387056 224653
rect 387280 224601 387286 224653
rect 387338 224641 387344 224653
rect 517648 224641 517654 224653
rect 387338 224613 517654 224641
rect 387338 224601 387344 224613
rect 517648 224601 517654 224613
rect 517706 224601 517712 224653
rect 322288 224527 322294 224579
rect 322346 224567 322352 224579
rect 453424 224567 453430 224579
rect 322346 224539 453430 224567
rect 322346 224527 322352 224539
rect 453424 224527 453430 224539
rect 453482 224527 453488 224579
rect 325072 224453 325078 224505
rect 325130 224493 325136 224505
rect 459568 224493 459574 224505
rect 325130 224465 459574 224493
rect 325130 224453 325136 224465
rect 459568 224453 459574 224465
rect 459626 224453 459632 224505
rect 331504 224379 331510 224431
rect 331562 224419 331568 224431
rect 471568 224419 471574 224431
rect 331562 224391 471574 224419
rect 331562 224379 331568 224391
rect 471568 224379 471574 224391
rect 471626 224379 471632 224431
rect 328240 224305 328246 224357
rect 328298 224345 328304 224357
rect 465616 224345 465622 224357
rect 328298 224317 465622 224345
rect 328298 224305 328304 224317
rect 465616 224305 465622 224317
rect 465674 224305 465680 224357
rect 661360 224305 661366 224357
rect 661418 224345 661424 224357
rect 676048 224345 676054 224357
rect 661418 224317 676054 224345
rect 661418 224305 661424 224317
rect 676048 224305 676054 224317
rect 676106 224305 676112 224357
rect 275632 224231 275638 224283
rect 275690 224271 275696 224283
rect 359920 224271 359926 224283
rect 275690 224243 359926 224271
rect 275690 224231 275696 224243
rect 359920 224231 359926 224243
rect 359978 224231 359984 224283
rect 362800 224231 362806 224283
rect 362858 224271 362864 224283
rect 498832 224271 498838 224283
rect 362858 224243 498838 224271
rect 362858 224231 362864 224243
rect 498832 224231 498838 224243
rect 498890 224231 498896 224283
rect 337168 224157 337174 224209
rect 337226 224197 337232 224209
rect 483760 224197 483766 224209
rect 337226 224169 483766 224197
rect 337226 224157 337232 224169
rect 483760 224157 483766 224169
rect 483818 224157 483824 224209
rect 334480 224083 334486 224135
rect 334538 224123 334544 224135
rect 477616 224123 477622 224135
rect 334538 224095 477622 224123
rect 334538 224083 334544 224095
rect 477616 224083 477622 224095
rect 477674 224083 477680 224135
rect 338128 224009 338134 224061
rect 338186 224049 338192 224061
rect 482896 224049 482902 224061
rect 338186 224021 482902 224049
rect 338186 224009 338192 224021
rect 482896 224009 482902 224021
rect 482954 224009 482960 224061
rect 340432 223935 340438 223987
rect 340490 223975 340496 223987
rect 489712 223975 489718 223987
rect 340490 223947 489718 223975
rect 340490 223935 340496 223947
rect 489712 223935 489718 223947
rect 489770 223935 489776 223987
rect 346672 223861 346678 223913
rect 346730 223901 346736 223913
rect 346730 223873 358718 223901
rect 346730 223861 346736 223873
rect 358690 223827 358718 223873
rect 358768 223861 358774 223913
rect 358826 223901 358832 223913
rect 497296 223901 497302 223913
rect 358826 223873 497302 223901
rect 358826 223861 358832 223873
rect 497296 223861 497302 223873
rect 497354 223861 497360 223913
rect 503344 223827 503350 223839
rect 358690 223799 503350 223827
rect 503344 223787 503350 223799
rect 503402 223787 503408 223839
rect 663856 223787 663862 223839
rect 663914 223827 663920 223839
rect 676048 223827 676054 223839
rect 663914 223799 676054 223827
rect 663914 223787 663920 223799
rect 676048 223787 676054 223799
rect 676106 223787 676112 223839
rect 347920 223713 347926 223765
rect 347978 223753 347984 223765
rect 347978 223725 348494 223753
rect 347978 223713 347984 223725
rect 266512 223639 266518 223691
rect 266570 223679 266576 223691
rect 341776 223679 341782 223691
rect 266570 223651 341782 223679
rect 266570 223639 266576 223651
rect 341776 223639 341782 223651
rect 341834 223639 341840 223691
rect 264592 223565 264598 223617
rect 264650 223605 264656 223617
rect 338704 223605 338710 223617
rect 264650 223577 338710 223605
rect 264650 223565 264656 223577
rect 338704 223565 338710 223577
rect 338762 223565 338768 223617
rect 348466 223605 348494 223725
rect 361648 223713 361654 223765
rect 361706 223753 361712 223765
rect 501808 223753 501814 223765
rect 361706 223725 501814 223753
rect 361706 223713 361712 223725
rect 501808 223713 501814 223725
rect 501866 223713 501872 223765
rect 349936 223639 349942 223691
rect 349994 223679 350000 223691
rect 509392 223679 509398 223691
rect 349994 223651 509398 223679
rect 349994 223639 350000 223651
rect 509392 223639 509398 223651
rect 509450 223639 509456 223691
rect 504784 223605 504790 223617
rect 348466 223577 504790 223605
rect 504784 223565 504790 223577
rect 504842 223565 504848 223617
rect 268048 223491 268054 223543
rect 268106 223531 268112 223543
rect 344848 223531 344854 223543
rect 268106 223503 344854 223531
rect 268106 223491 268112 223503
rect 344848 223491 344854 223503
rect 344906 223491 344912 223543
rect 350800 223491 350806 223543
rect 350858 223531 350864 223543
rect 364528 223531 364534 223543
rect 350858 223503 364534 223531
rect 350858 223491 350864 223503
rect 364528 223491 364534 223503
rect 364586 223491 364592 223543
rect 364624 223491 364630 223543
rect 364682 223531 364688 223543
rect 507856 223531 507862 223543
rect 364682 223503 507862 223531
rect 364682 223491 364688 223503
rect 507856 223491 507862 223503
rect 507914 223491 507920 223543
rect 269584 223417 269590 223469
rect 269642 223457 269648 223469
rect 347728 223457 347734 223469
rect 269642 223429 347734 223457
rect 269642 223417 269648 223429
rect 347728 223417 347734 223429
rect 347786 223417 347792 223469
rect 353008 223417 353014 223469
rect 353066 223457 353072 223469
rect 515344 223457 515350 223469
rect 353066 223429 515350 223457
rect 353066 223417 353072 223429
rect 515344 223417 515350 223429
rect 515402 223417 515408 223469
rect 270928 223343 270934 223395
rect 270986 223383 270992 223395
rect 350800 223383 350806 223395
rect 270986 223355 350806 223383
rect 270986 223343 270992 223355
rect 350800 223343 350806 223355
rect 350858 223343 350864 223395
rect 352528 223343 352534 223395
rect 352586 223383 352592 223395
rect 352586 223355 364478 223383
rect 352586 223343 352592 223355
rect 272560 223269 272566 223321
rect 272618 223309 272624 223321
rect 353872 223309 353878 223321
rect 272618 223281 353878 223309
rect 272618 223269 272624 223281
rect 353872 223269 353878 223281
rect 353930 223269 353936 223321
rect 355600 223269 355606 223321
rect 355658 223309 355664 223321
rect 364450 223309 364478 223355
rect 364528 223343 364534 223395
rect 364586 223383 364592 223395
rect 510832 223383 510838 223395
rect 364586 223355 510838 223383
rect 364586 223343 364592 223355
rect 510832 223343 510838 223355
rect 510890 223343 510896 223395
rect 513904 223309 513910 223321
rect 355658 223281 364382 223309
rect 364450 223281 513910 223309
rect 355658 223269 355664 223281
rect 274096 223195 274102 223247
rect 274154 223235 274160 223247
rect 356848 223235 356854 223247
rect 274154 223207 356854 223235
rect 274154 223195 274160 223207
rect 356848 223195 356854 223207
rect 356906 223195 356912 223247
rect 364354 223235 364382 223281
rect 513904 223269 513910 223281
rect 513962 223269 513968 223321
rect 519856 223235 519862 223247
rect 364354 223207 519862 223235
rect 519856 223195 519862 223207
rect 519914 223195 519920 223247
rect 321712 223121 321718 223173
rect 321770 223161 321776 223173
rect 449680 223161 449686 223173
rect 321770 223133 449686 223161
rect 321770 223121 321776 223133
rect 449680 223121 449686 223133
rect 449738 223121 449744 223173
rect 319408 223047 319414 223099
rect 319466 223087 319472 223099
rect 447472 223087 447478 223099
rect 319466 223059 447478 223087
rect 319466 223047 319472 223059
rect 447472 223047 447478 223059
rect 447530 223047 447536 223099
rect 316336 222973 316342 223025
rect 316394 223013 316400 223025
rect 441424 223013 441430 223025
rect 316394 222985 441430 223013
rect 316394 222973 316400 222985
rect 441424 222973 441430 222985
rect 441482 222973 441488 223025
rect 315280 222899 315286 222951
rect 315338 222939 315344 222951
rect 437680 222939 437686 222951
rect 315338 222911 437686 222939
rect 315338 222899 315344 222911
rect 437680 222899 437686 222911
rect 437738 222899 437744 222951
rect 310288 222825 310294 222877
rect 310346 222865 310352 222877
rect 429328 222865 429334 222877
rect 310346 222837 429334 222865
rect 310346 222825 310352 222837
rect 429328 222825 429334 222837
rect 429386 222825 429392 222877
rect 308848 222751 308854 222803
rect 308906 222791 308912 222803
rect 426352 222791 426358 222803
rect 308906 222763 426358 222791
rect 308906 222751 308912 222763
rect 426352 222751 426358 222763
rect 426410 222751 426416 222803
rect 312592 222677 312598 222729
rect 312650 222717 312656 222729
rect 431536 222717 431542 222729
rect 312650 222689 431542 222717
rect 312650 222677 312656 222689
rect 431536 222677 431542 222689
rect 431594 222677 431600 222729
rect 277072 222603 277078 222655
rect 277130 222643 277136 222655
rect 362896 222643 362902 222655
rect 277130 222615 362902 222643
rect 277130 222603 277136 222615
rect 362896 222603 362902 222615
rect 362954 222603 362960 222655
rect 363952 222603 363958 222655
rect 364010 222643 364016 222655
rect 479920 222643 479926 222655
rect 364010 222615 479926 222643
rect 364010 222603 364016 222615
rect 479920 222603 479926 222615
rect 479978 222603 479984 222655
rect 307888 222529 307894 222581
rect 307946 222569 307952 222581
rect 422512 222569 422518 222581
rect 307946 222541 422518 222569
rect 307946 222529 307952 222541
rect 422512 222529 422518 222541
rect 422570 222529 422576 222581
rect 306544 222455 306550 222507
rect 306602 222495 306608 222507
rect 419536 222495 419542 222507
rect 306602 222467 419542 222495
rect 306602 222455 306608 222467
rect 419536 222455 419542 222467
rect 419594 222455 419600 222507
rect 302800 222381 302806 222433
rect 302858 222421 302864 222433
rect 414256 222421 414262 222433
rect 302858 222393 414262 222421
rect 302858 222381 302864 222393
rect 414256 222381 414262 222393
rect 414314 222381 414320 222433
rect 305872 222307 305878 222359
rect 305930 222347 305936 222359
rect 420208 222347 420214 222359
rect 305930 222319 420214 222347
rect 305930 222307 305936 222319
rect 420208 222307 420214 222319
rect 420266 222307 420272 222359
rect 284656 222233 284662 222285
rect 284714 222273 284720 222285
rect 378064 222273 378070 222285
rect 284714 222245 378070 222273
rect 284714 222233 284720 222245
rect 378064 222233 378070 222245
rect 378122 222233 378128 222285
rect 398512 222233 398518 222285
rect 398570 222273 398576 222285
rect 502576 222273 502582 222285
rect 398570 222245 502582 222273
rect 398570 222233 398576 222245
rect 502576 222233 502582 222245
rect 502634 222233 502640 222285
rect 343600 222159 343606 222211
rect 343658 222199 343664 222211
rect 358768 222199 358774 222211
rect 343658 222171 358774 222199
rect 343658 222159 343664 222171
rect 358768 222159 358774 222171
rect 358826 222159 358832 222211
rect 374608 222159 374614 222211
rect 374666 222199 374672 222211
rect 458800 222199 458806 222211
rect 374666 222171 458806 222199
rect 374666 222159 374672 222171
rect 458800 222159 458806 222171
rect 458858 222159 458864 222211
rect 283120 222085 283126 222137
rect 283178 222125 283184 222137
rect 374992 222125 374998 222137
rect 283178 222097 374998 222125
rect 283178 222085 283184 222097
rect 374992 222085 374998 222097
rect 375050 222085 375056 222137
rect 349552 222011 349558 222063
rect 349610 222051 349616 222063
rect 364624 222051 364630 222063
rect 349610 222023 364630 222051
rect 349610 222011 349616 222023
rect 364624 222011 364630 222023
rect 364682 222011 364688 222063
rect 157072 221715 157078 221767
rect 157130 221755 157136 221767
rect 184336 221755 184342 221767
rect 157130 221727 184342 221755
rect 157130 221715 157136 221727
rect 184336 221715 184342 221727
rect 184394 221715 184400 221767
rect 498256 221715 498262 221767
rect 498314 221755 498320 221767
rect 499552 221755 499558 221767
rect 498314 221727 499558 221755
rect 498314 221715 498320 221727
rect 499552 221715 499558 221727
rect 499610 221715 499616 221767
rect 504208 221715 504214 221767
rect 504266 221755 504272 221767
rect 506368 221755 506374 221767
rect 504266 221727 506374 221755
rect 504266 221715 504272 221727
rect 506368 221715 506374 221727
rect 506426 221715 506432 221767
rect 541552 221715 541558 221767
rect 541610 221755 541616 221767
rect 544096 221755 544102 221767
rect 541610 221727 544102 221755
rect 541610 221715 541616 221727
rect 544096 221715 544102 221727
rect 544154 221715 544160 221767
rect 553216 221715 553222 221767
rect 553274 221755 553280 221767
rect 555280 221755 555286 221767
rect 553274 221727 555286 221755
rect 553274 221715 553280 221727
rect 555280 221715 555286 221727
rect 555338 221715 555344 221767
rect 576016 221715 576022 221767
rect 576074 221755 576080 221767
rect 577312 221755 577318 221767
rect 576074 221727 577318 221755
rect 576074 221715 576080 221727
rect 577312 221715 577318 221727
rect 577370 221715 577376 221767
rect 645136 221271 645142 221323
rect 645194 221311 645200 221323
rect 650032 221311 650038 221323
rect 645194 221283 650038 221311
rect 645194 221271 645200 221283
rect 650032 221271 650038 221283
rect 650090 221271 650096 221323
rect 149584 218903 149590 218955
rect 149642 218943 149648 218955
rect 165520 218943 165526 218955
rect 149642 218915 165526 218943
rect 149642 218903 149648 218915
rect 165520 218903 165526 218915
rect 165578 218903 165584 218955
rect 147376 216831 147382 216883
rect 147434 216871 147440 216883
rect 151504 216871 151510 216883
rect 147434 216843 151510 216871
rect 147434 216831 147440 216843
rect 151504 216831 151510 216843
rect 151562 216831 151568 216883
rect 645136 216831 645142 216883
rect 645194 216871 645200 216883
rect 649936 216871 649942 216883
rect 645194 216843 649942 216871
rect 645194 216831 645200 216843
rect 649936 216831 649942 216843
rect 649994 216831 650000 216883
rect 41584 216461 41590 216513
rect 41642 216501 41648 216513
rect 45136 216501 45142 216513
rect 41642 216473 45142 216501
rect 41642 216461 41648 216473
rect 45136 216461 45142 216473
rect 45194 216461 45200 216513
rect 674800 216387 674806 216439
rect 674858 216427 674864 216439
rect 676048 216427 676054 216439
rect 674858 216399 676054 216427
rect 674858 216387 674864 216399
rect 676048 216387 676054 216399
rect 676106 216387 676112 216439
rect 147280 216239 147286 216291
rect 147338 216279 147344 216291
rect 151216 216279 151222 216291
rect 147338 216251 151222 216279
rect 147338 216239 147344 216251
rect 151216 216239 151222 216251
rect 151274 216239 151280 216291
rect 41776 215721 41782 215773
rect 41834 215761 41840 215773
rect 44944 215761 44950 215773
rect 41834 215733 44950 215761
rect 41834 215721 41840 215733
rect 44944 215721 44950 215733
rect 45002 215721 45008 215773
rect 41776 215203 41782 215255
rect 41834 215243 41840 215255
rect 45232 215243 45238 215255
rect 41834 215215 45238 215243
rect 41834 215203 41840 215215
rect 45232 215203 45238 215215
rect 45290 215203 45296 215255
rect 41584 214981 41590 215033
rect 41642 215021 41648 215033
rect 43504 215021 43510 215033
rect 41642 214993 43510 215021
rect 41642 214981 41648 214993
rect 43504 214981 43510 214993
rect 43562 214981 43568 215033
rect 674416 214907 674422 214959
rect 674474 214947 674480 214959
rect 676048 214947 676054 214959
rect 674474 214919 676054 214947
rect 674474 214907 674480 214919
rect 676048 214907 676054 214919
rect 676106 214907 676112 214959
rect 41776 214241 41782 214293
rect 41834 214281 41840 214293
rect 45328 214281 45334 214293
rect 41834 214253 45334 214281
rect 41834 214241 41840 214253
rect 45328 214241 45334 214253
rect 45386 214241 45392 214293
rect 41776 213649 41782 213701
rect 41834 213689 41840 213701
rect 44656 213689 44662 213701
rect 41834 213661 44662 213689
rect 41834 213649 41840 213661
rect 44656 213649 44662 213661
rect 44714 213649 44720 213701
rect 41776 213279 41782 213331
rect 41834 213319 41840 213331
rect 43216 213319 43222 213331
rect 41834 213291 43222 213319
rect 41834 213279 41840 213291
rect 43216 213279 43222 213291
rect 43274 213279 43280 213331
rect 147376 213279 147382 213331
rect 147434 213319 147440 213331
rect 151408 213319 151414 213331
rect 147434 213291 151414 213319
rect 147434 213279 147440 213291
rect 151408 213279 151414 213291
rect 151466 213279 151472 213331
rect 674512 213279 674518 213331
rect 674570 213319 674576 213331
rect 675952 213319 675958 213331
rect 674570 213291 675958 213319
rect 674570 213279 674576 213291
rect 675952 213279 675958 213291
rect 676010 213279 676016 213331
rect 674608 213205 674614 213257
rect 674666 213245 674672 213257
rect 676240 213245 676246 213257
rect 674666 213217 676246 213245
rect 674666 213205 674672 213217
rect 676240 213205 676246 213217
rect 676298 213205 676304 213257
rect 149488 213131 149494 213183
rect 149546 213171 149552 213183
rect 182800 213171 182806 213183
rect 149546 213143 182806 213171
rect 149546 213131 149552 213143
rect 182800 213131 182806 213143
rect 182858 213131 182864 213183
rect 674704 213131 674710 213183
rect 674762 213171 674768 213183
rect 676048 213171 676054 213183
rect 674762 213143 676054 213171
rect 674762 213131 674768 213143
rect 676048 213131 676054 213143
rect 676106 213131 676112 213183
rect 41584 212909 41590 212961
rect 41642 212949 41648 212961
rect 44560 212949 44566 212961
rect 41642 212921 44566 212949
rect 41642 212909 41648 212921
rect 44560 212909 44566 212921
rect 44618 212909 44624 212961
rect 645136 212909 645142 212961
rect 645194 212949 645200 212961
rect 649840 212949 649846 212961
rect 645194 212921 649846 212949
rect 645194 212909 645200 212921
rect 649840 212909 649846 212921
rect 649898 212909 649904 212961
rect 147088 212465 147094 212517
rect 147146 212505 147152 212517
rect 151696 212505 151702 212517
rect 147146 212477 151702 212505
rect 147146 212465 147152 212477
rect 151696 212465 151702 212477
rect 151754 212465 151760 212517
rect 41776 212169 41782 212221
rect 41834 212209 41840 212221
rect 43408 212209 43414 212221
rect 41834 212181 43414 212209
rect 41834 212169 41840 212181
rect 43408 212169 43414 212181
rect 43466 212169 43472 212221
rect 147376 210319 147382 210371
rect 147434 210359 147440 210371
rect 151312 210359 151318 210371
rect 147434 210331 151318 210359
rect 147434 210319 147440 210331
rect 151312 210319 151318 210331
rect 151370 210319 151376 210371
rect 149488 210245 149494 210297
rect 149546 210285 149552 210297
rect 179920 210285 179926 210297
rect 149546 210257 179926 210285
rect 149546 210245 149552 210257
rect 179920 210245 179926 210257
rect 179978 210245 179984 210297
rect 646576 210245 646582 210297
rect 646634 210285 646640 210297
rect 679792 210285 679798 210297
rect 646634 210257 679798 210285
rect 646634 210245 646640 210257
rect 679792 210245 679798 210257
rect 679850 210245 679856 210297
rect 645136 209801 645142 209853
rect 645194 209841 645200 209853
rect 649744 209841 649750 209853
rect 645194 209813 649750 209841
rect 645194 209801 645200 209813
rect 649744 209801 649750 209813
rect 649802 209801 649808 209853
rect 147280 207433 147286 207485
rect 147338 207473 147344 207485
rect 151600 207473 151606 207485
rect 147338 207445 151606 207473
rect 147338 207433 147344 207445
rect 151600 207433 151606 207445
rect 151658 207433 151664 207485
rect 149488 207359 149494 207411
rect 149546 207399 149552 207411
rect 177040 207399 177046 207411
rect 149546 207371 177046 207399
rect 149546 207359 149552 207371
rect 177040 207359 177046 207371
rect 177098 207359 177104 207411
rect 41872 206175 41878 206227
rect 41930 206215 41936 206227
rect 42736 206215 42742 206227
rect 41930 206187 42742 206215
rect 41930 206175 41936 206187
rect 42736 206175 42742 206187
rect 42794 206175 42800 206227
rect 645136 206027 645142 206079
rect 645194 206067 645200 206079
rect 649648 206067 649654 206079
rect 645194 206039 649654 206067
rect 645194 206027 645200 206039
rect 649648 206027 649654 206039
rect 649706 206027 649712 206079
rect 675760 205953 675766 206005
rect 675818 205953 675824 206005
rect 41776 205879 41782 205931
rect 41834 205919 41840 205931
rect 43120 205919 43126 205931
rect 41834 205891 43126 205919
rect 41834 205879 41840 205891
rect 43120 205879 43126 205891
rect 43178 205879 43184 205931
rect 675778 205783 675806 205953
rect 675760 205731 675766 205783
rect 675818 205731 675824 205783
rect 41584 205139 41590 205191
rect 41642 205179 41648 205191
rect 42928 205179 42934 205191
rect 41642 205151 42934 205179
rect 41642 205139 41648 205151
rect 42928 205139 42934 205151
rect 42986 205139 42992 205191
rect 41680 204917 41686 204969
rect 41738 204957 41744 204969
rect 45040 204957 45046 204969
rect 41738 204929 45046 204957
rect 41738 204917 41744 204929
rect 45040 204917 45046 204929
rect 45098 204917 45104 204969
rect 41584 204843 41590 204895
rect 41642 204883 41648 204895
rect 42832 204883 42838 204895
rect 41642 204855 42838 204883
rect 41642 204843 41648 204855
rect 42832 204843 42838 204855
rect 42890 204843 42896 204895
rect 41776 204547 41782 204599
rect 41834 204587 41840 204599
rect 43024 204587 43030 204599
rect 41834 204559 43030 204587
rect 41834 204547 41840 204559
rect 43024 204547 43030 204559
rect 43082 204547 43088 204599
rect 149488 204547 149494 204599
rect 149546 204587 149552 204599
rect 168592 204587 168598 204599
rect 149546 204559 168598 204587
rect 149546 204547 149552 204559
rect 168592 204547 168598 204559
rect 168650 204547 168656 204599
rect 149296 204473 149302 204525
rect 149354 204513 149360 204525
rect 174256 204513 174262 204525
rect 149354 204485 174262 204513
rect 149354 204473 149360 204485
rect 174256 204473 174262 204485
rect 174314 204473 174320 204525
rect 41776 204325 41782 204377
rect 41834 204365 41840 204377
rect 44752 204365 44758 204377
rect 41834 204337 44758 204365
rect 41834 204325 41840 204337
rect 44752 204325 44758 204337
rect 44810 204325 44816 204377
rect 41776 203733 41782 203785
rect 41834 203773 41840 203785
rect 44848 203773 44854 203785
rect 41834 203745 44854 203773
rect 41834 203733 41840 203745
rect 44848 203733 44854 203745
rect 44906 203733 44912 203785
rect 674800 202031 674806 202083
rect 674858 202071 674864 202083
rect 675472 202071 675478 202083
rect 674858 202043 675478 202071
rect 674858 202031 674864 202043
rect 675472 202031 675478 202043
rect 675530 202031 675536 202083
rect 149680 201661 149686 201713
rect 149738 201701 149744 201713
rect 180016 201701 180022 201713
rect 149738 201673 180022 201701
rect 149738 201661 149744 201673
rect 180016 201661 180022 201673
rect 180074 201661 180080 201713
rect 149488 201587 149494 201639
rect 149546 201627 149552 201639
rect 182896 201627 182902 201639
rect 149546 201599 182902 201627
rect 149546 201587 149552 201599
rect 182896 201587 182902 201599
rect 182954 201587 182960 201639
rect 145744 201513 145750 201565
rect 145802 201553 145808 201565
rect 184336 201553 184342 201565
rect 145802 201525 184342 201553
rect 145802 201513 145808 201525
rect 184336 201513 184342 201525
rect 184394 201513 184400 201565
rect 645136 201513 645142 201565
rect 645194 201553 645200 201565
rect 649552 201553 649558 201565
rect 645194 201525 649558 201553
rect 645194 201513 645200 201525
rect 649552 201513 649558 201525
rect 649610 201513 649616 201565
rect 674704 200847 674710 200899
rect 674762 200887 674768 200899
rect 675376 200887 675382 200899
rect 674762 200859 675382 200887
rect 674762 200847 674768 200859
rect 675376 200847 675382 200859
rect 675434 200847 675440 200899
rect 149296 198775 149302 198827
rect 149354 198815 149360 198827
rect 159952 198815 159958 198827
rect 149354 198787 159958 198815
rect 149354 198775 149360 198787
rect 159952 198775 159958 198787
rect 160010 198775 160016 198827
rect 149488 198701 149494 198753
rect 149546 198741 149552 198753
rect 177136 198741 177142 198753
rect 149546 198713 177142 198741
rect 149546 198701 149552 198713
rect 177136 198701 177142 198713
rect 177194 198701 177200 198753
rect 181360 198627 181366 198679
rect 181418 198667 181424 198679
rect 184336 198667 184342 198679
rect 181418 198639 184342 198667
rect 181418 198627 181424 198639
rect 184336 198627 184342 198639
rect 184394 198627 184400 198679
rect 148912 198553 148918 198605
rect 148970 198593 148976 198605
rect 149488 198593 149494 198605
rect 148970 198565 149494 198593
rect 148970 198553 148976 198565
rect 149488 198553 149494 198565
rect 149546 198553 149552 198605
rect 178480 198553 178486 198605
rect 178538 198593 178544 198605
rect 184432 198593 184438 198605
rect 178538 198565 184438 198593
rect 178538 198553 178544 198565
rect 184432 198553 184438 198565
rect 184490 198553 184496 198605
rect 645136 198479 645142 198531
rect 645194 198519 645200 198531
rect 649456 198519 649462 198531
rect 645194 198491 649462 198519
rect 645194 198479 645200 198491
rect 649456 198479 649462 198491
rect 649514 198479 649520 198531
rect 148912 198405 148918 198457
rect 148970 198445 148976 198457
rect 149680 198445 149686 198457
rect 148970 198417 149686 198445
rect 148970 198405 148976 198417
rect 149680 198405 149686 198417
rect 149738 198405 149744 198457
rect 674608 197591 674614 197643
rect 674666 197631 674672 197643
rect 675376 197631 675382 197643
rect 674666 197603 675382 197631
rect 674666 197591 674672 197603
rect 675376 197591 675382 197603
rect 675434 197591 675440 197643
rect 42064 197369 42070 197421
rect 42122 197369 42128 197421
rect 42082 197199 42110 197369
rect 42064 197147 42070 197199
rect 42122 197147 42128 197199
rect 674416 196999 674422 197051
rect 674474 197039 674480 197051
rect 675472 197039 675478 197051
rect 674474 197011 675478 197039
rect 674474 196999 674480 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 42736 196851 42742 196903
rect 42794 196891 42800 196903
rect 43216 196891 43222 196903
rect 42794 196863 43222 196891
rect 42794 196851 42800 196863
rect 43216 196851 43222 196863
rect 43274 196851 43280 196903
rect 674512 196555 674518 196607
rect 674570 196595 674576 196607
rect 675376 196595 675382 196607
rect 674570 196567 675382 196595
rect 674570 196555 674576 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 149296 195889 149302 195941
rect 149354 195929 149360 195941
rect 162736 195929 162742 195941
rect 149354 195901 162742 195929
rect 149354 195889 149360 195901
rect 162736 195889 162742 195901
rect 162794 195889 162800 195941
rect 149680 195815 149686 195867
rect 149738 195855 149744 195867
rect 171280 195855 171286 195867
rect 149738 195827 171286 195855
rect 149738 195815 149744 195827
rect 171280 195815 171286 195827
rect 171338 195815 171344 195867
rect 166960 195741 166966 195793
rect 167018 195781 167024 195793
rect 184528 195781 184534 195793
rect 167018 195753 184534 195781
rect 167018 195741 167024 195753
rect 184528 195741 184534 195753
rect 184586 195741 184592 195793
rect 169840 195667 169846 195719
rect 169898 195707 169904 195719
rect 184432 195707 184438 195719
rect 169898 195679 184438 195707
rect 169898 195667 169904 195679
rect 184432 195667 184438 195679
rect 184490 195667 184496 195719
rect 172720 195593 172726 195645
rect 172778 195633 172784 195645
rect 184336 195633 184342 195645
rect 172778 195605 184342 195633
rect 172778 195593 172784 195605
rect 184336 195593 184342 195605
rect 184394 195593 184400 195645
rect 149392 194631 149398 194683
rect 149450 194671 149456 194683
rect 157072 194671 157078 194683
rect 149450 194643 157078 194671
rect 149450 194631 149456 194643
rect 157072 194631 157078 194643
rect 157130 194631 157136 194683
rect 645136 193965 645142 194017
rect 645194 194005 645200 194017
rect 649360 194005 649366 194017
rect 645194 193977 649366 194005
rect 645194 193965 645200 193977
rect 649360 193965 649366 193977
rect 649418 193965 649424 194017
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 42928 193487 42934 193499
rect 42122 193459 42934 193487
rect 42122 193447 42128 193459
rect 42928 193447 42934 193459
rect 42986 193447 42992 193499
rect 149392 193003 149398 193055
rect 149450 193043 149456 193055
rect 154096 193043 154102 193055
rect 149450 193015 154102 193043
rect 149450 193003 149456 193015
rect 154096 193003 154102 193015
rect 154154 193003 154160 193055
rect 152560 192929 152566 192981
rect 152618 192969 152624 192981
rect 184624 192969 184630 192981
rect 152618 192941 184630 192969
rect 152618 192929 152624 192941
rect 184624 192929 184630 192941
rect 184682 192929 184688 192981
rect 155440 192855 155446 192907
rect 155498 192895 155504 192907
rect 184528 192895 184534 192907
rect 155498 192867 184534 192895
rect 155498 192855 155504 192867
rect 184528 192855 184534 192867
rect 184586 192855 184592 192907
rect 158320 192781 158326 192833
rect 158378 192821 158384 192833
rect 184336 192821 184342 192833
rect 158378 192793 184342 192821
rect 158378 192781 158384 192793
rect 184336 192781 184342 192793
rect 184394 192781 184400 192833
rect 164080 192707 164086 192759
rect 164138 192747 164144 192759
rect 184432 192747 184438 192759
rect 164138 192719 184438 192747
rect 164138 192707 164144 192719
rect 184432 192707 184438 192719
rect 184490 192707 184496 192759
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 42832 192229 42838 192241
rect 42218 192201 42838 192229
rect 42218 192189 42224 192201
rect 42832 192189 42838 192201
rect 42890 192189 42896 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 43120 191489 43126 191501
rect 42122 191461 43126 191489
rect 42122 191449 42128 191461
rect 43120 191449 43126 191461
rect 43178 191449 43184 191501
rect 42160 191005 42166 191057
rect 42218 191045 42224 191057
rect 43024 191045 43030 191057
rect 42218 191017 43030 191045
rect 42218 191005 42224 191017
rect 43024 191005 43030 191017
rect 43082 191005 43088 191057
rect 645136 190413 645142 190465
rect 645194 190453 645200 190465
rect 653776 190453 653782 190465
rect 645194 190425 653782 190453
rect 645194 190413 645200 190425
rect 653776 190413 653782 190425
rect 653834 190413 653840 190465
rect 147568 190191 147574 190243
rect 147626 190231 147632 190243
rect 151792 190231 151798 190243
rect 147626 190203 151798 190231
rect 147626 190191 147632 190203
rect 151792 190191 151798 190203
rect 151850 190191 151856 190243
rect 143152 190043 143158 190095
rect 143210 190083 143216 190095
rect 184624 190083 184630 190095
rect 143210 190055 184630 190083
rect 143210 190043 143216 190055
rect 184624 190043 184630 190055
rect 184682 190043 184688 190095
rect 143248 189969 143254 190021
rect 143306 190009 143312 190021
rect 184528 190009 184534 190021
rect 143306 189981 184534 190009
rect 143306 189969 143312 189981
rect 184528 189969 184534 189981
rect 184586 189969 184592 190021
rect 145360 189895 145366 189947
rect 145418 189935 145424 189947
rect 184432 189935 184438 189947
rect 145418 189907 184438 189935
rect 145418 189895 145424 189907
rect 184432 189895 184438 189907
rect 184490 189895 184496 189947
rect 148912 189821 148918 189873
rect 148970 189861 148976 189873
rect 184336 189861 184342 189873
rect 148970 189833 184342 189861
rect 148970 189821 148976 189833
rect 184336 189821 184342 189833
rect 184394 189821 184400 189873
rect 146896 188785 146902 188837
rect 146954 188825 146960 188837
rect 147280 188825 147286 188837
rect 146954 188797 147286 188825
rect 146954 188785 146960 188797
rect 147280 188785 147286 188797
rect 147338 188785 147344 188837
rect 42160 187823 42166 187875
rect 42218 187863 42224 187875
rect 43216 187863 43222 187875
rect 42218 187835 43222 187863
rect 42218 187823 42224 187835
rect 43216 187823 43222 187835
rect 43274 187823 43280 187875
rect 149392 187231 149398 187283
rect 149450 187271 149456 187283
rect 165616 187271 165622 187283
rect 149450 187243 165622 187271
rect 149450 187231 149456 187243
rect 165616 187231 165622 187243
rect 165674 187231 165680 187283
rect 143152 187157 143158 187209
rect 143210 187197 143216 187209
rect 184432 187197 184438 187209
rect 143210 187169 184438 187197
rect 143210 187157 143216 187169
rect 184432 187157 184438 187169
rect 184490 187157 184496 187209
rect 143344 187083 143350 187135
rect 143402 187123 143408 187135
rect 184624 187123 184630 187135
rect 143402 187095 184630 187123
rect 143402 187083 143408 187095
rect 184624 187083 184630 187095
rect 184682 187083 184688 187135
rect 143248 187009 143254 187061
rect 143306 187049 143312 187061
rect 184336 187049 184342 187061
rect 143306 187021 184342 187049
rect 143306 187009 143312 187021
rect 184336 187009 184342 187021
rect 184394 187009 184400 187061
rect 168496 186935 168502 186987
rect 168554 186975 168560 186987
rect 184528 186975 184534 186987
rect 168554 186947 184534 186975
rect 168554 186935 168560 186947
rect 184528 186935 184534 186947
rect 184586 186935 184592 186987
rect 646192 184567 646198 184619
rect 646250 184607 646256 184619
rect 660880 184607 660886 184619
rect 646250 184579 660886 184607
rect 646250 184567 646256 184579
rect 660880 184567 660886 184579
rect 660938 184567 660944 184619
rect 149392 184345 149398 184397
rect 149450 184385 149456 184397
rect 168688 184385 168694 184397
rect 149450 184357 168694 184385
rect 149450 184345 149456 184357
rect 168688 184345 168694 184357
rect 168746 184345 168752 184397
rect 145648 184271 145654 184323
rect 145706 184311 145712 184323
rect 184528 184311 184534 184323
rect 145706 184283 184534 184311
rect 145706 184271 145712 184283
rect 184528 184271 184534 184283
rect 184586 184271 184592 184323
rect 145552 184197 145558 184249
rect 145610 184237 145616 184249
rect 184336 184237 184342 184249
rect 145610 184209 184342 184237
rect 145610 184197 145616 184209
rect 184336 184197 184342 184209
rect 184394 184197 184400 184249
rect 156880 184123 156886 184175
rect 156938 184163 156944 184175
rect 184624 184163 184630 184175
rect 156938 184135 184630 184163
rect 156938 184123 156944 184135
rect 184624 184123 184630 184135
rect 184682 184123 184688 184175
rect 162640 184049 162646 184101
rect 162698 184089 162704 184101
rect 184432 184089 184438 184101
rect 162698 184061 184438 184089
rect 162698 184049 162704 184061
rect 184432 184049 184438 184061
rect 184490 184049 184496 184101
rect 645904 183087 645910 183139
rect 645962 183127 645968 183139
rect 658288 183127 658294 183139
rect 645962 183099 658294 183127
rect 645962 183087 645968 183099
rect 658288 183087 658294 183099
rect 658346 183087 658352 183139
rect 149392 181459 149398 181511
rect 149450 181499 149456 181511
rect 171376 181499 171382 181511
rect 149450 181471 171382 181499
rect 149450 181459 149456 181471
rect 171376 181459 171382 181471
rect 171434 181459 171440 181511
rect 143056 181385 143062 181437
rect 143114 181425 143120 181437
rect 184624 181425 184630 181437
rect 143114 181397 184630 181425
rect 143114 181385 143120 181397
rect 184624 181385 184630 181397
rect 184682 181385 184688 181437
rect 151120 181311 151126 181363
rect 151178 181351 151184 181363
rect 184528 181351 184534 181363
rect 151178 181323 184534 181351
rect 151178 181311 151184 181323
rect 184528 181311 184534 181323
rect 184586 181311 184592 181363
rect 154000 181237 154006 181289
rect 154058 181277 154064 181289
rect 184336 181277 184342 181289
rect 154058 181249 184342 181277
rect 154058 181237 154064 181249
rect 184336 181237 184342 181249
rect 184394 181237 184400 181289
rect 159760 181163 159766 181215
rect 159818 181203 159824 181215
rect 184432 181203 184438 181215
rect 159818 181175 184438 181203
rect 159818 181163 159824 181175
rect 184432 181163 184438 181175
rect 184490 181163 184496 181215
rect 149392 179535 149398 179587
rect 149450 179575 149456 179587
rect 156880 179575 156886 179587
rect 149450 179547 156886 179575
rect 149450 179535 149456 179547
rect 156880 179535 156886 179547
rect 156938 179535 156944 179587
rect 646000 179387 646006 179439
rect 646058 179427 646064 179439
rect 658480 179427 658486 179439
rect 646058 179399 658486 179427
rect 646058 179387 646064 179399
rect 658480 179387 658486 179399
rect 658538 179387 658544 179439
rect 666640 179313 666646 179365
rect 666698 179353 666704 179365
rect 676048 179353 676054 179365
rect 666698 179325 676054 179353
rect 666698 179313 666704 179325
rect 676048 179313 676054 179325
rect 676106 179313 676112 179365
rect 147376 178795 147382 178847
rect 147434 178835 147440 178847
rect 154192 178835 154198 178847
rect 147434 178807 154198 178835
rect 147434 178795 147440 178807
rect 154192 178795 154198 178807
rect 154250 178795 154256 178847
rect 661456 178795 661462 178847
rect 661514 178835 661520 178847
rect 676048 178835 676054 178847
rect 661514 178807 676054 178835
rect 661514 178795 661520 178807
rect 676048 178795 676054 178807
rect 676106 178795 676112 178847
rect 655312 178647 655318 178699
rect 655370 178687 655376 178699
rect 676240 178687 676246 178699
rect 655370 178659 676246 178687
rect 655370 178647 655376 178659
rect 676240 178647 676246 178659
rect 676298 178647 676304 178699
rect 149680 178573 149686 178625
rect 149738 178613 149744 178625
rect 162640 178613 162646 178625
rect 149738 178585 162646 178613
rect 149738 178573 149744 178585
rect 162640 178573 162646 178585
rect 162698 178573 162704 178625
rect 143056 178499 143062 178551
rect 143114 178539 143120 178551
rect 184432 178539 184438 178551
rect 143114 178511 184438 178539
rect 143114 178499 143120 178511
rect 184432 178499 184438 178511
rect 184490 178499 184496 178551
rect 148912 178425 148918 178477
rect 148970 178465 148976 178477
rect 149680 178465 149686 178477
rect 148970 178437 149686 178465
rect 148970 178425 148976 178437
rect 149680 178425 149686 178437
rect 149738 178425 149744 178477
rect 184528 178465 184534 178477
rect 149890 178437 184534 178465
rect 143056 178351 143062 178403
rect 143114 178351 143120 178403
rect 143074 178243 143102 178351
rect 143152 178277 143158 178329
rect 143210 178317 143216 178329
rect 149890 178317 149918 178437
rect 184528 178425 184534 178437
rect 184586 178425 184592 178477
rect 184336 178391 184342 178403
rect 143210 178289 149918 178317
rect 155506 178363 184342 178391
rect 143210 178277 143216 178289
rect 155506 178243 155534 178363
rect 184336 178351 184342 178363
rect 184394 178351 184400 178403
rect 143074 178215 155534 178243
rect 147184 176723 147190 176775
rect 147242 176763 147248 176775
rect 151120 176763 151126 176775
rect 147242 176735 151126 176763
rect 147242 176723 147248 176735
rect 151120 176723 151126 176735
rect 151178 176723 151184 176775
rect 145456 175613 145462 175665
rect 145514 175653 145520 175665
rect 184336 175653 184342 175665
rect 145514 175625 184342 175653
rect 145514 175613 145520 175625
rect 184336 175613 184342 175625
rect 184394 175613 184400 175665
rect 156976 175539 156982 175591
rect 157034 175579 157040 175591
rect 184432 175579 184438 175591
rect 157034 175551 184438 175579
rect 157034 175539 157040 175551
rect 184432 175539 184438 175551
rect 184490 175539 184496 175591
rect 645136 174873 645142 174925
rect 645194 174913 645200 174925
rect 655216 174913 655222 174925
rect 645194 174885 655222 174913
rect 645194 174873 645200 174885
rect 655216 174873 655222 174885
rect 655274 174873 655280 174925
rect 674512 172875 674518 172927
rect 674570 172915 674576 172927
rect 676048 172915 676054 172927
rect 674570 172887 676054 172915
rect 674570 172875 674576 172887
rect 676048 172875 676054 172887
rect 676106 172875 676112 172927
rect 674800 172801 674806 172853
rect 674858 172841 674864 172853
rect 676240 172841 676246 172853
rect 674858 172813 676246 172841
rect 674858 172801 674864 172813
rect 676240 172801 676246 172813
rect 676298 172801 676304 172853
rect 148240 172727 148246 172779
rect 148298 172767 148304 172779
rect 184432 172767 184438 172779
rect 148298 172739 184438 172767
rect 148298 172727 148304 172739
rect 184432 172727 184438 172739
rect 184490 172727 184496 172779
rect 148720 172653 148726 172705
rect 148778 172693 148784 172705
rect 184528 172693 184534 172705
rect 148778 172665 184534 172693
rect 148778 172653 148784 172665
rect 184528 172653 184534 172665
rect 184586 172653 184592 172705
rect 168400 172579 168406 172631
rect 168458 172619 168464 172631
rect 184336 172619 184342 172631
rect 168458 172591 184342 172619
rect 168458 172579 168464 172591
rect 184336 172579 184342 172591
rect 184394 172579 184400 172631
rect 645136 171395 645142 171447
rect 645194 171435 645200 171447
rect 652336 171435 652342 171447
rect 645194 171407 652342 171435
rect 645194 171395 645200 171407
rect 652336 171395 652342 171407
rect 652394 171395 652400 171447
rect 147280 170359 147286 170411
rect 147338 170399 147344 170411
rect 148240 170399 148246 170411
rect 147338 170371 148246 170399
rect 147338 170359 147344 170371
rect 148240 170359 148246 170371
rect 148298 170359 148304 170411
rect 674608 169989 674614 170041
rect 674666 170029 674672 170041
rect 675952 170029 675958 170041
rect 674666 170001 675958 170029
rect 674666 169989 674672 170001
rect 675952 169989 675958 170001
rect 676010 169989 676016 170041
rect 149392 169915 149398 169967
rect 149450 169955 149456 169967
rect 180112 169955 180118 169967
rect 149450 169927 180118 169955
rect 149450 169915 149456 169927
rect 180112 169915 180118 169927
rect 180170 169915 180176 169967
rect 674704 169915 674710 169967
rect 674762 169955 674768 169967
rect 676048 169955 676054 169967
rect 674762 169927 676054 169955
rect 674762 169915 674768 169927
rect 676048 169915 676054 169927
rect 676106 169915 676112 169967
rect 148528 169841 148534 169893
rect 148586 169881 148592 169893
rect 184432 169881 184438 169893
rect 148586 169853 184438 169881
rect 148586 169841 148592 169853
rect 184432 169841 184438 169853
rect 184490 169841 184496 169893
rect 148336 169767 148342 169819
rect 148394 169807 148400 169819
rect 184528 169807 184534 169819
rect 148394 169779 184534 169807
rect 148394 169767 148400 169779
rect 184528 169767 184534 169779
rect 184586 169767 184592 169819
rect 149008 169693 149014 169745
rect 149066 169733 149072 169745
rect 184624 169733 184630 169745
rect 149066 169705 184630 169733
rect 149066 169693 149072 169705
rect 184624 169693 184630 169705
rect 184682 169693 184688 169745
rect 174160 169619 174166 169671
rect 174218 169659 174224 169671
rect 184336 169659 184342 169671
rect 174218 169631 184342 169659
rect 174218 169619 174224 169631
rect 184336 169619 184342 169631
rect 184394 169619 184400 169671
rect 645136 167991 645142 168043
rect 645194 168031 645200 168043
rect 652816 168031 652822 168043
rect 645194 168003 652822 168031
rect 645194 167991 645200 168003
rect 652816 167991 652822 168003
rect 652874 167991 652880 168043
rect 676240 167365 676246 167377
rect 659506 167337 676246 167365
rect 646672 167251 646678 167303
rect 646730 167291 646736 167303
rect 659506 167291 659534 167337
rect 676240 167325 676246 167337
rect 676298 167325 676304 167377
rect 646730 167263 659534 167291
rect 646730 167251 646736 167263
rect 646864 167177 646870 167229
rect 646922 167217 646928 167229
rect 676240 167217 676246 167229
rect 646922 167189 676246 167217
rect 646922 167177 646928 167189
rect 676240 167177 676246 167189
rect 676298 167177 676304 167229
rect 646768 167103 646774 167155
rect 646826 167143 646832 167155
rect 676144 167143 676150 167155
rect 646826 167115 676150 167143
rect 646826 167103 646832 167115
rect 676144 167103 676150 167115
rect 676202 167103 676208 167155
rect 149392 167029 149398 167081
rect 149450 167069 149456 167081
rect 182992 167069 182998 167081
rect 149450 167041 182998 167069
rect 149450 167029 149456 167041
rect 182992 167029 182998 167041
rect 183050 167029 183056 167081
rect 675184 167029 675190 167081
rect 675242 167069 675248 167081
rect 676048 167069 676054 167081
rect 675242 167041 676054 167069
rect 675242 167029 675248 167041
rect 676048 167029 676054 167041
rect 676106 167029 676112 167081
rect 148432 166955 148438 167007
rect 148490 166995 148496 167007
rect 184432 166995 184438 167007
rect 148490 166967 184438 166995
rect 148490 166955 148496 166967
rect 184432 166955 184438 166967
rect 184490 166955 184496 167007
rect 149200 166881 149206 166933
rect 149258 166921 149264 166933
rect 184528 166921 184534 166933
rect 149258 166893 184534 166921
rect 149258 166881 149264 166893
rect 184528 166881 184534 166893
rect 184586 166881 184592 166933
rect 159856 166807 159862 166859
rect 159914 166847 159920 166859
rect 184336 166847 184342 166859
rect 159914 166819 184342 166847
rect 159914 166807 159920 166819
rect 184336 166807 184342 166819
rect 184394 166807 184400 166859
rect 146992 164439 146998 164491
rect 147050 164439 147056 164491
rect 147010 163961 147038 164439
rect 148624 164069 148630 164121
rect 148682 164109 148688 164121
rect 184336 164109 184342 164121
rect 148682 164081 184342 164109
rect 148682 164069 148688 164081
rect 184336 164069 184342 164081
rect 184394 164069 184400 164121
rect 149296 163995 149302 164047
rect 149354 164035 149360 164047
rect 184528 164035 184534 164047
rect 149354 164007 184534 164035
rect 149354 163995 149360 164007
rect 184528 163995 184534 164007
rect 184586 163995 184592 164047
rect 184432 163961 184438 163973
rect 147010 163933 184438 163961
rect 184432 163921 184438 163933
rect 184490 163921 184496 163973
rect 149008 163847 149014 163899
rect 149066 163887 149072 163899
rect 149296 163887 149302 163899
rect 149066 163859 149302 163887
rect 149066 163847 149072 163859
rect 149296 163847 149302 163859
rect 149354 163847 149360 163899
rect 184336 163887 184342 163899
rect 155506 163859 184342 163887
rect 148240 163699 148246 163751
rect 148298 163739 148304 163751
rect 155506 163739 155534 163859
rect 184336 163847 184342 163859
rect 184394 163847 184400 163899
rect 148298 163711 155534 163739
rect 148298 163699 148304 163711
rect 645520 161775 645526 161827
rect 645578 161815 645584 161827
rect 661072 161815 661078 161827
rect 645578 161787 661078 161815
rect 645578 161775 645584 161787
rect 661072 161775 661078 161787
rect 661130 161775 661136 161827
rect 148144 161183 148150 161235
rect 148202 161223 148208 161235
rect 184624 161223 184630 161235
rect 148202 161195 184630 161223
rect 148202 161183 148208 161195
rect 184624 161183 184630 161195
rect 184682 161183 184688 161235
rect 148816 161109 148822 161161
rect 148874 161149 148880 161161
rect 184336 161149 184342 161161
rect 148874 161121 184342 161149
rect 148874 161109 148880 161121
rect 184336 161109 184342 161121
rect 184394 161109 184400 161161
rect 149104 161035 149110 161087
rect 149162 161075 149168 161087
rect 184432 161075 184438 161087
rect 149162 161047 184438 161075
rect 149162 161035 149168 161047
rect 184432 161035 184438 161047
rect 184490 161035 184496 161087
rect 149584 160961 149590 161013
rect 149642 161001 149648 161013
rect 184528 161001 184534 161013
rect 149642 160973 184534 161001
rect 149642 160961 149648 160973
rect 184528 160961 184534 160973
rect 184586 160961 184592 161013
rect 675376 160961 675382 161013
rect 675434 160961 675440 161013
rect 675664 160961 675670 161013
rect 675722 160961 675728 161013
rect 675394 160791 675422 160961
rect 675376 160739 675382 160791
rect 675434 160739 675440 160791
rect 675682 160051 675710 160961
rect 675664 159999 675670 160051
rect 675722 159999 675728 160051
rect 674512 159407 674518 159459
rect 674570 159447 674576 159459
rect 675376 159447 675382 159459
rect 674570 159419 675382 159447
rect 674570 159407 674576 159419
rect 675376 159407 675382 159419
rect 675434 159407 675440 159459
rect 645520 158445 645526 158497
rect 645578 158485 645584 158497
rect 661168 158485 661174 158497
rect 645578 158457 661174 158485
rect 645578 158445 645584 158457
rect 661168 158445 661174 158457
rect 661226 158445 661232 158497
rect 148048 158371 148054 158423
rect 148106 158411 148112 158423
rect 184432 158411 184438 158423
rect 148106 158383 184438 158411
rect 148106 158371 148112 158383
rect 184432 158371 184438 158383
rect 184490 158371 184496 158423
rect 149488 158297 149494 158349
rect 149546 158337 149552 158349
rect 184528 158337 184534 158349
rect 149546 158309 184534 158337
rect 149546 158297 149552 158309
rect 184528 158297 184534 158309
rect 184586 158297 184592 158349
rect 151504 158223 151510 158275
rect 151562 158263 151568 158275
rect 184624 158263 184630 158275
rect 151562 158235 184630 158263
rect 151562 158223 151568 158235
rect 184624 158223 184630 158235
rect 184682 158223 184688 158275
rect 165520 158149 165526 158201
rect 165578 158189 165584 158201
rect 184336 158189 184342 158201
rect 165578 158161 184342 158189
rect 165578 158149 165584 158161
rect 184336 158149 184342 158161
rect 184394 158149 184400 158201
rect 674800 157705 674806 157757
rect 674858 157745 674864 157757
rect 675472 157745 675478 157757
rect 674858 157717 675478 157745
rect 674858 157705 674864 157717
rect 675472 157705 675478 157717
rect 675530 157705 675536 157757
rect 674704 156891 674710 156943
rect 674762 156931 674768 156943
rect 675472 156931 675478 156943
rect 674762 156903 675478 156931
rect 674762 156891 674768 156903
rect 675472 156891 675478 156903
rect 675530 156891 675536 156943
rect 674608 156299 674614 156351
rect 674666 156339 674672 156351
rect 675376 156339 675382 156351
rect 674666 156311 675382 156339
rect 674666 156299 674672 156311
rect 675376 156299 675382 156311
rect 675434 156299 675440 156351
rect 645136 155855 645142 155907
rect 645194 155895 645200 155907
rect 661264 155895 661270 155907
rect 645194 155867 661270 155895
rect 645194 155855 645200 155867
rect 661264 155855 661270 155867
rect 661322 155855 661328 155907
rect 675184 155855 675190 155907
rect 675242 155895 675248 155907
rect 675376 155895 675382 155907
rect 675242 155867 675382 155895
rect 675242 155855 675248 155867
rect 675376 155855 675382 155867
rect 675434 155855 675440 155907
rect 151408 155411 151414 155463
rect 151466 155451 151472 155463
rect 184432 155451 184438 155463
rect 151466 155423 184438 155451
rect 151466 155411 151472 155423
rect 184432 155411 184438 155423
rect 184490 155411 184496 155463
rect 151696 155337 151702 155389
rect 151754 155377 151760 155389
rect 184528 155377 184534 155389
rect 151754 155349 184534 155377
rect 151754 155337 151760 155349
rect 184528 155337 184534 155349
rect 184586 155337 184592 155389
rect 151216 155263 151222 155315
rect 151274 155303 151280 155315
rect 184336 155303 184342 155315
rect 151274 155275 184342 155303
rect 151274 155263 151280 155275
rect 184336 155263 184342 155275
rect 184394 155263 184400 155315
rect 182800 154893 182806 154945
rect 182858 154933 182864 154945
rect 184720 154933 184726 154945
rect 182858 154905 184726 154933
rect 182858 154893 182864 154905
rect 184720 154893 184726 154905
rect 184778 154893 184784 154945
rect 151312 152599 151318 152651
rect 151370 152639 151376 152651
rect 184336 152639 184342 152651
rect 151370 152611 184342 152639
rect 151370 152599 151376 152611
rect 184336 152599 184342 152611
rect 184394 152599 184400 152651
rect 151600 152525 151606 152577
rect 151658 152565 151664 152577
rect 184432 152565 184438 152577
rect 151658 152537 184438 152565
rect 151658 152525 151664 152537
rect 184432 152525 184438 152537
rect 184490 152525 184496 152577
rect 646000 152525 646006 152577
rect 646058 152565 646064 152577
rect 658576 152565 658582 152577
rect 646058 152537 658582 152565
rect 646058 152525 646064 152537
rect 658576 152525 658582 152537
rect 658634 152525 658640 152577
rect 179920 152451 179926 152503
rect 179978 152491 179984 152503
rect 184528 152491 184534 152503
rect 179978 152463 184534 152491
rect 179978 152451 179984 152463
rect 184528 152451 184534 152463
rect 184586 152451 184592 152503
rect 149200 150157 149206 150209
rect 149258 150197 149264 150209
rect 149680 150197 149686 150209
rect 149258 150169 149686 150197
rect 149258 150157 149264 150169
rect 149680 150157 149686 150169
rect 149738 150157 149744 150209
rect 168592 149713 168598 149765
rect 168650 149753 168656 149765
rect 184432 149753 184438 149765
rect 168650 149725 184438 149753
rect 168650 149713 168656 149725
rect 184432 149713 184438 149725
rect 184490 149713 184496 149765
rect 174256 149639 174262 149691
rect 174314 149679 174320 149691
rect 184336 149679 184342 149691
rect 174314 149651 184342 149679
rect 174314 149639 174320 149651
rect 184336 149639 184342 149651
rect 184394 149639 184400 149691
rect 180016 149565 180022 149617
rect 180074 149605 180080 149617
rect 184528 149605 184534 149617
rect 180074 149577 184534 149605
rect 180074 149565 180080 149577
rect 184528 149565 184534 149577
rect 184586 149565 184592 149617
rect 177040 149491 177046 149543
rect 177098 149531 177104 149543
rect 184624 149531 184630 149543
rect 177098 149503 184630 149531
rect 177098 149491 177104 149503
rect 184624 149491 184630 149503
rect 184682 149491 184688 149543
rect 645136 149343 645142 149395
rect 645194 149383 645200 149395
rect 658672 149383 658678 149395
rect 645194 149355 658678 149383
rect 645194 149343 645200 149355
rect 658672 149343 658678 149355
rect 658730 149343 658736 149395
rect 148048 148011 148054 148063
rect 148106 148051 148112 148063
rect 151696 148051 151702 148063
rect 148106 148023 151702 148051
rect 148106 148011 148112 148023
rect 151696 148011 151702 148023
rect 151754 148011 151760 148063
rect 148048 146975 148054 147027
rect 148106 147015 148112 147027
rect 151216 147015 151222 147027
rect 148106 146987 151222 147015
rect 148106 146975 148112 146987
rect 151216 146975 151222 146987
rect 151274 146975 151280 147027
rect 182896 146827 182902 146879
rect 182954 146867 182960 146879
rect 185776 146867 185782 146879
rect 182954 146839 185782 146867
rect 182954 146827 182960 146839
rect 185776 146827 185782 146839
rect 185834 146827 185840 146879
rect 159952 146753 159958 146805
rect 160010 146793 160016 146805
rect 184432 146793 184438 146805
rect 160010 146765 184438 146793
rect 160010 146753 160016 146765
rect 184432 146753 184438 146765
rect 184490 146753 184496 146805
rect 177136 146679 177142 146731
rect 177194 146719 177200 146731
rect 184528 146719 184534 146731
rect 177194 146691 184534 146719
rect 177194 146679 177200 146691
rect 184528 146679 184534 146691
rect 184586 146679 184592 146731
rect 147952 146605 147958 146657
rect 148010 146645 148016 146657
rect 184336 146645 184342 146657
rect 148010 146617 184342 146645
rect 148010 146605 148016 146617
rect 184336 146605 184342 146617
rect 184394 146605 184400 146657
rect 147952 145791 147958 145843
rect 148010 145831 148016 145843
rect 151600 145831 151606 145843
rect 148010 145803 151606 145831
rect 148010 145791 148016 145803
rect 151600 145791 151606 145803
rect 151658 145791 151664 145843
rect 147952 144311 147958 144363
rect 148010 144351 148016 144363
rect 151312 144351 151318 144363
rect 148010 144323 151318 144351
rect 148010 144311 148016 144323
rect 151312 144311 151318 144323
rect 151370 144311 151376 144363
rect 147856 143941 147862 143993
rect 147914 143981 147920 143993
rect 184432 143981 184438 143993
rect 147914 143953 184438 143981
rect 147914 143941 147920 143953
rect 184432 143941 184438 143953
rect 184490 143941 184496 143993
rect 157072 143867 157078 143919
rect 157130 143907 157136 143919
rect 184624 143907 184630 143919
rect 157130 143879 184630 143907
rect 157130 143867 157136 143879
rect 184624 143867 184630 143879
rect 184682 143867 184688 143919
rect 162736 143793 162742 143845
rect 162794 143833 162800 143845
rect 184528 143833 184534 143845
rect 162794 143805 184534 143833
rect 162794 143793 162800 143805
rect 184528 143793 184534 143805
rect 184586 143793 184592 143845
rect 171280 143719 171286 143771
rect 171338 143759 171344 143771
rect 184336 143759 184342 143771
rect 171338 143731 184342 143759
rect 171338 143719 171344 143731
rect 184336 143719 184342 143731
rect 184394 143719 184400 143771
rect 147856 142535 147862 142587
rect 147914 142575 147920 142587
rect 151888 142575 151894 142587
rect 147914 142547 151894 142575
rect 147914 142535 147920 142547
rect 151888 142535 151894 142547
rect 151946 142535 151952 142587
rect 147856 141499 147862 141551
rect 147914 141539 147920 141551
rect 151504 141539 151510 141551
rect 147914 141511 151510 141539
rect 147914 141499 147920 141511
rect 151504 141499 151510 141511
rect 151562 141499 151568 141551
rect 147664 141203 147670 141255
rect 147722 141243 147728 141255
rect 151408 141243 151414 141255
rect 147722 141215 151414 141243
rect 147722 141203 147728 141215
rect 151408 141203 151414 141215
rect 151466 141203 151472 141255
rect 147952 141055 147958 141107
rect 148010 141095 148016 141107
rect 184528 141095 184534 141107
rect 148010 141067 184534 141095
rect 148010 141055 148016 141067
rect 184528 141055 184534 141067
rect 184586 141055 184592 141107
rect 147472 140981 147478 141033
rect 147530 141021 147536 141033
rect 184624 141021 184630 141033
rect 147530 140993 184630 141021
rect 147530 140981 147536 140993
rect 184624 140981 184630 140993
rect 184682 140981 184688 141033
rect 149200 140907 149206 140959
rect 149258 140947 149264 140959
rect 185680 140947 185686 140959
rect 149258 140919 185686 140947
rect 149258 140907 149264 140919
rect 185680 140907 185686 140919
rect 185738 140907 185744 140959
rect 151792 140833 151798 140885
rect 151850 140873 151856 140885
rect 184432 140873 184438 140885
rect 151850 140845 184438 140873
rect 151850 140833 151856 140845
rect 184432 140833 184438 140845
rect 184490 140833 184496 140885
rect 154096 140759 154102 140811
rect 154154 140799 154160 140811
rect 184336 140799 184342 140811
rect 154154 140771 184342 140799
rect 154154 140759 154160 140771
rect 184336 140759 184342 140771
rect 184394 140759 184400 140811
rect 147856 138169 147862 138221
rect 147914 138209 147920 138221
rect 184528 138209 184534 138221
rect 147914 138181 184534 138209
rect 147914 138169 147920 138181
rect 184528 138169 184534 138181
rect 184586 138169 184592 138221
rect 165616 138095 165622 138147
rect 165674 138135 165680 138147
rect 184336 138135 184342 138147
rect 165674 138107 184342 138135
rect 165674 138095 165680 138107
rect 184336 138095 184342 138107
rect 184394 138095 184400 138147
rect 168688 138021 168694 138073
rect 168746 138061 168752 138073
rect 184432 138061 184438 138073
rect 168746 138033 184438 138061
rect 168746 138021 168752 138033
rect 184432 138021 184438 138033
rect 184490 138021 184496 138073
rect 147568 135283 147574 135335
rect 147626 135323 147632 135335
rect 184432 135323 184438 135335
rect 147626 135295 184438 135323
rect 147626 135283 147632 135295
rect 184432 135283 184438 135295
rect 184490 135283 184496 135335
rect 149488 135209 149494 135261
rect 149546 135249 149552 135261
rect 184336 135249 184342 135261
rect 149546 135221 184342 135249
rect 149546 135209 149552 135221
rect 184336 135209 184342 135221
rect 184394 135209 184400 135261
rect 162640 135135 162646 135187
rect 162698 135175 162704 135187
rect 184528 135175 184534 135187
rect 162698 135147 184534 135175
rect 162698 135135 162704 135147
rect 184528 135135 184534 135147
rect 184586 135135 184592 135187
rect 171376 135061 171382 135113
rect 171434 135101 171440 135113
rect 184336 135101 184342 135113
rect 171434 135073 184342 135101
rect 171434 135061 171440 135073
rect 184336 135061 184342 135073
rect 184394 135061 184400 135113
rect 672400 134321 672406 134373
rect 672458 134361 672464 134373
rect 676240 134361 676246 134373
rect 672458 134333 676246 134361
rect 672458 134321 672464 134333
rect 676240 134321 676246 134333
rect 676298 134321 676304 134373
rect 655408 132767 655414 132819
rect 655466 132807 655472 132819
rect 676240 132807 676246 132819
rect 655466 132779 676246 132807
rect 655466 132767 655472 132779
rect 676240 132767 676246 132779
rect 676298 132767 676304 132819
rect 655120 132619 655126 132671
rect 655178 132659 655184 132671
rect 676144 132659 676150 132671
rect 655178 132631 676150 132659
rect 655178 132619 655184 132631
rect 676144 132619 676150 132631
rect 676202 132619 676208 132671
rect 646576 132471 646582 132523
rect 646634 132511 646640 132523
rect 676048 132511 676054 132523
rect 646634 132483 676054 132511
rect 646634 132471 646640 132483
rect 676048 132471 676054 132483
rect 676106 132471 676112 132523
rect 147184 132397 147190 132449
rect 147242 132437 147248 132449
rect 184624 132437 184630 132449
rect 147242 132409 184630 132437
rect 147242 132397 147248 132409
rect 184624 132397 184630 132409
rect 184682 132397 184688 132449
rect 151120 132323 151126 132375
rect 151178 132363 151184 132375
rect 184528 132363 184534 132375
rect 151178 132335 184534 132363
rect 151178 132323 151184 132335
rect 184528 132323 184534 132335
rect 184586 132323 184592 132375
rect 154192 132249 154198 132301
rect 154250 132289 154256 132301
rect 184432 132289 184438 132301
rect 154250 132261 184438 132289
rect 154250 132249 154256 132261
rect 184432 132249 184438 132261
rect 184490 132249 184496 132301
rect 156880 132175 156886 132227
rect 156938 132215 156944 132227
rect 184336 132215 184342 132227
rect 156938 132187 184342 132215
rect 156938 132175 156944 132187
rect 184336 132175 184342 132187
rect 184394 132175 184400 132227
rect 650992 129807 650998 129859
rect 651050 129847 651056 129859
rect 676048 129847 676054 129859
rect 651050 129819 676054 129847
rect 651050 129807 651056 129819
rect 676048 129807 676054 129819
rect 676106 129807 676112 129859
rect 647728 129659 647734 129711
rect 647786 129699 647792 129711
rect 650992 129699 650998 129711
rect 647786 129671 650998 129699
rect 647786 129659 647792 129671
rect 650992 129659 650998 129671
rect 651050 129659 651056 129711
rect 647920 129585 647926 129637
rect 647978 129625 647984 129637
rect 650896 129625 650902 129637
rect 647978 129597 650902 129625
rect 647978 129585 647984 129597
rect 650896 129585 650902 129597
rect 650954 129625 650960 129637
rect 676240 129625 676246 129637
rect 650954 129597 676246 129625
rect 650954 129585 650960 129597
rect 676240 129585 676246 129597
rect 676298 129585 676304 129637
rect 147088 129511 147094 129563
rect 147146 129551 147152 129563
rect 184336 129551 184342 129563
rect 147146 129523 184342 129551
rect 147146 129511 147152 129523
rect 184336 129511 184342 129523
rect 184394 129511 184400 129563
rect 147376 129437 147382 129489
rect 147434 129477 147440 129489
rect 184432 129477 184438 129489
rect 147434 129449 184438 129477
rect 147434 129437 147440 129449
rect 184432 129437 184438 129449
rect 184490 129437 184496 129489
rect 149296 129363 149302 129415
rect 149354 129403 149360 129415
rect 184528 129403 184534 129415
rect 149354 129375 184534 129403
rect 149354 129363 149360 129375
rect 184528 129363 184534 129375
rect 184586 129363 184592 129415
rect 180112 129289 180118 129341
rect 180170 129329 180176 129341
rect 184720 129329 184726 129341
rect 180170 129301 184726 129329
rect 180170 129289 180176 129301
rect 184720 129289 184726 129301
rect 184778 129289 184784 129341
rect 674512 126699 674518 126751
rect 674570 126739 674576 126751
rect 676048 126739 676054 126751
rect 674570 126711 676054 126739
rect 674570 126699 674576 126711
rect 676048 126699 676054 126711
rect 676106 126699 676112 126751
rect 147280 126625 147286 126677
rect 147338 126665 147344 126677
rect 184336 126665 184342 126677
rect 147338 126637 184342 126665
rect 147338 126625 147344 126637
rect 184336 126625 184342 126637
rect 184394 126625 184400 126677
rect 148912 126551 148918 126603
rect 148970 126591 148976 126603
rect 184432 126591 184438 126603
rect 148970 126563 184438 126591
rect 148970 126551 148976 126563
rect 184432 126551 184438 126563
rect 184490 126551 184496 126603
rect 182992 126477 182998 126529
rect 183050 126517 183056 126529
rect 186832 126517 186838 126529
rect 183050 126489 186838 126517
rect 183050 126477 183056 126489
rect 186832 126477 186838 126489
rect 186890 126477 186896 126529
rect 674224 124701 674230 124753
rect 674282 124741 674288 124753
rect 676048 124741 676054 124753
rect 674282 124713 676054 124741
rect 674282 124701 674288 124713
rect 676048 124701 676054 124713
rect 676106 124701 676112 124753
rect 674416 124035 674422 124087
rect 674474 124075 674480 124087
rect 676240 124075 676246 124087
rect 674474 124047 676246 124075
rect 674474 124035 674480 124047
rect 676240 124035 676246 124047
rect 676298 124035 676304 124087
rect 674032 123961 674038 124013
rect 674090 124001 674096 124013
rect 675952 124001 675958 124013
rect 674090 123973 675958 124001
rect 674090 123961 674096 123973
rect 675952 123961 675958 123973
rect 676010 123961 676016 124013
rect 674128 123887 674134 123939
rect 674186 123927 674192 123939
rect 676048 123927 676054 123939
rect 674186 123899 676054 123927
rect 674186 123887 674192 123899
rect 676048 123887 676054 123899
rect 676106 123887 676112 123939
rect 146896 123813 146902 123865
rect 146954 123853 146960 123865
rect 184624 123853 184630 123865
rect 146954 123825 184630 123853
rect 146954 123813 146960 123825
rect 184624 123813 184630 123825
rect 184682 123813 184688 123865
rect 146992 123739 146998 123791
rect 147050 123779 147056 123791
rect 184432 123779 184438 123791
rect 147050 123751 184438 123779
rect 147050 123739 147056 123751
rect 184432 123739 184438 123751
rect 184490 123739 184496 123791
rect 149488 123665 149494 123717
rect 149546 123705 149552 123717
rect 184528 123705 184534 123717
rect 149546 123677 184534 123705
rect 149546 123665 149552 123677
rect 184528 123665 184534 123677
rect 184586 123665 184592 123717
rect 149680 123591 149686 123643
rect 149738 123631 149744 123643
rect 184336 123631 184342 123643
rect 149738 123603 184342 123631
rect 149738 123591 149744 123603
rect 184336 123591 184342 123603
rect 184394 123591 184400 123643
rect 646672 121223 646678 121275
rect 646730 121263 646736 121275
rect 676336 121263 676342 121275
rect 646730 121235 676342 121263
rect 646730 121223 646736 121235
rect 676336 121223 676342 121235
rect 676394 121223 676400 121275
rect 647920 121149 647926 121201
rect 647978 121189 647984 121201
rect 676144 121189 676150 121201
rect 647978 121161 676150 121189
rect 647978 121149 647984 121161
rect 676144 121149 676150 121161
rect 676202 121149 676208 121201
rect 647824 121075 647830 121127
rect 647882 121115 647888 121127
rect 676240 121115 676246 121127
rect 647882 121087 676246 121115
rect 647882 121075 647888 121087
rect 676240 121075 676246 121087
rect 676298 121075 676304 121127
rect 674608 121001 674614 121053
rect 674666 121041 674672 121053
rect 676048 121041 676054 121053
rect 674666 121013 676054 121041
rect 674666 121001 674672 121013
rect 676048 121001 676054 121013
rect 676106 121001 676112 121053
rect 149104 120927 149110 120979
rect 149162 120967 149168 120979
rect 184528 120967 184534 120979
rect 149162 120939 184534 120967
rect 149162 120927 149168 120939
rect 184528 120927 184534 120939
rect 184586 120927 184592 120979
rect 149584 120853 149590 120905
rect 149642 120893 149648 120905
rect 184624 120893 184630 120905
rect 149642 120865 184630 120893
rect 149642 120853 149648 120865
rect 184624 120853 184630 120865
rect 184682 120853 184688 120905
rect 149008 120779 149014 120831
rect 149066 120819 149072 120831
rect 184336 120819 184342 120831
rect 149066 120791 184342 120819
rect 149066 120779 149072 120791
rect 184336 120779 184342 120791
rect 184394 120779 184400 120831
rect 151696 120705 151702 120757
rect 151754 120745 151760 120757
rect 184432 120745 184438 120757
rect 151754 120717 184438 120745
rect 151754 120705 151760 120717
rect 184432 120705 184438 120717
rect 184490 120705 184496 120757
rect 151312 118041 151318 118093
rect 151370 118081 151376 118093
rect 184624 118081 184630 118093
rect 151370 118053 184630 118081
rect 151370 118041 151376 118053
rect 184624 118041 184630 118053
rect 184682 118041 184688 118093
rect 151216 117967 151222 118019
rect 151274 118007 151280 118019
rect 184336 118007 184342 118019
rect 151274 117979 184342 118007
rect 151274 117967 151280 117979
rect 184336 117967 184342 117979
rect 184394 117967 184400 118019
rect 151600 117893 151606 117945
rect 151658 117933 151664 117945
rect 184432 117933 184438 117945
rect 151658 117905 184438 117933
rect 151658 117893 151664 117905
rect 184432 117893 184438 117905
rect 184490 117893 184496 117945
rect 151888 117819 151894 117871
rect 151946 117859 151952 117871
rect 184528 117859 184534 117871
rect 151946 117831 184534 117859
rect 151946 117819 151952 117831
rect 184528 117819 184534 117831
rect 184586 117819 184592 117871
rect 675472 115747 675478 115799
rect 675530 115747 675536 115799
rect 675490 115577 675518 115747
rect 675472 115525 675478 115577
rect 675530 115525 675536 115577
rect 647920 115229 647926 115281
rect 647978 115269 647984 115281
rect 665200 115269 665206 115281
rect 647978 115241 665206 115269
rect 647978 115229 647984 115241
rect 665200 115229 665206 115241
rect 665258 115229 665264 115281
rect 148336 115155 148342 115207
rect 148394 115195 148400 115207
rect 184528 115195 184534 115207
rect 148394 115167 184534 115195
rect 148394 115155 148400 115167
rect 184528 115155 184534 115167
rect 184586 115155 184592 115207
rect 148816 115081 148822 115133
rect 148874 115121 148880 115133
rect 184624 115121 184630 115133
rect 148874 115093 184630 115121
rect 148874 115081 148880 115093
rect 184624 115081 184630 115093
rect 184682 115081 184688 115133
rect 151408 115007 151414 115059
rect 151466 115047 151472 115059
rect 184432 115047 184438 115059
rect 151466 115019 184438 115047
rect 151466 115007 151472 115019
rect 184432 115007 184438 115019
rect 184490 115007 184496 115059
rect 151504 114933 151510 114985
rect 151562 114973 151568 114985
rect 184336 114973 184342 114985
rect 151562 114945 184342 114973
rect 151562 114933 151568 114945
rect 184336 114933 184342 114945
rect 184394 114933 184400 114985
rect 674512 114785 674518 114837
rect 674570 114825 674576 114837
rect 675376 114825 675382 114837
rect 674570 114797 675382 114825
rect 674570 114785 674576 114797
rect 675376 114785 675382 114797
rect 675434 114785 675440 114837
rect 148240 112269 148246 112321
rect 148298 112309 148304 112321
rect 184432 112309 184438 112321
rect 148298 112281 184438 112309
rect 148298 112269 148304 112281
rect 184432 112269 184438 112281
rect 184490 112269 184496 112321
rect 148624 112195 148630 112247
rect 148682 112235 148688 112247
rect 184528 112235 184534 112247
rect 148682 112207 184534 112235
rect 148682 112195 148688 112207
rect 184528 112195 184534 112207
rect 184586 112195 184592 112247
rect 148432 112121 148438 112173
rect 148490 112161 148496 112173
rect 184336 112161 184342 112173
rect 148490 112133 184342 112161
rect 148490 112121 148496 112133
rect 184336 112121 184342 112133
rect 184394 112121 184400 112173
rect 674416 111677 674422 111729
rect 674474 111717 674480 111729
rect 675376 111717 675382 111729
rect 674474 111689 675382 111717
rect 674474 111677 674480 111689
rect 675376 111677 675382 111689
rect 675434 111677 675440 111729
rect 674224 111159 674230 111211
rect 674282 111199 674288 111211
rect 675376 111199 675382 111211
rect 674282 111171 675382 111199
rect 674282 111159 674288 111171
rect 675376 111159 675382 111171
rect 675434 111159 675440 111211
rect 674128 110641 674134 110693
rect 674186 110681 674192 110693
rect 675376 110681 675382 110693
rect 674186 110653 675382 110681
rect 674186 110641 674192 110653
rect 675376 110641 675382 110653
rect 675434 110641 675440 110693
rect 147952 109383 147958 109435
rect 148010 109423 148016 109435
rect 184528 109423 184534 109435
rect 148010 109395 184534 109423
rect 148010 109383 148016 109395
rect 184528 109383 184534 109395
rect 184586 109383 184592 109435
rect 148720 109309 148726 109361
rect 148778 109349 148784 109361
rect 184432 109349 184438 109361
rect 148778 109321 184438 109349
rect 148778 109309 148784 109321
rect 184432 109309 184438 109321
rect 184490 109309 184496 109361
rect 148528 109235 148534 109287
rect 148586 109275 148592 109287
rect 184336 109275 184342 109287
rect 148586 109247 184342 109275
rect 148586 109235 148592 109247
rect 184336 109235 184342 109247
rect 184394 109235 184400 109287
rect 674032 107311 674038 107363
rect 674090 107351 674096 107363
rect 675376 107351 675382 107363
rect 674090 107323 675382 107351
rect 674090 107311 674096 107323
rect 675376 107311 675382 107323
rect 675434 107311 675440 107363
rect 147664 106497 147670 106549
rect 147722 106537 147728 106549
rect 184624 106537 184630 106549
rect 147722 106509 184630 106537
rect 147722 106497 147728 106509
rect 184624 106497 184630 106509
rect 184682 106497 184688 106549
rect 148048 106423 148054 106475
rect 148106 106463 148112 106475
rect 184432 106463 184438 106475
rect 148106 106435 184438 106463
rect 148106 106423 148112 106435
rect 184432 106423 184438 106435
rect 184490 106423 184496 106475
rect 147856 106349 147862 106401
rect 147914 106389 147920 106401
rect 184528 106389 184534 106401
rect 147914 106361 184534 106389
rect 147914 106349 147920 106361
rect 184528 106349 184534 106361
rect 184586 106349 184592 106401
rect 149392 106275 149398 106327
rect 149450 106315 149456 106327
rect 184336 106315 184342 106327
rect 149450 106287 184342 106315
rect 149450 106275 149456 106287
rect 184336 106275 184342 106287
rect 184394 106275 184400 106327
rect 674608 106127 674614 106179
rect 674666 106167 674672 106179
rect 675376 106167 675382 106179
rect 674666 106139 675382 106167
rect 674666 106127 674672 106139
rect 675376 106127 675382 106139
rect 675434 106127 675440 106179
rect 647920 103907 647926 103959
rect 647978 103947 647984 103959
rect 661168 103947 661174 103959
rect 647978 103919 661174 103947
rect 647978 103907 647984 103919
rect 661168 103907 661174 103919
rect 661226 103907 661232 103959
rect 645904 103685 645910 103737
rect 645962 103725 645968 103737
rect 657520 103725 657526 103737
rect 645962 103697 657526 103725
rect 645962 103685 645968 103697
rect 657520 103685 657526 103697
rect 657578 103685 657584 103737
rect 147568 103611 147574 103663
rect 147626 103651 147632 103663
rect 184528 103651 184534 103663
rect 147626 103623 184534 103651
rect 147626 103611 147632 103623
rect 184528 103611 184534 103623
rect 184586 103611 184592 103663
rect 147088 103537 147094 103589
rect 147146 103577 147152 103589
rect 184624 103577 184630 103589
rect 147146 103549 184630 103577
rect 147146 103537 147152 103549
rect 184624 103537 184630 103549
rect 184682 103537 184688 103589
rect 147760 103463 147766 103515
rect 147818 103503 147824 103515
rect 184432 103503 184438 103515
rect 147818 103475 184438 103503
rect 147818 103463 147824 103475
rect 184432 103463 184438 103475
rect 184490 103463 184496 103515
rect 148144 103389 148150 103441
rect 148202 103429 148208 103441
rect 184336 103429 184342 103441
rect 148202 103401 184342 103429
rect 148202 103389 148208 103401
rect 184336 103389 184342 103401
rect 184394 103389 184400 103441
rect 645136 102057 645142 102109
rect 645194 102097 645200 102109
rect 652432 102097 652438 102109
rect 645194 102069 652438 102097
rect 645194 102057 645200 102069
rect 652432 102057 652438 102069
rect 652490 102057 652496 102109
rect 147184 100725 147190 100777
rect 147242 100765 147248 100777
rect 184432 100765 184438 100777
rect 147242 100737 184438 100765
rect 147242 100725 147248 100737
rect 184432 100725 184438 100737
rect 184490 100725 184496 100777
rect 147280 100651 147286 100703
rect 147338 100691 147344 100703
rect 184528 100691 184534 100703
rect 147338 100663 184534 100691
rect 147338 100651 147344 100663
rect 184528 100651 184534 100663
rect 184586 100651 184592 100703
rect 147376 100577 147382 100629
rect 147434 100617 147440 100629
rect 184624 100617 184630 100629
rect 147434 100589 184630 100617
rect 147434 100577 147440 100589
rect 184624 100577 184630 100589
rect 184682 100577 184688 100629
rect 149776 100503 149782 100555
rect 149834 100543 149840 100555
rect 184336 100543 184342 100555
rect 149834 100515 184342 100543
rect 149834 100503 149840 100515
rect 184336 100503 184342 100515
rect 184394 100503 184400 100555
rect 647920 97913 647926 97965
rect 647978 97953 647984 97965
rect 662512 97953 662518 97965
rect 647978 97925 662518 97953
rect 647978 97913 647984 97925
rect 662512 97913 662518 97925
rect 662570 97913 662576 97965
rect 146992 97839 146998 97891
rect 147050 97879 147056 97891
rect 184528 97879 184534 97891
rect 147050 97851 184534 97879
rect 147050 97839 147056 97851
rect 184528 97839 184534 97851
rect 184586 97839 184592 97891
rect 147472 97765 147478 97817
rect 147530 97805 147536 97817
rect 184336 97805 184342 97817
rect 147530 97777 184342 97805
rect 147530 97765 147536 97777
rect 184336 97765 184342 97777
rect 184394 97765 184400 97817
rect 149296 97691 149302 97743
rect 149354 97731 149360 97743
rect 184432 97731 184438 97743
rect 149354 97703 184438 97731
rect 149354 97691 149360 97703
rect 184432 97691 184438 97703
rect 184490 97691 184496 97743
rect 645424 95915 645430 95967
rect 645482 95955 645488 95967
rect 653680 95955 653686 95967
rect 645482 95927 653686 95955
rect 645482 95915 645488 95927
rect 653680 95915 653686 95927
rect 653738 95915 653744 95967
rect 148912 94953 148918 95005
rect 148970 94993 148976 95005
rect 184528 94993 184534 95005
rect 148970 94965 184534 94993
rect 148970 94953 148976 94965
rect 184528 94953 184534 94965
rect 184586 94953 184592 95005
rect 149200 94879 149206 94931
rect 149258 94919 149264 94931
rect 184336 94919 184342 94931
rect 149258 94891 184342 94919
rect 149258 94879 149264 94891
rect 184336 94879 184342 94891
rect 184394 94879 184400 94931
rect 149104 94805 149110 94857
rect 149162 94845 149168 94857
rect 184432 94845 184438 94857
rect 149162 94817 184438 94845
rect 149162 94805 149168 94817
rect 184432 94805 184438 94817
rect 184490 94805 184496 94857
rect 149584 94731 149590 94783
rect 149642 94771 149648 94783
rect 184336 94771 184342 94783
rect 149642 94743 184342 94771
rect 149642 94731 149648 94743
rect 184336 94731 184342 94743
rect 184394 94731 184400 94783
rect 649552 93547 649558 93599
rect 649610 93587 649616 93599
rect 668176 93587 668182 93599
rect 649610 93559 668182 93587
rect 649610 93547 649616 93559
rect 668176 93547 668182 93559
rect 668234 93547 668240 93599
rect 646768 92659 646774 92711
rect 646826 92699 646832 92711
rect 663088 92699 663094 92711
rect 646826 92671 663094 92699
rect 646826 92659 646832 92671
rect 663088 92659 663094 92671
rect 663146 92659 663152 92711
rect 646480 92363 646486 92415
rect 646538 92403 646544 92415
rect 660688 92403 660694 92415
rect 646538 92375 660694 92403
rect 646538 92363 646544 92375
rect 660688 92363 660694 92375
rect 660746 92363 660752 92415
rect 645520 92289 645526 92341
rect 645578 92329 645584 92341
rect 661744 92329 661750 92341
rect 645578 92301 661750 92329
rect 645578 92289 645584 92301
rect 661744 92289 661750 92301
rect 661802 92289 661808 92341
rect 646864 92215 646870 92267
rect 646922 92255 646928 92267
rect 659824 92255 659830 92267
rect 646922 92227 659830 92255
rect 646922 92215 646928 92227
rect 659824 92215 659830 92227
rect 659882 92215 659888 92267
rect 647152 92141 647158 92193
rect 647210 92181 647216 92193
rect 658864 92181 658870 92193
rect 647210 92153 658870 92181
rect 647210 92141 647216 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 146896 92067 146902 92119
rect 146954 92107 146960 92119
rect 184528 92107 184534 92119
rect 146954 92079 184534 92107
rect 146954 92067 146960 92079
rect 184528 92067 184534 92079
rect 184586 92067 184592 92119
rect 148816 91993 148822 92045
rect 148874 92033 148880 92045
rect 184624 92033 184630 92045
rect 148874 92005 184630 92033
rect 148874 91993 148880 92005
rect 184624 91993 184630 92005
rect 184682 91993 184688 92045
rect 149392 91919 149398 91971
rect 149450 91959 149456 91971
rect 184432 91959 184438 91971
rect 149450 91931 184438 91959
rect 149450 91919 149456 91931
rect 184432 91919 184438 91931
rect 184490 91919 184496 91971
rect 149008 91845 149014 91897
rect 149066 91885 149072 91897
rect 184336 91885 184342 91897
rect 149066 91857 184342 91885
rect 149066 91845 149072 91857
rect 184336 91845 184342 91857
rect 184394 91845 184400 91897
rect 147952 89181 147958 89233
rect 148010 89221 148016 89233
rect 184624 89221 184630 89233
rect 148010 89193 184630 89221
rect 148010 89181 148016 89193
rect 184624 89181 184630 89193
rect 184682 89181 184688 89233
rect 148432 89107 148438 89159
rect 148490 89147 148496 89159
rect 184528 89147 184534 89159
rect 148490 89119 184534 89147
rect 148490 89107 148496 89119
rect 184528 89107 184534 89119
rect 184586 89107 184592 89159
rect 148336 89033 148342 89085
rect 148394 89073 148400 89085
rect 184336 89073 184342 89085
rect 148394 89045 184342 89073
rect 148394 89033 148400 89045
rect 184336 89033 184342 89045
rect 184394 89033 184400 89085
rect 148624 88959 148630 89011
rect 148682 88999 148688 89011
rect 184432 88999 184438 89011
rect 148682 88971 184438 88999
rect 148682 88959 148688 88971
rect 184432 88959 184438 88971
rect 184490 88959 184496 89011
rect 645904 87479 645910 87531
rect 645962 87519 645968 87531
rect 650896 87519 650902 87531
rect 645962 87491 650902 87519
rect 645962 87479 645968 87491
rect 650896 87479 650902 87491
rect 650954 87479 650960 87531
rect 647920 87257 647926 87309
rect 647978 87297 647984 87309
rect 658000 87297 658006 87309
rect 647978 87269 658006 87297
rect 647978 87257 647984 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 647056 87035 647062 87087
rect 647114 87075 647120 87087
rect 663280 87075 663286 87087
rect 647114 87047 663286 87075
rect 647114 87035 647120 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 148048 86369 148054 86421
rect 148106 86409 148112 86421
rect 184336 86409 184342 86421
rect 148106 86381 184342 86409
rect 148106 86369 148112 86381
rect 184336 86369 184342 86381
rect 184394 86369 184400 86421
rect 147664 86295 147670 86347
rect 147722 86335 147728 86347
rect 184432 86335 184438 86347
rect 147722 86307 184438 86335
rect 147722 86295 147728 86307
rect 184432 86295 184438 86307
rect 184490 86295 184496 86347
rect 148528 86221 148534 86273
rect 148586 86261 148592 86273
rect 184528 86261 184534 86273
rect 148586 86233 184534 86261
rect 148586 86221 148592 86233
rect 184528 86221 184534 86233
rect 184586 86221 184592 86273
rect 645904 84149 645910 84201
rect 645962 84189 645968 84201
rect 657040 84189 657046 84201
rect 645962 84161 657046 84189
rect 645962 84149 645968 84161
rect 657040 84149 657046 84161
rect 657098 84149 657104 84201
rect 640720 83631 640726 83683
rect 640778 83671 640784 83683
rect 649552 83671 649558 83683
rect 640778 83643 649558 83671
rect 640778 83631 640784 83643
rect 649552 83631 649558 83643
rect 649610 83631 649616 83683
rect 646768 83557 646774 83609
rect 646826 83597 646832 83609
rect 651760 83597 651766 83609
rect 646826 83569 651766 83597
rect 646826 83557 646832 83569
rect 651760 83557 651766 83569
rect 651818 83557 651824 83609
rect 148240 83483 148246 83535
rect 148298 83523 148304 83535
rect 184528 83523 184534 83535
rect 148298 83495 184534 83523
rect 148298 83483 148304 83495
rect 184528 83483 184534 83495
rect 184586 83483 184592 83535
rect 148720 83409 148726 83461
rect 148778 83449 148784 83461
rect 184624 83449 184630 83461
rect 148778 83421 184630 83449
rect 148778 83409 148784 83421
rect 184624 83409 184630 83421
rect 184682 83409 184688 83461
rect 149680 83335 149686 83387
rect 149738 83375 149744 83387
rect 184336 83375 184342 83387
rect 149738 83347 184342 83375
rect 149738 83335 149744 83347
rect 184336 83335 184342 83347
rect 184394 83335 184400 83387
rect 148144 83261 148150 83313
rect 148202 83301 148208 83313
rect 184432 83301 184438 83313
rect 148202 83273 184438 83301
rect 148202 83261 148208 83273
rect 184432 83261 184438 83273
rect 184490 83261 184496 83313
rect 647920 81855 647926 81907
rect 647978 81895 647984 81907
rect 663280 81895 663286 81907
rect 647978 81867 663286 81895
rect 647978 81855 647984 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 647824 81781 647830 81833
rect 647882 81821 647888 81833
rect 663376 81821 663382 81833
rect 647882 81793 663382 81821
rect 647882 81781 647888 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 657040 81633 657046 81685
rect 657098 81673 657104 81685
rect 658576 81673 658582 81685
rect 657098 81645 658582 81673
rect 657098 81633 657104 81645
rect 658576 81633 658582 81645
rect 658634 81633 658640 81685
rect 647728 81559 647734 81611
rect 647786 81599 647792 81611
rect 662416 81599 662422 81611
rect 647786 81571 662422 81599
rect 647786 81559 647792 81571
rect 662416 81559 662422 81571
rect 662474 81559 662480 81611
rect 647920 80745 647926 80797
rect 647978 80785 647984 80797
rect 662512 80785 662518 80797
rect 647978 80757 662518 80785
rect 647978 80745 647984 80757
rect 662512 80745 662518 80757
rect 662570 80745 662576 80797
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 149200 80597 149206 80649
rect 149258 80637 149264 80649
rect 184624 80637 184630 80649
rect 149258 80609 184630 80637
rect 149258 80597 149264 80609
rect 184624 80597 184630 80609
rect 184682 80597 184688 80649
rect 149488 80523 149494 80575
rect 149546 80563 149552 80575
rect 184336 80563 184342 80575
rect 149546 80535 184342 80563
rect 149546 80523 149552 80535
rect 184336 80523 184342 80535
rect 184394 80523 184400 80575
rect 147568 80449 147574 80501
rect 147626 80489 147632 80501
rect 184432 80489 184438 80501
rect 147626 80461 184438 80489
rect 147626 80449 147632 80461
rect 184432 80449 184438 80461
rect 184490 80449 184496 80501
rect 148912 80375 148918 80427
rect 148970 80415 148976 80427
rect 184528 80415 184534 80427
rect 148970 80387 184534 80415
rect 148970 80375 148976 80387
rect 184528 80375 184534 80387
rect 184586 80375 184592 80427
rect 149008 77711 149014 77763
rect 149066 77751 149072 77763
rect 184432 77751 184438 77763
rect 149066 77723 184438 77751
rect 149066 77711 149072 77723
rect 184432 77711 184438 77723
rect 184490 77711 184496 77763
rect 646960 77711 646966 77763
rect 647018 77751 647024 77763
rect 658288 77751 658294 77763
rect 647018 77723 658294 77751
rect 647018 77711 647024 77723
rect 658288 77711 658294 77723
rect 658346 77711 658352 77763
rect 149104 77637 149110 77689
rect 149162 77677 149168 77689
rect 184528 77677 184534 77689
rect 149162 77649 184534 77677
rect 149162 77637 149168 77649
rect 184528 77637 184534 77649
rect 184586 77637 184592 77689
rect 646576 77637 646582 77689
rect 646634 77677 646640 77689
rect 659440 77677 659446 77689
rect 646634 77649 659446 77677
rect 646634 77637 646640 77649
rect 659440 77637 659446 77649
rect 659498 77637 659504 77689
rect 149392 77563 149398 77615
rect 149450 77603 149456 77615
rect 184624 77603 184630 77615
rect 149450 77575 184630 77603
rect 149450 77563 149456 77575
rect 184624 77563 184630 77575
rect 184682 77563 184688 77615
rect 646672 77563 646678 77615
rect 646730 77603 646736 77615
rect 661744 77603 661750 77615
rect 646730 77575 661750 77603
rect 646730 77563 646736 77575
rect 661744 77563 661750 77575
rect 661802 77563 661808 77615
rect 149296 77489 149302 77541
rect 149354 77529 149360 77541
rect 184336 77529 184342 77541
rect 149354 77501 184342 77529
rect 149354 77489 149360 77501
rect 184336 77489 184342 77501
rect 184394 77489 184400 77541
rect 647920 77489 647926 77541
rect 647978 77529 647984 77541
rect 656944 77529 656950 77541
rect 647978 77501 656950 77529
rect 647978 77489 647984 77501
rect 656944 77489 656950 77501
rect 657002 77489 657008 77541
rect 646000 76083 646006 76135
rect 646058 76123 646064 76135
rect 657520 76123 657526 76135
rect 646058 76095 657526 76123
rect 646058 76083 646064 76095
rect 657520 76083 657526 76095
rect 657578 76083 657584 76135
rect 647056 74899 647062 74951
rect 647114 74939 647120 74951
rect 660112 74939 660118 74951
rect 647114 74911 660118 74939
rect 647114 74899 647120 74911
rect 660112 74899 660118 74911
rect 660170 74899 660176 74951
rect 148816 74825 148822 74877
rect 148874 74865 148880 74877
rect 184336 74865 184342 74877
rect 148874 74837 184342 74865
rect 148874 74825 148880 74837
rect 184336 74825 184342 74837
rect 184394 74825 184400 74877
rect 148336 74751 148342 74803
rect 148394 74791 148400 74803
rect 184432 74791 184438 74803
rect 148394 74763 184438 74791
rect 148394 74751 148400 74763
rect 184432 74751 184438 74763
rect 184490 74751 184496 74803
rect 148528 74677 148534 74729
rect 148586 74717 148592 74729
rect 184528 74717 184534 74729
rect 148586 74689 184534 74717
rect 148586 74677 148592 74689
rect 184528 74677 184534 74689
rect 184586 74677 184592 74729
rect 149584 74603 149590 74655
rect 149642 74643 149648 74655
rect 184624 74643 184630 74655
rect 149642 74615 184630 74643
rect 149642 74603 149648 74615
rect 184624 74603 184630 74615
rect 184682 74603 184688 74655
rect 647920 72087 647926 72139
rect 647978 72127 647984 72139
rect 660688 72127 660694 72139
rect 647978 72099 660694 72127
rect 647978 72087 647984 72099
rect 660688 72087 660694 72099
rect 660746 72087 660752 72139
rect 148432 71939 148438 71991
rect 148490 71979 148496 71991
rect 184336 71979 184342 71991
rect 148490 71951 184342 71979
rect 148490 71939 148496 71951
rect 184336 71939 184342 71951
rect 184394 71939 184400 71991
rect 148720 71865 148726 71917
rect 148778 71905 148784 71917
rect 184432 71905 184438 71917
rect 148778 71877 184438 71905
rect 148778 71865 148784 71877
rect 184432 71865 184438 71877
rect 184490 71865 184496 71917
rect 149680 71791 149686 71843
rect 149738 71831 149744 71843
rect 184528 71831 184534 71843
rect 149738 71803 184534 71831
rect 149738 71791 149744 71803
rect 184528 71791 184534 71803
rect 184586 71791 184592 71843
rect 647920 69571 647926 69623
rect 647978 69611 647984 69623
rect 661456 69611 661462 69623
rect 647978 69583 661462 69611
rect 647978 69571 647984 69583
rect 661456 69571 661462 69583
rect 661514 69571 661520 69623
rect 148624 69053 148630 69105
rect 148682 69093 148688 69105
rect 184336 69093 184342 69105
rect 148682 69065 184342 69093
rect 148682 69053 148688 69065
rect 184336 69053 184342 69065
rect 184394 69053 184400 69105
rect 149488 68979 149494 69031
rect 149546 69019 149552 69031
rect 184528 69019 184534 69031
rect 149546 68991 184534 69019
rect 149546 68979 149552 68991
rect 184528 68979 184534 68991
rect 184586 68979 184592 69031
rect 149104 68905 149110 68957
rect 149162 68945 149168 68957
rect 184336 68945 184342 68957
rect 149162 68917 184342 68945
rect 149162 68905 149168 68917
rect 184336 68905 184342 68917
rect 184394 68905 184400 68957
rect 149584 68831 149590 68883
rect 149642 68871 149648 68883
rect 184432 68871 184438 68883
rect 149642 68843 184438 68871
rect 149642 68831 149648 68843
rect 184432 68831 184438 68843
rect 184490 68831 184496 68883
rect 149392 66167 149398 66219
rect 149450 66207 149456 66219
rect 184624 66207 184630 66219
rect 149450 66179 184630 66207
rect 149450 66167 149456 66179
rect 184624 66167 184630 66179
rect 184682 66167 184688 66219
rect 646000 66167 646006 66219
rect 646058 66207 646064 66219
rect 652336 66207 652342 66219
rect 646058 66179 652342 66207
rect 646058 66167 646064 66179
rect 652336 66167 652342 66179
rect 652394 66167 652400 66219
rect 149200 66093 149206 66145
rect 149258 66133 149264 66145
rect 184528 66133 184534 66145
rect 149258 66105 184534 66133
rect 149258 66093 149264 66105
rect 184528 66093 184534 66105
rect 184586 66093 184592 66145
rect 149008 66019 149014 66071
rect 149066 66059 149072 66071
rect 184336 66059 184342 66071
rect 149066 66031 184342 66059
rect 149066 66019 149072 66031
rect 184336 66019 184342 66031
rect 184394 66019 184400 66071
rect 149296 65945 149302 65997
rect 149354 65985 149360 65997
rect 184432 65985 184438 65997
rect 149354 65957 184438 65985
rect 149354 65945 149360 65957
rect 184432 65945 184438 65957
rect 184490 65945 184496 65997
rect 647920 63577 647926 63629
rect 647978 63617 647984 63629
rect 663184 63617 663190 63629
rect 647978 63589 663190 63617
rect 647978 63577 647984 63589
rect 663184 63577 663190 63589
rect 663242 63577 663248 63629
rect 149680 63281 149686 63333
rect 149738 63321 149744 63333
rect 184624 63321 184630 63333
rect 149738 63293 184630 63321
rect 149738 63281 149744 63293
rect 184624 63281 184630 63293
rect 184682 63281 184688 63333
rect 149488 63207 149494 63259
rect 149546 63247 149552 63259
rect 184432 63247 184438 63259
rect 149546 63219 184438 63247
rect 149546 63207 149552 63219
rect 184432 63207 184438 63219
rect 184490 63207 184496 63259
rect 149584 63133 149590 63185
rect 149642 63173 149648 63185
rect 184336 63173 184342 63185
rect 149642 63145 184342 63173
rect 149642 63133 149648 63145
rect 184336 63133 184342 63145
rect 184394 63133 184400 63185
rect 149392 63059 149398 63111
rect 149450 63099 149456 63111
rect 184528 63099 184534 63111
rect 149450 63071 184534 63099
rect 149450 63059 149456 63071
rect 184528 63059 184534 63071
rect 184586 63059 184592 63111
rect 647920 60987 647926 61039
rect 647978 61027 647984 61039
rect 663472 61027 663478 61039
rect 647978 60999 663478 61027
rect 647978 60987 647984 60999
rect 663472 60987 663478 60999
rect 663530 60987 663536 61039
rect 149392 60395 149398 60447
rect 149450 60435 149456 60447
rect 184432 60435 184438 60447
rect 149450 60407 184438 60435
rect 149450 60395 149456 60407
rect 184432 60395 184438 60407
rect 184490 60395 184496 60447
rect 149488 60321 149494 60373
rect 149546 60361 149552 60373
rect 184528 60361 184534 60373
rect 149546 60333 184534 60361
rect 149546 60321 149552 60333
rect 184528 60321 184534 60333
rect 184586 60321 184592 60373
rect 149296 60247 149302 60299
rect 149354 60287 149360 60299
rect 184336 60287 184342 60299
rect 149354 60259 184342 60287
rect 149354 60247 149360 60259
rect 184336 60247 184342 60259
rect 184394 60247 184400 60299
rect 646000 59063 646006 59115
rect 646058 59103 646064 59115
rect 652240 59103 652246 59115
rect 646058 59075 652246 59103
rect 646058 59063 646064 59075
rect 652240 59063 652246 59075
rect 652298 59063 652304 59115
rect 149392 58989 149398 59041
rect 149450 59029 149456 59041
rect 184336 59029 184342 59041
rect 149450 59001 184342 59029
rect 149450 58989 149456 59001
rect 184336 58989 184342 59001
rect 184394 58989 184400 59041
rect 149392 57509 149398 57561
rect 149450 57549 149456 57561
rect 184336 57549 184342 57561
rect 149450 57521 184342 57549
rect 149450 57509 149456 57521
rect 184336 57509 184342 57521
rect 184394 57509 184400 57561
rect 149392 56177 149398 56229
rect 149450 56217 149456 56229
rect 184432 56217 184438 56229
rect 149450 56189 184438 56217
rect 149450 56177 149456 56189
rect 184432 56177 184438 56189
rect 184490 56177 184496 56229
rect 149488 56103 149494 56155
rect 149546 56143 149552 56155
rect 184336 56143 184342 56155
rect 149546 56115 184342 56143
rect 149546 56103 149552 56115
rect 184336 56103 184342 56115
rect 184394 56103 184400 56155
rect 149680 54623 149686 54675
rect 149738 54663 149744 54675
rect 184336 54663 184342 54675
rect 149738 54635 184342 54663
rect 149738 54623 149744 54635
rect 184336 54623 184342 54635
rect 184394 54623 184400 54675
rect 149392 53217 149398 53269
rect 149450 53257 149456 53269
rect 184336 53257 184342 53269
rect 149450 53229 184342 53257
rect 149450 53217 149456 53229
rect 184336 53217 184342 53229
rect 184394 53217 184400 53269
rect 331216 48037 331222 48089
rect 331274 48077 331280 48089
rect 354832 48077 354838 48089
rect 331274 48049 354838 48077
rect 331274 48037 331280 48049
rect 354832 48037 354838 48049
rect 354890 48037 354896 48089
rect 362032 48037 362038 48089
rect 362090 48077 362096 48089
rect 389200 48077 389206 48089
rect 362090 48049 389206 48077
rect 362090 48037 362096 48049
rect 389200 48037 389206 48049
rect 389258 48037 389264 48089
rect 411856 48037 411862 48089
rect 411914 48077 411920 48089
rect 424048 48077 424054 48089
rect 411914 48049 424054 48077
rect 411914 48037 411920 48049
rect 424048 48037 424054 48049
rect 424106 48037 424112 48089
rect 434896 48037 434902 48089
rect 434954 48077 434960 48089
rect 475696 48077 475702 48089
rect 434954 48049 475702 48077
rect 434954 48037 434960 48049
rect 475696 48037 475702 48049
rect 475754 48037 475760 48089
rect 311056 47963 311062 48015
rect 311114 48003 311120 48015
rect 371920 48003 371926 48015
rect 311114 47975 371926 48003
rect 311114 47963 311120 47975
rect 371920 47963 371926 47975
rect 371978 47963 371984 48015
rect 405520 47963 405526 48015
rect 405578 48003 405584 48015
rect 441328 48003 441334 48015
rect 405578 47975 441334 48003
rect 405578 47963 405584 47975
rect 441328 47963 441334 47975
rect 441386 47963 441392 48015
rect 460336 47963 460342 48015
rect 460394 48003 460400 48015
rect 510352 48003 510358 48015
rect 460394 47975 510358 48003
rect 460394 47963 460400 47975
rect 510352 47963 510358 47975
rect 510410 47963 510416 48015
rect 320176 47889 320182 47941
rect 320234 47929 320240 47941
rect 515536 47929 515542 47941
rect 320234 47901 515542 47929
rect 320234 47889 320240 47901
rect 515536 47889 515542 47901
rect 515594 47889 515600 47941
rect 285808 47815 285814 47867
rect 285866 47855 285872 47867
rect 493936 47855 493942 47867
rect 285866 47827 493942 47855
rect 285866 47815 285872 47827
rect 493936 47815 493942 47827
rect 493994 47815 494000 47867
rect 302896 47741 302902 47793
rect 302954 47781 302960 47793
rect 525904 47781 525910 47793
rect 302954 47753 525910 47781
rect 302954 47741 302960 47753
rect 525904 47741 525910 47753
rect 525962 47741 525968 47793
rect 268528 47667 268534 47719
rect 268586 47707 268592 47719
rect 503920 47707 503926 47719
rect 268586 47679 503926 47707
rect 268586 47667 268592 47679
rect 503920 47667 503926 47679
rect 503978 47667 503984 47719
rect 233680 47593 233686 47645
rect 233738 47633 233744 47645
rect 475600 47633 475606 47645
rect 233738 47605 475606 47633
rect 233738 47593 233744 47605
rect 475600 47593 475606 47605
rect 475658 47593 475664 47645
rect 250960 47519 250966 47571
rect 251018 47559 251024 47571
rect 521200 47559 521206 47571
rect 251018 47531 521206 47559
rect 251018 47519 251024 47531
rect 521200 47519 521206 47531
rect 521258 47519 521264 47571
rect 145360 47075 145366 47127
rect 145418 47115 145424 47127
rect 199120 47115 199126 47127
rect 145418 47087 199126 47115
rect 145418 47075 145424 47087
rect 199120 47075 199126 47087
rect 199178 47075 199184 47127
rect 455056 46927 455062 46979
rect 455114 46967 455120 46979
rect 458608 46967 458614 46979
rect 455114 46939 458614 46967
rect 455114 46927 455120 46939
rect 458608 46927 458614 46939
rect 458666 46927 458672 46979
rect 521488 46335 521494 46387
rect 521546 46375 521552 46387
rect 527920 46375 527926 46387
rect 521546 46347 527926 46375
rect 521546 46335 521552 46347
rect 527920 46335 527926 46347
rect 527978 46335 527984 46387
rect 515536 45077 515542 45129
rect 515594 45117 515600 45129
rect 529264 45117 529270 45129
rect 515594 45089 529270 45117
rect 515594 45077 515600 45089
rect 529264 45077 529270 45089
rect 529322 45077 529328 45129
rect 521488 43267 521494 43279
rect 518386 43239 521494 43267
rect 509776 43153 509782 43205
rect 509834 43193 509840 43205
rect 518386 43193 518414 43239
rect 521488 43227 521494 43239
rect 521546 43227 521552 43279
rect 633616 43227 633622 43279
rect 633674 43267 633680 43279
rect 640720 43267 640726 43279
rect 633674 43239 640726 43267
rect 633674 43227 633680 43239
rect 640720 43227 640726 43239
rect 640778 43227 640784 43279
rect 509834 43165 518414 43193
rect 509834 43153 509840 43165
rect 398896 42339 398902 42391
rect 398954 42379 398960 42391
rect 411856 42379 411862 42391
rect 398954 42351 411862 42379
rect 398954 42339 398960 42351
rect 411856 42339 411862 42351
rect 411914 42339 411920 42391
rect 471664 41747 471670 41799
rect 471722 41787 471728 41799
rect 475504 41787 475510 41799
rect 471722 41759 475510 41787
rect 471722 41747 471728 41759
rect 475504 41747 475510 41759
rect 475562 41747 475568 41799
rect 514000 41747 514006 41799
rect 514058 41787 514064 41799
rect 514864 41787 514870 41799
rect 514058 41759 514870 41787
rect 514058 41747 514064 41759
rect 514864 41747 514870 41759
rect 514922 41747 514928 41799
rect 503920 40267 503926 40319
rect 503978 40307 503984 40319
rect 506800 40307 506806 40319
rect 503978 40279 506806 40307
rect 503978 40267 503984 40279
rect 506800 40267 506806 40279
rect 506858 40267 506864 40319
rect 365902 37381 365908 37433
rect 365960 37421 365966 37433
rect 398896 37421 398902 37433
rect 365960 37393 398902 37421
rect 365960 37381 365966 37393
rect 398896 37381 398902 37393
rect 398954 37381 398960 37433
rect 420688 37381 420694 37433
rect 420746 37421 420752 37433
rect 455056 37421 455062 37433
rect 420746 37393 455062 37421
rect 420746 37381 420752 37393
rect 455056 37381 455062 37393
rect 455114 37381 455120 37433
rect 475504 37381 475510 37433
rect 475562 37421 475568 37433
rect 509776 37421 509782 37433
rect 475562 37393 509782 37421
rect 475562 37381 475568 37393
rect 509776 37381 509782 37393
rect 509834 37381 509840 37433
rect 475600 37307 475606 37359
rect 475658 37347 475664 37359
rect 514000 37347 514006 37359
rect 475658 37319 514006 37347
rect 475658 37307 475664 37319
rect 514000 37307 514006 37319
rect 514058 37307 514064 37359
<< via1 >>
rect 261334 1006411 261386 1006463
rect 276598 1006411 276650 1006463
rect 92854 1006115 92906 1006167
rect 102454 1006115 102506 1006167
rect 356374 1006041 356426 1006093
rect 371638 1006041 371690 1006093
rect 558166 1006041 558218 1006093
rect 574678 1006041 574730 1006093
rect 357910 1005967 357962 1006019
rect 377302 1005967 377354 1006019
rect 358774 1005893 358826 1005945
rect 378838 1005893 378890 1005945
rect 425686 1005893 425738 1005945
rect 471670 1005893 471722 1005945
rect 92566 1005819 92618 1005871
rect 101014 1005819 101066 1005871
rect 262294 1005819 262346 1005871
rect 276502 1005819 276554 1005871
rect 359350 1005819 359402 1005871
rect 380086 1005819 380138 1005871
rect 429718 1005819 429770 1005871
rect 466486 1005819 466538 1005871
rect 551638 1005819 551690 1005871
rect 571606 1005819 571658 1005871
rect 428278 1005745 428330 1005797
rect 460822 1005745 460874 1005797
rect 502294 1005745 502346 1005797
rect 518518 1005745 518570 1005797
rect 553654 1005745 553706 1005797
rect 571318 1005745 571370 1005797
rect 361846 1005671 361898 1005723
rect 383638 1005671 383690 1005723
rect 428662 1005671 428714 1005723
rect 469270 1005671 469322 1005723
rect 501718 1005671 501770 1005723
rect 523990 1005671 524042 1005723
rect 554614 1005671 554666 1005723
rect 573046 1005671 573098 1005723
rect 92950 1005597 93002 1005649
rect 109942 1005597 109994 1005649
rect 358294 1005597 358346 1005649
rect 379990 1005597 380042 1005649
rect 426742 1005597 426794 1005649
rect 472054 1005597 472106 1005649
rect 554038 1005597 554090 1005649
rect 572950 1005597 573002 1005649
rect 94102 1005523 94154 1005575
rect 110518 1005523 110570 1005575
rect 158518 1005523 158570 1005575
rect 172918 1005523 172970 1005575
rect 356758 1005523 356810 1005575
rect 371542 1005523 371594 1005575
rect 425302 1005523 425354 1005575
rect 471862 1005523 471914 1005575
rect 502678 1005523 502730 1005575
rect 92662 1005449 92714 1005501
rect 102070 1005449 102122 1005501
rect 151126 1005449 151178 1005501
rect 161398 1005449 161450 1005501
rect 197206 1005449 197258 1005501
rect 207382 1005449 207434 1005501
rect 357142 1005449 357194 1005501
rect 372022 1005449 372074 1005501
rect 423766 1005449 423818 1005501
rect 471766 1005449 471818 1005501
rect 500758 1005449 500810 1005501
rect 509686 1005449 509738 1005501
rect 518422 1005449 518474 1005501
rect 555190 1005449 555242 1005501
rect 571990 1005449 572042 1005501
rect 152662 1005375 152714 1005427
rect 161878 1005375 161930 1005427
rect 361270 1005375 361322 1005427
rect 374998 1005375 375050 1005427
rect 424726 1005375 424778 1005427
rect 472150 1005375 472202 1005427
rect 503734 1005375 503786 1005427
rect 520534 1005375 520586 1005427
rect 107062 1005301 107114 1005353
rect 124630 1005301 124682 1005353
rect 159478 1005301 159530 1005353
rect 172822 1005301 172874 1005353
rect 210838 1005301 210890 1005353
rect 227350 1005301 227402 1005353
rect 316438 1005301 316490 1005353
rect 331222 1005301 331274 1005353
rect 360886 1005301 360938 1005353
rect 374518 1005301 374570 1005353
rect 424150 1005301 424202 1005353
rect 471958 1005301 472010 1005353
rect 505270 1005301 505322 1005353
rect 520342 1005301 520394 1005353
rect 552598 1005301 552650 1005353
rect 561526 1005301 561578 1005353
rect 161494 1005227 161546 1005279
rect 169942 1005227 169994 1005279
rect 201622 1005227 201674 1005279
rect 212854 1005227 212906 1005279
rect 313846 1005227 313898 1005279
rect 329686 1005227 329738 1005279
rect 362326 1005227 362378 1005279
rect 374614 1005227 374666 1005279
rect 426166 1005227 426218 1005279
rect 472246 1005227 472298 1005279
rect 503254 1005227 503306 1005279
rect 521302 1005227 521354 1005279
rect 552214 1005227 552266 1005279
rect 561046 1005227 561098 1005279
rect 98038 1005153 98090 1005205
rect 105430 1005153 105482 1005205
rect 108022 1005153 108074 1005205
rect 126646 1005153 126698 1005205
rect 160918 1005153 160970 1005205
rect 166964 1005153 167016 1005205
rect 209878 1005153 209930 1005205
rect 225430 1005153 225482 1005205
rect 298486 1005153 298538 1005205
rect 308278 1005153 308330 1005205
rect 312886 1005153 312938 1005205
rect 329782 1005153 329834 1005205
rect 362806 1005153 362858 1005205
rect 374422 1005153 374474 1005205
rect 501142 1005153 501194 1005205
rect 506710 1005153 506762 1005205
rect 509782 1005079 509834 1005131
rect 552982 1005153 553034 1005205
rect 521494 1005079 521546 1005131
rect 564310 1005079 564362 1005131
rect 372022 1005005 372074 1005057
rect 380182 1005005 380234 1005057
rect 371542 1004931 371594 1004983
rect 380374 1004931 380426 1004983
rect 371638 1004857 371690 1004909
rect 380470 1004857 380522 1004909
rect 143830 1004783 143882 1004835
rect 156982 1004783 157034 1004835
rect 520342 1002711 520394 1002763
rect 521590 1002711 521642 1002763
rect 299542 1002637 299594 1002689
rect 306742 1002637 306794 1002689
rect 299734 1002563 299786 1002615
rect 307318 1002563 307370 1002615
rect 300118 1002489 300170 1002541
rect 307894 1002489 307946 1002541
rect 97846 1002415 97898 1002467
rect 103030 1002415 103082 1002467
rect 246934 1002415 246986 1002467
rect 255286 1002415 255338 1002467
rect 299638 1002415 299690 1002467
rect 305302 1002415 305354 1002467
rect 95062 1002341 95114 1002393
rect 101494 1002341 101546 1002393
rect 246550 1002341 246602 1002393
rect 253654 1002341 253706 1002393
rect 300022 1002341 300074 1002393
rect 306358 1002341 306410 1002393
rect 561046 1002341 561098 1002393
rect 564406 1002341 564458 1002393
rect 100534 1002267 100586 1002319
rect 103606 1002267 103658 1002319
rect 143926 1002267 143978 1002319
rect 153046 1002267 153098 1002319
rect 246838 1002267 246890 1002319
rect 254230 1002267 254282 1002319
rect 299830 1002267 299882 1002319
rect 305782 1002267 305834 1002319
rect 505654 1002267 505706 1002319
rect 521398 1002267 521450 1002319
rect 558550 1002267 558602 1002319
rect 567382 1002267 567434 1002319
rect 509686 1002193 509738 1002245
rect 515830 1002193 515882 1002245
rect 374422 1000935 374474 1000987
rect 383446 1000935 383498 1000987
rect 430198 1000935 430250 1000987
rect 472630 1000935 472682 1000987
rect 374998 1000861 375050 1000913
rect 383350 1000861 383402 1000913
rect 429238 1000861 429290 1000913
rect 472534 1000861 472586 1000913
rect 195190 1000787 195242 1000839
rect 208438 1000787 208490 1000839
rect 359734 1000787 359786 1000839
rect 383542 1000787 383594 1000839
rect 427126 1000787 427178 1000839
rect 472630 1000787 472682 1000839
rect 507190 1000787 507242 1000839
rect 517862 1000787 517914 1000839
rect 506230 1000639 506282 1000691
rect 518086 1000639 518138 1000691
rect 298238 1000121 298290 1000173
rect 299638 1000121 299690 1000173
rect 92470 999677 92522 999729
rect 95062 999677 95114 999729
rect 590710 999677 590762 999729
rect 625558 999677 625610 999729
rect 609046 999603 609098 999655
rect 625846 999603 625898 999655
rect 246646 999529 246698 999581
rect 259798 999529 259850 999581
rect 298142 999529 298194 999581
rect 311446 999529 311498 999581
rect 540310 999529 540362 999581
rect 572854 999529 572906 999581
rect 590614 999529 590666 999581
rect 625750 999529 625802 999581
rect 92298 999475 92350 999527
rect 100534 999455 100586 999507
rect 247030 999455 247082 999507
rect 256630 999455 256682 999507
rect 298334 999455 298386 999507
rect 299830 999455 299882 999507
rect 380182 999455 380234 999507
rect 382870 999455 382922 999507
rect 469270 999455 469322 999507
rect 472438 999455 472490 999507
rect 504214 999455 504266 999507
rect 518086 999455 518138 999507
rect 561622 999455 561674 999507
rect 574870 999455 574922 999507
rect 590518 999455 590570 999507
rect 625654 999455 625706 999507
rect 92374 999381 92426 999433
rect 98038 999381 98090 999433
rect 143734 999381 143786 999433
rect 154966 999381 155018 999433
rect 195094 999381 195146 999433
rect 206326 999381 206378 999433
rect 246550 999381 246602 999433
rect 257782 999381 257834 999433
rect 298142 999381 298194 999433
rect 309334 999381 309386 999433
rect 380278 999381 380330 999433
rect 382966 999381 383018 999433
rect 399922 999381 399974 999433
rect 446518 999381 446570 999433
rect 460822 999381 460874 999433
rect 469366 999381 469418 999433
rect 509782 999381 509834 999433
rect 517750 999381 517802 999433
rect 564310 999381 564362 999433
rect 573142 999307 573194 999359
rect 564502 998123 564554 998175
rect 573238 998123 573290 998175
rect 92758 997901 92810 997953
rect 106006 997901 106058 997953
rect 567382 997679 567434 997731
rect 590518 997679 590570 997731
rect 555574 997605 555626 997657
rect 625846 997605 625898 997657
rect 571990 997531 572042 997583
rect 609046 997531 609098 997583
rect 557590 997457 557642 997509
rect 590614 997457 590666 997509
rect 574870 997383 574922 997435
rect 590710 997383 590762 997435
rect 377302 997087 377354 997139
rect 382678 997087 382730 997139
rect 246742 996495 246794 996547
rect 256246 996495 256298 996547
rect 299446 996495 299498 996547
rect 309814 996495 309866 996547
rect 378838 996495 378890 996547
rect 382774 996495 382826 996547
rect 572854 996495 572906 996547
rect 576310 996495 576362 996547
rect 146902 996273 146954 996325
rect 154390 996273 154442 996325
rect 108502 996199 108554 996251
rect 112438 996199 112490 996251
rect 149686 996199 149738 996251
rect 153430 996199 153482 996251
rect 115222 996125 115274 996177
rect 159958 996199 160010 996251
rect 201526 996199 201578 996251
rect 204886 996199 204938 996251
rect 166966 996125 167018 996177
rect 211414 996125 211466 996177
rect 216022 996125 216074 996177
rect 262774 996125 262826 996177
rect 276502 996125 276554 996177
rect 314230 996125 314282 996177
rect 321622 996125 321674 996177
rect 374422 996125 374474 996177
rect 432790 996125 432842 996177
rect 440662 996125 440714 996177
rect 509782 996125 509834 996177
rect 510742 996125 510794 996177
rect 515734 996125 515786 996177
rect 126646 996051 126698 996103
rect 124630 995977 124682 996029
rect 92758 995903 92810 995955
rect 100534 995829 100586 995881
rect 146806 995977 146858 996029
rect 152374 995977 152426 996029
rect 146710 995903 146762 995955
rect 151990 995903 152042 995955
rect 158902 996051 158954 996103
rect 164278 996051 164330 996103
rect 172822 996051 172874 996103
rect 210838 996051 210890 996103
rect 212758 996051 212810 996103
rect 216118 996051 216170 996103
rect 227350 996051 227402 996103
rect 172918 995977 172970 996029
rect 159670 995903 159722 995955
rect 164182 995903 164234 995955
rect 198742 995903 198794 995955
rect 205942 995903 205994 995955
rect 263734 996051 263786 996103
rect 313846 996051 313898 996103
rect 366742 996051 366794 996103
rect 371638 996051 371690 996103
rect 434134 996051 434186 996103
rect 437782 996051 437834 996103
rect 512662 996051 512714 996103
rect 561142 996051 561194 996103
rect 561910 996051 561962 996103
rect 569974 996051 570026 996103
rect 262486 995977 262538 996029
rect 268054 995977 268106 996029
rect 276598 995977 276650 996029
rect 313078 995977 313130 996029
rect 317206 995977 317258 996029
rect 366262 995977 366314 996029
rect 371734 995977 371786 996029
rect 382678 995977 382730 996029
rect 216598 995903 216650 995955
rect 225430 995903 225482 995955
rect 261526 995903 261578 995955
rect 265174 995903 265226 995955
rect 382966 995903 383018 995955
rect 158902 995829 158954 995881
rect 203926 995829 203978 995881
rect 210166 995829 210218 995881
rect 213142 995829 213194 995881
rect 246454 995829 246506 995881
rect 78646 995755 78698 995807
rect 82294 995755 82346 995807
rect 86230 995755 86282 995807
rect 94966 995755 95018 995807
rect 142966 995755 143018 995807
rect 143734 995755 143786 995807
rect 146710 995755 146762 995807
rect 154006 995755 154058 995807
rect 188854 995755 188906 995807
rect 189430 995755 189482 995807
rect 202294 995755 202346 995807
rect 240886 995755 240938 995807
rect 245686 995755 245738 995807
rect 246550 995755 246602 995807
rect 292534 995755 292586 995807
rect 298238 995829 298290 995881
rect 383446 995829 383498 995881
rect 297334 995755 297386 995807
rect 298142 995755 298194 995807
rect 383638 995755 383690 995807
rect 384406 995755 384458 995807
rect 386038 995755 386090 995807
rect 433558 995977 433610 996029
rect 437878 995977 437930 996029
rect 511126 995977 511178 996029
rect 515638 995977 515690 996029
rect 471766 995903 471818 995955
rect 472246 995829 472298 995881
rect 388054 995755 388106 995807
rect 393046 995755 393098 995807
rect 396598 995755 396650 995807
rect 399862 995755 399914 995807
rect 472630 995755 472682 995807
rect 474070 995755 474122 995807
rect 477718 995755 477770 995807
rect 523702 995903 523754 995955
rect 523894 995829 523946 995881
rect 625558 995903 625610 995955
rect 625654 995829 625706 995881
rect 482710 995755 482762 995807
rect 524086 995755 524138 995807
rect 525334 995755 525386 995807
rect 526102 995755 526154 995807
rect 529078 995755 529130 995807
rect 537142 995755 537194 995807
rect 540310 995755 540362 995807
rect 625846 995755 625898 995807
rect 627094 995755 627146 995807
rect 627862 995755 627914 995807
rect 634582 995755 634634 995807
rect 91510 995681 91562 995733
rect 92278 995681 92330 995733
rect 141046 995681 141098 995733
rect 143830 995681 143882 995733
rect 194422 995681 194474 995733
rect 195094 995681 195146 995733
rect 243958 995681 244010 995733
rect 246646 995681 246698 995733
rect 295414 995681 295466 995733
rect 298046 995681 298098 995733
rect 383542 995681 383594 995733
rect 384982 995681 385034 995733
rect 472534 995681 472586 995733
rect 473302 995681 473354 995733
rect 523990 995681 524042 995733
rect 524758 995681 524810 995733
rect 625750 995681 625802 995733
rect 626518 995681 626570 995733
rect 89782 995607 89834 995659
rect 92374 995607 92426 995659
rect 139318 995607 139370 995659
rect 143926 995607 143978 995659
rect 192502 995607 192554 995659
rect 195190 995607 195242 995659
rect 235798 995607 235850 995659
rect 246742 995607 246794 995659
rect 290614 995607 290666 995659
rect 299446 995607 299498 995659
rect 383350 995607 383402 995659
rect 387478 995607 387530 995659
rect 472726 995607 472778 995659
rect 474646 995607 474698 995659
rect 523798 995607 523850 995659
rect 529750 995607 529802 995659
rect 625942 995607 625994 995659
rect 630166 995607 630218 995659
rect 85366 995533 85418 995585
rect 94966 995533 95018 995585
rect 236470 995533 236522 995585
rect 254806 995533 254858 995585
rect 291190 995533 291242 995585
rect 298334 995533 298386 995585
rect 382870 995533 382922 995585
rect 389398 995533 389450 995585
rect 472054 995533 472106 995585
rect 476950 995533 477002 995585
rect 87862 995459 87914 995511
rect 92470 995459 92522 995511
rect 183766 995459 183818 995511
rect 205270 995459 205322 995511
rect 239542 995459 239594 995511
rect 246838 995459 246890 995511
rect 287926 995459 287978 995511
rect 300022 995459 300074 995511
rect 380374 995459 380426 995511
rect 392374 995459 392426 995511
rect 472438 995459 472490 995511
rect 476374 995459 476426 995511
rect 380470 995385 380522 995437
rect 393718 995385 393770 995437
rect 469366 995385 469418 995437
rect 480982 995533 481034 995585
rect 523606 995533 523658 995585
rect 528406 995533 528458 995585
rect 140374 995089 140426 995141
rect 186934 995015 186986 995067
rect 517750 994127 517802 994179
rect 532822 994127 532874 994179
rect 515830 993979 515882 994031
rect 534358 993979 534410 994031
rect 571318 993905 571370 993957
rect 635254 993905 635306 993957
rect 129334 993831 129386 993883
rect 146902 993831 146954 993883
rect 180502 993831 180554 993883
rect 198742 993831 198794 993883
rect 77686 993757 77738 993809
rect 97846 993757 97898 993809
rect 131830 993757 131882 993809
rect 156214 993757 156266 993809
rect 179830 993757 179882 993809
rect 207862 993757 207914 993809
rect 561622 993757 561674 993809
rect 634294 993757 634346 993809
rect 77302 993683 77354 993735
rect 103606 993683 103658 993735
rect 128470 993683 128522 993735
rect 156502 993683 156554 993735
rect 181366 993683 181418 993735
rect 209110 993683 209162 993735
rect 232534 993683 232586 993735
rect 260374 993683 260426 993735
rect 360022 993683 360074 993735
rect 398806 993683 398858 993735
rect 427414 993683 427466 993735
rect 487798 993683 487850 993735
rect 504406 993683 504458 993735
rect 538966 993683 539018 993735
rect 555958 993683 556010 993735
rect 641014 993683 641066 993735
rect 362902 993165 362954 993217
rect 430870 993165 430922 993217
rect 363862 993091 363914 993143
rect 431830 993091 431882 993143
rect 434902 993091 434954 993143
rect 507862 993091 507914 993143
rect 431254 993017 431306 993069
rect 508822 993017 508874 993069
rect 430198 992943 430250 992995
rect 434902 992943 434954 992995
rect 507286 992943 507338 992995
rect 559126 993091 559178 993143
rect 508438 992869 508490 992921
rect 560182 993017 560234 993069
rect 331222 992573 331274 992625
rect 332566 992573 332618 992625
rect 105814 990649 105866 990701
rect 109558 990649 109610 990701
rect 373942 990649 373994 990701
rect 381622 990649 381674 990701
rect 89590 989983 89642 990035
rect 94102 989983 94154 990035
rect 569782 989761 569834 989813
rect 592438 989761 592490 989813
rect 138262 989687 138314 989739
rect 151126 989687 151178 989739
rect 371638 989687 371690 989739
rect 397846 989687 397898 989739
rect 437782 989687 437834 989739
rect 462742 989687 462794 989739
rect 515638 989687 515690 989739
rect 527638 989687 527690 989739
rect 569878 989687 569930 989739
rect 608758 989687 608810 989739
rect 371542 989613 371594 989665
rect 414070 989613 414122 989665
rect 437974 989613 438026 989665
rect 478966 989613 479018 989665
rect 491830 989613 491882 989665
rect 511414 989613 511466 989665
rect 515542 989613 515594 989665
rect 543766 989613 543818 989665
rect 569974 989613 570026 989665
rect 624982 989613 625034 989665
rect 319702 989539 319754 989591
rect 365398 989539 365450 989591
rect 371734 989539 371786 989591
rect 430294 989539 430346 989591
rect 437878 989539 437930 989591
rect 495190 989539 495242 989591
rect 515734 989539 515786 989591
rect 560086 989539 560138 989591
rect 567190 989539 567242 989591
rect 660886 989539 660938 989591
rect 216118 989465 216170 989517
rect 235606 989465 235658 989517
rect 267958 989465 268010 989517
rect 300502 989465 300554 989517
rect 319606 989465 319658 989517
rect 349174 989465 349226 989517
rect 351286 989465 351338 989517
rect 649558 989465 649610 989517
rect 110326 989391 110378 989443
rect 122038 989391 122090 989443
rect 270742 989391 270794 989443
rect 284278 989391 284330 989443
rect 305302 989391 305354 989443
rect 649654 989391 649706 989443
rect 73462 989317 73514 989369
rect 92950 989317 93002 989369
rect 265174 989317 265226 989369
rect 658006 989317 658058 989369
rect 45046 989243 45098 989295
rect 108598 989243 108650 989295
rect 250486 989243 250538 989295
rect 649750 989243 649802 989295
rect 152662 989169 152714 989221
rect 154486 989169 154538 989221
rect 201622 988799 201674 988851
rect 203158 988799 203210 988851
rect 329686 987763 329738 987815
rect 650902 987763 650954 987815
rect 329782 987689 329834 987741
rect 650998 987689 651050 987741
rect 44662 987615 44714 987667
rect 364438 987615 364490 987667
rect 44566 987541 44618 987593
rect 363478 987541 363530 987593
rect 44854 987467 44906 987519
rect 363862 987467 363914 987519
rect 44758 987393 44810 987445
rect 362902 987393 362954 987445
rect 417526 987393 417578 987445
rect 649462 987393 649514 987445
rect 321622 987319 321674 987371
rect 652246 987319 652298 987371
rect 317206 987245 317258 987297
rect 652438 987245 652490 987297
rect 268054 987171 268106 987223
rect 658102 987171 658154 987223
rect 45142 987097 45194 987149
rect 431254 987097 431306 987149
rect 44950 987023 45002 987075
rect 430198 987023 430250 987075
rect 495286 987023 495338 987075
rect 649366 987023 649418 987075
rect 216598 986949 216650 987001
rect 658198 986949 658250 987001
rect 213142 986875 213194 986927
rect 658390 986875 658442 986927
rect 198646 986801 198698 986853
rect 649846 986801 649898 986853
rect 45238 986727 45290 986779
rect 507286 986727 507338 986779
rect 45334 986653 45386 986705
rect 508438 986653 508490 986705
rect 571606 986653 571658 986705
rect 653782 986653 653834 986705
rect 164182 986579 164234 986631
rect 655126 986579 655178 986631
rect 146614 986505 146666 986557
rect 649942 986505 649994 986557
rect 62038 986431 62090 986483
rect 112342 986431 112394 986483
rect 669622 986431 669674 986483
rect 62134 986357 62186 986409
rect 112438 986357 112490 986409
rect 669814 986357 669866 986409
rect 565462 985025 565514 985077
rect 566038 985025 566090 985077
rect 669718 985025 669770 985077
rect 565846 984951 565898 985003
rect 566326 984951 566378 985003
rect 669910 984951 669962 985003
rect 164278 983693 164330 983745
rect 660982 983693 661034 983745
rect 61942 983619 61994 983671
rect 566326 983619 566378 983671
rect 61846 983545 61898 983597
rect 565462 983545 565514 983597
rect 94870 983471 94922 983523
rect 650038 983471 650090 983523
rect 65110 983397 65162 983449
rect 652630 983397 652682 983449
rect 63382 983323 63434 983375
rect 652918 983323 652970 983375
rect 63190 983249 63242 983301
rect 652534 983249 652586 983301
rect 62902 983175 62954 983227
rect 652822 983175 652874 983227
rect 63094 983101 63146 983153
rect 653014 983101 653066 983153
rect 60982 983027 61034 983079
rect 655414 983027 655466 983079
rect 63286 982953 63338 983005
rect 655318 982953 655370 983005
rect 57622 982879 57674 982931
rect 652726 982879 652778 982931
rect 48982 982805 49034 982857
rect 652342 982805 652394 982857
rect 58198 979253 58250 979305
rect 63190 979253 63242 979305
rect 55414 979179 55466 979231
rect 60982 979179 61034 979231
rect 52054 977699 52106 977751
rect 63094 977699 63146 977751
rect 58870 976441 58922 976493
rect 63286 976441 63338 976493
rect 58966 976367 59018 976419
rect 65110 976367 65162 976419
rect 51958 974887 52010 974939
rect 62902 974887 62954 974939
rect 56278 973555 56330 973607
rect 58198 973555 58250 973607
rect 51862 973481 51914 973533
rect 58966 973481 59018 973533
rect 56086 973407 56138 973459
rect 63382 973481 63434 973533
rect 45622 972001 45674 972053
rect 48886 972001 48938 972053
rect 42358 970669 42410 970721
rect 59542 970669 59594 970721
rect 44374 970521 44426 970573
rect 52054 970595 52106 970647
rect 48982 969189 49034 969241
rect 57526 969189 57578 969241
rect 50326 969115 50378 969167
rect 58870 969115 58922 969167
rect 46678 968449 46730 968501
rect 51958 968449 52010 968501
rect 45526 967709 45578 967761
rect 51862 967709 51914 967761
rect 42166 967265 42218 967317
rect 42358 967265 42410 967317
rect 44278 966081 44330 966133
rect 46678 966081 46730 966133
rect 46006 964971 46058 965023
rect 55414 964971 55466 965023
rect 51862 964897 51914 964949
rect 56278 964897 56330 964949
rect 45718 964749 45770 964801
rect 48982 964823 49034 964875
rect 52438 964823 52490 964875
rect 56086 964823 56138 964875
rect 47542 961937 47594 961989
rect 59542 961937 59594 961989
rect 674710 961271 674762 961323
rect 675382 961271 675434 961323
rect 655606 959125 655658 959177
rect 674806 959125 674858 959177
rect 45910 959051 45962 959103
rect 50326 959051 50378 959103
rect 674806 955425 674858 955477
rect 675382 955425 675434 955477
rect 48982 953279 49034 953331
rect 52438 953279 52490 953331
rect 47446 951873 47498 951925
rect 51766 951873 51818 951925
rect 38806 950393 38858 950445
rect 42358 950393 42410 950445
rect 34486 947507 34538 947559
rect 59542 947507 59594 947559
rect 44470 945805 44522 945857
rect 48982 945805 49034 945857
rect 41782 943807 41834 943859
rect 47542 943807 47594 943859
rect 41590 943585 41642 943637
rect 45046 943585 45098 943637
rect 40246 941735 40298 941787
rect 62134 941735 62186 941787
rect 660886 939737 660938 939789
rect 676054 939737 676106 939789
rect 655702 939367 655754 939419
rect 676246 939367 676298 939419
rect 655510 939219 655562 939271
rect 676150 939219 676202 939271
rect 670774 939145 670826 939197
rect 676054 939145 676106 939197
rect 655222 939071 655274 939123
rect 676342 939071 676394 939123
rect 41590 938923 41642 938975
rect 62038 938923 62090 938975
rect 39766 938849 39818 938901
rect 59542 938849 59594 938901
rect 669910 938849 669962 938901
rect 676246 938849 676298 938901
rect 670870 938035 670922 938087
rect 676246 938035 676298 938087
rect 669718 937739 669770 937791
rect 676054 937739 676106 937791
rect 670966 937147 671018 937199
rect 676054 937147 676106 937199
rect 41590 932115 41642 932167
rect 45046 932115 45098 932167
rect 660886 927379 660938 927431
rect 679798 927379 679850 927431
rect 43126 921607 43178 921659
rect 58582 921607 58634 921659
rect 656374 921607 656426 921659
rect 666646 921607 666698 921659
rect 50422 910063 50474 910115
rect 59542 910063 59594 910115
rect 654454 908731 654506 908783
rect 661078 908731 661130 908783
rect 47638 895707 47690 895759
rect 59542 895707 59594 895759
rect 654454 895707 654506 895759
rect 672598 895707 672650 895759
rect 53398 884163 53450 884215
rect 58006 884163 58058 884215
rect 673750 876541 673802 876593
rect 675382 876541 675434 876593
rect 673558 873433 673610 873485
rect 675382 873433 675434 873485
rect 673846 872619 673898 872671
rect 675382 872619 675434 872671
rect 672790 872101 672842 872153
rect 675478 872101 675530 872153
rect 656566 871139 656618 871191
rect 674710 871139 674762 871191
rect 47542 869807 47594 869859
rect 59542 869807 59594 869859
rect 654454 869289 654506 869341
rect 663766 869289 663818 869341
rect 673462 869141 673514 869193
rect 675478 869141 675530 869193
rect 674614 868327 674666 868379
rect 675382 868327 675434 868379
rect 673366 867809 673418 867861
rect 675382 867809 675434 867861
rect 669526 866921 669578 866973
rect 675208 866921 675260 866973
rect 674230 866477 674282 866529
rect 675382 866477 675434 866529
rect 674710 866255 674762 866307
rect 675382 866255 675434 866307
rect 53206 858263 53258 858315
rect 58390 858263 58442 858315
rect 654454 855377 654506 855429
rect 672502 855377 672554 855429
rect 53302 843833 53354 843885
rect 59542 843833 59594 843885
rect 654454 840947 654506 840999
rect 666742 840947 666794 840999
rect 50518 832363 50570 832415
rect 59542 832363 59594 832415
rect 654742 829477 654794 829529
rect 661270 829477 661322 829529
rect 41686 823705 41738 823757
rect 62038 823705 62090 823757
rect 39958 820819 40010 820871
rect 41686 820819 41738 820871
rect 41590 819265 41642 819317
rect 47638 819265 47690 819317
rect 41782 818525 41834 818577
rect 53398 818525 53450 818577
rect 41782 818007 41834 818059
rect 50422 818007 50474 818059
rect 50326 817933 50378 817985
rect 59542 817933 59594 817985
rect 41782 816971 41834 817023
rect 43222 816971 43274 817023
rect 655510 815047 655562 815099
rect 661174 815047 661226 815099
rect 41590 812679 41642 812731
rect 43030 812679 43082 812731
rect 41782 812235 41834 812287
rect 42646 812235 42698 812287
rect 42070 810089 42122 810141
rect 43030 810089 43082 810141
rect 41590 806759 41642 806811
rect 42742 806759 42794 806811
rect 47638 806463 47690 806515
rect 59542 806463 59594 806515
rect 41590 806389 41642 806441
rect 45430 806389 45482 806441
rect 42358 802023 42410 802075
rect 42838 802023 42890 802075
rect 654454 800617 654506 800669
rect 670006 800617 670058 800669
rect 41494 800469 41546 800521
rect 43510 800469 43562 800521
rect 42070 800247 42122 800299
rect 43414 800247 43466 800299
rect 41878 800173 41930 800225
rect 42166 800173 42218 800225
rect 43318 800173 43370 800225
rect 41878 799951 41930 800003
rect 42166 798101 42218 798153
rect 42646 798101 42698 798153
rect 653014 797805 653066 797857
rect 657910 797731 657962 797783
rect 42070 797287 42122 797339
rect 43126 797287 43178 797339
rect 43222 797287 43274 797339
rect 43222 797065 43274 797117
rect 42166 794993 42218 795045
rect 42742 794993 42794 795045
rect 42742 794845 42794 794897
rect 43126 794845 43178 794897
rect 43126 794697 43178 794749
rect 43414 794697 43466 794749
rect 42166 793809 42218 793861
rect 42454 793809 42506 793861
rect 42166 793143 42218 793195
rect 42838 793143 42890 793195
rect 42838 792995 42890 793047
rect 43126 792995 43178 793047
rect 43126 792847 43178 792899
rect 43510 792847 43562 792899
rect 47830 792033 47882 792085
rect 59542 792033 59594 792085
rect 42166 790627 42218 790679
rect 42742 790627 42794 790679
rect 42166 789887 42218 789939
rect 43126 789887 43178 789939
rect 42166 789443 42218 789495
rect 42838 789443 42890 789495
rect 655606 789147 655658 789199
rect 663862 789147 663914 789199
rect 652918 789073 652970 789125
rect 655510 789073 655562 789125
rect 657910 789073 657962 789125
rect 662326 789073 662378 789125
rect 42166 788777 42218 788829
rect 42934 788777 42986 788829
rect 673270 787297 673322 787349
rect 675478 787297 675530 787349
rect 42166 787001 42218 787053
rect 43030 787001 43082 787053
rect 42166 786409 42218 786461
rect 42742 786409 42794 786461
rect 42070 785743 42122 785795
rect 42454 785743 42506 785795
rect 42166 784559 42218 784611
rect 45526 784559 45578 784611
rect 42070 784263 42122 784315
rect 45718 784263 45770 784315
rect 673174 784263 673226 784315
rect 675478 784263 675530 784315
rect 662326 783671 662378 783723
rect 666838 783671 666890 783723
rect 673078 783449 673130 783501
rect 675382 783449 675434 783501
rect 661270 783301 661322 783353
rect 674710 783301 674762 783353
rect 672982 782931 673034 782983
rect 675478 782931 675530 782983
rect 673654 779897 673706 779949
rect 675382 779897 675434 779949
rect 672886 778565 672938 778617
rect 675382 778565 675434 778617
rect 53398 777603 53450 777655
rect 59542 777603 59594 777655
rect 674710 777011 674762 777063
rect 675382 777011 675434 777063
rect 41590 776049 41642 776101
rect 53302 776049 53354 776101
rect 41782 775309 41834 775361
rect 50518 775309 50570 775361
rect 41782 774791 41834 774843
rect 53206 774791 53258 774843
rect 41590 774569 41642 774621
rect 43222 774569 43274 774621
rect 41590 773607 41642 773659
rect 43222 773607 43274 773659
rect 41782 769981 41834 770033
rect 42934 769981 42986 770033
rect 41782 769463 41834 769515
rect 43030 769463 43082 769515
rect 41878 766355 41930 766407
rect 43126 766355 43178 766407
rect 41590 766059 41642 766111
rect 42838 766059 42890 766111
rect 53206 766059 53258 766111
rect 59542 766059 59594 766111
rect 41590 763247 41642 763299
rect 45526 763247 45578 763299
rect 654454 763247 654506 763299
rect 672406 763247 672458 763299
rect 661078 762877 661130 762929
rect 676054 762877 676106 762929
rect 666646 762285 666698 762337
rect 676054 762285 676106 762337
rect 672598 761989 672650 762041
rect 676246 761989 676298 762041
rect 655510 761767 655562 761819
rect 666358 761767 666410 761819
rect 670774 761545 670826 761597
rect 676246 761545 676298 761597
rect 672598 760583 672650 760635
rect 676246 760583 676298 760635
rect 670870 760287 670922 760339
rect 676054 760287 676106 760339
rect 670678 759843 670730 759895
rect 676054 759843 676106 759895
rect 670966 759325 671018 759377
rect 676054 759325 676106 759377
rect 666358 758807 666410 758859
rect 670774 758807 670826 758859
rect 676054 758807 676106 758859
rect 669718 757549 669770 757601
rect 670870 757549 670922 757601
rect 42070 757475 42122 757527
rect 40438 757401 40490 757453
rect 42454 757401 42506 757453
rect 43126 757475 43178 757527
rect 43606 757475 43658 757527
rect 43702 757475 43754 757527
rect 47542 757475 47594 757527
rect 669910 757475 669962 757527
rect 670966 757475 671018 757527
rect 45814 757401 45866 757453
rect 40342 757327 40394 757379
rect 41554 757327 41606 757379
rect 43126 757327 43178 757379
rect 41686 757253 41738 757305
rect 42838 757253 42890 757305
rect 43030 757253 43082 757305
rect 43510 757253 43562 757305
rect 42166 757179 42218 757231
rect 43414 757179 43466 757231
rect 41974 757105 42026 757157
rect 43318 757105 43370 757157
rect 41782 757031 41834 757083
rect 43030 757031 43082 757083
rect 41878 756957 41930 757009
rect 42934 756957 42986 757009
rect 41878 756735 41930 756787
rect 42166 755477 42218 755529
rect 42454 755477 42506 755529
rect 673750 755403 673802 755455
rect 676054 755403 676106 755455
rect 42166 755181 42218 755233
rect 673558 755033 673610 755085
rect 676246 755033 676298 755085
rect 42070 754885 42122 754937
rect 673846 754293 673898 754345
rect 676054 754293 676106 754345
rect 42166 754071 42218 754123
rect 43702 754071 43754 754123
rect 42070 753035 42122 753087
rect 42838 753035 42890 753087
rect 42838 752887 42890 752939
rect 43318 752887 43370 752939
rect 672790 752813 672842 752865
rect 676054 752813 676106 752865
rect 673462 752369 673514 752421
rect 676054 752369 676106 752421
rect 673366 751851 673418 751903
rect 676054 751851 676106 751903
rect 42070 751777 42122 751829
rect 42934 751777 42986 751829
rect 47734 751703 47786 751755
rect 59542 751703 59594 751755
rect 652534 751703 652586 751755
rect 655510 751703 655562 751755
rect 42934 751629 42986 751681
rect 43414 751629 43466 751681
rect 42166 750593 42218 750645
rect 43126 750593 43178 750645
rect 43126 750445 43178 750497
rect 43510 750445 43562 750497
rect 42070 749927 42122 749979
rect 43030 749927 43082 749979
rect 654454 748891 654506 748943
rect 666646 748891 666698 748943
rect 658294 748817 658346 748869
rect 679798 748817 679850 748869
rect 42166 746893 42218 746945
rect 42838 746893 42890 746945
rect 42070 746819 42122 746871
rect 42934 746819 42986 746871
rect 42070 746079 42122 746131
rect 43606 746079 43658 746131
rect 42166 745635 42218 745687
rect 43126 745635 43178 745687
rect 42166 743711 42218 743763
rect 43030 743711 43082 743763
rect 42070 743193 42122 743245
rect 42646 743193 42698 743245
rect 42166 742379 42218 742431
rect 42742 742379 42794 742431
rect 42070 741343 42122 741395
rect 45622 741343 45674 741395
rect 41686 741121 41738 741173
rect 44278 741121 44330 741173
rect 47926 740159 47978 740211
rect 58582 740159 58634 740211
rect 673846 739123 673898 739175
rect 675478 739123 675530 739175
rect 655222 738679 655274 738731
rect 674710 738679 674762 738731
rect 673462 738457 673514 738509
rect 675382 738457 675434 738509
rect 673366 737865 673418 737917
rect 675382 737865 675434 737917
rect 654454 735867 654506 735919
rect 661270 735867 661322 735919
rect 673750 734905 673802 734957
rect 675382 734905 675434 734957
rect 672790 733573 672842 733625
rect 675478 733573 675530 733625
rect 41590 732833 41642 732885
rect 47830 732833 47882 732885
rect 672694 732315 672746 732367
rect 675478 732315 675530 732367
rect 41782 732093 41834 732145
rect 53398 732093 53450 732145
rect 674710 732019 674762 732071
rect 675382 732019 675434 732071
rect 655510 731871 655562 731923
rect 658870 731871 658922 731923
rect 41590 731797 41642 731849
rect 47638 731797 47690 731849
rect 41590 731353 41642 731405
rect 43222 731353 43274 731405
rect 666838 731205 666890 731257
rect 670102 731205 670154 731257
rect 674326 730465 674378 730517
rect 675478 730465 675530 730517
rect 41590 730391 41642 730443
rect 43222 730391 43274 730443
rect 674518 728615 674570 728667
rect 675478 728615 675530 728667
rect 658870 728541 658922 728593
rect 662134 728541 662186 728593
rect 50518 725803 50570 725855
rect 59158 725803 59210 725855
rect 41782 723287 41834 723339
rect 42934 723287 42986 723339
rect 41782 723139 41834 723191
rect 43030 723139 43082 723191
rect 41590 722991 41642 723043
rect 42838 722991 42890 723043
rect 672598 722917 672650 722969
rect 679702 722917 679754 722969
rect 662134 720919 662186 720971
rect 663382 720919 663434 720971
rect 41782 720179 41834 720231
rect 45622 720179 45674 720231
rect 41590 720105 41642 720157
rect 43126 720105 43178 720157
rect 672502 718033 672554 718085
rect 676246 718033 676298 718085
rect 663766 717293 663818 717345
rect 676054 717293 676106 717345
rect 663382 717145 663434 717197
rect 670390 717145 670442 717197
rect 666742 716997 666794 717049
rect 676246 716997 676298 717049
rect 652534 715665 652586 715717
rect 670678 715665 670730 715717
rect 670678 715295 670730 715347
rect 676054 715295 676106 715347
rect 670102 714851 670154 714903
rect 670966 714851 671018 714903
rect 676054 714851 676106 714903
rect 43702 714333 43754 714385
rect 50326 714333 50378 714385
rect 670774 714333 670826 714385
rect 676054 714333 676106 714385
rect 47542 714259 47594 714311
rect 59542 714259 59594 714311
rect 41494 714049 41546 714101
rect 43606 714037 43658 714089
rect 41878 713815 41930 713867
rect 42070 713815 42122 713867
rect 43414 713815 43466 713867
rect 670390 713741 670442 713793
rect 670870 713741 670922 713793
rect 676054 713741 676106 713793
rect 41878 713519 41930 713571
rect 42454 713223 42506 713275
rect 43510 713223 43562 713275
rect 42166 710855 42218 710907
rect 43702 710855 43754 710907
rect 673270 710411 673322 710463
rect 676054 710411 676106 710463
rect 654454 710263 654506 710315
rect 663766 710263 663818 710315
rect 673174 710041 673226 710093
rect 676246 710041 676298 710093
rect 42166 709893 42218 709945
rect 42934 709893 42986 709945
rect 673078 709301 673130 709353
rect 676054 709301 676106 709353
rect 42070 708561 42122 708613
rect 43510 708561 43562 708613
rect 42166 708043 42218 708095
rect 43030 708043 43082 708095
rect 672982 707969 673034 708021
rect 676246 707969 676298 708021
rect 43030 707895 43082 707947
rect 43414 707895 43466 707947
rect 42166 707377 42218 707429
rect 43126 707377 43178 707429
rect 673654 707377 673706 707429
rect 676054 707377 676106 707429
rect 672886 706859 672938 706911
rect 676054 706859 676106 706911
rect 42166 706563 42218 706615
rect 43030 706563 43082 706615
rect 43030 706415 43082 706467
rect 43606 706415 43658 706467
rect 42262 704787 42314 704839
rect 42454 704787 42506 704839
rect 42262 703677 42314 703729
rect 42934 703677 42986 703729
rect 42070 703529 42122 703581
rect 42838 703529 42890 703581
rect 658486 702715 658538 702767
rect 679990 702715 680042 702767
rect 42166 702271 42218 702323
rect 43030 702271 43082 702323
rect 42070 700347 42122 700399
rect 43126 700347 43178 700399
rect 42166 700051 42218 700103
rect 42838 700051 42890 700103
rect 47638 699829 47690 699881
rect 59542 699829 59594 699881
rect 673174 699829 673226 699881
rect 679702 699829 679754 699881
rect 42166 699385 42218 699437
rect 42454 699385 42506 699437
rect 654454 696943 654506 696995
rect 670102 696943 670154 696995
rect 41878 694649 41930 694701
rect 46006 694649 46058 694701
rect 673654 693465 673706 693517
rect 675478 693465 675530 693517
rect 673558 692873 673610 692925
rect 675478 692873 675530 692925
rect 655222 692577 655274 692629
rect 674710 692577 674762 692629
rect 672886 689765 672938 689817
rect 675382 689765 675434 689817
rect 41782 689469 41834 689521
rect 47926 689469 47978 689521
rect 673270 689099 673322 689151
rect 675382 689099 675434 689151
rect 41782 688877 41834 688929
rect 50518 688877 50570 688929
rect 41590 688581 41642 688633
rect 47734 688581 47786 688633
rect 672982 688581 673034 688633
rect 675478 688581 675530 688633
rect 50422 688359 50474 688411
rect 59542 688359 59594 688411
rect 41590 688137 41642 688189
rect 43222 688137 43274 688189
rect 41590 687175 41642 687227
rect 43222 687175 43274 687227
rect 674710 687027 674762 687079
rect 675478 687027 675530 687079
rect 41782 685917 41834 685969
rect 45910 685917 45962 685969
rect 674230 685473 674282 685525
rect 675478 685473 675530 685525
rect 674422 683623 674474 683675
rect 675478 683623 675530 683675
rect 41590 682809 41642 682861
rect 42742 682809 42794 682861
rect 654454 682587 654506 682639
rect 666742 682587 666794 682639
rect 41590 680219 41642 680271
rect 42934 680219 42986 680271
rect 41590 679183 41642 679235
rect 42742 679183 42794 679235
rect 41686 678887 41738 678939
rect 42454 678887 42506 678939
rect 42454 678739 42506 678791
rect 42934 678739 42986 678791
rect 41782 678443 41834 678495
rect 42838 678443 42890 678495
rect 41590 676963 41642 677015
rect 43126 676963 43178 677015
rect 41782 676889 41834 676941
rect 45910 676889 45962 676941
rect 53302 673929 53354 673981
rect 59062 673929 59114 673981
rect 670006 672671 670058 672723
rect 676054 672671 676106 672723
rect 661174 672301 661226 672353
rect 676246 672301 676298 672353
rect 41974 671931 42026 671983
rect 42934 671931 42986 671983
rect 663862 671561 663914 671613
rect 676054 671561 676106 671613
rect 673174 671191 673226 671243
rect 676054 671191 676106 671243
rect 43606 671043 43658 671095
rect 53206 671043 53258 671095
rect 41398 670925 41450 670977
rect 43510 670925 43562 670977
rect 41494 670851 41546 670903
rect 43414 670851 43466 670903
rect 42742 670777 42794 670829
rect 43318 670777 43370 670829
rect 41878 670599 41930 670651
rect 42166 670599 42218 670651
rect 42742 670599 42794 670651
rect 672310 670599 672362 670651
rect 676054 670599 676106 670651
rect 41878 670303 41930 670355
rect 670966 670081 671018 670133
rect 676054 670081 676106 670133
rect 667990 669563 668042 669615
rect 676054 669563 676106 669615
rect 670870 669341 670922 669393
rect 676246 669341 676298 669393
rect 42166 668379 42218 668431
rect 43030 668379 43082 668431
rect 43030 668231 43082 668283
rect 43318 668231 43370 668283
rect 674326 668083 674378 668135
rect 676054 668083 676106 668135
rect 674518 668009 674570 668061
rect 676246 668009 676298 668061
rect 42166 667861 42218 667913
rect 43606 667861 43658 667913
rect 42166 665345 42218 665397
rect 42838 665345 42890 665397
rect 42166 664827 42218 664879
rect 42934 664827 42986 664879
rect 42934 664679 42986 664731
rect 43414 664679 43466 664731
rect 673846 664605 673898 664657
rect 676054 664605 676106 664657
rect 673462 664309 673514 664361
rect 676246 664309 676298 664361
rect 42070 663939 42122 663991
rect 43126 663939 43178 663991
rect 672694 663865 672746 663917
rect 676246 663865 676298 663917
rect 43126 663791 43178 663843
rect 43510 663791 43562 663843
rect 673366 662607 673418 662659
rect 676054 662607 676106 662659
rect 50326 662385 50378 662437
rect 58102 662385 58154 662437
rect 655414 662311 655466 662363
rect 659062 662311 659114 662363
rect 673750 662237 673802 662289
rect 676054 662237 676106 662289
rect 672790 661645 672842 661697
rect 676054 661645 676106 661697
rect 42070 661053 42122 661105
rect 43030 661053 43082 661105
rect 42070 660387 42122 660439
rect 42838 660387 42890 660439
rect 42166 659869 42218 659921
rect 42742 659869 42794 659921
rect 42742 659721 42794 659773
rect 42934 659721 42986 659773
rect 42934 659573 42986 659625
rect 43126 659573 43178 659625
rect 655222 659499 655274 659551
rect 679798 659499 679850 659551
rect 42070 659055 42122 659107
rect 42934 659055 42986 659107
rect 42070 657205 42122 657257
rect 42838 657205 42890 657257
rect 42166 656687 42218 656739
rect 42934 656687 42986 656739
rect 654454 656687 654506 656739
rect 661078 656687 661130 656739
rect 672502 656687 672554 656739
rect 679894 656687 679946 656739
rect 42166 656169 42218 656221
rect 43030 656169 43082 656221
rect 659062 653801 659114 653853
rect 665014 653727 665066 653779
rect 673750 652099 673802 652151
rect 675478 652099 675530 652151
rect 673078 649065 673130 649117
rect 675478 649065 675530 649117
rect 673174 648251 673226 648303
rect 675382 648251 675434 648303
rect 53206 648029 53258 648081
rect 59542 648029 59594 648081
rect 673846 647881 673898 647933
rect 675478 647881 675530 647933
rect 655510 646549 655562 646601
rect 674710 646549 674762 646601
rect 41782 646253 41834 646305
rect 50422 646253 50474 646305
rect 41782 645735 41834 645787
rect 53302 645735 53354 645787
rect 41590 645365 41642 645417
rect 47638 645365 47690 645417
rect 41782 644773 41834 644825
rect 43222 644773 43274 644825
rect 672790 644773 672842 644825
rect 675382 644773 675434 644825
rect 673462 643959 673514 644011
rect 675478 643959 675530 644011
rect 672694 643367 672746 643419
rect 675382 643367 675434 643419
rect 654454 642257 654506 642309
rect 672598 642257 672650 642309
rect 673366 642257 673418 642309
rect 675478 642257 675530 642309
rect 674710 641813 674762 641865
rect 675382 641813 675434 641865
rect 665014 640407 665066 640459
rect 668086 640407 668138 640459
rect 41782 639519 41834 639571
rect 43126 639519 43178 639571
rect 41686 637003 41738 637055
rect 43030 637003 43082 637055
rect 47734 636485 47786 636537
rect 59542 636485 59594 636537
rect 672310 635597 672362 635649
rect 679702 635597 679754 635649
rect 41686 634931 41738 634983
rect 42838 634931 42890 634983
rect 41686 633895 41738 633947
rect 46006 633895 46058 633947
rect 42934 629677 42986 629729
rect 43414 629677 43466 629729
rect 25846 629233 25898 629285
rect 43702 629233 43754 629285
rect 42838 627827 42890 627879
rect 47542 627827 47594 627879
rect 654454 627827 654506 627879
rect 663958 627827 664010 627879
rect 655318 627753 655370 627805
rect 665206 627753 665258 627805
rect 668086 627753 668138 627805
rect 670870 627753 670922 627805
rect 43030 627679 43082 627731
rect 43510 627679 43562 627731
rect 666646 627679 666698 627731
rect 676054 627679 676106 627731
rect 42070 627531 42122 627583
rect 43126 627531 43178 627583
rect 41974 627457 42026 627509
rect 43030 627457 43082 627509
rect 41782 627383 41834 627435
rect 41878 627383 41930 627435
rect 42934 627383 42986 627435
rect 672406 627309 672458 627361
rect 676246 627309 676298 627361
rect 41782 627013 41834 627065
rect 661270 626569 661322 626621
rect 676054 626569 676106 626621
rect 672022 625607 672074 625659
rect 676054 625607 676106 625659
rect 42166 625311 42218 625363
rect 43222 625311 43274 625363
rect 674230 624867 674282 624919
rect 676054 624867 676106 624919
rect 42166 624645 42218 624697
rect 42838 624645 42890 624697
rect 670870 624645 670922 624697
rect 675958 624645 676010 624697
rect 42838 624497 42890 624549
rect 43414 624497 43466 624549
rect 665206 623535 665258 623587
rect 670966 623535 671018 623587
rect 675958 623535 676010 623587
rect 42166 623461 42218 623513
rect 43510 623461 43562 623513
rect 47542 622055 47594 622107
rect 59542 622055 59594 622107
rect 674422 621981 674474 622033
rect 676246 621981 676298 622033
rect 42166 621611 42218 621663
rect 42838 621611 42890 621663
rect 42166 620353 42218 620405
rect 42934 620353 42986 620405
rect 673654 619169 673706 619221
rect 676054 619169 676106 619221
rect 42262 619021 42314 619073
rect 43030 619021 43082 619073
rect 673270 618133 673322 618185
rect 676054 618133 676106 618185
rect 42070 617837 42122 617889
rect 43126 617837 43178 617889
rect 673558 617615 673610 617667
rect 676054 617615 676106 617667
rect 672886 617393 672938 617445
rect 676246 617393 676298 617445
rect 42262 616653 42314 616705
rect 42934 616653 42986 616705
rect 672982 616653 673034 616705
rect 676054 616653 676106 616705
rect 652342 616357 652394 616409
rect 655318 616357 655370 616409
rect 653878 614507 653930 614559
rect 661174 614507 661226 614559
rect 42166 614137 42218 614189
rect 42838 614137 42890 614189
rect 42166 613619 42218 613671
rect 42934 613619 42986 613671
rect 652342 613471 652394 613523
rect 679798 613471 679850 613523
rect 42070 612805 42122 612857
rect 43030 612805 43082 612857
rect 47638 610585 47690 610637
rect 59254 610585 59306 610637
rect 660598 607921 660650 607973
rect 666838 607921 666890 607973
rect 652918 607699 652970 607751
rect 653878 607699 653930 607751
rect 672214 607033 672266 607085
rect 675478 607033 675530 607085
rect 673558 603925 673610 603977
rect 675478 603925 675530 603977
rect 654550 603333 654602 603385
rect 674614 603333 674666 603385
rect 673270 603259 673322 603311
rect 675382 603259 675434 603311
rect 41782 603037 41834 603089
rect 47734 603037 47786 603089
rect 41590 602741 41642 602793
rect 47542 602741 47594 602793
rect 672310 602667 672362 602719
rect 675382 602667 675434 602719
rect 41590 602149 41642 602201
rect 53206 602149 53258 602201
rect 653014 602001 653066 602053
rect 660598 602001 660650 602053
rect 654454 601927 654506 601979
rect 672502 601927 672554 601979
rect 41782 601557 41834 601609
rect 43510 601557 43562 601609
rect 41782 600965 41834 601017
rect 43222 600965 43274 601017
rect 41590 599855 41642 599907
rect 43318 599855 43370 599907
rect 44374 599855 44426 599907
rect 672118 599781 672170 599833
rect 675382 599781 675434 599833
rect 672886 599263 672938 599315
rect 675382 599263 675434 599315
rect 41782 598967 41834 599019
rect 43510 598967 43562 599019
rect 672982 598375 673034 598427
rect 675478 598375 675530 598427
rect 41590 597709 41642 597761
rect 42934 597709 42986 597761
rect 672406 597117 672458 597169
rect 675478 597117 675530 597169
rect 674614 596821 674666 596873
rect 675382 596821 675434 596873
rect 43510 596155 43562 596207
rect 47542 596155 47594 596207
rect 53206 596155 53258 596207
rect 59350 596155 59402 596207
rect 41782 593935 41834 593987
rect 42742 593935 42794 593987
rect 41782 593491 41834 593543
rect 43126 593491 43178 593543
rect 41782 592529 41834 592581
rect 43030 592529 43082 592581
rect 41782 591197 41834 591249
rect 42838 591197 42890 591249
rect 41590 590679 41642 590731
rect 47446 590679 47498 590731
rect 654454 590383 654506 590435
rect 666838 590383 666890 590435
rect 655318 588607 655370 588659
rect 658870 588607 658922 588659
rect 658870 586017 658922 586069
rect 668086 586017 668138 586069
rect 43510 584685 43562 584737
rect 50326 584685 50378 584737
rect 50422 584685 50474 584737
rect 59542 584685 59594 584737
rect 41782 584315 41834 584367
rect 43702 584315 43754 584367
rect 41974 584241 42026 584293
rect 43798 584241 43850 584293
rect 41878 584167 41930 584219
rect 42166 584167 42218 584219
rect 43414 584167 43466 584219
rect 41878 583945 41930 583997
rect 42454 583649 42506 583701
rect 43318 583649 43370 583701
rect 670102 582465 670154 582517
rect 676054 582465 676106 582517
rect 42166 582095 42218 582147
rect 42934 582095 42986 582147
rect 652822 581947 652874 581999
rect 43030 581873 43082 581925
rect 43318 581873 43370 581925
rect 663766 581947 663818 581999
rect 676054 581947 676106 581999
rect 668086 581799 668138 581851
rect 670774 581799 670826 581851
rect 665878 581725 665930 581777
rect 666742 581577 666794 581629
rect 676246 581577 676298 581629
rect 42070 581355 42122 581407
rect 43510 581355 43562 581407
rect 672022 580985 672074 581037
rect 676054 580985 676106 581037
rect 42070 580245 42122 580297
rect 42742 580245 42794 580297
rect 670582 580171 670634 580223
rect 676246 580171 676298 580223
rect 42742 580097 42794 580149
rect 43126 580097 43178 580149
rect 670870 579949 670922 580001
rect 676054 579949 676106 580001
rect 43030 579801 43082 579853
rect 43414 579801 43466 579853
rect 670774 579431 670826 579483
rect 676054 579431 676106 579483
rect 42166 578987 42218 579039
rect 42838 578987 42890 579039
rect 670966 578913 671018 578965
rect 676054 578913 676106 578965
rect 665878 578395 665930 578447
rect 670678 578395 670730 578447
rect 676054 578395 676106 578447
rect 42070 578247 42122 578299
rect 42742 578247 42794 578299
rect 42166 577655 42218 577707
rect 42934 577655 42986 577707
rect 654454 577285 654506 577337
rect 661174 577285 661226 577337
rect 42166 577137 42218 577189
rect 43510 577137 43562 577189
rect 673750 574991 673802 575043
rect 676054 574991 676106 575043
rect 42166 574621 42218 574673
rect 43126 574621 43178 574673
rect 673078 574621 673130 574673
rect 676246 574621 676298 574673
rect 42166 574103 42218 574155
rect 43030 574103 43082 574155
rect 673174 573881 673226 573933
rect 676054 573881 676106 573933
rect 673366 573511 673418 573563
rect 676054 573511 676106 573563
rect 42166 573437 42218 573489
rect 43606 573437 43658 573489
rect 673462 572993 673514 573045
rect 676054 572993 676106 573045
rect 42166 572771 42218 572823
rect 42838 572771 42890 572823
rect 673846 572401 673898 572453
rect 676054 572401 676106 572453
rect 672790 571957 672842 572009
rect 676054 571957 676106 572009
rect 672694 571661 672746 571713
rect 676246 571661 676298 571713
rect 42166 570847 42218 570899
rect 42934 570847 42986 570899
rect 42166 570403 42218 570455
rect 42358 570403 42410 570455
rect 42358 570255 42410 570307
rect 59542 570255 59594 570307
rect 42070 569663 42122 569715
rect 42742 569663 42794 569715
rect 652822 567369 652874 567421
rect 679990 567369 680042 567421
rect 41782 559821 41834 559873
rect 50422 559821 50474 559873
rect 652726 559821 652778 559873
rect 663766 559821 663818 559873
rect 674614 559377 674666 559429
rect 675382 559377 675434 559429
rect 674518 558933 674570 558985
rect 675478 558933 675530 558985
rect 41782 558785 41834 558837
rect 53206 558785 53258 558837
rect 50326 558711 50378 558763
rect 59542 558711 59594 558763
rect 41782 558341 41834 558393
rect 43222 558341 43274 558393
rect 673846 558045 673898 558097
rect 675382 558045 675434 558097
rect 41782 557823 41834 557875
rect 43606 557823 43658 557875
rect 656566 557231 656618 557283
rect 675286 557231 675338 557283
rect 674710 555233 674762 555285
rect 675478 555233 675530 555285
rect 673750 554345 673802 554397
rect 675382 554345 675434 554397
rect 673078 553901 673130 553953
rect 675478 553901 675530 553953
rect 41590 553161 41642 553213
rect 42838 553161 42890 553213
rect 673174 553161 673226 553213
rect 675382 553161 675434 553213
rect 673654 551903 673706 551955
rect 675478 551903 675530 551955
rect 41878 550423 41930 550475
rect 43126 550423 43178 550475
rect 652630 550201 652682 550253
rect 656566 550201 656618 550253
rect 41590 550127 41642 550179
rect 42742 550127 42794 550179
rect 654838 550127 654890 550179
rect 666646 550127 666698 550179
rect 674422 548869 674474 548921
rect 675286 548869 675338 548921
rect 41878 548795 41930 548847
rect 42838 548795 42890 548847
rect 674326 548203 674378 548255
rect 675286 548203 675338 548255
rect 41878 547315 41930 547367
rect 44470 547315 44522 547367
rect 670774 547167 670826 547219
rect 679702 547167 679754 547219
rect 53302 544355 53354 544407
rect 59542 544355 59594 544407
rect 42262 542801 42314 542853
rect 43030 542801 43082 542853
rect 42070 541765 42122 541817
rect 43126 541765 43178 541817
rect 656662 541543 656714 541595
rect 42742 541469 42794 541521
rect 47638 541469 47690 541521
rect 670774 541395 670826 541447
rect 41398 541321 41450 541373
rect 43222 541321 43274 541373
rect 663766 541321 663818 541373
rect 676726 541321 676778 541373
rect 41494 541247 41546 541299
rect 43414 541247 43466 541299
rect 41782 540951 41834 541003
rect 41782 540729 41834 540781
rect 42070 538879 42122 538931
rect 42934 538879 42986 538931
rect 42934 538731 42986 538783
rect 43222 538731 43274 538783
rect 42166 538287 42218 538339
rect 42742 538287 42794 538339
rect 654454 537473 654506 537525
rect 663862 537473 663914 537525
rect 672598 537473 672650 537525
rect 676054 537473 676106 537525
rect 670774 537325 670826 537377
rect 676630 537325 676682 537377
rect 42070 537029 42122 537081
rect 43318 537029 43370 537081
rect 661078 536881 661130 536933
rect 676054 536881 676106 536933
rect 663958 536585 664010 536637
rect 676246 536585 676298 536637
rect 42070 535771 42122 535823
rect 42838 535771 42890 535823
rect 670966 534883 671018 534935
rect 676054 534883 676106 534935
rect 42166 534439 42218 534491
rect 42934 534439 42986 534491
rect 42166 533921 42218 533973
rect 43126 533921 43178 533973
rect 670870 533921 670922 533973
rect 676054 533921 676106 533973
rect 47638 532811 47690 532863
rect 59542 532811 59594 532863
rect 42166 531479 42218 531531
rect 42838 531479 42890 531531
rect 42070 530147 42122 530199
rect 43126 530147 43178 530199
rect 672214 529999 672266 530051
rect 676054 529999 676106 530051
rect 673558 529629 673610 529681
rect 676246 529629 676298 529681
rect 673270 528889 673322 528941
rect 676054 528889 676106 528941
rect 674710 528519 674762 528571
rect 674998 528519 675050 528571
rect 672406 528445 672458 528497
rect 676054 528445 676106 528497
rect 672886 528149 672938 528201
rect 676246 528149 676298 528201
rect 672310 527409 672362 527461
rect 676054 527409 676106 527461
rect 42166 527187 42218 527239
rect 43030 527187 43082 527239
rect 42070 527039 42122 527091
rect 42838 527039 42890 527091
rect 672118 526965 672170 527017
rect 676054 526965 676106 527017
rect 672982 526669 673034 526721
rect 676246 526669 676298 526721
rect 654454 524227 654506 524279
rect 663958 524227 664010 524279
rect 661078 524153 661130 524205
rect 679798 524153 679850 524205
rect 47830 518381 47882 518433
rect 59542 518381 59594 518433
rect 654454 509797 654506 509849
rect 672406 509797 672458 509849
rect 47734 504025 47786 504077
rect 59542 504025 59594 504077
rect 676534 498253 676586 498305
rect 679702 498253 679754 498305
rect 654454 495367 654506 495419
rect 670102 495367 670154 495419
rect 666838 493665 666890 493717
rect 676246 493665 676298 493717
rect 672502 492925 672554 492977
rect 676054 492925 676106 492977
rect 50422 492481 50474 492533
rect 59542 492481 59594 492533
rect 661174 492333 661226 492385
rect 676054 492333 676106 492385
rect 674998 489521 675050 489573
rect 676246 489521 676298 489573
rect 674614 489447 674666 489499
rect 676054 489447 676106 489499
rect 674422 489373 674474 489425
rect 676150 489373 676202 489425
rect 674518 486635 674570 486687
rect 676054 486635 676106 486687
rect 674326 486561 674378 486613
rect 676246 486561 676298 486613
rect 673846 485081 673898 485133
rect 676246 485081 676298 485133
rect 673654 484489 673706 484541
rect 676054 484489 676106 484541
rect 654454 484045 654506 484097
rect 661462 484045 661514 484097
rect 673078 483971 673130 484023
rect 676054 483971 676106 484023
rect 673750 483009 673802 483061
rect 676054 483009 676106 483061
rect 673174 482417 673226 482469
rect 676054 482417 676106 482469
rect 661174 479457 661226 479509
rect 679990 479457 680042 479509
rect 48022 478125 48074 478177
rect 59542 478125 59594 478177
rect 654454 469467 654506 469519
rect 666742 469467 666794 469519
rect 53494 466581 53546 466633
rect 57814 466581 57866 466633
rect 654454 455037 654506 455089
rect 661558 455037 661610 455089
rect 53206 452151 53258 452203
rect 59542 452151 59594 452203
rect 654454 443567 654506 443619
rect 672598 443567 672650 443619
rect 47926 440681 47978 440733
rect 57814 440681 57866 440733
rect 41782 432245 41834 432297
rect 47638 432245 47690 432297
rect 41782 431727 41834 431779
rect 47830 431727 47882 431779
rect 41590 431357 41642 431409
rect 53302 431357 53354 431409
rect 41782 430765 41834 430817
rect 43222 430765 43274 430817
rect 41782 430173 41834 430225
rect 43318 430173 43370 430225
rect 654454 429137 654506 429189
rect 663766 429137 663818 429189
rect 41590 428471 41642 428523
rect 43222 428471 43274 428523
rect 53398 426251 53450 426303
rect 59542 426251 59594 426303
rect 41590 421071 41642 421123
rect 43030 421071 43082 421123
rect 41590 420923 41642 420975
rect 42934 420923 42986 420975
rect 41974 420701 42026 420753
rect 43126 420701 43178 420753
rect 41782 420479 41834 420531
rect 42838 420479 42890 420531
rect 41782 419739 41834 419791
rect 47638 419739 47690 419791
rect 654454 417593 654506 417645
rect 672502 417593 672554 417645
rect 40726 417519 40778 417571
rect 44278 417519 44330 417571
rect 50614 414707 50666 414759
rect 59542 414707 59594 414759
rect 41878 413375 41930 413427
rect 41878 413153 41930 413205
rect 42070 410489 42122 410541
rect 50326 410489 50378 410541
rect 42166 409453 42218 409505
rect 42838 409453 42890 409505
rect 42166 408195 42218 408247
rect 42934 408195 42986 408247
rect 42070 407455 42122 407507
rect 43126 407455 43178 407507
rect 42166 406863 42218 406915
rect 43030 406863 43082 406915
rect 663862 405457 663914 405509
rect 676246 405457 676298 405509
rect 666646 404717 666698 404769
rect 676054 404717 676106 404769
rect 663958 404199 664010 404251
rect 676054 404199 676106 404251
rect 654454 403237 654506 403289
rect 666838 403237 666890 403289
rect 673846 403237 673898 403289
rect 676054 403237 676106 403289
rect 670870 402201 670922 402253
rect 676054 402201 676106 402253
rect 676054 402053 676106 402105
rect 676630 402053 676682 402105
rect 666646 401239 666698 401291
rect 676054 401239 676106 401291
rect 670966 400943 671018 400995
rect 676246 400943 676298 400995
rect 50326 400351 50378 400403
rect 59542 400351 59594 400403
rect 674326 400351 674378 400403
rect 676726 400351 676778 400403
rect 673750 395689 673802 395741
rect 676054 395689 676106 395741
rect 673654 393987 673706 394039
rect 676246 393987 676298 394039
rect 661270 391693 661322 391745
rect 679798 391693 679850 391745
rect 654838 390731 654890 390783
rect 661366 390731 661418 390783
rect 41782 389029 41834 389081
rect 48022 389029 48074 389081
rect 53302 388807 53354 388859
rect 59542 388807 59594 388859
rect 41590 388733 41642 388785
rect 53494 388733 53546 388785
rect 41782 387993 41834 388045
rect 50422 387993 50474 388045
rect 41782 387549 41834 387601
rect 43318 387549 43370 387601
rect 41782 386957 41834 387009
rect 43510 386957 43562 387009
rect 670198 385847 670250 385899
rect 674326 385847 674378 385899
rect 41590 385181 41642 385233
rect 43222 385181 43274 385233
rect 44182 385181 44234 385233
rect 34486 381555 34538 381607
rect 43318 381555 43370 381607
rect 61846 381555 61898 381607
rect 41782 380075 41834 380127
rect 42838 380075 42890 380127
rect 655318 378669 655370 378721
rect 666646 378669 666698 378721
rect 41590 378447 41642 378499
rect 43126 378447 43178 378499
rect 41782 378299 41834 378351
rect 42742 378299 42794 378351
rect 41590 378225 41642 378277
rect 43030 378225 43082 378277
rect 41782 377559 41834 377611
rect 42934 377559 42986 377611
rect 654454 377263 654506 377315
rect 670006 377263 670058 377315
rect 673750 377189 673802 377241
rect 675382 377189 675434 377241
rect 673654 376819 673706 376871
rect 675286 376819 675338 376871
rect 40246 376523 40298 376575
rect 41782 376523 41834 376575
rect 47830 376523 47882 376575
rect 50518 374377 50570 374429
rect 59446 374377 59498 374429
rect 41878 370159 41930 370211
rect 652630 370085 652682 370137
rect 670198 370085 670250 370137
rect 41878 369937 41930 369989
rect 42070 367347 42122 367399
rect 47734 367347 47786 367399
rect 42070 366237 42122 366289
rect 42838 366237 42890 366289
rect 42166 364979 42218 365031
rect 42934 364979 42986 365031
rect 654454 364831 654506 364883
rect 663862 364831 663914 364883
rect 42070 364387 42122 364439
rect 42742 364387 42794 364439
rect 42166 363647 42218 363699
rect 43030 363647 43082 363699
rect 48022 362907 48074 362959
rect 58390 362907 58442 362959
rect 652726 362833 652778 362885
rect 655318 362833 655370 362885
rect 42166 360613 42218 360665
rect 43126 360613 43178 360665
rect 670102 360021 670154 360073
rect 676054 360021 676106 360073
rect 672406 359725 672458 359777
rect 676246 359725 676298 359777
rect 661462 358985 661514 359037
rect 676054 358985 676106 359037
rect 673846 358541 673898 358593
rect 676054 358541 676106 358593
rect 670102 357727 670154 357779
rect 670870 357727 670922 357779
rect 676246 357727 676298 357779
rect 670966 356543 671018 356595
rect 676054 356543 676106 356595
rect 670294 354249 670346 354301
rect 670966 354249 671018 354301
rect 654454 351363 654506 351415
rect 666646 351363 666698 351415
rect 674806 351363 674858 351415
rect 676054 351363 676106 351415
rect 673942 349883 673994 349935
rect 676246 349883 676298 349935
rect 674038 349143 674090 349195
rect 676054 349143 676106 349195
rect 674230 348551 674282 348603
rect 676246 348551 676298 348603
rect 47734 348477 47786 348529
rect 59542 348477 59594 348529
rect 674710 348477 674762 348529
rect 676054 348477 676106 348529
rect 41782 345887 41834 345939
rect 53398 345887 53450 345939
rect 658582 345591 658634 345643
rect 679798 345591 679850 345643
rect 41590 345517 41642 345569
rect 50614 345517 50666 345569
rect 41782 344777 41834 344829
rect 47926 344777 47978 344829
rect 41782 344333 41834 344385
rect 43510 344333 43562 344385
rect 41782 343815 41834 343867
rect 43222 343815 43274 343867
rect 41782 343297 41834 343349
rect 43414 343297 43466 343349
rect 45334 343297 45386 343349
rect 41782 342335 41834 342387
rect 43510 342335 43562 342387
rect 45238 342335 45290 342387
rect 41590 341965 41642 342017
rect 43318 341965 43370 342017
rect 675766 341151 675818 341203
rect 675766 340929 675818 340981
rect 674806 337895 674858 337947
rect 675478 337895 675530 337947
rect 50422 337007 50474 337059
rect 59542 337007 59594 337059
rect 674230 336045 674282 336097
rect 675382 336045 675434 336097
rect 41590 335231 41642 335283
rect 43126 335231 43178 335283
rect 41782 334935 41834 334987
rect 42934 334935 42986 334987
rect 41590 334639 41642 334691
rect 43030 334639 43082 334691
rect 41782 334491 41834 334543
rect 42838 334491 42890 334543
rect 41782 333307 41834 333359
rect 47926 333307 47978 333359
rect 674038 332715 674090 332767
rect 675382 332715 675434 332767
rect 673942 332197 673994 332249
rect 675478 332197 675530 332249
rect 674710 331753 674762 331805
rect 675382 331753 675434 331805
rect 41878 327017 41930 327069
rect 41878 326721 41930 326773
rect 43030 326647 43082 326699
rect 43318 326647 43370 326699
rect 42454 326499 42506 326551
rect 43030 326499 43082 326551
rect 42166 324131 42218 324183
rect 53206 324131 53258 324183
rect 654838 323243 654890 323295
rect 661462 323243 661514 323295
rect 42166 323095 42218 323147
rect 42934 323095 42986 323147
rect 42934 322947 42986 322999
rect 43318 322947 43370 322999
rect 53398 322577 53450 322629
rect 59542 322577 59594 322629
rect 42070 321763 42122 321815
rect 42838 321763 42890 321815
rect 42166 321023 42218 321075
rect 43126 321023 43178 321075
rect 42166 320579 42218 320631
rect 42934 320579 42986 320631
rect 43414 318359 43466 318411
rect 43414 318137 43466 318189
rect 42166 317471 42218 317523
rect 43030 317471 43082 317523
rect 45718 316065 45770 316117
rect 49270 316065 49322 316117
rect 661558 315029 661610 315081
rect 676054 315029 676106 315081
rect 666742 314733 666794 314785
rect 676246 314733 676298 314785
rect 672598 313993 672650 314045
rect 676054 313993 676106 314045
rect 45238 311033 45290 311085
rect 58582 311033 58634 311085
rect 654454 311033 654506 311085
rect 672406 311033 672458 311085
rect 674326 309627 674378 309679
rect 676054 309627 676106 309679
rect 674230 308147 674282 308199
rect 676054 308147 676106 308199
rect 674134 306371 674186 306423
rect 676246 306371 676298 306423
rect 674038 305335 674090 305387
rect 676246 305335 676298 305387
rect 45814 305261 45866 305313
rect 49270 305187 49322 305239
rect 53206 305187 53258 305239
rect 674518 305261 674570 305313
rect 676054 305261 676106 305313
rect 58966 305187 59018 305239
rect 41782 302671 41834 302723
rect 50518 302671 50570 302723
rect 44374 302523 44426 302575
rect 53686 302523 53738 302575
rect 658678 302523 658730 302575
rect 679894 302523 679946 302575
rect 673942 302449 673994 302501
rect 676054 302449 676106 302501
rect 674422 302375 674474 302427
rect 676246 302375 676298 302427
rect 41590 302301 41642 302353
rect 48022 302301 48074 302353
rect 41782 301561 41834 301613
rect 53302 301561 53354 301613
rect 41782 301191 41834 301243
rect 43222 301191 43274 301243
rect 53686 301117 53738 301169
rect 55318 301117 55370 301169
rect 41782 300599 41834 300651
rect 43606 300599 43658 300651
rect 41782 300081 41834 300133
rect 43510 300081 43562 300133
rect 45142 300081 45194 300133
rect 41782 299637 41834 299689
rect 43414 299637 43466 299689
rect 41590 299341 41642 299393
rect 43222 299341 43274 299393
rect 44950 299341 45002 299393
rect 41782 298601 41834 298653
rect 43318 298601 43370 298653
rect 45142 296677 45194 296729
rect 59542 296677 59594 296729
rect 674230 295937 674282 295989
rect 675382 295937 675434 295989
rect 674518 295345 674570 295397
rect 675478 295345 675530 295397
rect 674326 294531 674378 294583
rect 675382 294531 675434 294583
rect 44278 293791 44330 293843
rect 55318 293791 55370 293843
rect 60310 293791 60362 293843
rect 60406 293717 60458 293769
rect 41878 292311 41930 292363
rect 43126 292311 43178 292363
rect 674134 292015 674186 292067
rect 675478 292015 675530 292067
rect 41590 291571 41642 291623
rect 43030 291571 43082 291623
rect 674038 291571 674090 291623
rect 675382 291571 675434 291623
rect 41590 291127 41642 291179
rect 42742 291127 42794 291179
rect 41878 291053 41930 291105
rect 42934 291053 42986 291105
rect 674422 291053 674474 291105
rect 675382 291053 675434 291105
rect 41782 290905 41834 290957
rect 42838 290905 42890 290957
rect 53206 290905 53258 290957
rect 57526 290905 57578 290957
rect 41782 290091 41834 290143
rect 48022 290091 48074 290143
rect 673942 286539 673994 286591
rect 675382 286539 675434 286591
rect 57526 285207 57578 285259
rect 63286 285207 63338 285259
rect 44950 285133 45002 285185
rect 59542 285133 59594 285185
rect 47542 285059 47594 285111
rect 60406 285059 60458 285111
rect 41974 283801 42026 283853
rect 41974 283505 42026 283557
rect 42166 281063 42218 281115
rect 50326 281063 50378 281115
rect 42166 279879 42218 279931
rect 42838 279879 42890 279931
rect 60310 278621 60362 278673
rect 652918 278621 652970 278673
rect 42166 278547 42218 278599
rect 42742 278547 42794 278599
rect 58966 278547 59018 278599
rect 652726 278547 652778 278599
rect 60502 278473 60554 278525
rect 653014 278473 653066 278525
rect 60598 278399 60650 278451
rect 652534 278399 652586 278451
rect 320950 278029 321002 278081
rect 422518 278029 422570 278081
rect 317878 277955 317930 278007
rect 415414 277955 415466 278007
rect 319510 277881 319562 277933
rect 419062 277881 419114 277933
rect 42166 277807 42218 277859
rect 43030 277807 43082 277859
rect 322102 277807 322154 277859
rect 426262 277807 426314 277859
rect 323830 277733 323882 277785
rect 429622 277733 429674 277785
rect 324982 277659 325034 277711
rect 433462 277659 433514 277711
rect 328054 277585 328106 277637
rect 440566 277585 440618 277637
rect 408022 277511 408074 277563
rect 546646 277511 546698 277563
rect 316630 277437 316682 277489
rect 412246 277437 412298 277489
rect 42070 277363 42122 277415
rect 42934 277363 42986 277415
rect 326422 277363 326474 277415
rect 437014 277363 437066 277415
rect 329302 277289 329354 277341
rect 444214 277289 444266 277341
rect 332374 277215 332426 277267
rect 451222 277215 451274 277267
rect 330742 277141 330794 277193
rect 447670 277141 447722 277193
rect 333622 277067 333674 277119
rect 454774 277067 454826 277119
rect 336694 276993 336746 277045
rect 461878 276993 461930 277045
rect 405430 276919 405482 276971
rect 612982 276919 613034 276971
rect 393910 276845 393962 276897
rect 603670 276845 603722 276897
rect 396790 276771 396842 276823
rect 610774 276771 610826 276823
rect 398230 276697 398282 276749
rect 614422 276697 614474 276749
rect 401110 276623 401162 276675
rect 621430 276623 621482 276675
rect 399382 276549 399434 276601
rect 617974 276549 618026 276601
rect 402550 276475 402602 276527
rect 625078 276475 625130 276527
rect 350230 276401 350282 276453
rect 496150 276401 496202 276453
rect 353398 276327 353450 276379
rect 503254 276327 503306 276379
rect 357430 276253 357482 276305
rect 513910 276253 513962 276305
rect 293014 276179 293066 276231
rect 354262 276179 354314 276231
rect 356182 276179 356234 276231
rect 510358 276179 510410 276231
rect 294646 276105 294698 276157
rect 357910 276105 357962 276157
rect 360310 276105 360362 276157
rect 521014 276105 521066 276157
rect 295894 276031 295946 276083
rect 361366 276031 361418 276083
rect 363382 276031 363434 276083
rect 528118 276031 528170 276083
rect 297334 275957 297386 276009
rect 364918 275957 364970 276009
rect 365974 275957 366026 276009
rect 535126 275957 535178 276009
rect 298966 275883 299018 275935
rect 368470 275883 368522 275935
rect 372502 275883 372554 275935
rect 550486 275883 550538 275935
rect 300214 275809 300266 275861
rect 372022 275809 372074 275861
rect 375094 275809 375146 275861
rect 557590 275809 557642 275861
rect 301750 275735 301802 275787
rect 375574 275735 375626 275787
rect 380566 275735 380618 275787
rect 303286 275661 303338 275713
rect 379126 275661 379178 275713
rect 381046 275661 381098 275713
rect 399094 275735 399146 275787
rect 564694 275735 564746 275787
rect 303766 275587 303818 275639
rect 380374 275587 380426 275639
rect 383446 275587 383498 275639
rect 570646 275661 570698 275713
rect 304438 275513 304490 275565
rect 382582 275513 382634 275565
rect 386518 275513 386570 275565
rect 571798 275587 571850 275639
rect 305014 275439 305066 275491
rect 383830 275439 383882 275491
rect 577750 275513 577802 275565
rect 586006 275439 586058 275491
rect 306358 275365 306410 275417
rect 387382 275365 387434 275417
rect 306166 275291 306218 275343
rect 386230 275291 386282 275343
rect 386326 275291 386378 275343
rect 584854 275365 584906 275417
rect 390358 275291 390410 275343
rect 308086 275217 308138 275269
rect 390934 275217 390986 275269
rect 395158 275217 395210 275269
rect 407926 275291 407978 275343
rect 591958 275291 592010 275343
rect 310390 275143 310442 275195
rect 396886 275143 396938 275195
rect 404950 275143 405002 275195
rect 595414 275217 595466 275269
rect 314710 275069 314762 275121
rect 407446 275069 407498 275121
rect 313558 274995 313610 275047
rect 405142 274995 405194 275047
rect 607318 275143 607370 275195
rect 407734 275069 407786 275121
rect 634390 275069 634442 275121
rect 630934 274995 630986 275047
rect 347638 274921 347690 274973
rect 489046 274921 489098 274973
rect 344566 274847 344618 274899
rect 481942 274847 481994 274899
rect 341686 274773 341738 274825
rect 474934 274773 474986 274825
rect 339094 274699 339146 274751
rect 467830 274699 467882 274751
rect 336022 274625 336074 274677
rect 460630 274625 460682 274677
rect 333142 274551 333194 274603
rect 453526 274551 453578 274603
rect 330454 274477 330506 274529
rect 446518 274477 446570 274529
rect 327574 274403 327626 274455
rect 439414 274403 439466 274455
rect 325942 274329 325994 274381
rect 435862 274329 435914 274381
rect 42166 274255 42218 274307
rect 43126 274255 43178 274307
rect 321622 274255 321674 274307
rect 425206 274255 425258 274307
rect 320182 274181 320234 274233
rect 421654 274181 421706 274233
rect 317302 274107 317354 274159
rect 414550 274107 414602 274159
rect 315958 274033 316010 274085
rect 411094 274033 411146 274085
rect 311638 273959 311690 274011
rect 400342 273959 400394 274011
rect 307318 273885 307370 273937
rect 389686 273885 389738 273937
rect 378262 273811 378314 273863
rect 399094 273811 399146 273863
rect 388918 273737 388970 273789
rect 407926 273737 407978 273789
rect 406102 273663 406154 273715
rect 407734 273663 407786 273715
rect 409654 273663 409706 273715
rect 480886 273663 480938 273715
rect 403702 273589 403754 273641
rect 506806 273589 506858 273641
rect 84790 273515 84842 273567
rect 142390 273515 142442 273567
rect 149782 273515 149834 273567
rect 207670 273515 207722 273567
rect 277750 273515 277802 273567
rect 316438 273515 316490 273567
rect 342166 273515 342218 273567
rect 476086 273515 476138 273567
rect 480886 273515 480938 273567
rect 642742 273515 642794 273567
rect 80086 273441 80138 273493
rect 142486 273441 142538 273493
rect 146230 273441 146282 273493
rect 210166 273441 210218 273493
rect 275350 273441 275402 273493
rect 310486 273441 310538 273493
rect 312790 273441 312842 273493
rect 402742 273441 402794 273493
rect 402838 273441 402890 273493
rect 545878 273441 545930 273493
rect 546646 273441 546698 273493
rect 639190 273441 639242 273493
rect 139126 273367 139178 273419
rect 207286 273367 207338 273419
rect 276310 273367 276362 273419
rect 312886 273367 312938 273419
rect 313942 273367 313994 273419
rect 329494 273367 329546 273419
rect 350998 273367 351050 273419
rect 497398 273367 497450 273419
rect 506806 273367 506858 273419
rect 628534 273367 628586 273419
rect 119062 273293 119114 273345
rect 120886 273293 120938 273345
rect 132022 273293 132074 273345
rect 206998 273293 207050 273345
rect 278230 273293 278282 273345
rect 317686 273293 317738 273345
rect 352630 273293 352682 273345
rect 502006 273293 502058 273345
rect 612982 273293 613034 273345
rect 632086 273293 632138 273345
rect 127318 273219 127370 273271
rect 209974 273219 210026 273271
rect 219574 273219 219626 273271
rect 238678 273219 238730 273271
rect 281302 273219 281354 273271
rect 324790 273219 324842 273271
rect 353686 273219 353738 273271
rect 504406 273219 504458 273271
rect 123766 273145 123818 273197
rect 209014 273145 209066 273197
rect 279670 273145 279722 273197
rect 321142 273145 321194 273197
rect 355798 273145 355850 273197
rect 509110 273145 509162 273197
rect 509206 273145 509258 273197
rect 635638 273145 635690 273197
rect 116662 273071 116714 273123
rect 207094 273071 207146 273123
rect 217174 273071 217226 273123
rect 237622 273071 237674 273123
rect 280630 273071 280682 273123
rect 323542 273071 323594 273123
rect 356758 273071 356810 273123
rect 511510 273071 511562 273123
rect 113206 272997 113258 273049
rect 205942 272997 205994 273049
rect 218326 272997 218378 273049
rect 238102 272997 238154 273049
rect 279286 272997 279338 273049
rect 319990 272997 320042 273049
rect 359350 272997 359402 273049
rect 120214 272923 120266 272975
rect 207958 272923 208010 272975
rect 220726 272923 220778 272975
rect 239158 272923 239210 272975
rect 288502 272923 288554 272975
rect 342454 272923 342506 272975
rect 361270 272923 361322 272975
rect 376054 272997 376106 273049
rect 516214 272997 516266 273049
rect 109558 272849 109610 272901
rect 205270 272849 205322 272901
rect 214870 272849 214922 272901
rect 236470 272849 236522 272901
rect 284950 272849 285002 272901
rect 334102 272849 334154 272901
rect 362230 272849 362282 272901
rect 518614 272923 518666 272975
rect 107158 272775 107210 272827
rect 204694 272775 204746 272827
rect 213622 272775 213674 272827
rect 236278 272775 236330 272827
rect 287926 272775 287978 272827
rect 341302 272775 341354 272827
rect 364150 272775 364202 272827
rect 523414 272849 523466 272901
rect 102550 272701 102602 272753
rect 203350 272701 203402 272753
rect 215926 272701 215978 272753
rect 236950 272701 237002 272753
rect 271030 272701 271082 272753
rect 299926 272701 299978 272753
rect 301846 272701 301898 272753
rect 358966 272701 359018 272753
rect 365302 272701 365354 272753
rect 375574 272701 375626 272753
rect 525718 272775 525770 272827
rect 530518 272701 530570 272753
rect 95446 272627 95498 272679
rect 201142 272627 201194 272679
rect 233686 272627 233738 272679
rect 244054 272627 244106 272679
rect 292726 272627 292778 272679
rect 353110 272627 353162 272679
rect 367030 272627 367082 272679
rect 537526 272627 537578 272679
rect 100150 272553 100202 272605
rect 202870 272553 202922 272605
rect 212470 272553 212522 272605
rect 235702 272553 235754 272605
rect 295414 272553 295466 272605
rect 360214 272553 360266 272605
rect 367894 272553 367946 272605
rect 93046 272479 93098 272531
rect 200950 272479 201002 272531
rect 208822 272479 208874 272531
rect 234358 272479 234410 272531
rect 270262 272479 270314 272531
rect 297526 272479 297578 272531
rect 298294 272479 298346 272531
rect 367222 272479 367274 272531
rect 374134 272479 374186 272531
rect 375574 272553 375626 272605
rect 532822 272553 532874 272605
rect 90646 272405 90698 272457
rect 199702 272405 199754 272457
rect 232534 272405 232586 272457
rect 243670 272405 243722 272457
rect 271798 272405 271850 272457
rect 301078 272405 301130 272457
rect 301366 272405 301418 272457
rect 374326 272405 374378 272457
rect 539830 272479 539882 272531
rect 555190 272405 555242 272457
rect 87094 272331 87146 272383
rect 199030 272331 199082 272383
rect 207766 272331 207818 272383
rect 233878 272331 233930 272383
rect 236086 272331 236138 272383
rect 245302 272331 245354 272383
rect 272758 272331 272810 272383
rect 303382 272331 303434 272383
rect 303958 272331 304010 272383
rect 381526 272331 381578 272383
rect 382966 272331 383018 272383
rect 576598 272331 576650 272383
rect 81238 272257 81290 272309
rect 196822 272257 196874 272309
rect 210070 272257 210122 272309
rect 234550 272257 234602 272309
rect 234934 272257 234986 272309
rect 244822 272257 244874 272309
rect 273430 272257 273482 272309
rect 305782 272257 305834 272309
rect 306838 272257 306890 272309
rect 388630 272257 388682 272309
rect 388726 272257 388778 272309
rect 590710 272257 590762 272309
rect 82390 272183 82442 272235
rect 197398 272183 197450 272235
rect 228982 272183 229034 272235
rect 242422 272183 242474 272235
rect 275158 272183 275210 272235
rect 309430 272183 309482 272235
rect 309910 272183 309962 272235
rect 395734 272183 395786 272235
rect 397078 272183 397130 272235
rect 612022 272183 612074 272235
rect 72982 272109 73034 272161
rect 194422 272109 194474 272161
rect 194710 272109 194762 272161
rect 224566 272109 224618 272161
rect 227830 272109 227882 272161
rect 242134 272109 242186 272161
rect 277078 272109 277130 272161
rect 314134 272109 314186 272161
rect 315478 272109 315530 272161
rect 409846 272109 409898 272161
rect 410902 272109 410954 272161
rect 646294 272109 646346 272161
rect 101302 272035 101354 272087
rect 159766 272035 159818 272087
rect 163990 272035 164042 272087
rect 207862 272035 207914 272087
rect 230230 272035 230282 272087
rect 242902 272035 242954 272087
rect 273910 272035 273962 272087
rect 307030 272035 307082 272087
rect 348118 272035 348170 272087
rect 490294 272035 490346 272087
rect 97750 271961 97802 272013
rect 151126 271961 151178 272013
rect 156886 271961 156938 272013
rect 207766 271961 207818 272013
rect 231382 271961 231434 272013
rect 243094 271961 243146 272013
rect 272950 271961 273002 272013
rect 304630 271961 304682 272013
rect 350038 271961 350090 272013
rect 494998 271961 495050 272013
rect 89494 271887 89546 271939
rect 142582 271887 142634 271939
rect 168694 271887 168746 271939
rect 169846 271887 169898 271939
rect 179350 271887 179402 271939
rect 181366 271887 181418 271939
rect 182902 271887 182954 271939
rect 184246 271887 184298 271939
rect 111958 271813 112010 271865
rect 162646 271813 162698 271865
rect 170998 271813 171050 271865
rect 207478 271887 207530 271939
rect 211222 271887 211274 271939
rect 235030 271887 235082 271939
rect 270550 271887 270602 271939
rect 298678 271887 298730 271939
rect 299446 271887 299498 271939
rect 327094 271887 327146 271939
rect 346966 271887 347018 271939
rect 487894 271887 487946 271939
rect 191158 271813 191210 271865
rect 227158 271813 227210 271865
rect 272278 271813 272330 271865
rect 302326 271813 302378 271865
rect 345238 271813 345290 271865
rect 483190 271813 483242 271865
rect 94198 271739 94250 271791
rect 142774 271739 142826 271791
rect 155638 271739 155690 271791
rect 104854 271665 104906 271717
rect 154006 271665 154058 271717
rect 108406 271591 108458 271643
rect 156886 271591 156938 271643
rect 126166 271517 126218 271569
rect 143062 271517 143114 271569
rect 162742 271739 162794 271791
rect 192982 271739 193034 271791
rect 195862 271739 195914 271791
rect 221590 271739 221642 271791
rect 344086 271739 344138 271791
rect 480790 271739 480842 271791
rect 178102 271665 178154 271717
rect 207382 271665 207434 271717
rect 341494 271665 341546 271717
rect 473686 271665 473738 271717
rect 161590 271591 161642 271643
rect 164086 271591 164138 271643
rect 185398 271591 185450 271643
rect 186358 271591 186410 271643
rect 193174 271591 193226 271643
rect 201814 271591 201866 271643
rect 224278 271591 224330 271643
rect 338614 271591 338666 271643
rect 466582 271591 466634 271643
rect 192310 271517 192362 271569
rect 221974 271517 222026 271569
rect 335446 271517 335498 271569
rect 459574 271517 459626 271569
rect 129622 271443 129674 271495
rect 142966 271443 143018 271495
rect 181750 271443 181802 271495
rect 210454 271443 210506 271495
rect 332566 271443 332618 271495
rect 452470 271443 452522 271495
rect 133270 271369 133322 271421
rect 142870 271369 142922 271421
rect 169750 271369 169802 271421
rect 198646 271369 198698 271421
rect 199510 271369 199562 271421
rect 221494 271369 221546 271421
rect 329974 271369 330026 271421
rect 445270 271369 445322 271421
rect 185206 271295 185258 271347
rect 210358 271295 210410 271347
rect 237238 271295 237290 271347
rect 245494 271295 245546 271347
rect 326902 271295 326954 271347
rect 438166 271295 438218 271347
rect 136822 271221 136874 271273
rect 143158 271221 143210 271273
rect 193462 271221 193514 271273
rect 221686 271221 221738 271273
rect 238486 271221 238538 271273
rect 246070 271221 246122 271273
rect 324022 271221 324074 271273
rect 431158 271221 431210 271273
rect 75286 271147 75338 271199
rect 77494 271147 77546 271199
rect 176950 271147 177002 271199
rect 204022 271147 204074 271199
rect 205366 271147 205418 271199
rect 232630 271147 232682 271199
rect 239542 271147 239594 271199
rect 246454 271147 246506 271199
rect 321430 271147 321482 271199
rect 424054 271147 424106 271199
rect 140278 271073 140330 271125
rect 143254 271073 143306 271125
rect 175798 271073 175850 271125
rect 178486 271073 178538 271125
rect 188758 271073 188810 271125
rect 210262 271073 210314 271125
rect 240790 271073 240842 271125
rect 247222 271073 247274 271125
rect 318358 271073 318410 271125
rect 416950 271073 417002 271125
rect 187606 270999 187658 271051
rect 205846 270999 205898 271051
rect 221878 270999 221930 271051
rect 239350 270999 239402 271051
rect 241942 270999 241994 271051
rect 247702 270999 247754 271051
rect 358582 270999 358634 271051
rect 376054 270999 376106 271051
rect 198262 270925 198314 270977
rect 68182 270703 68234 270755
rect 69046 270703 69098 270755
rect 115510 270703 115562 270755
rect 118006 270703 118058 270755
rect 122518 270703 122570 270755
rect 123766 270703 123818 270755
rect 143926 270703 143978 270755
rect 145366 270703 145418 270755
rect 147382 270703 147434 270755
rect 149686 270703 149738 270755
rect 151030 270703 151082 270755
rect 152566 270703 152618 270755
rect 154486 270703 154538 270755
rect 155446 270703 155498 270755
rect 165142 270703 165194 270755
rect 166966 270703 167018 270755
rect 223126 270925 223178 270977
rect 240022 270925 240074 270977
rect 243190 270925 243242 270977
rect 247990 270925 248042 270977
rect 224182 270851 224234 270903
rect 240502 270851 240554 270903
rect 244342 270851 244394 270903
rect 248662 270851 248714 270903
rect 225430 270777 225482 270829
rect 241078 270777 241130 270829
rect 245590 270777 245642 270829
rect 249142 270777 249194 270829
rect 340534 270777 340586 270829
rect 348406 270777 348458 270829
rect 142678 270629 142730 270681
rect 214294 270629 214346 270681
rect 226582 270703 226634 270755
rect 241270 270703 241322 270755
rect 246742 270703 246794 270755
rect 249622 270703 249674 270755
rect 230038 270629 230090 270681
rect 262006 270629 262058 270681
rect 137878 270555 137930 270607
rect 212662 270555 212714 270607
rect 262966 270555 263018 270607
rect 134422 270481 134474 270533
rect 211894 270481 211946 270533
rect 124918 270407 124970 270459
rect 209494 270407 209546 270459
rect 262486 270407 262538 270459
rect 121366 270333 121418 270385
rect 208342 270333 208394 270385
rect 117910 270259 117962 270311
rect 207574 270259 207626 270311
rect 207670 270259 207722 270311
rect 216214 270259 216266 270311
rect 253942 270259 253994 270311
rect 257302 270259 257354 270311
rect 264886 270259 264938 270311
rect 269878 270259 269930 270311
rect 283702 270629 283754 270681
rect 330646 270629 330698 270681
rect 284182 270555 284234 270607
rect 331798 270555 331850 270607
rect 285622 270481 285674 270533
rect 335350 270481 335402 270533
rect 277462 270407 277514 270459
rect 286294 270407 286346 270459
rect 337750 270703 337802 270755
rect 348406 270629 348458 270681
rect 491446 270629 491498 270681
rect 349462 270555 349514 270607
rect 493750 270555 493802 270607
rect 352438 270481 352490 270533
rect 500854 270481 500906 270533
rect 351286 270407 351338 270459
rect 498550 270407 498602 270459
rect 279766 270333 279818 270385
rect 286774 270333 286826 270385
rect 338902 270333 338954 270385
rect 355030 270333 355082 270385
rect 507958 270333 508010 270385
rect 278710 270259 278762 270311
rect 290614 270259 290666 270311
rect 340534 270259 340586 270311
rect 354070 270259 354122 270311
rect 505654 270259 505706 270311
rect 114262 270185 114314 270237
rect 206422 270185 206474 270237
rect 210166 270185 210218 270237
rect 214966 270185 215018 270237
rect 255286 270185 255338 270237
rect 260950 270185 261002 270237
rect 266038 270185 266090 270237
rect 286870 270185 286922 270237
rect 289174 270185 289226 270237
rect 344854 270185 344906 270237
rect 357910 270185 357962 270237
rect 515062 270185 515114 270237
rect 110806 270111 110858 270163
rect 205750 270111 205802 270163
rect 207382 270111 207434 270163
rect 223606 270111 223658 270163
rect 264694 270111 264746 270163
rect 103702 270037 103754 270089
rect 203542 270037 203594 270089
rect 210454 270037 210506 270089
rect 224758 270037 224810 270089
rect 265366 270037 265418 270089
rect 269878 270111 269930 270163
rect 284566 270111 284618 270163
rect 289942 270111 289994 270163
rect 346006 270111 346058 270163
rect 356950 270111 357002 270163
rect 512758 270111 512810 270163
rect 106006 269963 106058 270015
rect 204214 269963 204266 270015
rect 210358 269963 210410 270015
rect 225526 269963 225578 270015
rect 266518 269963 266570 270015
rect 283318 270037 283370 270089
rect 291094 270037 291146 270089
rect 349558 270037 349610 270089
rect 359830 270037 359882 270089
rect 519766 270037 519818 270089
rect 672502 270037 672554 270089
rect 676054 270037 676106 270089
rect 98902 269889 98954 269941
rect 202294 269889 202346 269941
rect 207478 269889 207530 269941
rect 221782 269889 221834 269941
rect 96598 269815 96650 269867
rect 201622 269815 201674 269867
rect 210262 269815 210314 269867
rect 226678 269815 226730 269867
rect 258646 269815 258698 269867
rect 269206 269815 269258 269867
rect 285718 269963 285770 270015
rect 293974 269963 294026 270015
rect 356662 269963 356714 270015
rect 360982 269963 361034 270015
rect 522166 269963 522218 270015
rect 269494 269889 269546 269941
rect 289270 269889 289322 269941
rect 292246 269889 292298 269941
rect 351862 269889 351914 269941
rect 363574 269889 363626 269941
rect 529270 269889 529322 269941
rect 288022 269815 288074 269867
rect 293494 269815 293546 269867
rect 355510 269815 355562 269867
rect 362806 269815 362858 269867
rect 526870 269815 526922 269867
rect 91798 269741 91850 269793
rect 177046 269741 177098 269793
rect 204022 269741 204074 269793
rect 223414 269741 223466 269793
rect 268438 269741 268490 269793
rect 292822 269741 292874 269793
rect 296470 269741 296522 269793
rect 362614 269741 362666 269793
rect 365686 269741 365738 269793
rect 533974 269741 534026 269793
rect 663766 269741 663818 269793
rect 676246 269741 676298 269793
rect 88342 269667 88394 269719
rect 199222 269667 199274 269719
rect 205846 269667 205898 269719
rect 226006 269667 226058 269719
rect 255766 269667 255818 269719
rect 262102 269667 262154 269719
rect 267286 269667 267338 269719
rect 290422 269667 290474 269719
rect 297046 269667 297098 269719
rect 363766 269667 363818 269719
rect 366550 269667 366602 269719
rect 536374 269667 536426 269719
rect 85942 269593 85994 269645
rect 198550 269593 198602 269645
rect 198646 269593 198698 269645
rect 221206 269593 221258 269645
rect 249046 269593 249098 269645
rect 250294 269593 250346 269645
rect 269206 269593 269258 269645
rect 295126 269593 295178 269645
rect 299638 269593 299690 269645
rect 83542 269519 83594 269571
rect 198070 269519 198122 269571
rect 206518 269519 206570 269571
rect 233398 269519 233450 269571
rect 253366 269519 253418 269571
rect 256150 269519 256202 269571
rect 267094 269519 267146 269571
rect 269494 269519 269546 269571
rect 269686 269519 269738 269571
rect 296374 269519 296426 269571
rect 302614 269519 302666 269571
rect 367126 269519 367178 269571
rect 369622 269593 369674 269645
rect 543478 269593 543530 269645
rect 370870 269519 370922 269571
rect 76438 269445 76490 269497
rect 195670 269445 195722 269497
rect 204118 269445 204170 269497
rect 232150 269445 232202 269497
rect 256246 269445 256298 269497
rect 263254 269445 263306 269497
rect 267766 269445 267818 269497
rect 291670 269445 291722 269497
rect 305686 269445 305738 269497
rect 384982 269519 385034 269571
rect 78838 269371 78890 269423
rect 196630 269371 196682 269423
rect 202966 269371 203018 269423
rect 231958 269371 232010 269423
rect 268630 269371 268682 269423
rect 294070 269371 294122 269423
rect 308278 269371 308330 269423
rect 74038 269297 74090 269349
rect 194998 269297 195050 269349
rect 200566 269297 200618 269349
rect 230998 269297 231050 269349
rect 258166 269297 258218 269349
rect 267958 269297 268010 269349
rect 274678 269297 274730 269349
rect 308182 269297 308234 269349
rect 367126 269297 367178 269349
rect 377974 269297 378026 269349
rect 379126 269371 379178 269423
rect 567094 269519 567146 269571
rect 392086 269297 392138 269349
rect 77686 269223 77738 269275
rect 196150 269223 196202 269275
rect 197110 269223 197162 269275
rect 229558 269223 229610 269275
rect 260086 269223 260138 269275
rect 272662 269223 272714 269275
rect 384118 269223 384170 269275
rect 580054 269445 580106 269497
rect 392758 269371 392810 269423
rect 601366 269371 601418 269423
rect 398998 269297 399050 269349
rect 615574 269297 615626 269349
rect 407254 269223 407306 269275
rect 636790 269223 636842 269275
rect 135670 269149 135722 269201
rect 212374 269149 212426 269201
rect 260566 269149 260618 269201
rect 273814 269149 273866 269201
rect 281782 269149 281834 269201
rect 325366 269149 325418 269201
rect 345430 269149 345482 269201
rect 484246 269149 484298 269201
rect 666838 269149 666890 269201
rect 676246 269149 676298 269201
rect 141526 269075 141578 269127
rect 213814 269075 213866 269127
rect 259894 269075 259946 269127
rect 271510 269075 271562 269127
rect 282550 269075 282602 269127
rect 328246 269075 328298 269127
rect 346486 269075 346538 269127
rect 486646 269075 486698 269127
rect 144982 269001 145034 269053
rect 214486 269001 214538 269053
rect 261814 269001 261866 269053
rect 276214 269001 276266 269053
rect 280150 269001 280202 269053
rect 322390 269001 322442 269053
rect 343606 269001 343658 269053
rect 479638 269001 479690 269053
rect 148630 268927 148682 268979
rect 215734 268927 215786 268979
rect 278902 268927 278954 268979
rect 318742 268927 318794 268979
rect 342646 268927 342698 268979
rect 477238 268927 477290 268979
rect 152182 268853 152234 268905
rect 216694 268853 216746 268905
rect 264118 268853 264170 268905
rect 153334 268779 153386 268831
rect 216886 268779 216938 268831
rect 257014 268779 257066 268831
rect 264406 268779 264458 268831
rect 277558 268853 277610 268905
rect 315286 268853 315338 268905
rect 339766 268853 339818 268905
rect 470134 268853 470186 268905
rect 282166 268779 282218 268831
rect 283030 268779 283082 268831
rect 313942 268779 313994 268831
rect 341014 268779 341066 268831
rect 472534 268779 472586 268831
rect 160438 268705 160490 268757
rect 218902 268705 218954 268757
rect 257686 268705 257738 268757
rect 266806 268705 266858 268757
rect 282070 268705 282122 268757
rect 299446 268705 299498 268757
rect 336886 268705 336938 268757
rect 463030 268705 463082 268757
rect 159286 268631 159338 268683
rect 218614 268631 218666 268683
rect 275830 268631 275882 268683
rect 311734 268631 311786 268683
rect 334294 268631 334346 268683
rect 455926 268631 455978 268683
rect 166390 268557 166442 268609
rect 220534 268557 220586 268609
rect 331222 268557 331274 268609
rect 448822 268557 448874 268609
rect 167542 268483 167594 268535
rect 221014 268483 221066 268535
rect 253174 268483 253226 268535
rect 254998 268483 255050 268535
rect 259414 268483 259466 268535
rect 270358 268483 270410 268535
rect 328342 268483 328394 268535
rect 441814 268483 441866 268535
rect 173398 268409 173450 268461
rect 222358 268409 222410 268461
rect 325750 268409 325802 268461
rect 434710 268409 434762 268461
rect 174646 268335 174698 268387
rect 222838 268335 222890 268387
rect 247894 268335 247946 268387
rect 249814 268335 249866 268387
rect 252694 268335 252746 268387
rect 253846 268335 253898 268387
rect 261238 268335 261290 268387
rect 275062 268335 275114 268387
rect 322582 268335 322634 268387
rect 427606 268335 427658 268387
rect 177046 268261 177098 268313
rect 200470 268261 200522 268313
rect 205366 268261 205418 268313
rect 225238 268261 225290 268313
rect 257494 268261 257546 268313
rect 265558 268261 265610 268313
rect 319702 268261 319754 268313
rect 420502 268261 420554 268313
rect 180502 268187 180554 268239
rect 205462 268187 205514 268239
rect 205654 268187 205706 268239
rect 224086 268187 224138 268239
rect 224278 268187 224330 268239
rect 231478 268187 231530 268239
rect 254614 268187 254666 268239
rect 258550 268187 258602 268239
rect 263638 268187 263690 268239
rect 281014 268187 281066 268239
rect 317110 268187 317162 268239
rect 413398 268187 413450 268239
rect 184150 268113 184202 268165
rect 205366 268113 205418 268165
rect 192982 268039 193034 268091
rect 219286 268113 219338 268165
rect 224566 268113 224618 268165
rect 228406 268113 228458 268165
rect 311158 268113 311210 268165
rect 399190 268113 399242 268165
rect 207286 268039 207338 268091
rect 213334 268039 213386 268091
rect 221494 268039 221546 268091
rect 230422 268039 230474 268091
rect 314230 268039 314282 268091
rect 406294 268039 406346 268091
rect 193174 267965 193226 268017
rect 217366 267965 217418 268017
rect 221590 267965 221642 268017
rect 229078 267965 229130 268017
rect 334966 267965 335018 268017
rect 346870 267965 346922 268017
rect 207862 267891 207914 267943
rect 219958 267891 220010 267943
rect 221974 267891 222026 267943
rect 227638 267891 227690 267943
rect 255094 267891 255146 267943
rect 259702 267891 259754 267943
rect 337846 267891 337898 267943
rect 207766 267817 207818 267869
rect 218134 267817 218186 267869
rect 221686 267817 221738 267869
rect 227830 267817 227882 267869
rect 295222 267817 295274 267869
rect 301846 267817 301898 267869
rect 339286 267817 339338 267869
rect 354262 267817 354314 267869
rect 359926 267817 359978 267869
rect 359158 267743 359210 267795
rect 517366 267743 517418 267795
rect 361750 267669 361802 267721
rect 524470 267669 524522 267721
rect 364630 267595 364682 267647
rect 531574 267595 531626 267647
rect 367702 267521 367754 267573
rect 538774 267521 538826 267573
rect 370774 267447 370826 267499
rect 547030 267447 547082 267499
rect 286102 267373 286154 267425
rect 336502 267373 336554 267425
rect 372022 267373 372074 267425
rect 549334 267373 549386 267425
rect 284470 267299 284522 267351
rect 333046 267299 333098 267351
rect 373174 267299 373226 267351
rect 552886 267299 552938 267351
rect 288694 267225 288746 267277
rect 343318 267225 343370 267277
rect 373846 267225 373898 267277
rect 554134 267225 554186 267277
rect 287350 267151 287402 267203
rect 340150 267151 340202 267203
rect 374614 267151 374666 267203
rect 556438 267151 556490 267203
rect 291574 267077 291626 267129
rect 350710 267077 350762 267129
rect 377494 267077 377546 267129
rect 563542 267077 563594 267129
rect 290422 267003 290474 267055
rect 347254 267003 347306 267055
rect 376822 267003 376874 267055
rect 561238 267003 561290 267055
rect 297814 266929 297866 266981
rect 366070 266929 366122 266981
rect 376246 266929 376298 266981
rect 559990 266929 560042 266981
rect 300694 266855 300746 266907
rect 373270 266855 373322 266907
rect 379414 266855 379466 266907
rect 568246 266855 568298 266907
rect 299446 266781 299498 266833
rect 369334 266781 369386 266833
rect 382294 266781 382346 266833
rect 575350 266781 575402 266833
rect 302038 266707 302090 266759
rect 376726 266707 376778 266759
rect 385366 266707 385418 266759
rect 582454 266707 582506 266759
rect 308758 266633 308810 266685
rect 309238 266559 309290 266611
rect 392278 266633 392330 266685
rect 600214 266633 600266 266685
rect 310678 266485 310730 266537
rect 393334 266559 393386 266611
rect 394678 266559 394730 266611
rect 606070 266559 606122 266611
rect 394486 266485 394538 266537
rect 398902 266485 398954 266537
rect 616726 266485 616778 266537
rect 398038 266411 398090 266463
rect 400630 266411 400682 266463
rect 620278 266411 620330 266463
rect 187222 266337 187274 266389
rect 189718 266337 189770 266389
rect 312310 266337 312362 266389
rect 401590 266337 401642 266389
rect 403222 266337 403274 266389
rect 627382 266337 627434 266389
rect 354838 266263 354890 266315
rect 506518 266263 506570 266315
rect 351958 266189 352010 266241
rect 499702 266189 499754 266241
rect 348886 266115 348938 266167
rect 492598 266115 492650 266167
rect 346006 266041 346058 266093
rect 485494 266041 485546 266093
rect 343318 265967 343370 266019
rect 478390 265967 478442 266019
rect 340246 265893 340298 265945
rect 471286 265893 471338 265945
rect 337366 265819 337418 265871
rect 464278 265819 464330 265871
rect 334774 265745 334826 265797
rect 457174 265745 457226 265797
rect 331894 265671 331946 265723
rect 450070 265671 450122 265723
rect 328822 265597 328874 265649
rect 442966 265597 443018 265649
rect 324502 265523 324554 265575
rect 432310 265523 432362 265575
rect 323350 265449 323402 265501
rect 428854 265449 428906 265501
rect 313078 265375 313130 265427
rect 403990 265375 404042 265427
rect 406582 265375 406634 265427
rect 509206 265375 509258 265427
rect 319030 265301 319082 265353
rect 418102 265301 418154 265353
rect 314902 265227 314954 265279
rect 408694 265227 408746 265279
rect 354262 264931 354314 264983
rect 468886 264931 468938 264983
rect 346870 264857 346922 264909
rect 458326 264857 458378 264909
rect 359926 264783 359978 264835
rect 465430 264783 465482 264835
rect 142390 262415 142442 262467
rect 142678 262415 142730 262467
rect 420406 262119 420458 262171
rect 606166 262119 606218 262171
rect 674614 261379 674666 261431
rect 676246 261379 676298 261431
rect 41590 259677 41642 259729
rect 50422 259677 50474 259729
rect 674710 259307 674762 259359
rect 676054 259307 676106 259359
rect 420406 259233 420458 259285
rect 603286 259233 603338 259285
rect 43222 259159 43274 259211
rect 44854 259159 44906 259211
rect 41782 258937 41834 258989
rect 53398 258937 53450 258989
rect 41782 258345 41834 258397
rect 47734 258345 47786 258397
rect 41782 257975 41834 258027
rect 43606 257975 43658 258027
rect 41782 257383 41834 257435
rect 43510 257383 43562 257435
rect 41782 256865 41834 256917
rect 43222 256865 43274 256917
rect 41782 256495 41834 256547
rect 43414 256495 43466 256547
rect 674038 256421 674090 256473
rect 676054 256421 676106 256473
rect 420406 256347 420458 256399
rect 603382 256347 603434 256399
rect 646486 256347 646538 256399
rect 679702 256347 679754 256399
rect 41782 255903 41834 255955
rect 43414 255903 43466 255955
rect 41782 255385 41834 255437
rect 43318 255385 43370 255437
rect 43414 255385 43466 255437
rect 44758 255385 44810 255437
rect 420406 253461 420458 253513
rect 603478 253461 603530 253513
rect 675670 251167 675722 251219
rect 675766 251167 675818 251219
rect 675670 250945 675722 250997
rect 420406 250575 420458 250627
rect 603574 250575 603626 250627
rect 675766 250205 675818 250257
rect 120886 249465 120938 249517
rect 145558 249465 145610 249517
rect 48022 249391 48074 249443
rect 186838 249391 186890 249443
rect 47638 249317 47690 249369
rect 186742 249317 186794 249369
rect 41590 249243 41642 249295
rect 43126 249243 43178 249295
rect 47830 249243 47882 249295
rect 186934 249243 186986 249295
rect 47926 249169 47978 249221
rect 187030 249169 187082 249221
rect 44470 249095 44522 249147
rect 186454 249095 186506 249147
rect 41590 248355 41642 248407
rect 42838 248355 42890 248407
rect 41590 248059 41642 248111
rect 42934 248059 42986 248111
rect 41782 247911 41834 247963
rect 42742 247911 42794 247963
rect 41974 247837 42026 247889
rect 43030 247837 43082 247889
rect 420310 247763 420362 247815
rect 600406 247763 600458 247815
rect 41590 247689 41642 247741
rect 157078 247689 157130 247741
rect 420406 247689 420458 247741
rect 626326 247689 626378 247741
rect 674614 247023 674666 247075
rect 675478 247023 675530 247075
rect 118006 246949 118058 247001
rect 145654 246949 145706 247001
rect 123766 246875 123818 246927
rect 168502 246875 168554 246927
rect 77494 246801 77546 246853
rect 145462 246801 145514 246853
rect 69046 246727 69098 246779
rect 145750 246727 145802 246779
rect 47446 246653 47498 246705
rect 186646 246653 186698 246705
rect 45910 246579 45962 246631
rect 186166 246579 186218 246631
rect 46006 246505 46058 246557
rect 186550 246505 186602 246557
rect 45430 246431 45482 246483
rect 186070 246431 186122 246483
rect 45622 246357 45674 246409
rect 186358 246357 186410 246409
rect 45526 246283 45578 246335
rect 186262 246283 186314 246335
rect 45046 246209 45098 246261
rect 185878 246209 185930 246261
rect 41590 244803 41642 244855
rect 156982 244803 157034 244855
rect 420406 244803 420458 244855
rect 629206 244803 629258 244855
rect 41686 243323 41738 243375
rect 185590 243323 185642 243375
rect 674710 242953 674762 243005
rect 675382 242953 675434 243005
rect 45046 242805 45098 242857
rect 185302 242805 185354 242857
rect 45334 242731 45386 242783
rect 185974 242731 186026 242783
rect 44854 242657 44906 242709
rect 185494 242657 185546 242709
rect 44758 242583 44810 242635
rect 185782 242583 185834 242635
rect 149398 241917 149450 241969
rect 168406 241917 168458 241969
rect 420406 241917 420458 241969
rect 600502 241917 600554 241969
rect 674038 241769 674090 241821
rect 675286 241769 675338 241821
rect 41878 240585 41930 240637
rect 41878 240363 41930 240415
rect 383062 239623 383114 239675
rect 464758 239623 464810 239675
rect 352822 239549 352874 239601
rect 439126 239549 439178 239601
rect 363238 239475 363290 239527
rect 378838 239475 378890 239527
rect 383158 239475 383210 239527
rect 473878 239475 473930 239527
rect 369286 239401 369338 239453
rect 376150 239401 376202 239453
rect 394486 239401 394538 239453
rect 496534 239401 496586 239453
rect 365014 239327 365066 239379
rect 505654 239327 505706 239379
rect 372118 239253 372170 239305
rect 523798 239253 523850 239305
rect 388534 239179 388586 239231
rect 413398 239179 413450 239231
rect 420406 239179 420458 239231
rect 596182 239179 596234 239231
rect 367222 239105 367274 239157
rect 542614 239105 542666 239157
rect 149398 239031 149450 239083
rect 174166 239031 174218 239083
rect 377590 239031 377642 239083
rect 561718 239031 561770 239083
rect 323926 238957 323978 239009
rect 455062 238957 455114 239009
rect 327670 238883 327722 238935
rect 461878 238883 461930 238935
rect 326710 238809 326762 238861
rect 462550 238809 462602 238861
rect 329878 238735 329930 238787
rect 468598 238735 468650 238787
rect 332662 238661 332714 238713
rect 474646 238661 474698 238713
rect 335734 238587 335786 238639
rect 480694 238587 480746 238639
rect 338998 238513 339050 238565
rect 486742 238513 486794 238565
rect 341782 238439 341834 238491
rect 492790 238439 492842 238491
rect 345910 238365 345962 238417
rect 498262 238365 498314 238417
rect 345334 238291 345386 238343
rect 500278 238291 500330 238343
rect 348118 238217 348170 238269
rect 504118 238217 504170 238269
rect 351190 238143 351242 238195
rect 512374 238143 512426 238195
rect 354166 238069 354218 238121
rect 518518 238069 518570 238121
rect 361366 237995 361418 238047
rect 532054 237995 532106 238047
rect 363094 237921 363146 237973
rect 535126 237921 535178 237973
rect 360310 237847 360362 237899
rect 530518 237847 530570 237899
rect 364438 237773 364490 237825
rect 538006 237773 538058 237825
rect 365878 237699 365930 237751
rect 538582 237699 538634 237751
rect 367606 237625 367658 237677
rect 541558 237625 541610 237677
rect 370390 237551 370442 237603
rect 550870 237551 550922 237603
rect 323158 237477 323210 237529
rect 452758 237477 452810 237529
rect 320854 237403 320906 237455
rect 450454 237403 450506 237455
rect 317590 237329 317642 237381
rect 444502 237329 444554 237381
rect 314806 237255 314858 237307
rect 438358 237255 438410 237307
rect 313846 237181 313898 237233
rect 434614 237181 434666 237233
rect 310774 237107 310826 237159
rect 428662 237107 428714 237159
rect 307030 237033 307082 237085
rect 423286 237033 423338 237085
rect 304822 236959 304874 237011
rect 301750 236885 301802 236937
rect 409654 236885 409706 236937
rect 286198 236811 286250 236863
rect 381046 236811 381098 236863
rect 411574 236959 411626 237011
rect 413974 236959 414026 237011
rect 410710 236885 410762 236937
rect 413686 236885 413738 236937
rect 416470 236811 416522 236863
rect 281590 236737 281642 236789
rect 372406 236737 372458 236789
rect 42166 236663 42218 236715
rect 42742 236663 42794 236715
rect 278422 236663 278474 236715
rect 366742 236663 366794 236715
rect 388822 236663 388874 236715
rect 390358 236663 390410 236715
rect 279862 236589 279914 236641
rect 368950 236589 369002 236641
rect 388630 236589 388682 236641
rect 389014 236589 389066 236641
rect 390358 236515 390410 236567
rect 476950 236515 477002 236567
rect 42838 236441 42890 236493
rect 43126 236441 43178 236493
rect 397366 236441 397418 236493
rect 483862 236441 483914 236493
rect 363574 236293 363626 236345
rect 381430 236293 381482 236345
rect 346294 236145 346346 236197
rect 361654 236145 361706 236197
rect 383830 236145 383882 236197
rect 388726 236145 388778 236197
rect 231190 236071 231242 236123
rect 253558 236071 253610 236123
rect 255286 236071 255338 236123
rect 273718 236071 273770 236123
rect 285142 236071 285194 236123
rect 326806 236071 326858 236123
rect 350422 236071 350474 236123
rect 508630 236367 508682 236419
rect 403318 236293 403370 236345
rect 520726 236293 520778 236345
rect 403222 236219 403274 236271
rect 526678 236219 526730 236271
rect 411670 236145 411722 236197
rect 544342 236145 544394 236197
rect 400246 236071 400298 236123
rect 485590 236071 485642 236123
rect 250486 235997 250538 236049
rect 272374 235997 272426 236049
rect 282166 235997 282218 236049
rect 325366 235997 325418 236049
rect 333814 235997 333866 236049
rect 466486 235997 466538 236049
rect 211222 235923 211274 235975
rect 229270 235923 229322 235975
rect 241654 235923 241706 235975
rect 266326 235923 266378 235975
rect 286678 235923 286730 235975
rect 331126 235923 331178 235975
rect 339862 235923 339914 235975
rect 475222 235923 475274 235975
rect 210646 235849 210698 235901
rect 230038 235849 230090 235901
rect 244342 235849 244394 235901
rect 268150 235849 268202 235901
rect 271990 235849 272042 235901
rect 282358 235849 282410 235901
rect 287446 235849 287498 235901
rect 341974 235849 342026 235901
rect 343126 235849 343178 235901
rect 483766 235849 483818 235901
rect 212950 235775 213002 235827
rect 232342 235775 232394 235827
rect 233494 235775 233546 235827
rect 211990 235701 212042 235753
rect 233014 235701 233066 235753
rect 211606 235627 211658 235679
rect 230710 235627 230762 235679
rect 238006 235775 238058 235827
rect 264694 235775 264746 235827
rect 265750 235775 265802 235827
rect 290998 235775 291050 235827
rect 294454 235775 294506 235827
rect 338518 235775 338570 235827
rect 339478 235775 339530 235827
rect 397366 235775 397418 235827
rect 398230 235775 398282 235827
rect 400246 235775 400298 235827
rect 400342 235775 400394 235827
rect 559222 235775 559274 235827
rect 257974 235701 258026 235753
rect 279190 235701 279242 235753
rect 283894 235701 283946 235753
rect 325846 235701 325898 235753
rect 328918 235701 328970 235753
rect 262006 235627 262058 235679
rect 279286 235627 279338 235679
rect 322486 235627 322538 235679
rect 348886 235627 348938 235679
rect 365014 235627 365066 235679
rect 214198 235553 214250 235605
rect 235318 235553 235370 235605
rect 249718 235553 249770 235605
rect 293782 235553 293834 235605
rect 298006 235553 298058 235605
rect 338326 235553 338378 235605
rect 358006 235553 358058 235605
rect 372118 235553 372170 235605
rect 378646 235701 378698 235753
rect 398518 235701 398570 235753
rect 398614 235701 398666 235753
rect 564310 235701 564362 235753
rect 374518 235627 374570 235679
rect 410710 235627 410762 235679
rect 410806 235627 410858 235679
rect 585238 235627 585290 235679
rect 383062 235553 383114 235605
rect 211030 235479 211082 235531
rect 231574 235479 231626 235531
rect 234262 235479 234314 235531
rect 264886 235479 264938 235531
rect 273430 235479 273482 235531
rect 336502 235479 336554 235531
rect 341206 235479 341258 235531
rect 42166 235405 42218 235457
rect 42934 235405 42986 235457
rect 220630 235405 220682 235457
rect 235894 235405 235946 235457
rect 235990 235405 236042 235457
rect 240694 235405 240746 235457
rect 245206 235405 245258 235457
rect 278230 235405 278282 235457
rect 284758 235405 284810 235457
rect 345622 235405 345674 235457
rect 347638 235405 347690 235457
rect 378646 235405 378698 235457
rect 383062 235405 383114 235457
rect 219382 235331 219434 235383
rect 244534 235331 244586 235383
rect 251158 235331 251210 235383
rect 299254 235331 299306 235383
rect 311542 235331 311594 235383
rect 325270 235331 325322 235383
rect 332182 235331 332234 235383
rect 372886 235331 372938 235383
rect 373078 235331 373130 235383
rect 411574 235553 411626 235605
rect 397654 235479 397706 235531
rect 400246 235479 400298 235531
rect 401782 235479 401834 235531
rect 410614 235479 410666 235531
rect 411766 235479 411818 235531
rect 587446 235479 587498 235531
rect 409174 235405 409226 235457
rect 588886 235405 588938 235457
rect 384406 235331 384458 235383
rect 398806 235331 398858 235383
rect 403606 235331 403658 235383
rect 585142 235331 585194 235383
rect 210070 235257 210122 235309
rect 227830 235257 227882 235309
rect 228406 235257 228458 235309
rect 264022 235257 264074 235309
rect 267478 235257 267530 235309
rect 328342 235257 328394 235309
rect 330454 235257 330506 235309
rect 392854 235257 392906 235309
rect 396310 235257 396362 235309
rect 587350 235257 587402 235309
rect 213430 235183 213482 235235
rect 209302 235109 209354 235161
rect 228502 235109 228554 235161
rect 208918 235035 208970 235087
rect 226966 235035 227018 235087
rect 235702 235183 235754 235235
rect 271126 235183 271178 235235
rect 275254 235183 275306 235235
rect 291094 235183 291146 235235
rect 293494 235183 293546 235235
rect 359926 235183 359978 235235
rect 390838 235183 390890 235235
rect 590134 235183 590186 235235
rect 232918 235109 232970 235161
rect 259030 235109 259082 235161
rect 290710 235109 290762 235161
rect 354358 235109 354410 235161
rect 389782 235109 389834 235161
rect 587926 235109 587978 235161
rect 235798 235035 235850 235087
rect 235894 235035 235946 235087
rect 245014 235035 245066 235087
rect 246646 235035 246698 235087
rect 290902 235035 290954 235087
rect 296086 235035 296138 235087
rect 362710 235035 362762 235087
rect 372886 235035 372938 235087
rect 392086 235035 392138 235087
rect 392278 235035 392330 235087
rect 593110 235035 593162 235087
rect 225142 234961 225194 235013
rect 250582 234961 250634 235013
rect 254230 234961 254282 235013
rect 305110 234961 305162 235013
rect 318358 234961 318410 235013
rect 393910 234961 393962 235013
rect 396694 234961 396746 235013
rect 408310 234961 408362 235013
rect 410422 234961 410474 235013
rect 609046 234961 609098 235013
rect 204406 234887 204458 234939
rect 217942 234887 217994 234939
rect 225526 234887 225578 234939
rect 260182 234887 260234 234939
rect 261910 234887 261962 234939
rect 311062 234887 311114 234939
rect 313078 234887 313130 234939
rect 323446 234887 323498 234939
rect 324406 234887 324458 234939
rect 391414 234887 391466 234939
rect 393046 234887 393098 234939
rect 594646 234887 594698 234939
rect 42166 234813 42218 234865
rect 42838 234813 42890 234865
rect 203254 234813 203306 234865
rect 216502 234813 216554 234865
rect 222358 234813 222410 234865
rect 250486 234813 250538 234865
rect 258742 234813 258794 234865
rect 308182 234813 308234 234865
rect 317110 234813 317162 234865
rect 391510 234813 391562 234865
rect 392662 234813 392714 234865
rect 593974 234813 594026 234865
rect 206998 234739 207050 234791
rect 221782 234739 221834 234791
rect 223894 234739 223946 234791
rect 250774 234739 250826 234791
rect 255766 234739 255818 234791
rect 305782 234739 305834 234791
rect 309334 234739 309386 234791
rect 394198 234739 394250 234791
rect 394390 234739 394442 234791
rect 596950 234739 597002 234791
rect 206518 234665 206570 234717
rect 222454 234665 222506 234717
rect 227062 234665 227114 234717
rect 263254 234665 263306 234717
rect 264406 234665 264458 234717
rect 319606 234665 319658 234717
rect 319894 234665 319946 234717
rect 403414 234665 403466 234717
rect 407734 234665 407786 234717
rect 624118 234665 624170 234717
rect 204790 234591 204842 234643
rect 207286 234591 207338 234643
rect 207862 234591 207914 234643
rect 225526 234591 225578 234643
rect 202870 234517 202922 234569
rect 214870 234517 214922 234569
rect 217846 234517 217898 234569
rect 235990 234591 236042 234643
rect 246550 234591 246602 234643
rect 267958 234591 268010 234643
rect 277558 234591 277610 234643
rect 318166 234591 318218 234643
rect 326230 234591 326282 234643
rect 449302 234591 449354 234643
rect 228790 234517 228842 234569
rect 266230 234517 266282 234569
rect 267094 234517 267146 234569
rect 298198 234517 298250 234569
rect 303478 234517 303530 234569
rect 354262 234517 354314 234569
rect 391222 234517 391274 234569
rect 512662 234517 512714 234569
rect 202006 234443 202058 234495
rect 213430 234443 213482 234495
rect 249334 234443 249386 234495
rect 271030 234443 271082 234495
rect 280630 234443 280682 234495
rect 322198 234443 322250 234495
rect 323542 234443 323594 234495
rect 446326 234443 446378 234495
rect 149398 234369 149450 234421
rect 159862 234369 159914 234421
rect 206134 234369 206186 234421
rect 220918 234369 220970 234421
rect 252598 234369 252650 234421
rect 273622 234369 273674 234421
rect 276118 234369 276170 234421
rect 313942 234369 313994 234421
rect 320278 234369 320330 234421
rect 443446 234369 443498 234421
rect 207382 234295 207434 234347
rect 219382 234295 219434 234347
rect 247414 234295 247466 234347
rect 269398 234295 269450 234347
rect 270262 234295 270314 234347
rect 304342 234295 304394 234347
rect 314422 234295 314474 234347
rect 436150 234295 436202 234347
rect 200278 234221 200330 234273
rect 210358 234221 210410 234273
rect 253462 234221 253514 234273
rect 270838 234221 270890 234273
rect 273046 234221 273098 234273
rect 306646 234221 306698 234273
rect 317206 234221 317258 234273
rect 434902 234221 434954 234273
rect 200182 234147 200234 234199
rect 208822 234147 208874 234199
rect 209686 234147 209738 234199
rect 226294 234147 226346 234199
rect 268534 234147 268586 234199
rect 293974 234147 294026 234199
rect 295702 234147 295754 234199
rect 303574 234147 303626 234199
rect 308470 234147 308522 234199
rect 424054 234147 424106 234199
rect 198742 234073 198794 234125
rect 207382 234073 207434 234125
rect 207478 234073 207530 234125
rect 223990 234073 224042 234125
rect 264310 234073 264362 234125
rect 289846 234073 289898 234125
rect 298966 234073 299018 234125
rect 348502 234073 348554 234125
rect 352150 234073 352202 234125
rect 400438 234073 400490 234125
rect 403510 234073 403562 234125
rect 509782 234073 509834 234125
rect 42070 233999 42122 234051
rect 43030 233999 43082 234051
rect 198358 233999 198410 234051
rect 205942 233999 205994 234051
rect 206902 233999 206954 234051
rect 220246 233999 220298 234051
rect 261238 233999 261290 234051
rect 279670 233999 279722 234051
rect 281206 233999 281258 234051
rect 300790 233999 300842 234051
rect 311158 233999 311210 234051
rect 420406 233999 420458 234051
rect 197494 233925 197546 233977
rect 204310 233925 204362 233977
rect 205174 233925 205226 233977
rect 207286 233925 207338 233977
rect 208726 233925 208778 233977
rect 224758 233925 224810 233977
rect 258358 233925 258410 233977
rect 278134 233925 278186 233977
rect 287062 233925 287114 233977
rect 321142 233925 321194 233977
rect 326134 233925 326186 233977
rect 374614 233925 374666 233977
rect 199126 233851 199178 233903
rect 205078 233851 205130 233903
rect 205558 233851 205610 233903
rect 218710 233851 218762 233903
rect 299350 233851 299402 233903
rect 344662 233851 344714 233903
rect 354934 233851 354986 233903
rect 387190 233925 387242 233977
rect 403318 233925 403370 233977
rect 196918 233777 196970 233829
rect 202870 233777 202922 233829
rect 204214 233777 204266 233829
rect 215542 233777 215594 233829
rect 261622 233777 261674 233829
rect 279286 233777 279338 233829
rect 292918 233777 292970 233829
rect 325462 233777 325514 233829
rect 196534 233703 196586 233755
rect 200566 233703 200618 233755
rect 201526 233703 201578 233755
rect 211894 233703 211946 233755
rect 299830 233703 299882 233755
rect 339862 233777 339914 233829
rect 356758 233777 356810 233829
rect 392086 233851 392138 233903
rect 396982 233851 397034 233903
rect 401206 233851 401258 233903
rect 492502 233925 492554 233977
rect 406198 233851 406250 233903
rect 489622 233851 489674 233903
rect 385366 233777 385418 233829
rect 334966 233703 335018 233755
rect 390358 233703 390410 233755
rect 399478 233703 399530 233755
rect 406198 233703 406250 233755
rect 409558 233777 409610 233829
rect 582550 233777 582602 233829
rect 455254 233703 455306 233755
rect 195670 233629 195722 233681
rect 201334 233629 201386 233681
rect 202486 233629 202538 233681
rect 212566 233629 212618 233681
rect 305206 233629 305258 233681
rect 192886 233555 192938 233607
rect 195286 233555 195338 233607
rect 195574 233555 195626 233607
rect 199798 233555 199850 233607
rect 201046 233555 201098 233607
rect 209686 233555 209738 233607
rect 290326 233555 290378 233607
rect 325174 233555 325226 233607
rect 325462 233555 325514 233607
rect 336310 233555 336362 233607
rect 338326 233629 338378 233681
rect 358486 233629 358538 233681
rect 358582 233629 358634 233681
rect 429142 233629 429194 233681
rect 342934 233555 342986 233607
rect 343510 233555 343562 233607
rect 348694 233555 348746 233607
rect 365686 233555 365738 233607
rect 408982 233555 409034 233607
rect 194230 233481 194282 233533
rect 198358 233481 198410 233533
rect 200662 233481 200714 233533
rect 208150 233481 208202 233533
rect 208438 233481 208490 233533
rect 223222 233481 223274 233533
rect 256534 233481 256586 233533
rect 274678 233481 274730 233533
rect 304438 233481 304490 233533
rect 334006 233481 334058 233533
rect 336694 233481 336746 233533
rect 363958 233481 364010 233533
rect 364054 233481 364106 233533
rect 406102 233481 406154 233533
rect 194614 233407 194666 233459
rect 196054 233407 196106 233459
rect 196150 233407 196202 233459
rect 199126 233407 199178 233459
rect 199702 233407 199754 233459
rect 206614 233407 206666 233459
rect 207286 233407 207338 233459
rect 217174 233407 217226 233459
rect 268918 233407 268970 233459
rect 273430 233407 273482 233459
rect 277942 233407 277994 233459
rect 294454 233407 294506 233459
rect 315766 233407 315818 233459
rect 352822 233407 352874 233459
rect 361270 233407 361322 233459
rect 400342 233407 400394 233459
rect 410038 233407 410090 233459
rect 411670 233407 411722 233459
rect 192406 233333 192458 233385
rect 193750 233333 193802 233385
rect 193846 233333 193898 233385
rect 196822 233333 196874 233385
rect 197974 233333 198026 233385
rect 203638 233333 203690 233385
rect 203926 233333 203978 233385
rect 214198 233333 214250 233385
rect 262870 233333 262922 233385
rect 281206 233333 281258 233385
rect 285718 233333 285770 233385
rect 290710 233333 290762 233385
rect 291574 233333 291626 233385
rect 193462 233259 193514 233311
rect 194614 233259 194666 233311
rect 195190 233259 195242 233311
rect 197494 233259 197546 233311
rect 197878 233259 197930 233311
rect 202102 233259 202154 233311
rect 202390 233259 202442 233311
rect 211126 233259 211178 233311
rect 266134 233259 266186 233311
rect 280918 233259 280970 233311
rect 288502 233259 288554 233311
rect 292822 233259 292874 233311
rect 297238 233333 297290 233385
rect 312694 233333 312746 233385
rect 321718 233333 321770 233385
rect 332086 233333 332138 233385
rect 333430 233333 333482 233385
rect 383158 233333 383210 233385
rect 406294 233333 406346 233385
rect 409174 233333 409226 233385
rect 409942 233333 409994 233385
rect 411766 233333 411818 233385
rect 301558 233259 301610 233311
rect 301654 233259 301706 233311
rect 310198 233259 310250 233311
rect 325174 233259 325226 233311
rect 326902 233259 326954 233311
rect 329302 233259 329354 233311
rect 460726 233259 460778 233311
rect 259126 233185 259178 233237
rect 328150 233185 328202 233237
rect 331606 233185 331658 233237
rect 343414 233185 343466 233237
rect 350326 233185 350378 233237
rect 263542 233111 263594 233163
rect 335734 233111 335786 233163
rect 337942 233111 337994 233163
rect 355318 233111 355370 233163
rect 367222 233185 367274 233237
rect 497974 233185 498026 233237
rect 507094 233111 507146 233163
rect 262102 233037 262154 233089
rect 334198 233037 334250 233089
rect 334294 233037 334346 233089
rect 346294 233037 346346 233089
rect 353110 233037 353162 233089
rect 513142 233111 513194 233163
rect 512662 233037 512714 233089
rect 590902 233037 590954 233089
rect 325366 232963 325418 233015
rect 265174 232889 265226 232941
rect 335446 232889 335498 232941
rect 338038 232889 338090 232941
rect 352342 232889 352394 232941
rect 360790 232963 360842 233015
rect 360886 232963 360938 233015
rect 378934 232963 378986 233015
rect 522166 232963 522218 233015
rect 528310 232889 528362 232941
rect 277462 232815 277514 232867
rect 295606 232815 295658 232867
rect 322486 232815 322538 232867
rect 268438 232741 268490 232793
rect 334294 232741 334346 232793
rect 363382 232815 363434 232867
rect 375382 232815 375434 232867
rect 378454 232815 378506 232867
rect 381430 232815 381482 232867
rect 534262 232815 534314 232867
rect 345526 232741 345578 232793
rect 367222 232741 367274 232793
rect 378838 232741 378890 232793
rect 536566 232741 536618 232793
rect 266614 232667 266666 232719
rect 338230 232667 338282 232719
rect 338326 232667 338378 232719
rect 356086 232667 356138 232719
rect 366646 232667 366698 232719
rect 540310 232667 540362 232719
rect 271606 232593 271658 232645
rect 350038 232593 350090 232645
rect 360790 232593 360842 232645
rect 371254 232593 371306 232645
rect 371830 232593 371882 232645
rect 380182 232593 380234 232645
rect 380278 232593 380330 232645
rect 546358 232593 546410 232645
rect 219766 232519 219818 232571
rect 248086 232519 248138 232571
rect 274870 232519 274922 232571
rect 338326 232519 338378 232571
rect 338422 232519 338474 232571
rect 358294 232519 358346 232571
rect 364918 232519 364970 232571
rect 539542 232519 539594 232571
rect 218230 232445 218282 232497
rect 245110 232445 245162 232497
rect 271222 232445 271274 232497
rect 338038 232445 338090 232497
rect 338710 232445 338762 232497
rect 361270 232445 361322 232497
rect 366262 232445 366314 232497
rect 542614 232445 542666 232497
rect 221014 232371 221066 232423
rect 251158 232371 251210 232423
rect 269686 232371 269738 232423
rect 222550 232297 222602 232349
rect 254230 232297 254282 232349
rect 272950 232297 273002 232349
rect 337942 232297 337994 232349
rect 345622 232371 345674 232423
rect 379510 232371 379562 232423
rect 349366 232297 349418 232349
rect 357622 232297 357674 232349
rect 378934 232297 378986 232349
rect 380182 232297 380234 232349
rect 550870 232297 550922 232349
rect 224278 232223 224330 232275
rect 257206 232223 257258 232275
rect 274198 232223 274250 232275
rect 338326 232223 338378 232275
rect 338422 232223 338474 232275
rect 362038 232223 362090 232275
rect 363190 232223 363242 232275
rect 224374 232149 224426 232201
rect 258742 232149 258794 232201
rect 278998 232149 279050 232201
rect 295510 232149 295562 232201
rect 295606 232149 295658 232201
rect 364438 232149 364490 232201
rect 227446 232075 227498 232127
rect 264790 232075 264842 232127
rect 275734 232075 275786 232127
rect 338710 232075 338762 232127
rect 354262 232075 354314 232127
rect 367126 232075 367178 232127
rect 368086 232223 368138 232275
rect 545590 232223 545642 232275
rect 369910 232149 369962 232201
rect 380278 232149 380330 232201
rect 376438 232075 376490 232127
rect 554710 232149 554762 232201
rect 233206 232001 233258 232053
rect 275350 232001 275402 232053
rect 280246 232001 280298 232053
rect 370390 232001 370442 232053
rect 372310 232001 372362 232053
rect 380662 232075 380714 232127
rect 551638 232075 551690 232127
rect 378454 232001 378506 232053
rect 560758 232001 560810 232053
rect 234838 231927 234890 231979
rect 278326 231927 278378 231979
rect 283510 231927 283562 231979
rect 237622 231853 237674 231905
rect 284374 231853 284426 231905
rect 295510 231927 295562 231979
rect 367414 231927 367466 231979
rect 377206 231927 377258 231979
rect 561430 231927 561482 231979
rect 363190 231853 363242 231905
rect 236086 231779 236138 231831
rect 281302 231779 281354 231831
rect 281974 231779 282026 231831
rect 363382 231779 363434 231831
rect 365110 231779 365162 231831
rect 366934 231853 366986 231905
rect 377110 231853 377162 231905
rect 378550 231853 378602 231905
rect 566710 231853 566762 231905
rect 373462 231779 373514 231831
rect 376822 231779 376874 231831
rect 563638 231779 563690 231831
rect 260278 231705 260330 231757
rect 329590 231705 329642 231757
rect 338230 231705 338282 231757
rect 343222 231705 343274 231757
rect 257494 231631 257546 231683
rect 323638 231631 323690 231683
rect 334870 231631 334922 231683
rect 479158 231705 479210 231757
rect 343414 231631 343466 231683
rect 473110 231631 473162 231683
rect 243862 231557 243914 231609
rect 289750 231557 289802 231609
rect 240598 231483 240650 231535
rect 290422 231557 290474 231609
rect 297142 231557 297194 231609
rect 400246 231557 400298 231609
rect 408982 231557 409034 231609
rect 538870 231557 538922 231609
rect 289942 231483 289994 231535
rect 386326 231483 386378 231535
rect 400342 231483 400394 231535
rect 529750 231483 529802 231535
rect 248374 231409 248426 231461
rect 305494 231409 305546 231461
rect 312214 231409 312266 231461
rect 433846 231409 433898 231461
rect 242134 231335 242186 231387
rect 239350 231261 239402 231313
rect 287446 231261 287498 231313
rect 290902 231335 290954 231387
rect 302518 231335 302570 231387
rect 307606 231335 307658 231387
rect 424726 231335 424778 231387
rect 290806 231261 290858 231313
rect 374518 231261 374570 231313
rect 383062 231261 383114 231313
rect 293494 231187 293546 231239
rect 293878 231187 293930 231239
rect 379990 231187 380042 231239
rect 387766 231187 387818 231239
rect 392566 231187 392618 231239
rect 392854 231187 392906 231239
rect 403222 231261 403274 231313
rect 514678 231261 514730 231313
rect 252982 231113 253034 231165
rect 314518 231113 314570 231165
rect 334006 231113 334058 231165
rect 42070 231039 42122 231091
rect 42742 231039 42794 231091
rect 278230 231039 278282 231091
rect 299446 231039 299498 231091
rect 299542 231039 299594 231091
rect 368662 231039 368714 231091
rect 370774 231039 370826 231091
rect 380662 231039 380714 231091
rect 289750 230965 289802 231017
rect 296470 230965 296522 231017
rect 311062 230965 311114 231017
rect 332662 230965 332714 231017
rect 339862 230965 339914 231017
rect 398710 230965 398762 231017
rect 488950 231187 489002 231239
rect 467830 231039 467882 231091
rect 418774 230965 418826 231017
rect 293782 230891 293834 230943
rect 308182 230891 308234 230943
rect 326710 230891 326762 230943
rect 326806 230891 326858 230943
rect 338326 230891 338378 230943
rect 338518 230891 338570 230943
rect 395350 230891 395402 230943
rect 403414 230891 403466 230943
rect 446614 230891 446666 230943
rect 305782 230817 305834 230869
rect 320662 230817 320714 230869
rect 336310 230817 336362 230869
rect 392374 230817 392426 230869
rect 393910 230817 393962 230869
rect 443734 230817 443786 230869
rect 308566 230743 308618 230795
rect 325846 230743 325898 230795
rect 374230 230743 374282 230795
rect 376150 230743 376202 230795
rect 548566 230743 548618 230795
rect 299254 230669 299306 230721
rect 311638 230669 311690 230721
rect 318166 230669 318218 230721
rect 338422 230669 338474 230721
rect 348502 230669 348554 230721
rect 263926 230595 263978 230647
rect 337270 230595 337322 230647
rect 260662 230521 260714 230573
rect 331222 230521 331274 230573
rect 331318 230521 331370 230573
rect 380278 230595 380330 230647
rect 398710 230669 398762 230721
rect 409654 230669 409706 230721
rect 404470 230595 404522 230647
rect 338326 230521 338378 230573
rect 366934 230521 366986 230573
rect 305110 230447 305162 230499
rect 317590 230447 317642 230499
rect 322198 230447 322250 230499
rect 368086 230521 368138 230573
rect 394198 230521 394250 230573
rect 425590 230595 425642 230647
rect 367126 230447 367178 230499
rect 413494 230447 413546 230499
rect 420406 230447 420458 230499
rect 430102 230447 430154 230499
rect 246166 230373 246218 230425
rect 298678 230373 298730 230425
rect 300214 230373 300266 230425
rect 313270 230373 313322 230425
rect 325750 230373 325802 230425
rect 461014 230373 461066 230425
rect 471286 230373 471338 230425
rect 481462 230373 481514 230425
rect 248950 230299 249002 230351
rect 304822 230299 304874 230351
rect 330262 230299 330314 230351
rect 251926 230225 251978 230277
rect 310774 230225 310826 230277
rect 336214 230225 336266 230277
rect 343702 230299 343754 230351
rect 467062 230299 467114 230351
rect 475222 230299 475274 230351
rect 487510 230299 487562 230351
rect 298198 230151 298250 230203
rect 341014 230151 341066 230203
rect 470134 230225 470186 230277
rect 352726 230151 352778 230203
rect 492502 230151 492554 230203
rect 610486 230151 610538 230203
rect 290998 230077 291050 230129
rect 338038 230077 338090 230129
rect 250294 230003 250346 230055
rect 310006 230003 310058 230055
rect 313942 230003 313994 230055
rect 321622 230003 321674 230055
rect 337558 230003 337610 230055
rect 485206 230077 485258 230129
rect 501046 230077 501098 230129
rect 613558 230077 613610 230129
rect 352726 230003 352778 230055
rect 482134 230003 482186 230055
rect 485590 230003 485642 230055
rect 604534 230003 604586 230055
rect 247030 229929 247082 229981
rect 303958 229929 304010 229981
rect 304342 229929 304394 229981
rect 347158 229929 347210 229981
rect 357238 229929 357290 229981
rect 378934 229929 378986 229981
rect 489622 229929 489674 229981
rect 607510 229929 607562 229981
rect 255190 229855 255242 229907
rect 316822 229855 316874 229907
rect 317974 229855 318026 229907
rect 338518 229855 338570 229907
rect 343990 229855 344042 229907
rect 495094 229855 495146 229907
rect 254806 229781 254858 229833
rect 319126 229781 319178 229833
rect 323446 229781 323498 229833
rect 338422 229781 338474 229833
rect 347062 229781 347114 229833
rect 501046 229781 501098 229833
rect 506134 229781 506186 229833
rect 516118 229781 516170 229833
rect 245686 229707 245738 229759
rect 300982 229707 301034 229759
rect 306646 229707 306698 229759
rect 251542 229633 251594 229685
rect 313078 229633 313130 229685
rect 313270 229707 313322 229759
rect 407446 229707 407498 229759
rect 416950 229707 417002 229759
rect 572086 229707 572138 229759
rect 220150 229559 220202 229611
rect 249718 229559 249770 229611
rect 257590 229559 257642 229611
rect 325174 229559 325226 229611
rect 325270 229559 325322 229611
rect 338326 229559 338378 229611
rect 351766 229633 351818 229685
rect 353110 229559 353162 229611
rect 354838 229559 354890 229611
rect 506134 229559 506186 229611
rect 509782 229633 509834 229685
rect 614998 229633 615050 229685
rect 510166 229559 510218 229611
rect 516214 229559 516266 229611
rect 618070 229559 618122 229611
rect 222934 229485 222986 229537
rect 255670 229485 255722 229537
rect 259798 229485 259850 229537
rect 321430 229485 321482 229537
rect 221590 229411 221642 229463
rect 252598 229411 252650 229463
rect 256150 229411 256202 229463
rect 322102 229485 322154 229537
rect 328534 229485 328586 229537
rect 343702 229485 343754 229537
rect 362134 229485 362186 229537
rect 321622 229411 321674 229463
rect 359158 229411 359210 229463
rect 365398 229411 365450 229463
rect 378934 229485 378986 229537
rect 524470 229485 524522 229537
rect 216694 229337 216746 229389
rect 242134 229337 242186 229389
rect 242806 229337 242858 229389
rect 294934 229337 294986 229389
rect 296566 229337 296618 229389
rect 361366 229337 361418 229389
rect 368182 229337 368234 229389
rect 531286 229411 531338 229463
rect 226198 229263 226250 229315
rect 261718 229263 261770 229315
rect 262774 229263 262826 229315
rect 321334 229263 321386 229315
rect 321430 229263 321482 229315
rect 325846 229263 325898 229315
rect 333046 229263 333098 229315
rect 344758 229263 344810 229315
rect 231958 229189 232010 229241
rect 273814 229189 273866 229241
rect 287926 229189 287978 229241
rect 235222 229115 235274 229167
rect 279862 229115 279914 229167
rect 286294 229115 286346 229167
rect 239734 229041 239786 229093
rect 288886 229041 288938 229093
rect 289366 229115 289418 229167
rect 306646 229189 306698 229241
rect 367030 229189 367082 229241
rect 371542 229263 371594 229315
rect 537238 229337 537290 229389
rect 543382 229263 543434 229315
rect 564406 229263 564458 229315
rect 606742 229263 606794 229315
rect 372694 229189 372746 229241
rect 552406 229189 552458 229241
rect 559222 229189 559274 229241
rect 603670 229189 603722 229241
rect 374422 229115 374474 229167
rect 375766 229115 375818 229167
rect 558454 229115 558506 229167
rect 564310 229115 564362 229167
rect 605302 229115 605354 229167
rect 215254 228967 215306 229019
rect 239062 228967 239114 229019
rect 244150 228967 244202 229019
rect 298006 228967 298058 229019
rect 378742 229041 378794 229093
rect 564502 229041 564554 229093
rect 306646 228967 306698 229019
rect 312694 228967 312746 229019
rect 316246 228967 316298 229019
rect 241078 228893 241130 228945
rect 291958 228893 292010 228945
rect 298390 228893 298442 228945
rect 406006 228967 406058 229019
rect 408310 228967 408362 229019
rect 601462 228967 601514 229019
rect 321334 228893 321386 228945
rect 331894 228893 331946 228945
rect 243190 228819 243242 228871
rect 292630 228819 292682 228871
rect 295318 228819 295370 228871
rect 332470 228819 332522 228871
rect 228886 228745 228938 228797
rect 267862 228745 267914 228797
rect 274678 228745 274730 228797
rect 319894 228745 319946 228797
rect 322390 228745 322442 228797
rect 455158 228893 455210 228945
rect 455254 228893 455306 228945
rect 578038 228893 578090 228945
rect 338710 228819 338762 228871
rect 394582 228819 394634 228871
rect 406102 228819 406154 228871
rect 535798 228819 535850 228871
rect 230806 228671 230858 228723
rect 270742 228671 270794 228723
rect 270838 228671 270890 228723
rect 313846 228671 313898 228723
rect 321238 228671 321290 228723
rect 451990 228745 452042 228797
rect 338518 228671 338570 228723
rect 445942 228671 445994 228723
rect 231670 228597 231722 228649
rect 272278 228597 272330 228649
rect 272374 228597 272426 228649
rect 307702 228597 307754 228649
rect 313462 228597 313514 228649
rect 436918 228597 436970 228649
rect 230326 228523 230378 228575
rect 269302 228523 269354 228575
rect 269398 228523 269450 228575
rect 301750 228523 301802 228575
rect 308950 228523 309002 228575
rect 427798 228523 427850 228575
rect 429142 228523 429194 228575
rect 526006 228523 526058 228575
rect 538582 228523 538634 228575
rect 541078 228523 541130 228575
rect 561718 228523 561770 228575
rect 562966 228523 563018 228575
rect 567382 228523 567434 228575
rect 569014 228523 569066 228575
rect 268150 228449 268202 228501
rect 295702 228449 295754 228501
rect 306166 228449 306218 228501
rect 421846 228449 421898 228501
rect 455062 228449 455114 228501
rect 456502 228449 456554 228501
rect 466486 228449 466538 228501
rect 475318 228449 475370 228501
rect 483862 228449 483914 228501
rect 485974 228449 486026 228501
rect 266326 228375 266378 228427
rect 289750 228375 289802 228427
rect 289846 228375 289898 228427
rect 334966 228375 335018 228427
rect 340822 228375 340874 228427
rect 344566 228375 344618 228427
rect 344758 228375 344810 228427
rect 476182 228375 476234 228427
rect 483766 228375 483818 228427
rect 493462 228375 493514 228427
rect 262006 228301 262058 228353
rect 276790 228301 276842 228353
rect 279190 228301 279242 228353
rect 322966 228301 323018 228353
rect 338326 228301 338378 228353
rect 432406 228301 432458 228353
rect 449302 228301 449354 228353
rect 460246 228301 460298 228353
rect 264694 228227 264746 228279
rect 285910 228227 285962 228279
rect 291478 228227 291530 228279
rect 389302 228227 389354 228279
rect 400438 228227 400490 228279
rect 511606 228227 511658 228279
rect 248758 228153 248810 228205
rect 307030 228153 307082 228205
rect 310198 228153 310250 228205
rect 412726 228153 412778 228205
rect 303574 228079 303626 228131
rect 398326 228079 398378 228131
rect 400630 228079 400682 228131
rect 492022 228079 492074 228131
rect 288406 228005 288458 228057
rect 383254 228005 383306 228057
rect 396982 228005 397034 228057
rect 470902 228005 470954 228057
rect 253078 227931 253130 227983
rect 316150 227931 316202 227983
rect 316246 227931 316298 227983
rect 401398 227931 401450 227983
rect 434902 227931 434954 227983
rect 442198 227931 442250 227983
rect 292534 227857 292586 227909
rect 380086 227857 380138 227909
rect 391414 227857 391466 227909
rect 455734 227857 455786 227909
rect 301174 227783 301226 227835
rect 363286 227783 363338 227835
rect 391510 227783 391562 227835
rect 440662 227783 440714 227835
rect 292150 227709 292202 227761
rect 354262 227709 354314 227761
rect 385846 227709 385898 227761
rect 401974 227709 402026 227761
rect 407158 227709 407210 227761
rect 413206 227709 413258 227761
rect 446326 227709 446378 227761
rect 454294 227709 454346 227761
rect 293974 227635 294026 227687
rect 343990 227635 344042 227687
rect 344566 227635 344618 227687
rect 491254 227635 491306 227687
rect 279670 227561 279722 227613
rect 328918 227561 328970 227613
rect 338422 227561 338474 227613
rect 435382 227561 435434 227613
rect 443446 227561 443498 227613
rect 448246 227561 448298 227613
rect 460726 227561 460778 227613
rect 466390 227561 466442 227613
rect 190006 227487 190058 227539
rect 191542 227487 191594 227539
rect 228022 227487 228074 227539
rect 262486 227487 262538 227539
rect 291094 227487 291146 227539
rect 357622 227487 357674 227539
rect 392182 227487 392234 227539
rect 226582 227413 226634 227465
rect 259414 227413 259466 227465
rect 282358 227413 282410 227465
rect 351574 227413 351626 227465
rect 354262 227413 354314 227465
rect 393142 227413 393194 227465
rect 395062 227487 395114 227539
rect 584854 227487 584906 227539
rect 585238 227487 585290 227539
rect 630166 227487 630218 227539
rect 592342 227413 592394 227465
rect 606166 227413 606218 227465
rect 232918 227339 232970 227391
rect 261046 227339 261098 227391
rect 294454 227339 294506 227391
rect 363670 227339 363722 227391
rect 390070 227339 390122 227391
rect 390454 227339 390506 227391
rect 407638 227339 407690 227391
rect 407830 227339 407882 227391
rect 585622 227339 585674 227391
rect 588982 227339 589034 227391
rect 599158 227339 599210 227391
rect 639958 227339 640010 227391
rect 229558 227265 229610 227317
rect 265558 227265 265610 227317
rect 267958 227265 268010 227317
rect 300214 227265 300266 227317
rect 300790 227265 300842 227317
rect 369622 227265 369674 227317
rect 371542 227265 371594 227317
rect 385558 227265 385610 227317
rect 407158 227265 407210 227317
rect 413206 227265 413258 227317
rect 588598 227265 588650 227317
rect 600502 227265 600554 227317
rect 634678 227265 634730 227317
rect 229750 227191 229802 227243
rect 266998 227191 267050 227243
rect 273430 227191 273482 227243
rect 345526 227191 345578 227243
rect 354358 227191 354410 227243
rect 390070 227191 390122 227243
rect 394966 227191 395018 227243
rect 231094 227117 231146 227169
rect 268534 227117 268586 227169
rect 270646 227117 270698 227169
rect 348598 227117 348650 227169
rect 359926 227117 359978 227169
rect 396118 227117 396170 227169
rect 399958 227191 400010 227243
rect 407350 227191 407402 227243
rect 407638 227191 407690 227243
rect 589366 227191 589418 227243
rect 596182 227191 596234 227243
rect 633142 227191 633194 227243
rect 598486 227117 598538 227169
rect 603382 227117 603434 227169
rect 638518 227117 638570 227169
rect 233878 227043 233930 227095
rect 274486 227043 274538 227095
rect 276694 227043 276746 227095
rect 360598 227043 360650 227095
rect 394870 227043 394922 227095
rect 597718 227043 597770 227095
rect 232534 226969 232586 227021
rect 271606 226969 271658 227021
rect 279766 226969 279818 227021
rect 366742 226969 366794 227021
rect 368662 226969 368714 227021
rect 408214 226969 408266 227021
rect 410614 226969 410666 227021
rect 612118 226969 612170 227021
rect 235606 226895 235658 226947
rect 277558 226895 277610 226947
rect 282550 226895 282602 226947
rect 372694 226895 372746 226947
rect 374518 226895 374570 226947
rect 390742 226895 390794 226947
rect 401974 226895 402026 226947
rect 406486 226895 406538 226947
rect 407350 226895 407402 226947
rect 418966 226895 419018 226947
rect 419254 226895 419306 226947
rect 609814 226895 609866 226947
rect 213046 226821 213098 226873
rect 233782 226821 233834 226873
rect 237430 226821 237482 226873
rect 282070 226821 282122 226873
rect 301558 226821 301610 226873
rect 390838 226821 390890 226873
rect 401686 226821 401738 226873
rect 213814 226747 213866 226799
rect 237526 226747 237578 226799
rect 238390 226747 238442 226799
rect 252214 226747 252266 226799
rect 214582 226673 214634 226725
rect 236854 226673 236906 226725
rect 280630 226747 280682 226799
rect 290710 226747 290762 226799
rect 216118 226599 216170 226651
rect 239830 226599 239882 226651
rect 240118 226599 240170 226651
rect 247702 226599 247754 226651
rect 212374 226525 212426 226577
rect 234550 226525 234602 226577
rect 237046 226525 237098 226577
rect 252406 226673 252458 226725
rect 282934 226673 282986 226725
rect 283990 226673 284042 226725
rect 358486 226673 358538 226725
rect 388150 226747 388202 226799
rect 395062 226747 395114 226799
rect 400822 226747 400874 226799
rect 413206 226747 413258 226799
rect 611254 226821 611306 226873
rect 419158 226747 419210 226799
rect 608950 226747 609002 226799
rect 609046 226747 609098 226799
rect 629398 226747 629450 226799
rect 378742 226673 378794 226725
rect 379990 226673 380042 226725
rect 397654 226673 397706 226725
rect 402838 226673 402890 226725
rect 247894 226599 247946 226651
rect 286678 226599 286730 226651
rect 292822 226599 292874 226651
rect 384790 226599 384842 226651
rect 388534 226599 388586 226651
rect 407638 226599 407690 226651
rect 407734 226599 407786 226651
rect 418870 226599 418922 226651
rect 419062 226673 419114 226725
rect 608278 226673 608330 226725
rect 609142 226673 609194 226725
rect 630934 226673 630986 226725
rect 614326 226599 614378 226651
rect 247990 226525 248042 226577
rect 221686 226451 221738 226503
rect 250390 226451 250442 226503
rect 252214 226525 252266 226577
rect 283606 226525 283658 226577
rect 293110 226525 293162 226577
rect 393814 226525 393866 226577
rect 406678 226525 406730 226577
rect 621814 226525 621866 226577
rect 303190 226451 303242 226503
rect 304246 226451 304298 226503
rect 409558 226451 409610 226503
rect 217462 226377 217514 226429
rect 215734 226303 215786 226355
rect 238390 226303 238442 226355
rect 240214 226377 240266 226429
rect 288118 226377 288170 226429
rect 294838 226377 294890 226429
rect 396886 226377 396938 226429
rect 397558 226377 397610 226429
rect 411958 226451 412010 226503
rect 413206 226451 413258 226503
rect 419254 226451 419306 226503
rect 588886 226451 588938 226503
rect 626422 226451 626474 226503
rect 629206 226451 629258 226503
rect 634006 226451 634058 226503
rect 409750 226377 409802 226429
rect 619606 226377 619658 226429
rect 241270 226303 241322 226355
rect 243286 226303 243338 226355
rect 217078 226229 217130 226281
rect 243574 226229 243626 226281
rect 244918 226229 244970 226281
rect 250870 226303 250922 226355
rect 285142 226303 285194 226355
rect 297622 226303 297674 226355
rect 402838 226303 402890 226355
rect 407254 226303 407306 226355
rect 622678 226303 622730 226355
rect 218326 226155 218378 226207
rect 246646 226155 246698 226207
rect 294262 226229 294314 226281
rect 295222 226229 295274 226281
rect 399094 226229 399146 226281
rect 400246 226229 400298 226281
rect 403702 226229 403754 226281
rect 297238 226155 297290 226207
rect 302134 226155 302186 226207
rect 397558 226155 397610 226207
rect 215638 226081 215690 226133
rect 240598 226081 240650 226133
rect 241846 226081 241898 226133
rect 291190 226081 291242 226133
rect 300886 226081 300938 226133
rect 408982 226155 409034 226207
rect 397750 226081 397802 226133
rect 415030 226229 415082 226281
rect 418870 226229 418922 226281
rect 623350 226229 623402 226281
rect 412150 226155 412202 226207
rect 632374 226155 632426 226207
rect 411766 226081 411818 226133
rect 627862 226081 627914 226133
rect 226678 226007 226730 226059
rect 232918 226007 232970 226059
rect 250774 226007 250826 226059
rect 254902 226007 254954 226059
rect 264886 226007 264938 226059
rect 276118 226007 276170 226059
rect 224950 225933 225002 225985
rect 256438 225933 256490 225985
rect 257110 225933 257162 225985
rect 321334 226007 321386 226059
rect 326902 226007 326954 226059
rect 387766 226007 387818 226059
rect 321142 225933 321194 225985
rect 381814 225933 381866 225985
rect 387670 225933 387722 225985
rect 583414 226007 583466 226059
rect 587446 226007 587498 226059
rect 631702 226007 631754 226059
rect 389494 225933 389546 225985
rect 587158 225933 587210 225985
rect 600406 225933 600458 225985
rect 636214 225933 636266 225985
rect 218806 225859 218858 225911
rect 244342 225859 244394 225911
rect 253846 225859 253898 225911
rect 315382 225859 315434 225911
rect 335446 225859 335498 225911
rect 340246 225859 340298 225911
rect 341974 225859 342026 225911
rect 384022 225859 384074 225911
rect 387382 225859 387434 225911
rect 220342 225785 220394 225837
rect 247414 225785 247466 225837
rect 238774 225711 238826 225763
rect 250870 225785 250922 225837
rect 251062 225785 251114 225837
rect 250582 225711 250634 225763
rect 257974 225711 258026 225763
rect 271126 225785 271178 225837
rect 279094 225785 279146 225837
rect 280918 225785 280970 225837
rect 339478 225785 339530 225837
rect 374422 225785 374474 225837
rect 388630 225785 388682 225837
rect 388918 225859 388970 225911
rect 586390 225859 586442 225911
rect 603286 225859 603338 225911
rect 639190 225859 639242 225911
rect 582646 225785 582698 225837
rect 603574 225785 603626 225837
rect 636886 225785 636938 225837
rect 309334 225711 309386 225763
rect 319606 225711 319658 225763
rect 336406 225711 336458 225763
rect 336502 225711 336554 225763
rect 354550 225711 354602 225763
rect 358486 225711 358538 225763
rect 375766 225711 375818 225763
rect 390742 225711 390794 225763
rect 391510 225711 391562 225763
rect 392566 225711 392618 225763
rect 223318 225637 223370 225689
rect 253462 225637 253514 225689
rect 253558 225637 253610 225689
rect 269974 225637 270026 225689
rect 281206 225637 281258 225689
rect 333526 225637 333578 225689
rect 380086 225637 380138 225689
rect 394390 225637 394442 225689
rect 394870 225711 394922 225763
rect 406486 225711 406538 225763
rect 580342 225711 580394 225763
rect 603478 225711 603530 225763
rect 236470 225563 236522 225615
rect 252406 225563 252458 225615
rect 259030 225563 259082 225615
rect 273046 225563 273098 225615
rect 279286 225563 279338 225615
rect 330454 225563 330506 225615
rect 367030 225563 367082 225615
rect 382582 225563 382634 225615
rect 386614 225563 386666 225615
rect 394486 225563 394538 225615
rect 394582 225563 394634 225615
rect 397846 225563 397898 225615
rect 581110 225637 581162 225689
rect 585142 225637 585194 225689
rect 615862 225637 615914 225689
rect 626326 225711 626378 225763
rect 635446 225711 635498 225763
rect 637750 225637 637802 225689
rect 584086 225563 584138 225615
rect 587350 225563 587402 225615
rect 600790 225563 600842 225615
rect 273718 225489 273770 225541
rect 318358 225489 318410 225541
rect 318934 225489 318986 225541
rect 445174 225489 445226 225541
rect 582550 225489 582602 225541
rect 627190 225489 627242 225541
rect 273622 225415 273674 225467
rect 312310 225415 312362 225467
rect 312982 225415 313034 225467
rect 433174 225415 433226 225467
rect 278134 225341 278186 225393
rect 324406 225341 324458 225393
rect 332086 225341 332138 225393
rect 451222 225341 451274 225393
rect 271030 225267 271082 225319
rect 306262 225267 306314 225319
rect 309910 225267 309962 225319
rect 427030 225267 427082 225319
rect 306742 225193 306794 225245
rect 420982 225193 421034 225245
rect 303862 225119 303914 225171
rect 397750 225119 397802 225171
rect 397846 225119 397898 225171
rect 400630 225119 400682 225171
rect 415414 225119 415466 225171
rect 628630 225119 628682 225171
rect 259894 225045 259946 225097
rect 327382 225045 327434 225097
rect 328342 225045 328394 225097
rect 342550 225045 342602 225097
rect 342934 225045 342986 225097
rect 418006 225045 418058 225097
rect 670006 225045 670058 225097
rect 676246 225045 676298 225097
rect 344662 224971 344714 225023
rect 405910 224971 405962 225023
rect 406006 224971 406058 225023
rect 406774 224971 406826 225023
rect 409558 224971 409610 225023
rect 417238 224971 417290 225023
rect 189910 224897 189962 224949
rect 192310 224897 192362 224949
rect 363286 224897 363338 224949
rect 411286 224897 411338 224949
rect 250486 224823 250538 224875
rect 251926 224823 251978 224875
rect 358582 224823 358634 224875
rect 405142 224823 405194 224875
rect 405526 224823 405578 224875
rect 409750 224823 409802 224875
rect 245014 224749 245066 224801
rect 248854 224749 248906 224801
rect 361366 224749 361418 224801
rect 402166 224749 402218 224801
rect 185686 224675 185738 224727
rect 187126 224675 187178 224727
rect 190774 224675 190826 224727
rect 240694 224675 240746 224727
rect 242902 224675 242954 224727
rect 244534 224675 244586 224727
rect 245878 224675 245930 224727
rect 362710 224675 362762 224727
rect 399958 224675 400010 224727
rect 400054 224675 400106 224727
rect 419062 224675 419114 224727
rect 289078 224601 289130 224653
rect 386998 224601 387050 224653
rect 387286 224601 387338 224653
rect 517654 224601 517706 224653
rect 322294 224527 322346 224579
rect 453430 224527 453482 224579
rect 325078 224453 325130 224505
rect 459574 224453 459626 224505
rect 331510 224379 331562 224431
rect 471574 224379 471626 224431
rect 328246 224305 328298 224357
rect 465622 224305 465674 224357
rect 661366 224305 661418 224357
rect 676054 224305 676106 224357
rect 275638 224231 275690 224283
rect 359926 224231 359978 224283
rect 362806 224231 362858 224283
rect 498838 224231 498890 224283
rect 337174 224157 337226 224209
rect 483766 224157 483818 224209
rect 334486 224083 334538 224135
rect 477622 224083 477674 224135
rect 338134 224009 338186 224061
rect 482902 224009 482954 224061
rect 340438 223935 340490 223987
rect 489718 223935 489770 223987
rect 346678 223861 346730 223913
rect 358774 223861 358826 223913
rect 497302 223861 497354 223913
rect 503350 223787 503402 223839
rect 663862 223787 663914 223839
rect 676054 223787 676106 223839
rect 347926 223713 347978 223765
rect 266518 223639 266570 223691
rect 341782 223639 341834 223691
rect 264598 223565 264650 223617
rect 338710 223565 338762 223617
rect 361654 223713 361706 223765
rect 501814 223713 501866 223765
rect 349942 223639 349994 223691
rect 509398 223639 509450 223691
rect 504790 223565 504842 223617
rect 268054 223491 268106 223543
rect 344854 223491 344906 223543
rect 350806 223491 350858 223543
rect 364534 223491 364586 223543
rect 364630 223491 364682 223543
rect 507862 223491 507914 223543
rect 269590 223417 269642 223469
rect 347734 223417 347786 223469
rect 353014 223417 353066 223469
rect 515350 223417 515402 223469
rect 270934 223343 270986 223395
rect 350806 223343 350858 223395
rect 352534 223343 352586 223395
rect 272566 223269 272618 223321
rect 353878 223269 353930 223321
rect 355606 223269 355658 223321
rect 364534 223343 364586 223395
rect 510838 223343 510890 223395
rect 274102 223195 274154 223247
rect 356854 223195 356906 223247
rect 513910 223269 513962 223321
rect 519862 223195 519914 223247
rect 321718 223121 321770 223173
rect 449686 223121 449738 223173
rect 319414 223047 319466 223099
rect 447478 223047 447530 223099
rect 316342 222973 316394 223025
rect 441430 222973 441482 223025
rect 315286 222899 315338 222951
rect 437686 222899 437738 222951
rect 310294 222825 310346 222877
rect 429334 222825 429386 222877
rect 308854 222751 308906 222803
rect 426358 222751 426410 222803
rect 312598 222677 312650 222729
rect 431542 222677 431594 222729
rect 277078 222603 277130 222655
rect 362902 222603 362954 222655
rect 363958 222603 364010 222655
rect 479926 222603 479978 222655
rect 307894 222529 307946 222581
rect 422518 222529 422570 222581
rect 306550 222455 306602 222507
rect 419542 222455 419594 222507
rect 302806 222381 302858 222433
rect 414262 222381 414314 222433
rect 305878 222307 305930 222359
rect 420214 222307 420266 222359
rect 284662 222233 284714 222285
rect 378070 222233 378122 222285
rect 398518 222233 398570 222285
rect 502582 222233 502634 222285
rect 343606 222159 343658 222211
rect 358774 222159 358826 222211
rect 374614 222159 374666 222211
rect 458806 222159 458858 222211
rect 283126 222085 283178 222137
rect 374998 222085 375050 222137
rect 349558 222011 349610 222063
rect 364630 222011 364682 222063
rect 157078 221715 157130 221767
rect 184342 221715 184394 221767
rect 498262 221715 498314 221767
rect 499558 221715 499610 221767
rect 504214 221715 504266 221767
rect 506374 221715 506426 221767
rect 541558 221715 541610 221767
rect 544102 221715 544154 221767
rect 553222 221715 553274 221767
rect 555286 221715 555338 221767
rect 576022 221715 576074 221767
rect 577318 221715 577370 221767
rect 645142 221271 645194 221323
rect 650038 221271 650090 221323
rect 149590 218903 149642 218955
rect 165526 218903 165578 218955
rect 147382 216831 147434 216883
rect 151510 216831 151562 216883
rect 645142 216831 645194 216883
rect 649942 216831 649994 216883
rect 41590 216461 41642 216513
rect 45142 216461 45194 216513
rect 674806 216387 674858 216439
rect 676054 216387 676106 216439
rect 147286 216239 147338 216291
rect 151222 216239 151274 216291
rect 41782 215721 41834 215773
rect 44950 215721 45002 215773
rect 41782 215203 41834 215255
rect 45238 215203 45290 215255
rect 41590 214981 41642 215033
rect 43510 214981 43562 215033
rect 674422 214907 674474 214959
rect 676054 214907 676106 214959
rect 41782 214241 41834 214293
rect 45334 214241 45386 214293
rect 41782 213649 41834 213701
rect 44662 213649 44714 213701
rect 41782 213279 41834 213331
rect 43222 213279 43274 213331
rect 147382 213279 147434 213331
rect 151414 213279 151466 213331
rect 674518 213279 674570 213331
rect 675958 213279 676010 213331
rect 674614 213205 674666 213257
rect 676246 213205 676298 213257
rect 149494 213131 149546 213183
rect 182806 213131 182858 213183
rect 674710 213131 674762 213183
rect 676054 213131 676106 213183
rect 41590 212909 41642 212961
rect 44566 212909 44618 212961
rect 645142 212909 645194 212961
rect 649846 212909 649898 212961
rect 147094 212465 147146 212517
rect 151702 212465 151754 212517
rect 41782 212169 41834 212221
rect 43414 212169 43466 212221
rect 147382 210319 147434 210371
rect 151318 210319 151370 210371
rect 149494 210245 149546 210297
rect 179926 210245 179978 210297
rect 646582 210245 646634 210297
rect 679798 210245 679850 210297
rect 645142 209801 645194 209853
rect 649750 209801 649802 209853
rect 147286 207433 147338 207485
rect 151606 207433 151658 207485
rect 149494 207359 149546 207411
rect 177046 207359 177098 207411
rect 41878 206175 41930 206227
rect 42742 206175 42794 206227
rect 645142 206027 645194 206079
rect 649654 206027 649706 206079
rect 675766 205953 675818 206005
rect 41782 205879 41834 205931
rect 43126 205879 43178 205931
rect 675766 205731 675818 205783
rect 41590 205139 41642 205191
rect 42934 205139 42986 205191
rect 41686 204917 41738 204969
rect 45046 204917 45098 204969
rect 41590 204843 41642 204895
rect 42838 204843 42890 204895
rect 41782 204547 41834 204599
rect 43030 204547 43082 204599
rect 149494 204547 149546 204599
rect 168598 204547 168650 204599
rect 149302 204473 149354 204525
rect 174262 204473 174314 204525
rect 41782 204325 41834 204377
rect 44758 204325 44810 204377
rect 41782 203733 41834 203785
rect 44854 203733 44906 203785
rect 674806 202031 674858 202083
rect 675478 202031 675530 202083
rect 149686 201661 149738 201713
rect 180022 201661 180074 201713
rect 149494 201587 149546 201639
rect 182902 201587 182954 201639
rect 145750 201513 145802 201565
rect 184342 201513 184394 201565
rect 645142 201513 645194 201565
rect 649558 201513 649610 201565
rect 674710 200847 674762 200899
rect 675382 200847 675434 200899
rect 149302 198775 149354 198827
rect 159958 198775 160010 198827
rect 149494 198701 149546 198753
rect 177142 198701 177194 198753
rect 181366 198627 181418 198679
rect 184342 198627 184394 198679
rect 148918 198553 148970 198605
rect 149494 198553 149546 198605
rect 178486 198553 178538 198605
rect 184438 198553 184490 198605
rect 645142 198479 645194 198531
rect 649462 198479 649514 198531
rect 148918 198405 148970 198457
rect 149686 198405 149738 198457
rect 674614 197591 674666 197643
rect 675382 197591 675434 197643
rect 42070 197369 42122 197421
rect 42070 197147 42122 197199
rect 674422 196999 674474 197051
rect 675478 196999 675530 197051
rect 42742 196851 42794 196903
rect 43222 196851 43274 196903
rect 674518 196555 674570 196607
rect 675382 196555 675434 196607
rect 149302 195889 149354 195941
rect 162742 195889 162794 195941
rect 149686 195815 149738 195867
rect 171286 195815 171338 195867
rect 166966 195741 167018 195793
rect 184534 195741 184586 195793
rect 169846 195667 169898 195719
rect 184438 195667 184490 195719
rect 172726 195593 172778 195645
rect 184342 195593 184394 195645
rect 149398 194631 149450 194683
rect 157078 194631 157130 194683
rect 645142 193965 645194 194017
rect 649366 193965 649418 194017
rect 42070 193447 42122 193499
rect 42934 193447 42986 193499
rect 149398 193003 149450 193055
rect 154102 193003 154154 193055
rect 152566 192929 152618 192981
rect 184630 192929 184682 192981
rect 155446 192855 155498 192907
rect 184534 192855 184586 192907
rect 158326 192781 158378 192833
rect 184342 192781 184394 192833
rect 164086 192707 164138 192759
rect 184438 192707 184490 192759
rect 42166 192189 42218 192241
rect 42838 192189 42890 192241
rect 42070 191449 42122 191501
rect 43126 191449 43178 191501
rect 42166 191005 42218 191057
rect 43030 191005 43082 191057
rect 645142 190413 645194 190465
rect 653782 190413 653834 190465
rect 147574 190191 147626 190243
rect 151798 190191 151850 190243
rect 143158 190043 143210 190095
rect 184630 190043 184682 190095
rect 143254 189969 143306 190021
rect 184534 189969 184586 190021
rect 145366 189895 145418 189947
rect 184438 189895 184490 189947
rect 148918 189821 148970 189873
rect 184342 189821 184394 189873
rect 146902 188785 146954 188837
rect 147286 188785 147338 188837
rect 42166 187823 42218 187875
rect 43222 187823 43274 187875
rect 149398 187231 149450 187283
rect 165622 187231 165674 187283
rect 143158 187157 143210 187209
rect 184438 187157 184490 187209
rect 143350 187083 143402 187135
rect 184630 187083 184682 187135
rect 143254 187009 143306 187061
rect 184342 187009 184394 187061
rect 168502 186935 168554 186987
rect 184534 186935 184586 186987
rect 646198 184567 646250 184619
rect 660886 184567 660938 184619
rect 149398 184345 149450 184397
rect 168694 184345 168746 184397
rect 145654 184271 145706 184323
rect 184534 184271 184586 184323
rect 145558 184197 145610 184249
rect 184342 184197 184394 184249
rect 156886 184123 156938 184175
rect 184630 184123 184682 184175
rect 162646 184049 162698 184101
rect 184438 184049 184490 184101
rect 645910 183087 645962 183139
rect 658294 183087 658346 183139
rect 149398 181459 149450 181511
rect 171382 181459 171434 181511
rect 143062 181385 143114 181437
rect 184630 181385 184682 181437
rect 151126 181311 151178 181363
rect 184534 181311 184586 181363
rect 154006 181237 154058 181289
rect 184342 181237 184394 181289
rect 159766 181163 159818 181215
rect 184438 181163 184490 181215
rect 149398 179535 149450 179587
rect 156886 179535 156938 179587
rect 646006 179387 646058 179439
rect 658486 179387 658538 179439
rect 666646 179313 666698 179365
rect 676054 179313 676106 179365
rect 147382 178795 147434 178847
rect 154198 178795 154250 178847
rect 661462 178795 661514 178847
rect 676054 178795 676106 178847
rect 655318 178647 655370 178699
rect 676246 178647 676298 178699
rect 149686 178573 149738 178625
rect 162646 178573 162698 178625
rect 143062 178499 143114 178551
rect 184438 178499 184490 178551
rect 148918 178425 148970 178477
rect 149686 178425 149738 178477
rect 143062 178351 143114 178403
rect 143158 178277 143210 178329
rect 184534 178425 184586 178477
rect 184342 178351 184394 178403
rect 147190 176723 147242 176775
rect 151126 176723 151178 176775
rect 145462 175613 145514 175665
rect 184342 175613 184394 175665
rect 156982 175539 157034 175591
rect 184438 175539 184490 175591
rect 645142 174873 645194 174925
rect 655222 174873 655274 174925
rect 674518 172875 674570 172927
rect 676054 172875 676106 172927
rect 674806 172801 674858 172853
rect 676246 172801 676298 172853
rect 148246 172727 148298 172779
rect 184438 172727 184490 172779
rect 148726 172653 148778 172705
rect 184534 172653 184586 172705
rect 168406 172579 168458 172631
rect 184342 172579 184394 172631
rect 645142 171395 645194 171447
rect 652342 171395 652394 171447
rect 147286 170359 147338 170411
rect 148246 170359 148298 170411
rect 674614 169989 674666 170041
rect 675958 169989 676010 170041
rect 149398 169915 149450 169967
rect 180118 169915 180170 169967
rect 674710 169915 674762 169967
rect 676054 169915 676106 169967
rect 148534 169841 148586 169893
rect 184438 169841 184490 169893
rect 148342 169767 148394 169819
rect 184534 169767 184586 169819
rect 149014 169693 149066 169745
rect 184630 169693 184682 169745
rect 174166 169619 174218 169671
rect 184342 169619 184394 169671
rect 645142 167991 645194 168043
rect 652822 167991 652874 168043
rect 646678 167251 646730 167303
rect 676246 167325 676298 167377
rect 646870 167177 646922 167229
rect 676246 167177 676298 167229
rect 646774 167103 646826 167155
rect 676150 167103 676202 167155
rect 149398 167029 149450 167081
rect 182998 167029 183050 167081
rect 675190 167029 675242 167081
rect 676054 167029 676106 167081
rect 148438 166955 148490 167007
rect 184438 166955 184490 167007
rect 149206 166881 149258 166933
rect 184534 166881 184586 166933
rect 159862 166807 159914 166859
rect 184342 166807 184394 166859
rect 146998 164439 147050 164491
rect 148630 164069 148682 164121
rect 184342 164069 184394 164121
rect 149302 163995 149354 164047
rect 184534 163995 184586 164047
rect 184438 163921 184490 163973
rect 149014 163847 149066 163899
rect 149302 163847 149354 163899
rect 148246 163699 148298 163751
rect 184342 163847 184394 163899
rect 645526 161775 645578 161827
rect 661078 161775 661130 161827
rect 148150 161183 148202 161235
rect 184630 161183 184682 161235
rect 148822 161109 148874 161161
rect 184342 161109 184394 161161
rect 149110 161035 149162 161087
rect 184438 161035 184490 161087
rect 149590 160961 149642 161013
rect 184534 160961 184586 161013
rect 675382 160961 675434 161013
rect 675670 160961 675722 161013
rect 675382 160739 675434 160791
rect 675670 159999 675722 160051
rect 674518 159407 674570 159459
rect 675382 159407 675434 159459
rect 645526 158445 645578 158497
rect 661174 158445 661226 158497
rect 148054 158371 148106 158423
rect 184438 158371 184490 158423
rect 149494 158297 149546 158349
rect 184534 158297 184586 158349
rect 151510 158223 151562 158275
rect 184630 158223 184682 158275
rect 165526 158149 165578 158201
rect 184342 158149 184394 158201
rect 674806 157705 674858 157757
rect 675478 157705 675530 157757
rect 674710 156891 674762 156943
rect 675478 156891 675530 156943
rect 674614 156299 674666 156351
rect 675382 156299 675434 156351
rect 645142 155855 645194 155907
rect 661270 155855 661322 155907
rect 675190 155855 675242 155907
rect 675382 155855 675434 155907
rect 151414 155411 151466 155463
rect 184438 155411 184490 155463
rect 151702 155337 151754 155389
rect 184534 155337 184586 155389
rect 151222 155263 151274 155315
rect 184342 155263 184394 155315
rect 182806 154893 182858 154945
rect 184726 154893 184778 154945
rect 151318 152599 151370 152651
rect 184342 152599 184394 152651
rect 151606 152525 151658 152577
rect 184438 152525 184490 152577
rect 646006 152525 646058 152577
rect 658582 152525 658634 152577
rect 179926 152451 179978 152503
rect 184534 152451 184586 152503
rect 149206 150157 149258 150209
rect 149686 150157 149738 150209
rect 168598 149713 168650 149765
rect 184438 149713 184490 149765
rect 174262 149639 174314 149691
rect 184342 149639 184394 149691
rect 180022 149565 180074 149617
rect 184534 149565 184586 149617
rect 177046 149491 177098 149543
rect 184630 149491 184682 149543
rect 645142 149343 645194 149395
rect 658678 149343 658730 149395
rect 148054 148011 148106 148063
rect 151702 148011 151754 148063
rect 148054 146975 148106 147027
rect 151222 146975 151274 147027
rect 182902 146827 182954 146879
rect 185782 146827 185834 146879
rect 159958 146753 160010 146805
rect 184438 146753 184490 146805
rect 177142 146679 177194 146731
rect 184534 146679 184586 146731
rect 147958 146605 148010 146657
rect 184342 146605 184394 146657
rect 147958 145791 148010 145843
rect 151606 145791 151658 145843
rect 147958 144311 148010 144363
rect 151318 144311 151370 144363
rect 147862 143941 147914 143993
rect 184438 143941 184490 143993
rect 157078 143867 157130 143919
rect 184630 143867 184682 143919
rect 162742 143793 162794 143845
rect 184534 143793 184586 143845
rect 171286 143719 171338 143771
rect 184342 143719 184394 143771
rect 147862 142535 147914 142587
rect 151894 142535 151946 142587
rect 147862 141499 147914 141551
rect 151510 141499 151562 141551
rect 147670 141203 147722 141255
rect 151414 141203 151466 141255
rect 147958 141055 148010 141107
rect 184534 141055 184586 141107
rect 147478 140981 147530 141033
rect 184630 140981 184682 141033
rect 149206 140907 149258 140959
rect 185686 140907 185738 140959
rect 151798 140833 151850 140885
rect 184438 140833 184490 140885
rect 154102 140759 154154 140811
rect 184342 140759 184394 140811
rect 147862 138169 147914 138221
rect 184534 138169 184586 138221
rect 165622 138095 165674 138147
rect 184342 138095 184394 138147
rect 168694 138021 168746 138073
rect 184438 138021 184490 138073
rect 147574 135283 147626 135335
rect 184438 135283 184490 135335
rect 149494 135209 149546 135261
rect 184342 135209 184394 135261
rect 162646 135135 162698 135187
rect 184534 135135 184586 135187
rect 171382 135061 171434 135113
rect 184342 135061 184394 135113
rect 672406 134321 672458 134373
rect 676246 134321 676298 134373
rect 655414 132767 655466 132819
rect 676246 132767 676298 132819
rect 655126 132619 655178 132671
rect 676150 132619 676202 132671
rect 646582 132471 646634 132523
rect 676054 132471 676106 132523
rect 147190 132397 147242 132449
rect 184630 132397 184682 132449
rect 151126 132323 151178 132375
rect 184534 132323 184586 132375
rect 154198 132249 154250 132301
rect 184438 132249 184490 132301
rect 156886 132175 156938 132227
rect 184342 132175 184394 132227
rect 650998 129807 651050 129859
rect 676054 129807 676106 129859
rect 647734 129659 647786 129711
rect 650998 129659 651050 129711
rect 647926 129585 647978 129637
rect 650902 129585 650954 129637
rect 676246 129585 676298 129637
rect 147094 129511 147146 129563
rect 184342 129511 184394 129563
rect 147382 129437 147434 129489
rect 184438 129437 184490 129489
rect 149302 129363 149354 129415
rect 184534 129363 184586 129415
rect 180118 129289 180170 129341
rect 184726 129289 184778 129341
rect 674518 126699 674570 126751
rect 676054 126699 676106 126751
rect 147286 126625 147338 126677
rect 184342 126625 184394 126677
rect 148918 126551 148970 126603
rect 184438 126551 184490 126603
rect 182998 126477 183050 126529
rect 186838 126477 186890 126529
rect 674230 124701 674282 124753
rect 676054 124701 676106 124753
rect 674422 124035 674474 124087
rect 676246 124035 676298 124087
rect 674038 123961 674090 124013
rect 675958 123961 676010 124013
rect 674134 123887 674186 123939
rect 676054 123887 676106 123939
rect 146902 123813 146954 123865
rect 184630 123813 184682 123865
rect 146998 123739 147050 123791
rect 184438 123739 184490 123791
rect 149494 123665 149546 123717
rect 184534 123665 184586 123717
rect 149686 123591 149738 123643
rect 184342 123591 184394 123643
rect 646678 121223 646730 121275
rect 676342 121223 676394 121275
rect 647926 121149 647978 121201
rect 676150 121149 676202 121201
rect 647830 121075 647882 121127
rect 676246 121075 676298 121127
rect 674614 121001 674666 121053
rect 676054 121001 676106 121053
rect 149110 120927 149162 120979
rect 184534 120927 184586 120979
rect 149590 120853 149642 120905
rect 184630 120853 184682 120905
rect 149014 120779 149066 120831
rect 184342 120779 184394 120831
rect 151702 120705 151754 120757
rect 184438 120705 184490 120757
rect 151318 118041 151370 118093
rect 184630 118041 184682 118093
rect 151222 117967 151274 118019
rect 184342 117967 184394 118019
rect 151606 117893 151658 117945
rect 184438 117893 184490 117945
rect 151894 117819 151946 117871
rect 184534 117819 184586 117871
rect 675478 115747 675530 115799
rect 675478 115525 675530 115577
rect 647926 115229 647978 115281
rect 665206 115229 665258 115281
rect 148342 115155 148394 115207
rect 184534 115155 184586 115207
rect 148822 115081 148874 115133
rect 184630 115081 184682 115133
rect 151414 115007 151466 115059
rect 184438 115007 184490 115059
rect 151510 114933 151562 114985
rect 184342 114933 184394 114985
rect 674518 114785 674570 114837
rect 675382 114785 675434 114837
rect 148246 112269 148298 112321
rect 184438 112269 184490 112321
rect 148630 112195 148682 112247
rect 184534 112195 184586 112247
rect 148438 112121 148490 112173
rect 184342 112121 184394 112173
rect 674422 111677 674474 111729
rect 675382 111677 675434 111729
rect 674230 111159 674282 111211
rect 675382 111159 675434 111211
rect 674134 110641 674186 110693
rect 675382 110641 675434 110693
rect 147958 109383 148010 109435
rect 184534 109383 184586 109435
rect 148726 109309 148778 109361
rect 184438 109309 184490 109361
rect 148534 109235 148586 109287
rect 184342 109235 184394 109287
rect 674038 107311 674090 107363
rect 675382 107311 675434 107363
rect 147670 106497 147722 106549
rect 184630 106497 184682 106549
rect 148054 106423 148106 106475
rect 184438 106423 184490 106475
rect 147862 106349 147914 106401
rect 184534 106349 184586 106401
rect 149398 106275 149450 106327
rect 184342 106275 184394 106327
rect 674614 106127 674666 106179
rect 675382 106127 675434 106179
rect 647926 103907 647978 103959
rect 661174 103907 661226 103959
rect 645910 103685 645962 103737
rect 657526 103685 657578 103737
rect 147574 103611 147626 103663
rect 184534 103611 184586 103663
rect 147094 103537 147146 103589
rect 184630 103537 184682 103589
rect 147766 103463 147818 103515
rect 184438 103463 184490 103515
rect 148150 103389 148202 103441
rect 184342 103389 184394 103441
rect 645142 102057 645194 102109
rect 652438 102057 652490 102109
rect 147190 100725 147242 100777
rect 184438 100725 184490 100777
rect 147286 100651 147338 100703
rect 184534 100651 184586 100703
rect 147382 100577 147434 100629
rect 184630 100577 184682 100629
rect 149782 100503 149834 100555
rect 184342 100503 184394 100555
rect 647926 97913 647978 97965
rect 662518 97913 662570 97965
rect 146998 97839 147050 97891
rect 184534 97839 184586 97891
rect 147478 97765 147530 97817
rect 184342 97765 184394 97817
rect 149302 97691 149354 97743
rect 184438 97691 184490 97743
rect 645430 95915 645482 95967
rect 653686 95915 653738 95967
rect 148918 94953 148970 95005
rect 184534 94953 184586 95005
rect 149206 94879 149258 94931
rect 184342 94879 184394 94931
rect 149110 94805 149162 94857
rect 184438 94805 184490 94857
rect 149590 94731 149642 94783
rect 184342 94731 184394 94783
rect 649558 93547 649610 93599
rect 668182 93547 668234 93599
rect 646774 92659 646826 92711
rect 663094 92659 663146 92711
rect 646486 92363 646538 92415
rect 660694 92363 660746 92415
rect 645526 92289 645578 92341
rect 661750 92289 661802 92341
rect 646870 92215 646922 92267
rect 659830 92215 659882 92267
rect 647158 92141 647210 92193
rect 658870 92141 658922 92193
rect 146902 92067 146954 92119
rect 184534 92067 184586 92119
rect 148822 91993 148874 92045
rect 184630 91993 184682 92045
rect 149398 91919 149450 91971
rect 184438 91919 184490 91971
rect 149014 91845 149066 91897
rect 184342 91845 184394 91897
rect 147958 89181 148010 89233
rect 184630 89181 184682 89233
rect 148438 89107 148490 89159
rect 184534 89107 184586 89159
rect 148342 89033 148394 89085
rect 184342 89033 184394 89085
rect 148630 88959 148682 89011
rect 184438 88959 184490 89011
rect 645910 87479 645962 87531
rect 650902 87479 650954 87531
rect 647926 87257 647978 87309
rect 658006 87257 658058 87309
rect 647062 87035 647114 87087
rect 663286 87035 663338 87087
rect 148054 86369 148106 86421
rect 184342 86369 184394 86421
rect 147670 86295 147722 86347
rect 184438 86295 184490 86347
rect 148534 86221 148586 86273
rect 184534 86221 184586 86273
rect 645910 84149 645962 84201
rect 657046 84149 657098 84201
rect 640726 83631 640778 83683
rect 649558 83631 649610 83683
rect 646774 83557 646826 83609
rect 651766 83557 651818 83609
rect 148246 83483 148298 83535
rect 184534 83483 184586 83535
rect 148726 83409 148778 83461
rect 184630 83409 184682 83461
rect 149686 83335 149738 83387
rect 184342 83335 184394 83387
rect 148150 83261 148202 83313
rect 184438 83261 184490 83313
rect 647926 81855 647978 81907
rect 663286 81855 663338 81907
rect 647830 81781 647882 81833
rect 663382 81781 663434 81833
rect 657046 81633 657098 81685
rect 658582 81633 658634 81685
rect 647734 81559 647786 81611
rect 662422 81559 662474 81611
rect 647926 80745 647978 80797
rect 662518 80745 662570 80797
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 149206 80597 149258 80649
rect 184630 80597 184682 80649
rect 149494 80523 149546 80575
rect 184342 80523 184394 80575
rect 147574 80449 147626 80501
rect 184438 80449 184490 80501
rect 148918 80375 148970 80427
rect 184534 80375 184586 80427
rect 149014 77711 149066 77763
rect 184438 77711 184490 77763
rect 646966 77711 647018 77763
rect 658294 77711 658346 77763
rect 149110 77637 149162 77689
rect 184534 77637 184586 77689
rect 646582 77637 646634 77689
rect 659446 77637 659498 77689
rect 149398 77563 149450 77615
rect 184630 77563 184682 77615
rect 646678 77563 646730 77615
rect 661750 77563 661802 77615
rect 149302 77489 149354 77541
rect 184342 77489 184394 77541
rect 647926 77489 647978 77541
rect 656950 77489 657002 77541
rect 646006 76083 646058 76135
rect 657526 76083 657578 76135
rect 647062 74899 647114 74951
rect 660118 74899 660170 74951
rect 148822 74825 148874 74877
rect 184342 74825 184394 74877
rect 148342 74751 148394 74803
rect 184438 74751 184490 74803
rect 148534 74677 148586 74729
rect 184534 74677 184586 74729
rect 149590 74603 149642 74655
rect 184630 74603 184682 74655
rect 647926 72087 647978 72139
rect 660694 72087 660746 72139
rect 148438 71939 148490 71991
rect 184342 71939 184394 71991
rect 148726 71865 148778 71917
rect 184438 71865 184490 71917
rect 149686 71791 149738 71843
rect 184534 71791 184586 71843
rect 647926 69571 647978 69623
rect 661462 69571 661514 69623
rect 148630 69053 148682 69105
rect 184342 69053 184394 69105
rect 149494 68979 149546 69031
rect 184534 68979 184586 69031
rect 149110 68905 149162 68957
rect 184342 68905 184394 68957
rect 149590 68831 149642 68883
rect 184438 68831 184490 68883
rect 149398 66167 149450 66219
rect 184630 66167 184682 66219
rect 646006 66167 646058 66219
rect 652342 66167 652394 66219
rect 149206 66093 149258 66145
rect 184534 66093 184586 66145
rect 149014 66019 149066 66071
rect 184342 66019 184394 66071
rect 149302 65945 149354 65997
rect 184438 65945 184490 65997
rect 647926 63577 647978 63629
rect 663190 63577 663242 63629
rect 149686 63281 149738 63333
rect 184630 63281 184682 63333
rect 149494 63207 149546 63259
rect 184438 63207 184490 63259
rect 149590 63133 149642 63185
rect 184342 63133 184394 63185
rect 149398 63059 149450 63111
rect 184534 63059 184586 63111
rect 647926 60987 647978 61039
rect 663478 60987 663530 61039
rect 149398 60395 149450 60447
rect 184438 60395 184490 60447
rect 149494 60321 149546 60373
rect 184534 60321 184586 60373
rect 149302 60247 149354 60299
rect 184342 60247 184394 60299
rect 646006 59063 646058 59115
rect 652246 59063 652298 59115
rect 149398 58989 149450 59041
rect 184342 58989 184394 59041
rect 149398 57509 149450 57561
rect 184342 57509 184394 57561
rect 149398 56177 149450 56229
rect 184438 56177 184490 56229
rect 149494 56103 149546 56155
rect 184342 56103 184394 56155
rect 149686 54623 149738 54675
rect 184342 54623 184394 54675
rect 149398 53217 149450 53269
rect 184342 53217 184394 53269
rect 331222 48037 331274 48089
rect 354838 48037 354890 48089
rect 362038 48037 362090 48089
rect 389206 48037 389258 48089
rect 411862 48037 411914 48089
rect 424054 48037 424106 48089
rect 434902 48037 434954 48089
rect 475702 48037 475754 48089
rect 311062 47963 311114 48015
rect 371926 47963 371978 48015
rect 405526 47963 405578 48015
rect 441334 47963 441386 48015
rect 460342 47963 460394 48015
rect 510358 47963 510410 48015
rect 320182 47889 320234 47941
rect 515542 47889 515594 47941
rect 285814 47815 285866 47867
rect 493942 47815 493994 47867
rect 302902 47741 302954 47793
rect 525910 47741 525962 47793
rect 268534 47667 268586 47719
rect 503926 47667 503978 47719
rect 233686 47593 233738 47645
rect 475606 47593 475658 47645
rect 250966 47519 251018 47571
rect 521206 47519 521258 47571
rect 145366 47075 145418 47127
rect 199126 47075 199178 47127
rect 455062 46927 455114 46979
rect 458614 46927 458666 46979
rect 521494 46335 521546 46387
rect 527926 46335 527978 46387
rect 515542 45077 515594 45129
rect 529270 45077 529322 45129
rect 509782 43153 509834 43205
rect 521494 43227 521546 43279
rect 633622 43227 633674 43279
rect 640726 43227 640778 43279
rect 398902 42339 398954 42391
rect 411862 42339 411914 42391
rect 471670 41747 471722 41799
rect 475510 41747 475562 41799
rect 514006 41747 514058 41799
rect 514870 41747 514922 41799
rect 503926 40267 503978 40319
rect 506806 40267 506858 40319
rect 365908 37381 365960 37433
rect 398902 37381 398954 37433
rect 420694 37381 420746 37433
rect 455062 37381 455114 37433
rect 475510 37381 475562 37433
rect 509782 37381 509834 37433
rect 475606 37307 475658 37359
rect 514006 37307 514058 37359
<< metal2 >>
rect 148532 1016270 148588 1016279
rect 148532 1016205 148588 1016214
rect 250484 1016270 250540 1016279
rect 250484 1016205 250540 1016214
rect 353396 1016270 353452 1016279
rect 353396 1016205 353452 1016214
rect 148546 1007991 148574 1016205
rect 146612 1007982 146668 1007991
rect 146612 1007917 146668 1007926
rect 148532 1007982 148588 1007991
rect 148532 1007917 148588 1007926
rect 102452 1006206 102508 1006215
rect 92854 1006167 92906 1006173
rect 102452 1006141 102454 1006150
rect 92854 1006109 92906 1006115
rect 102506 1006141 102508 1006150
rect 102454 1006109 102506 1006115
rect 92566 1005871 92618 1005877
rect 92566 1005813 92618 1005819
rect 92470 999729 92522 999735
rect 92470 999671 92522 999677
rect 92290 999527 92350 999533
rect 92290 999475 92298 999527
rect 92290 999469 92350 999475
rect 92290 999468 92338 999469
rect 85940 995846 85996 995855
rect 78384 995813 78686 995832
rect 82032 995813 82334 995832
rect 78384 995807 78698 995813
rect 78384 995804 78646 995807
rect 82032 995807 82346 995813
rect 82032 995804 82294 995807
rect 78646 995749 78698 995755
rect 85728 995804 85940 995832
rect 86242 995813 86352 995832
rect 85940 995781 85996 995790
rect 86230 995807 86352 995813
rect 82294 995749 82346 995755
rect 86282 995804 86352 995807
rect 86230 995749 86282 995755
rect 92290 995739 92318 999468
rect 92374 999433 92426 999439
rect 92374 999375 92426 999381
rect 91510 995733 91562 995739
rect 81620 995698 81676 995707
rect 81408 995656 81620 995684
rect 89424 995665 89822 995684
rect 91248 995681 91510 995684
rect 91248 995675 91562 995681
rect 92278 995733 92330 995739
rect 92278 995675 92330 995681
rect 89424 995659 89834 995665
rect 89424 995656 89782 995659
rect 81620 995633 81676 995642
rect 91248 995656 91550 995675
rect 92386 995665 92414 999375
rect 92374 995659 92426 995665
rect 89782 995601 89834 995607
rect 92374 995601 92426 995607
rect 85366 995585 85418 995591
rect 81044 995550 81100 995559
rect 77088 995508 77342 995536
rect 77314 993741 77342 995508
rect 77698 993815 77726 995522
rect 77686 993809 77738 993815
rect 80194 993783 80222 995522
rect 80784 995508 81044 995536
rect 85104 995533 85366 995536
rect 85104 995527 85418 995533
rect 81044 995485 81100 995494
rect 84514 994079 84542 995522
rect 85104 995508 85406 995527
rect 87552 995517 87902 995536
rect 87552 995511 87914 995517
rect 87552 995508 87862 995511
rect 87862 995453 87914 995459
rect 84500 994070 84556 994079
rect 84500 994005 84556 994014
rect 88738 993931 88766 995522
rect 92482 995517 92510 999671
rect 92578 995855 92606 1005813
rect 92662 1005501 92714 1005507
rect 92662 1005443 92714 1005449
rect 92564 995846 92620 995855
rect 92564 995781 92620 995790
rect 92674 995707 92702 1005443
rect 92758 997953 92810 997959
rect 92758 997895 92810 997901
rect 92770 995961 92798 997895
rect 92758 995955 92810 995961
rect 92758 995897 92810 995903
rect 92660 995698 92716 995707
rect 92660 995633 92716 995642
rect 92866 995559 92894 1006109
rect 101012 1005910 101068 1005919
rect 101012 1005845 101014 1005854
rect 101066 1005845 101068 1005854
rect 101014 1005813 101066 1005819
rect 92950 1005649 93002 1005655
rect 109942 1005649 109994 1005655
rect 92950 1005591 93002 1005597
rect 109940 1005614 109942 1005623
rect 109994 1005614 109996 1005623
rect 92852 995550 92908 995559
rect 92470 995511 92522 995517
rect 92852 995485 92908 995494
rect 92470 995453 92522 995459
rect 88724 993922 88780 993931
rect 88724 993857 88780 993866
rect 77686 993751 77738 993757
rect 80180 993774 80236 993783
rect 77302 993735 77354 993741
rect 80180 993709 80236 993718
rect 77302 993677 77354 993683
rect 89590 990035 89642 990041
rect 89590 989977 89642 989983
rect 73462 989369 73514 989375
rect 73462 989311 73514 989317
rect 45046 989295 45098 989301
rect 45046 989237 45098 989243
rect 44662 987667 44714 987673
rect 44662 987609 44714 987615
rect 44566 987593 44618 987599
rect 44566 987535 44618 987541
rect 42358 970721 42410 970727
rect 42358 970663 42410 970669
rect 42178 968771 42206 969252
rect 42164 968762 42220 968771
rect 42164 968697 42220 968706
rect 41794 967143 41822 967402
rect 42370 967323 42398 970663
rect 44374 970573 44426 970579
rect 44374 970515 44426 970521
rect 42166 967317 42218 967323
rect 42166 967259 42218 967265
rect 42358 967317 42410 967323
rect 42358 967259 42410 967265
rect 41780 967134 41836 967143
rect 41780 967069 41836 967078
rect 42178 966736 42206 967259
rect 44278 966133 44330 966139
rect 44278 966075 44330 966081
rect 41794 965071 41822 965552
rect 41780 965062 41836 965071
rect 41780 964997 41836 965006
rect 41794 964035 41822 964368
rect 41780 964026 41836 964035
rect 41780 963961 41836 963970
rect 41794 963443 41822 963702
rect 41780 963434 41836 963443
rect 41780 963369 41836 963378
rect 41794 962851 41822 963081
rect 41780 962842 41836 962851
rect 41780 962777 41836 962786
rect 41794 962259 41822 962518
rect 41780 962250 41836 962259
rect 41780 962185 41836 962194
rect 41794 959595 41822 960045
rect 41780 959586 41836 959595
rect 41780 959521 41836 959530
rect 41794 959151 41822 959410
rect 41780 959142 41836 959151
rect 41780 959077 41836 959086
rect 42192 958730 42302 958758
rect 41890 957819 41918 958226
rect 41876 957810 41932 957819
rect 41876 957745 41932 957754
rect 42274 957523 42302 958730
rect 42260 957514 42316 957523
rect 42260 957449 42316 957458
rect 42178 956316 42206 956376
rect 42260 956330 42316 956339
rect 42178 956288 42260 956316
rect 42260 956265 42316 956274
rect 42192 955696 42398 955724
rect 42192 955063 42302 955091
rect 38806 950445 38858 950451
rect 38806 950387 38858 950393
rect 34486 947559 34538 947565
rect 34486 947501 34538 947507
rect 34498 945091 34526 947501
rect 34484 945082 34540 945091
rect 34484 945017 34540 945026
rect 38818 937691 38846 950387
rect 39764 944046 39820 944055
rect 39764 943981 39820 943990
rect 39778 938907 39806 943981
rect 41782 943859 41834 943865
rect 41780 943824 41782 943833
rect 41834 943824 41836 943833
rect 41780 943759 41836 943768
rect 41590 943637 41642 943643
rect 41588 943602 41590 943611
rect 41642 943602 41644 943611
rect 41588 943537 41644 943546
rect 40436 942714 40492 942723
rect 40436 942649 40492 942658
rect 40246 941787 40298 941793
rect 40246 941729 40298 941735
rect 40258 941687 40286 941729
rect 40244 941678 40300 941687
rect 40244 941613 40300 941622
rect 40340 941086 40396 941095
rect 40340 941021 40396 941030
rect 39766 938901 39818 938907
rect 39766 938843 39818 938849
rect 38804 937682 38860 937691
rect 38804 937617 38860 937626
rect 28820 932650 28876 932659
rect 28820 932585 28876 932594
rect 28834 932215 28862 932585
rect 28820 932206 28876 932215
rect 28820 932141 28876 932150
rect 39958 820871 40010 820877
rect 39958 820813 40010 820819
rect 39970 816331 39998 820813
rect 39956 816322 40012 816331
rect 39956 816257 40012 816266
rect 40354 814851 40382 941021
rect 40450 817811 40478 942649
rect 41684 942122 41740 942131
rect 41684 942057 41740 942066
rect 41588 940642 41644 940651
rect 41588 940577 41644 940586
rect 41602 938981 41630 940577
rect 41590 938975 41642 938981
rect 41590 938917 41642 938923
rect 41588 932206 41644 932215
rect 41588 932141 41590 932150
rect 41642 932141 41644 932150
rect 41590 932109 41642 932115
rect 41698 823763 41726 942057
rect 42274 939319 42302 955063
rect 42370 950451 42398 955696
rect 42358 950445 42410 950451
rect 42358 950387 42410 950393
rect 42260 939310 42316 939319
rect 42260 939245 42316 939254
rect 43126 921659 43178 921665
rect 43126 921601 43178 921607
rect 41686 823757 41738 823763
rect 41686 823699 41738 823705
rect 41698 820877 41726 823699
rect 41686 820871 41738 820877
rect 41686 820813 41738 820819
rect 41590 819317 41642 819323
rect 41588 819282 41590 819291
rect 41642 819282 41644 819291
rect 41588 819217 41644 819226
rect 41782 818577 41834 818583
rect 41780 818542 41782 818551
rect 41834 818542 41836 818551
rect 41780 818477 41836 818486
rect 41782 818059 41834 818065
rect 41782 818001 41834 818007
rect 41794 817959 41822 818001
rect 41780 817950 41836 817959
rect 41780 817885 41836 817894
rect 40436 817802 40492 817811
rect 40436 817737 40492 817746
rect 41780 817062 41836 817071
rect 41780 816997 41782 817006
rect 41834 816997 41836 817006
rect 41782 816965 41834 816971
rect 40340 814842 40396 814851
rect 40340 814777 40396 814786
rect 42068 814620 42124 814629
rect 42068 814555 42124 814564
rect 41780 814102 41836 814111
rect 41780 814037 41836 814046
rect 34388 813362 34444 813371
rect 34388 813297 34444 813306
rect 23060 806850 23116 806859
rect 23060 806785 23116 806794
rect 23074 806415 23102 806785
rect 23060 806406 23116 806415
rect 23060 806341 23116 806350
rect 34402 802123 34430 813297
rect 41588 812918 41644 812927
rect 41588 812853 41644 812862
rect 41602 812737 41630 812853
rect 41590 812731 41642 812737
rect 41590 812673 41642 812679
rect 41794 812293 41822 814037
rect 41782 812287 41834 812293
rect 41782 812229 41834 812235
rect 41876 812030 41932 812039
rect 41876 811965 41932 811974
rect 34484 811438 34540 811447
rect 34484 811373 34540 811382
rect 34388 802114 34444 802123
rect 34388 802049 34444 802058
rect 34498 801827 34526 811373
rect 41492 810698 41548 810707
rect 41492 810633 41548 810642
rect 34484 801818 34540 801827
rect 34484 801753 34540 801762
rect 41506 800527 41534 810633
rect 41780 810106 41836 810115
rect 41780 810041 41836 810050
rect 41684 809366 41740 809375
rect 41684 809301 41740 809310
rect 41588 807886 41644 807895
rect 41588 807821 41644 807830
rect 41602 806817 41630 807821
rect 41590 806811 41642 806817
rect 41590 806753 41642 806759
rect 41590 806441 41642 806447
rect 41588 806406 41590 806415
rect 41642 806406 41644 806415
rect 41588 806341 41644 806350
rect 41698 800615 41726 809301
rect 41684 800606 41740 800615
rect 41684 800541 41740 800550
rect 41494 800521 41546 800527
rect 41494 800463 41546 800469
rect 41794 800347 41822 810041
rect 41780 800338 41836 800347
rect 41780 800273 41836 800282
rect 41890 800231 41918 811965
rect 41972 811068 42028 811077
rect 41972 811003 42028 811012
rect 41986 809944 42014 811003
rect 42082 810147 42110 814555
rect 43030 812731 43082 812737
rect 43030 812673 43082 812679
rect 42356 812622 42412 812631
rect 42356 812557 42412 812566
rect 42070 810141 42122 810147
rect 42070 810083 42122 810089
rect 41986 809916 42110 809944
rect 41972 808626 42028 808635
rect 41972 808561 42028 808570
rect 41986 800347 42014 808561
rect 41972 800338 42028 800347
rect 42082 800305 42110 809916
rect 42164 809070 42220 809079
rect 42164 809005 42220 809014
rect 41972 800273 42028 800282
rect 42070 800299 42122 800305
rect 42070 800241 42122 800247
rect 42178 800231 42206 809005
rect 42370 802081 42398 812557
rect 42646 812287 42698 812293
rect 42646 812229 42698 812235
rect 42358 802075 42410 802081
rect 42358 802017 42410 802023
rect 41878 800225 41930 800231
rect 41878 800167 41930 800173
rect 42166 800225 42218 800231
rect 42166 800167 42218 800173
rect 41878 800003 41930 800009
rect 41878 799945 41930 799951
rect 41890 799422 41918 799945
rect 42658 798159 42686 812229
rect 43042 812174 43070 812673
rect 42946 812146 43070 812174
rect 42742 806811 42794 806817
rect 42742 806753 42794 806759
rect 42166 798153 42218 798159
rect 42166 798095 42218 798101
rect 42646 798153 42698 798159
rect 42646 798095 42698 798101
rect 42178 797605 42206 798095
rect 42452 797526 42508 797535
rect 42452 797461 42508 797470
rect 42070 797339 42122 797345
rect 42070 797281 42122 797287
rect 42082 796980 42110 797281
rect 41780 796342 41836 796351
rect 41780 796277 41836 796286
rect 41794 795765 41822 796277
rect 42166 795045 42218 795051
rect 42166 794987 42218 794993
rect 42178 794569 42206 794987
rect 41876 794270 41932 794279
rect 41876 794205 41932 794214
rect 41890 793946 41918 794205
rect 42466 793867 42494 797461
rect 42754 795051 42782 806753
rect 42838 802075 42890 802081
rect 42838 802017 42890 802023
rect 42742 795045 42794 795051
rect 42742 794987 42794 794993
rect 42742 794897 42794 794903
rect 42742 794839 42794 794845
rect 42166 793861 42218 793867
rect 42166 793803 42218 793809
rect 42454 793861 42506 793867
rect 42454 793803 42506 793809
rect 42178 793280 42206 793803
rect 42166 793195 42218 793201
rect 42166 793137 42218 793143
rect 42178 792729 42206 793137
rect 42754 790685 42782 794839
rect 42850 793201 42878 802017
rect 42838 793195 42890 793201
rect 42838 793137 42890 793143
rect 42838 793047 42890 793053
rect 42838 792989 42890 792995
rect 42166 790679 42218 790685
rect 42166 790621 42218 790627
rect 42742 790679 42794 790685
rect 42742 790621 42794 790627
rect 42178 790246 42206 790621
rect 42740 790570 42796 790579
rect 42740 790505 42796 790514
rect 42166 789939 42218 789945
rect 42166 789881 42218 789887
rect 42178 789580 42206 789881
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42178 788957 42206 789437
rect 42452 789238 42508 789247
rect 42452 789173 42508 789182
rect 42166 788829 42218 788835
rect 42166 788771 42218 788777
rect 42178 788396 42206 788771
rect 42166 787053 42218 787059
rect 42166 786995 42218 787001
rect 42178 786546 42206 786995
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42178 785921 42206 786403
rect 42466 785801 42494 789173
rect 42754 786467 42782 790505
rect 42850 789501 42878 792989
rect 42838 789495 42890 789501
rect 42838 789437 42890 789443
rect 42946 788835 42974 812146
rect 43030 810141 43082 810147
rect 43030 810083 43082 810089
rect 42934 788829 42986 788835
rect 42934 788771 42986 788777
rect 43042 787059 43070 810083
rect 43138 797345 43166 921601
rect 43222 817023 43274 817029
rect 43222 816965 43274 816971
rect 43234 797345 43262 816965
rect 43510 800521 43562 800527
rect 43510 800463 43562 800469
rect 43414 800299 43466 800305
rect 43414 800241 43466 800247
rect 43318 800225 43370 800231
rect 43318 800167 43370 800173
rect 43126 797339 43178 797345
rect 43126 797281 43178 797287
rect 43222 797339 43274 797345
rect 43222 797281 43274 797287
rect 43330 797216 43358 800167
rect 43138 797188 43358 797216
rect 43138 794903 43166 797188
rect 43222 797117 43274 797123
rect 43222 797059 43274 797065
rect 43126 794897 43178 794903
rect 43126 794839 43178 794845
rect 43126 794749 43178 794755
rect 43126 794691 43178 794697
rect 43138 793053 43166 794691
rect 43126 793047 43178 793053
rect 43126 792989 43178 792995
rect 43126 792899 43178 792905
rect 43126 792841 43178 792847
rect 43138 789945 43166 792841
rect 43126 789939 43178 789945
rect 43126 789881 43178 789887
rect 43030 787053 43082 787059
rect 43030 786995 43082 787001
rect 42742 786461 42794 786467
rect 42742 786403 42794 786409
rect 42070 785795 42122 785801
rect 42070 785737 42122 785743
rect 42454 785795 42506 785801
rect 42454 785737 42506 785743
rect 42082 785288 42110 785737
rect 42166 784611 42218 784617
rect 42166 784553 42218 784559
rect 42070 784315 42122 784321
rect 42070 784257 42122 784263
rect 41590 776101 41642 776107
rect 41588 776066 41590 776075
rect 41642 776066 41644 776075
rect 41588 776001 41644 776010
rect 41782 775361 41834 775367
rect 41780 775326 41782 775335
rect 41834 775326 41836 775335
rect 41780 775261 41836 775270
rect 41782 774843 41834 774849
rect 41780 774808 41782 774817
rect 41834 774808 41836 774817
rect 41780 774743 41836 774752
rect 41590 774621 41642 774627
rect 41588 774586 41590 774595
rect 41642 774586 41644 774595
rect 41588 774521 41644 774530
rect 41588 773698 41644 773707
rect 41588 773633 41590 773642
rect 41642 773633 41644 773642
rect 41590 773601 41642 773607
rect 42082 772375 42110 784257
rect 42178 773263 42206 784553
rect 43234 774627 43262 797059
rect 43426 794755 43454 800241
rect 43414 794749 43466 794755
rect 43414 794691 43466 794697
rect 43522 792905 43550 800463
rect 43510 792899 43562 792905
rect 43510 792841 43562 792847
rect 43222 774621 43274 774627
rect 43222 774563 43274 774569
rect 43222 773659 43274 773665
rect 43222 773601 43274 773607
rect 42164 773254 42220 773263
rect 42164 773189 42220 773198
rect 42068 772366 42124 772375
rect 42068 772301 42124 772310
rect 42068 771922 42124 771931
rect 42068 771857 42124 771866
rect 41780 771404 41836 771413
rect 41780 771339 41836 771348
rect 40436 770590 40492 770599
rect 40436 770525 40492 770534
rect 33044 770146 33100 770155
rect 33044 770081 33100 770090
rect 23060 763634 23116 763643
rect 23060 763569 23116 763578
rect 23074 763199 23102 763569
rect 23060 763190 23116 763199
rect 23060 763125 23116 763134
rect 33058 758107 33086 770081
rect 40340 768666 40396 768675
rect 40340 768601 40396 768610
rect 33236 768222 33292 768231
rect 33236 768157 33292 768166
rect 33250 758255 33278 768157
rect 33236 758246 33292 758255
rect 33236 758181 33292 758190
rect 33044 758098 33100 758107
rect 33044 758033 33100 758042
rect 40354 757385 40382 768601
rect 40450 757459 40478 770525
rect 41794 770039 41822 771339
rect 41782 770033 41834 770039
rect 41782 769975 41834 769981
rect 41780 769924 41836 769933
rect 41780 769859 41836 769868
rect 41794 769521 41822 769859
rect 41782 769515 41834 769521
rect 41782 769457 41834 769463
rect 41780 769406 41836 769415
rect 41780 769341 41836 769350
rect 41684 766742 41740 766751
rect 41684 766677 41740 766686
rect 41588 766150 41644 766159
rect 41588 766085 41590 766094
rect 41642 766085 41644 766094
rect 41590 766053 41642 766059
rect 41492 765262 41548 765271
rect 41492 765197 41548 765206
rect 41506 757541 41534 765197
rect 41590 763299 41642 763305
rect 41590 763241 41642 763247
rect 41602 763199 41630 763241
rect 41588 763190 41644 763199
rect 41588 763125 41644 763134
rect 41506 757513 41594 757541
rect 40438 757453 40490 757459
rect 40438 757395 40490 757401
rect 41566 757385 41594 757513
rect 40342 757379 40394 757385
rect 40342 757321 40394 757327
rect 41554 757379 41606 757385
rect 41554 757321 41606 757327
rect 41698 757311 41726 766677
rect 41686 757305 41738 757311
rect 41686 757247 41738 757253
rect 41794 757089 41822 769341
rect 41876 767926 41932 767935
rect 41876 767861 41932 767870
rect 41890 766413 41918 767861
rect 41972 767334 42028 767343
rect 41972 767269 42028 767278
rect 41878 766407 41930 766413
rect 41878 766349 41930 766355
rect 41876 764892 41932 764901
rect 41876 764827 41932 764836
rect 41782 757083 41834 757089
rect 41782 757025 41834 757031
rect 41890 757015 41918 764827
rect 41986 757163 42014 767269
rect 42082 757533 42110 771857
rect 42934 770033 42986 770039
rect 42934 769975 42986 769981
rect 42838 766111 42890 766117
rect 42838 766053 42890 766059
rect 42164 765854 42220 765863
rect 42164 765789 42220 765798
rect 42070 757527 42122 757533
rect 42070 757469 42122 757475
rect 42178 757237 42206 765789
rect 42850 760334 42878 766053
rect 42754 760306 42878 760334
rect 42454 757453 42506 757459
rect 42454 757395 42506 757401
rect 42166 757231 42218 757237
rect 42166 757173 42218 757179
rect 41974 757157 42026 757163
rect 41974 757099 42026 757105
rect 41878 757009 41930 757015
rect 41878 756951 41930 756957
rect 41878 756787 41930 756793
rect 41878 756729 41930 756735
rect 41890 756245 41918 756729
rect 42466 755535 42494 757395
rect 42754 756539 42782 760306
rect 42838 757305 42890 757311
rect 42838 757247 42890 757253
rect 42740 756530 42796 756539
rect 42740 756465 42796 756474
rect 42166 755529 42218 755535
rect 42166 755471 42218 755477
rect 42454 755529 42506 755535
rect 42454 755471 42506 755477
rect 42178 755239 42206 755471
rect 42166 755233 42218 755239
rect 42166 755175 42218 755181
rect 42070 754937 42122 754943
rect 42070 754879 42122 754885
rect 42082 754430 42110 754879
rect 42166 754123 42218 754129
rect 42166 754065 42218 754071
rect 42178 753764 42206 754065
rect 42850 753093 42878 757247
rect 42946 757131 42974 769975
rect 43030 769515 43082 769521
rect 43030 769457 43082 769463
rect 43042 757311 43070 769457
rect 43126 766407 43178 766413
rect 43126 766349 43178 766355
rect 43138 757533 43166 766349
rect 43126 757527 43178 757533
rect 43126 757469 43178 757475
rect 43126 757379 43178 757385
rect 43126 757321 43178 757327
rect 43030 757305 43082 757311
rect 43030 757247 43082 757253
rect 42932 757122 42988 757131
rect 42932 757057 42988 757066
rect 43030 757083 43082 757089
rect 43030 757025 43082 757031
rect 42934 757009 42986 757015
rect 42934 756951 42986 756957
rect 42070 753087 42122 753093
rect 42070 753029 42122 753035
rect 42838 753087 42890 753093
rect 42838 753029 42890 753035
rect 42082 752580 42110 753029
rect 42838 752939 42890 752945
rect 42838 752881 42890 752887
rect 42070 751829 42122 751835
rect 42070 751771 42122 751777
rect 42082 751396 42110 751771
rect 42068 751054 42124 751063
rect 42068 750989 42124 750998
rect 42082 750730 42110 750989
rect 42166 750645 42218 750651
rect 42166 750587 42218 750593
rect 42178 750064 42206 750587
rect 42070 749979 42122 749985
rect 42070 749921 42122 749927
rect 42082 749546 42110 749921
rect 42644 748686 42700 748695
rect 42644 748621 42700 748630
rect 42082 746877 42110 747030
rect 42166 746945 42218 746951
rect 42166 746887 42218 746893
rect 42070 746871 42122 746877
rect 42070 746813 42122 746819
rect 42178 746401 42206 746887
rect 42070 746131 42122 746137
rect 42070 746073 42122 746079
rect 42082 745772 42110 746073
rect 42166 745687 42218 745693
rect 42166 745629 42218 745635
rect 42178 745180 42206 745629
rect 42166 743763 42218 743769
rect 42166 743705 42218 743711
rect 42178 743365 42206 743705
rect 42658 743251 42686 748621
rect 42740 748538 42796 748547
rect 42740 748473 42796 748482
rect 42070 743245 42122 743251
rect 42070 743187 42122 743193
rect 42646 743245 42698 743251
rect 42646 743187 42698 743193
rect 42082 742738 42110 743187
rect 42754 742437 42782 748473
rect 42850 746951 42878 752881
rect 42946 751835 42974 756951
rect 42934 751829 42986 751835
rect 42934 751771 42986 751777
rect 42934 751681 42986 751687
rect 42934 751623 42986 751629
rect 42838 746945 42890 746951
rect 42838 746887 42890 746893
rect 42946 746877 42974 751623
rect 43042 749985 43070 757025
rect 43138 750651 43166 757321
rect 43126 750645 43178 750651
rect 43126 750587 43178 750593
rect 43126 750497 43178 750503
rect 43126 750439 43178 750445
rect 43030 749979 43082 749985
rect 43030 749921 43082 749927
rect 43028 749870 43084 749879
rect 43028 749805 43084 749814
rect 42934 746871 42986 746877
rect 42934 746813 42986 746819
rect 43042 743769 43070 749805
rect 43138 745693 43166 750439
rect 43126 745687 43178 745693
rect 43126 745629 43178 745635
rect 43030 743763 43082 743769
rect 43030 743705 43082 743711
rect 42166 742431 42218 742437
rect 42166 742373 42218 742379
rect 42742 742431 42794 742437
rect 42742 742373 42794 742379
rect 42178 742072 42206 742373
rect 42070 741395 42122 741401
rect 42070 741337 42122 741343
rect 41686 741173 41738 741179
rect 41686 741115 41738 741121
rect 41590 732885 41642 732891
rect 41588 732850 41590 732859
rect 41642 732850 41644 732859
rect 41588 732785 41644 732794
rect 41590 731849 41642 731855
rect 41588 731814 41590 731823
rect 41642 731814 41644 731823
rect 41588 731749 41644 731758
rect 41590 731405 41642 731411
rect 41588 731370 41590 731379
rect 41642 731370 41644 731379
rect 41588 731305 41644 731314
rect 41588 730482 41644 730491
rect 41588 730417 41590 730426
rect 41642 730417 41644 730426
rect 41590 730385 41642 730391
rect 41698 729455 41726 741115
rect 41782 732145 41834 732151
rect 41780 732110 41782 732119
rect 41834 732110 41836 732119
rect 41780 732045 41836 732054
rect 42082 730121 42110 741337
rect 43234 731411 43262 773601
rect 43606 757527 43658 757533
rect 43606 757469 43658 757475
rect 43702 757527 43754 757533
rect 43702 757469 43754 757475
rect 43510 757305 43562 757311
rect 43510 757247 43562 757253
rect 43414 757231 43466 757237
rect 43414 757173 43466 757179
rect 43318 757157 43370 757163
rect 43318 757099 43370 757105
rect 43330 752945 43358 757099
rect 43318 752939 43370 752945
rect 43318 752881 43370 752887
rect 43426 751687 43454 757173
rect 43414 751681 43466 751687
rect 43414 751623 43466 751629
rect 43522 750503 43550 757247
rect 43510 750497 43562 750503
rect 43510 750439 43562 750445
rect 43618 746137 43646 757469
rect 43714 754129 43742 757469
rect 43702 754123 43754 754129
rect 43702 754065 43754 754071
rect 43606 746131 43658 746137
rect 43606 746073 43658 746079
rect 44290 741179 44318 966075
rect 44278 741173 44330 741179
rect 44278 741115 44330 741121
rect 43222 731405 43274 731411
rect 43222 731347 43274 731353
rect 43222 730443 43274 730449
rect 43222 730385 43274 730391
rect 42068 730112 42124 730121
rect 42068 730047 42124 730056
rect 41684 729446 41740 729455
rect 41684 729381 41740 729390
rect 41684 727966 41740 727975
rect 41684 727901 41740 727910
rect 34388 726930 34444 726939
rect 34388 726865 34444 726874
rect 23060 720418 23116 720427
rect 23060 720353 23116 720362
rect 23074 719835 23102 720353
rect 23060 719826 23116 719835
rect 23060 719761 23116 719770
rect 34402 717023 34430 726865
rect 41492 726486 41548 726495
rect 41492 726421 41548 726430
rect 34484 725006 34540 725015
rect 34484 724941 34540 724950
rect 34388 717014 34444 717023
rect 34388 716949 34444 716958
rect 34498 716579 34526 724941
rect 34484 716570 34540 716579
rect 34484 716505 34540 716514
rect 41506 714107 41534 726421
rect 41588 723970 41644 723979
rect 41588 723905 41644 723914
rect 41602 723049 41630 723905
rect 41590 723043 41642 723049
rect 41590 722985 41642 722991
rect 41588 722046 41644 722055
rect 41588 721981 41644 721990
rect 41602 720163 41630 721981
rect 41590 720157 41642 720163
rect 41590 720099 41642 720105
rect 41494 714101 41546 714107
rect 41494 714043 41546 714049
rect 41698 714070 41726 727901
rect 41972 727670 42028 727679
rect 41972 727605 42028 727614
rect 41876 725598 41932 725607
rect 41876 725533 41932 725542
rect 41780 723674 41836 723683
rect 41780 723609 41836 723618
rect 41794 723345 41822 723609
rect 41782 723339 41834 723345
rect 41782 723281 41834 723287
rect 41780 723230 41836 723239
rect 41780 723165 41782 723174
rect 41834 723165 41836 723174
rect 41782 723133 41834 723139
rect 41780 721158 41836 721167
rect 41780 721093 41836 721102
rect 41794 720237 41822 721093
rect 41782 720231 41834 720237
rect 41780 720196 41782 720205
rect 41834 720196 41836 720205
rect 41780 720131 41836 720140
rect 41698 714054 41836 714070
rect 41698 714042 41780 714054
rect 41780 713989 41836 713998
rect 41890 713873 41918 725533
rect 41986 713915 42014 727605
rect 42068 726190 42124 726199
rect 42068 726125 42124 726134
rect 41972 713906 42028 713915
rect 41878 713867 41930 713873
rect 42082 713873 42110 726125
rect 42164 724710 42220 724719
rect 42164 724645 42220 724654
rect 42178 713915 42206 724645
rect 42934 723339 42986 723345
rect 42934 723281 42986 723287
rect 42838 723043 42890 723049
rect 42838 722985 42890 722991
rect 42452 721602 42508 721611
rect 42452 721537 42508 721546
rect 42164 713906 42220 713915
rect 41972 713841 42028 713850
rect 42070 713867 42122 713873
rect 41878 713809 41930 713815
rect 42164 713841 42220 713850
rect 42070 713809 42122 713815
rect 41878 713571 41930 713577
rect 41878 713513 41930 713519
rect 41890 713064 41918 713513
rect 42466 713281 42494 721537
rect 42454 713275 42506 713281
rect 42454 713217 42506 713223
rect 42068 711686 42124 711695
rect 42068 711621 42124 711630
rect 42082 711214 42110 711621
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42178 710548 42206 710849
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42178 709364 42206 709887
rect 42070 708613 42122 708619
rect 42070 708555 42122 708561
rect 42082 708180 42110 708555
rect 42166 708095 42218 708101
rect 42166 708037 42218 708043
rect 42178 707514 42206 708037
rect 42166 707429 42218 707435
rect 42166 707371 42218 707377
rect 42178 706881 42206 707371
rect 42166 706615 42218 706621
rect 42166 706557 42218 706563
rect 42178 706330 42206 706557
rect 42452 706062 42508 706071
rect 42452 705997 42508 706006
rect 42466 705614 42494 705997
rect 42466 705586 42590 705614
rect 42562 705012 42590 705586
rect 42466 704984 42590 705012
rect 42466 704845 42494 704984
rect 42262 704839 42314 704845
rect 42262 704781 42314 704787
rect 42454 704839 42506 704845
rect 42454 704781 42506 704787
rect 42274 703859 42302 704781
rect 42192 703831 42302 703859
rect 42262 703729 42314 703735
rect 42262 703671 42314 703677
rect 42452 703694 42508 703703
rect 42070 703581 42122 703587
rect 42070 703523 42122 703529
rect 42082 703222 42110 703523
rect 42274 702570 42302 703671
rect 42452 703629 42508 703638
rect 42192 702542 42302 702570
rect 42166 702323 42218 702329
rect 42166 702265 42218 702271
rect 42178 702005 42206 702265
rect 42070 700399 42122 700405
rect 42070 700341 42122 700347
rect 42082 700188 42110 700341
rect 42166 700103 42218 700109
rect 42166 700045 42218 700051
rect 42178 699522 42206 700045
rect 42466 699443 42494 703629
rect 42850 703587 42878 722985
rect 42946 709951 42974 723281
rect 43030 723191 43082 723197
rect 43030 723133 43082 723139
rect 42934 709945 42986 709951
rect 42934 709887 42986 709893
rect 42932 709762 42988 709771
rect 42932 709697 42988 709706
rect 42946 703735 42974 709697
rect 43042 708101 43070 723133
rect 43126 720157 43178 720163
rect 43126 720099 43178 720105
rect 43030 708095 43082 708101
rect 43030 708037 43082 708043
rect 43030 707947 43082 707953
rect 43030 707889 43082 707895
rect 43042 706621 43070 707889
rect 43138 707435 43166 720099
rect 43126 707429 43178 707435
rect 43126 707371 43178 707377
rect 43124 707246 43180 707255
rect 43124 707181 43180 707190
rect 43030 706615 43082 706621
rect 43030 706557 43082 706563
rect 43030 706467 43082 706473
rect 43030 706409 43082 706415
rect 42934 703729 42986 703735
rect 42934 703671 42986 703677
rect 42838 703581 42890 703587
rect 42838 703523 42890 703529
rect 42836 703398 42892 703407
rect 42836 703333 42892 703342
rect 42850 700109 42878 703333
rect 43042 702329 43070 706409
rect 43030 702323 43082 702329
rect 43030 702265 43082 702271
rect 43138 700405 43166 707181
rect 43126 700399 43178 700405
rect 43126 700341 43178 700347
rect 42838 700103 42890 700109
rect 42838 700045 42890 700051
rect 42166 699437 42218 699443
rect 42166 699379 42218 699385
rect 42454 699437 42506 699443
rect 42454 699379 42506 699385
rect 42178 698856 42206 699379
rect 41878 694701 41930 694707
rect 41878 694643 41930 694649
rect 41782 689521 41834 689527
rect 41780 689486 41782 689495
rect 41834 689486 41836 689495
rect 41780 689421 41836 689430
rect 41782 688929 41834 688935
rect 41780 688894 41782 688903
rect 41834 688894 41836 688903
rect 41780 688829 41836 688838
rect 41590 688633 41642 688639
rect 41588 688598 41590 688607
rect 41642 688598 41644 688607
rect 41588 688533 41644 688542
rect 41590 688189 41642 688195
rect 41588 688154 41590 688163
rect 41642 688154 41644 688163
rect 41588 688089 41644 688098
rect 41588 687266 41644 687275
rect 41588 687201 41590 687210
rect 41642 687201 41644 687210
rect 41590 687169 41642 687175
rect 41890 686979 41918 694643
rect 43234 688195 43262 730385
rect 43702 714385 43754 714391
rect 43702 714327 43754 714333
rect 43606 714089 43658 714095
rect 43606 714031 43658 714037
rect 43414 713867 43466 713873
rect 43414 713809 43466 713815
rect 43426 707953 43454 713809
rect 43510 713275 43562 713281
rect 43510 713217 43562 713223
rect 43522 708619 43550 713217
rect 43510 708613 43562 708619
rect 43510 708555 43562 708561
rect 43414 707947 43466 707953
rect 43414 707889 43466 707895
rect 43618 706473 43646 714031
rect 43714 710913 43742 714327
rect 43702 710907 43754 710913
rect 43702 710849 43754 710855
rect 43606 706467 43658 706473
rect 43606 706409 43658 706415
rect 43222 688189 43274 688195
rect 43222 688131 43274 688137
rect 43222 687227 43274 687233
rect 43222 687169 43274 687175
rect 41876 686970 41932 686979
rect 41876 686905 41932 686914
rect 41782 685969 41834 685975
rect 41780 685934 41782 685943
rect 41834 685934 41836 685943
rect 41780 685869 41836 685878
rect 41780 685046 41836 685055
rect 41780 684981 41836 684990
rect 41588 684306 41644 684315
rect 41588 684241 41644 684250
rect 34388 683714 34444 683723
rect 34388 683649 34444 683658
rect 23060 677202 23116 677211
rect 23060 677137 23116 677146
rect 23074 676767 23102 677137
rect 23060 676758 23116 676767
rect 23060 676693 23116 676702
rect 34402 672623 34430 683649
rect 41602 682867 41630 684241
rect 41684 683270 41740 683279
rect 41684 683205 41740 683214
rect 41590 682861 41642 682867
rect 41590 682803 41642 682809
rect 34484 681790 34540 681799
rect 34484 681725 34540 681734
rect 34388 672614 34444 672623
rect 34388 672549 34444 672558
rect 34498 672475 34526 681725
rect 41588 680310 41644 680319
rect 41588 680245 41590 680254
rect 41642 680245 41644 680254
rect 41590 680213 41642 680219
rect 41698 679694 41726 683205
rect 41410 679666 41726 679694
rect 34484 672466 34540 672475
rect 34484 672401 34540 672410
rect 41410 670983 41438 679666
rect 41588 679274 41644 679283
rect 41588 679209 41590 679218
rect 41642 679209 41644 679218
rect 41590 679177 41642 679183
rect 41794 679112 41822 684981
rect 42452 682974 42508 682983
rect 42452 682909 42508 682918
rect 41876 682382 41932 682391
rect 41876 682317 41932 682326
rect 41506 679084 41822 679112
rect 41398 670977 41450 670983
rect 41398 670919 41450 670925
rect 41506 670909 41534 679084
rect 41686 678939 41738 678945
rect 41686 678881 41738 678887
rect 41588 678830 41644 678839
rect 41588 678765 41644 678774
rect 41602 677021 41630 678765
rect 41590 677015 41642 677021
rect 41590 676957 41642 676963
rect 41698 671416 41726 678881
rect 41780 678534 41836 678543
rect 41780 678469 41782 678478
rect 41834 678469 41836 678478
rect 41782 678437 41834 678443
rect 41780 677942 41836 677951
rect 41780 677877 41836 677886
rect 41794 676989 41822 677877
rect 41780 676980 41836 676989
rect 41780 676915 41782 676924
rect 41834 676915 41836 676924
rect 41782 676883 41834 676889
rect 41698 671388 41822 671416
rect 41494 670903 41546 670909
rect 41494 670845 41546 670851
rect 41794 670699 41822 671388
rect 41780 670690 41836 670699
rect 41890 670657 41918 682317
rect 42164 681494 42220 681503
rect 42164 681429 42220 681438
rect 42068 680902 42124 680911
rect 42068 680837 42124 680846
rect 41972 680014 42028 680023
rect 41972 679949 42028 679958
rect 41986 671989 42014 679949
rect 41974 671983 42026 671989
rect 41974 671925 42026 671931
rect 42082 670699 42110 680837
rect 42068 670690 42124 670699
rect 41780 670625 41836 670634
rect 41878 670651 41930 670657
rect 42178 670657 42206 681429
rect 42466 678945 42494 682909
rect 42742 682861 42794 682867
rect 42742 682803 42794 682809
rect 42754 679694 42782 682803
rect 42934 680271 42986 680277
rect 42934 680213 42986 680219
rect 42754 679666 42878 679694
rect 42742 679235 42794 679241
rect 42742 679177 42794 679183
rect 42454 678939 42506 678945
rect 42454 678881 42506 678887
rect 42454 678791 42506 678797
rect 42454 678733 42506 678739
rect 42068 670625 42124 670634
rect 42166 670651 42218 670657
rect 41878 670593 41930 670599
rect 42166 670593 42218 670599
rect 41878 670355 41930 670361
rect 41878 670297 41930 670303
rect 41890 669848 41918 670297
rect 42466 670107 42494 678733
rect 42754 670835 42782 679177
rect 42850 678668 42878 679666
rect 42946 678797 42974 680213
rect 42934 678791 42986 678797
rect 42934 678733 42986 678739
rect 42850 678640 43070 678668
rect 42838 678495 42890 678501
rect 42838 678437 42890 678443
rect 42742 670829 42794 670835
rect 42742 670771 42794 670777
rect 42742 670651 42794 670657
rect 42742 670593 42794 670599
rect 42452 670098 42508 670107
rect 42452 670033 42508 670042
rect 42166 668431 42218 668437
rect 42166 668373 42218 668379
rect 42178 667998 42206 668373
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42178 667361 42206 667855
rect 42164 666694 42220 666703
rect 42164 666629 42220 666638
rect 42178 666148 42206 666629
rect 42166 665397 42218 665403
rect 42166 665339 42218 665345
rect 42178 664964 42206 665339
rect 42166 664879 42218 664885
rect 42166 664821 42218 664827
rect 42178 664298 42206 664821
rect 42070 663991 42122 663997
rect 42070 663933 42122 663939
rect 42082 663706 42110 663933
rect 41780 663438 41836 663447
rect 41780 663373 41836 663382
rect 41794 663114 41822 663373
rect 42070 661105 42122 661111
rect 42070 661047 42122 661053
rect 42082 660672 42110 661047
rect 42070 660439 42122 660445
rect 42070 660381 42122 660387
rect 42082 660006 42110 660381
rect 42754 659927 42782 670593
rect 42850 665403 42878 678437
rect 42934 671983 42986 671989
rect 42934 671925 42986 671931
rect 42838 665397 42890 665403
rect 42838 665339 42890 665345
rect 42836 665214 42892 665223
rect 42836 665149 42892 665158
rect 42850 660445 42878 665149
rect 42946 664885 42974 671925
rect 43042 668437 43070 678640
rect 43126 677015 43178 677021
rect 43126 676957 43178 676963
rect 43030 668431 43082 668437
rect 43030 668373 43082 668379
rect 43030 668283 43082 668289
rect 43030 668225 43082 668231
rect 42934 664879 42986 664885
rect 42934 664821 42986 664827
rect 42934 664731 42986 664737
rect 42934 664673 42986 664679
rect 42838 660439 42890 660445
rect 42838 660381 42890 660387
rect 42836 660330 42892 660339
rect 42836 660265 42892 660274
rect 42166 659921 42218 659927
rect 42166 659863 42218 659869
rect 42742 659921 42794 659927
rect 42742 659863 42794 659869
rect 42178 659340 42206 659863
rect 42742 659773 42794 659779
rect 42742 659715 42794 659721
rect 42070 659107 42122 659113
rect 42070 659049 42122 659055
rect 42082 658822 42110 659049
rect 42754 658836 42782 659715
rect 42850 658984 42878 660265
rect 42946 659779 42974 664673
rect 43042 661111 43070 668225
rect 43138 663997 43166 676957
rect 43126 663991 43178 663997
rect 43126 663933 43178 663939
rect 43126 663843 43178 663849
rect 43126 663785 43178 663791
rect 43030 661105 43082 661111
rect 43030 661047 43082 661053
rect 43028 660922 43084 660931
rect 43028 660857 43084 660866
rect 42934 659773 42986 659779
rect 42934 659715 42986 659721
rect 42934 659625 42986 659631
rect 42934 659567 42986 659573
rect 42946 659113 42974 659567
rect 42934 659107 42986 659113
rect 42934 659049 42986 659055
rect 42850 658956 42974 658984
rect 42754 658808 42878 658836
rect 42850 657263 42878 658808
rect 42070 657257 42122 657263
rect 42070 657199 42122 657205
rect 42838 657257 42890 657263
rect 42838 657199 42890 657205
rect 42082 656972 42110 657199
rect 42946 656745 42974 658956
rect 42166 656739 42218 656745
rect 42166 656681 42218 656687
rect 42934 656739 42986 656745
rect 42934 656681 42986 656687
rect 42178 656306 42206 656681
rect 43042 656227 43070 660857
rect 43138 659631 43166 663785
rect 43126 659625 43178 659631
rect 43126 659567 43178 659573
rect 42166 656221 42218 656227
rect 42166 656163 42218 656169
rect 43030 656221 43082 656227
rect 43030 656163 43082 656169
rect 42178 655677 42206 656163
rect 41782 646305 41834 646311
rect 41780 646270 41782 646279
rect 41834 646270 41836 646279
rect 41780 646205 41836 646214
rect 41782 645787 41834 645793
rect 41780 645752 41782 645761
rect 41834 645752 41836 645761
rect 41780 645687 41836 645696
rect 41590 645417 41642 645423
rect 41588 645382 41590 645391
rect 41642 645382 41644 645391
rect 41588 645317 41644 645326
rect 43234 644831 43262 687169
rect 43606 671095 43658 671101
rect 43606 671037 43658 671043
rect 43510 670977 43562 670983
rect 43510 670919 43562 670925
rect 43414 670903 43466 670909
rect 43414 670845 43466 670851
rect 43318 670829 43370 670835
rect 43318 670771 43370 670777
rect 43330 668289 43358 670771
rect 43318 668283 43370 668289
rect 43318 668225 43370 668231
rect 43426 664737 43454 670845
rect 43414 664731 43466 664737
rect 43414 664673 43466 664679
rect 43522 663849 43550 670919
rect 43618 667919 43646 671037
rect 43606 667913 43658 667919
rect 43606 667855 43658 667861
rect 43510 663843 43562 663849
rect 43510 663785 43562 663791
rect 41782 644825 41834 644831
rect 41780 644790 41782 644799
rect 43222 644825 43274 644831
rect 41834 644790 41836 644799
rect 43222 644767 43274 644773
rect 41780 644725 41836 644734
rect 43796 644198 43852 644207
rect 43796 644133 43852 644142
rect 43316 643754 43372 643763
rect 43316 643689 43372 643698
rect 25844 642422 25900 642431
rect 25844 642357 25900 642366
rect 23156 633986 23212 633995
rect 23156 633921 23212 633930
rect 23170 633551 23198 633921
rect 23156 633542 23212 633551
rect 23156 633477 23212 633486
rect 25858 629291 25886 642357
rect 41588 641534 41644 641543
rect 41588 641469 41644 641478
rect 34388 640498 34444 640507
rect 34388 640433 34444 640442
rect 25846 629285 25898 629291
rect 25846 629227 25898 629233
rect 34402 627927 34430 640433
rect 41492 640054 41548 640063
rect 41492 639989 41548 639998
rect 34484 638574 34540 638583
rect 34484 638509 34540 638518
rect 34498 629111 34526 638509
rect 34484 629102 34540 629111
rect 34484 629037 34540 629046
rect 41506 627927 41534 639989
rect 34388 627918 34444 627927
rect 34388 627853 34444 627862
rect 41492 627918 41548 627927
rect 41492 627853 41548 627862
rect 41602 627779 41630 641469
rect 41780 641238 41836 641247
rect 41780 641173 41836 641182
rect 41794 639577 41822 641173
rect 41876 639758 41932 639767
rect 41876 639693 41932 639702
rect 41782 639571 41834 639577
rect 41782 639513 41834 639519
rect 41780 639166 41836 639175
rect 41780 639101 41836 639110
rect 41684 637094 41740 637103
rect 41684 637029 41686 637038
rect 41738 637029 41740 637038
rect 41686 636997 41738 637003
rect 41684 635022 41740 635031
rect 41684 634957 41686 634966
rect 41738 634957 41740 634966
rect 41686 634925 41738 634931
rect 41684 634578 41740 634587
rect 41684 634513 41740 634522
rect 41698 633995 41726 634513
rect 41684 633986 41740 633995
rect 41684 633921 41686 633930
rect 41738 633921 41740 633930
rect 41686 633889 41738 633895
rect 41588 627770 41644 627779
rect 41588 627705 41644 627714
rect 41794 627441 41822 639101
rect 41890 627441 41918 639693
rect 43126 639571 43178 639577
rect 43126 639513 43178 639519
rect 42164 638278 42220 638287
rect 42164 638213 42220 638222
rect 41972 637686 42028 637695
rect 41972 637621 42028 637630
rect 41986 627515 42014 637621
rect 42068 636206 42124 636215
rect 42068 636141 42124 636150
rect 42082 627589 42110 636141
rect 42070 627583 42122 627589
rect 42070 627525 42122 627531
rect 41974 627509 42026 627515
rect 42178 627483 42206 638213
rect 43030 637055 43082 637061
rect 43030 636997 43082 637003
rect 42932 636798 42988 636807
rect 42932 636733 42988 636742
rect 42838 634983 42890 634989
rect 42838 634925 42890 634931
rect 42850 628075 42878 634925
rect 42946 629735 42974 636733
rect 42934 629729 42986 629735
rect 42934 629671 42986 629677
rect 42836 628066 42892 628075
rect 42836 628001 42892 628010
rect 42838 627879 42890 627885
rect 42838 627821 42890 627827
rect 41974 627451 42026 627457
rect 42164 627474 42220 627483
rect 41782 627435 41834 627441
rect 41782 627377 41834 627383
rect 41878 627435 41930 627441
rect 42164 627409 42220 627418
rect 41878 627377 41930 627383
rect 41782 627065 41834 627071
rect 41782 627007 41834 627013
rect 41794 626632 41822 627007
rect 42166 625363 42218 625369
rect 42166 625305 42218 625311
rect 42178 624782 42206 625305
rect 42850 624703 42878 627821
rect 43042 627737 43070 636997
rect 43138 627756 43166 639513
rect 43030 627731 43082 627737
rect 43138 627728 43262 627756
rect 43030 627673 43082 627679
rect 43126 627583 43178 627589
rect 43126 627525 43178 627531
rect 43030 627509 43082 627515
rect 43030 627451 43082 627457
rect 42934 627435 42986 627441
rect 42934 627377 42986 627383
rect 42166 624697 42218 624703
rect 42166 624639 42218 624645
rect 42838 624697 42890 624703
rect 42838 624639 42890 624645
rect 42178 624161 42206 624639
rect 42838 624549 42890 624555
rect 42838 624491 42890 624497
rect 42166 623513 42218 623519
rect 42166 623455 42218 623461
rect 42178 622965 42206 623455
rect 42164 622146 42220 622155
rect 42164 622081 42220 622090
rect 42178 621748 42206 622081
rect 42850 621669 42878 624491
rect 42166 621663 42218 621669
rect 42166 621605 42218 621611
rect 42838 621663 42890 621669
rect 42838 621605 42890 621611
rect 42178 621125 42206 621605
rect 42836 621554 42892 621563
rect 42836 621489 42892 621498
rect 41780 620962 41836 620971
rect 41780 620897 41836 620906
rect 41794 620490 41822 620897
rect 42166 620405 42218 620411
rect 42166 620347 42218 620353
rect 42178 619929 42206 620347
rect 42262 619073 42314 619079
rect 42262 619015 42314 619021
rect 42070 617889 42122 617895
rect 42070 617831 42122 617837
rect 42082 617456 42110 617831
rect 42274 616804 42302 619015
rect 42192 616776 42302 616804
rect 42262 616705 42314 616711
rect 42262 616647 42314 616653
rect 42274 616171 42302 616647
rect 42192 616143 42302 616171
rect 41780 616078 41836 616087
rect 41780 616013 41836 616022
rect 41794 615606 41822 616013
rect 42850 614195 42878 621489
rect 42946 620411 42974 627377
rect 42934 620405 42986 620411
rect 42934 620347 42986 620353
rect 42932 620222 42988 620231
rect 42932 620157 42988 620166
rect 42946 616711 42974 620157
rect 43042 619079 43070 627451
rect 43030 619073 43082 619079
rect 43030 619015 43082 619021
rect 43028 618890 43084 618899
rect 43028 618825 43084 618834
rect 42934 616705 42986 616711
rect 42934 616647 42986 616653
rect 42932 616522 42988 616531
rect 42932 616457 42988 616466
rect 42166 614189 42218 614195
rect 42166 614131 42218 614137
rect 42838 614189 42890 614195
rect 42838 614131 42890 614137
rect 42178 613756 42206 614131
rect 42946 613677 42974 616457
rect 42166 613671 42218 613677
rect 42166 613613 42218 613619
rect 42934 613671 42986 613677
rect 42934 613613 42986 613619
rect 42178 613121 42206 613613
rect 43042 612863 43070 618825
rect 43138 617895 43166 627525
rect 43234 625369 43262 627728
rect 43222 625363 43274 625369
rect 43222 625305 43274 625311
rect 43126 617889 43178 617895
rect 43126 617831 43178 617837
rect 42070 612857 42122 612863
rect 42070 612799 42122 612805
rect 43030 612857 43082 612863
rect 43030 612799 43082 612805
rect 42082 612498 42110 612799
rect 41782 603089 41834 603095
rect 41780 603054 41782 603063
rect 41834 603054 41836 603063
rect 41780 602989 41836 602998
rect 41590 602793 41642 602799
rect 41588 602758 41590 602767
rect 41642 602758 41644 602767
rect 41588 602693 41644 602702
rect 41590 602201 41642 602207
rect 41588 602166 41590 602175
rect 41642 602166 41644 602175
rect 41588 602101 41644 602110
rect 41782 601609 41834 601615
rect 41780 601574 41782 601583
rect 41834 601574 41836 601583
rect 41780 601509 41836 601518
rect 41780 601056 41836 601065
rect 41780 600991 41782 601000
rect 41834 600991 41836 601000
rect 43222 601017 43274 601023
rect 41782 600959 41834 600965
rect 43222 600959 43274 600965
rect 41588 599946 41644 599955
rect 41588 599881 41590 599890
rect 41642 599881 41644 599890
rect 41590 599849 41642 599855
rect 41780 599058 41836 599067
rect 41780 598993 41782 599002
rect 41834 598993 41836 599002
rect 41782 598961 41834 598967
rect 41492 598318 41548 598327
rect 41492 598253 41548 598262
rect 34388 597282 34444 597291
rect 34388 597217 34444 597226
rect 23060 590770 23116 590779
rect 23060 590705 23116 590714
rect 23074 590335 23102 590705
rect 23060 590326 23116 590335
rect 23060 590261 23116 590270
rect 34402 585591 34430 597217
rect 34484 595358 34540 595367
rect 34484 595293 34540 595302
rect 34388 585582 34444 585591
rect 34388 585517 34444 585526
rect 34498 585443 34526 595293
rect 34484 585434 34540 585443
rect 34484 585369 34540 585378
rect 41506 584563 41534 598253
rect 41588 597874 41644 597883
rect 41588 597809 41644 597818
rect 41602 597767 41630 597809
rect 41590 597761 41642 597767
rect 41590 597703 41642 597709
rect 42934 597761 42986 597767
rect 42934 597703 42986 597709
rect 42068 597134 42124 597143
rect 42068 597069 42124 597078
rect 41684 596394 41740 596403
rect 41684 596329 41740 596338
rect 41588 591362 41644 591371
rect 41588 591297 41644 591306
rect 41602 590779 41630 591297
rect 41588 590770 41644 590779
rect 41588 590705 41590 590714
rect 41642 590705 41644 590714
rect 41590 590673 41642 590679
rect 41698 590414 41726 596329
rect 41876 596024 41932 596033
rect 41876 595959 41932 595968
rect 41780 594174 41836 594183
rect 41780 594109 41836 594118
rect 41794 593993 41822 594109
rect 41782 593987 41834 593993
rect 41782 593929 41834 593935
rect 41780 593582 41836 593591
rect 41780 593517 41782 593526
rect 41834 593517 41836 593526
rect 41782 593485 41834 593491
rect 41780 592620 41836 592629
rect 41780 592555 41782 592564
rect 41834 592555 41836 592564
rect 41782 592523 41834 592529
rect 41780 592102 41836 592111
rect 41780 592037 41836 592046
rect 41794 591255 41822 592037
rect 41782 591249 41834 591255
rect 41782 591191 41834 591197
rect 41698 590386 41822 590414
rect 41492 584554 41548 584563
rect 41492 584489 41548 584498
rect 41794 584373 41822 590386
rect 41782 584367 41834 584373
rect 41782 584309 41834 584315
rect 41890 584225 41918 595959
rect 41972 595062 42028 595071
rect 41972 594997 42028 595006
rect 41986 584299 42014 594997
rect 41974 584293 42026 584299
rect 42082 584267 42110 597069
rect 42164 594470 42220 594479
rect 42164 594405 42220 594414
rect 41974 584235 42026 584241
rect 42068 584258 42124 584267
rect 41878 584219 41930 584225
rect 42178 584225 42206 594405
rect 42742 593987 42794 593993
rect 42742 593929 42794 593935
rect 42452 592990 42508 592999
rect 42452 592925 42508 592934
rect 42068 584193 42124 584202
rect 42166 584219 42218 584225
rect 41878 584161 41930 584167
rect 42166 584161 42218 584167
rect 41878 583997 41930 584003
rect 41878 583939 41930 583945
rect 41890 583445 41918 583939
rect 42466 583707 42494 592925
rect 42454 583701 42506 583707
rect 42454 583643 42506 583649
rect 42166 582147 42218 582153
rect 42166 582089 42218 582095
rect 42178 581605 42206 582089
rect 42070 581407 42122 581413
rect 42070 581349 42122 581355
rect 42082 580974 42110 581349
rect 42754 580303 42782 593929
rect 42838 591249 42890 591255
rect 42838 591191 42890 591197
rect 42070 580297 42122 580303
rect 42070 580239 42122 580245
rect 42742 580297 42794 580303
rect 42742 580239 42794 580245
rect 42082 579790 42110 580239
rect 42742 580149 42794 580155
rect 42742 580091 42794 580097
rect 42166 579039 42218 579045
rect 42166 578981 42218 578987
rect 42178 578569 42206 578981
rect 42754 578305 42782 580091
rect 42850 579045 42878 591191
rect 42946 582153 42974 597703
rect 43126 593543 43178 593549
rect 43126 593485 43178 593491
rect 43030 592581 43082 592587
rect 43030 592523 43082 592529
rect 42934 582147 42986 582153
rect 42934 582089 42986 582095
rect 43042 582024 43070 592523
rect 42946 581996 43070 582024
rect 42838 579039 42890 579045
rect 42838 578981 42890 578987
rect 42836 578782 42892 578791
rect 42836 578717 42892 578726
rect 42070 578299 42122 578305
rect 42070 578241 42122 578247
rect 42742 578299 42794 578305
rect 42742 578241 42794 578247
rect 42082 577940 42110 578241
rect 42166 577707 42218 577713
rect 42166 577649 42218 577655
rect 42178 577274 42206 577649
rect 42166 577189 42218 577195
rect 42166 577131 42218 577137
rect 42178 576992 42206 577131
rect 42082 576964 42206 576992
rect 42082 576756 42110 576964
rect 42166 574673 42218 574679
rect 42166 574615 42218 574621
rect 42178 574240 42206 574615
rect 42356 574490 42412 574499
rect 42356 574425 42412 574434
rect 42166 574155 42218 574161
rect 42166 574097 42218 574103
rect 42178 573574 42206 574097
rect 42166 573489 42218 573495
rect 42166 573431 42218 573437
rect 42178 573292 42206 573431
rect 42082 573264 42206 573292
rect 42082 572982 42110 573264
rect 42166 572823 42218 572829
rect 42166 572765 42218 572771
rect 42178 572390 42206 572765
rect 42166 570899 42218 570905
rect 42166 570841 42218 570847
rect 42178 570540 42206 570841
rect 42370 570461 42398 574425
rect 42740 574046 42796 574055
rect 42740 573981 42796 573990
rect 42166 570455 42218 570461
rect 42166 570397 42218 570403
rect 42358 570455 42410 570461
rect 42358 570397 42410 570403
rect 42178 570254 42206 570397
rect 42082 570226 42206 570254
rect 42358 570307 42410 570313
rect 42358 570249 42410 570255
rect 42082 569948 42110 570226
rect 42070 569715 42122 569721
rect 42070 569657 42122 569663
rect 42082 569282 42110 569657
rect 41782 559873 41834 559879
rect 41780 559838 41782 559847
rect 41834 559838 41836 559847
rect 41780 559773 41836 559782
rect 42370 559403 42398 570249
rect 42754 569721 42782 573981
rect 42850 572829 42878 578717
rect 42946 577713 42974 581996
rect 43030 581925 43082 581931
rect 43030 581867 43082 581873
rect 43042 579952 43070 581867
rect 43138 580155 43166 593485
rect 43126 580149 43178 580155
rect 43126 580091 43178 580097
rect 43042 579924 43166 579952
rect 43030 579853 43082 579859
rect 43030 579795 43082 579801
rect 42934 577707 42986 577713
rect 42934 577649 42986 577655
rect 42932 577598 42988 577607
rect 42932 577533 42988 577542
rect 42838 572823 42890 572829
rect 42838 572765 42890 572771
rect 42946 570905 42974 577533
rect 43042 574161 43070 579795
rect 43138 574679 43166 579924
rect 43126 574673 43178 574679
rect 43126 574615 43178 574621
rect 43030 574155 43082 574161
rect 43030 574097 43082 574103
rect 42934 570899 42986 570905
rect 42934 570841 42986 570847
rect 42742 569715 42794 569721
rect 42742 569657 42794 569663
rect 42356 559394 42412 559403
rect 42356 559329 42412 559338
rect 41782 558837 41834 558843
rect 41780 558802 41782 558811
rect 41834 558802 41836 558811
rect 41780 558737 41836 558746
rect 43234 558399 43262 600959
rect 43330 599913 43358 643689
rect 43414 629729 43466 629735
rect 43414 629671 43466 629677
rect 43426 624555 43454 629671
rect 43702 629285 43754 629291
rect 43702 629227 43754 629233
rect 43510 627731 43562 627737
rect 43510 627673 43562 627679
rect 43414 624549 43466 624555
rect 43414 624491 43466 624497
rect 43522 623519 43550 627673
rect 43510 623513 43562 623519
rect 43510 623455 43562 623461
rect 43714 619912 43742 629227
rect 43426 619884 43742 619912
rect 43426 601412 43454 619884
rect 43810 610574 43838 644133
rect 44386 619195 44414 970515
rect 44470 945857 44522 945863
rect 44470 945799 44522 945805
rect 44372 619186 44428 619195
rect 44372 619121 44428 619130
rect 43522 610546 43838 610574
rect 43522 601615 43550 610546
rect 43510 601609 43562 601615
rect 43510 601551 43562 601557
rect 43426 601384 43550 601412
rect 43318 599907 43370 599913
rect 43318 599849 43370 599855
rect 43522 599025 43550 601384
rect 44374 599907 44426 599913
rect 44374 599849 44426 599855
rect 43510 599019 43562 599025
rect 43510 598961 43562 598967
rect 43522 596213 43550 598961
rect 43510 596207 43562 596213
rect 43510 596149 43562 596155
rect 43510 584737 43562 584743
rect 43510 584679 43562 584685
rect 43414 584219 43466 584225
rect 43414 584161 43466 584167
rect 43318 583701 43370 583707
rect 43318 583643 43370 583649
rect 43330 581931 43358 583643
rect 43318 581925 43370 581931
rect 43318 581867 43370 581873
rect 43426 579859 43454 584161
rect 43522 581413 43550 584679
rect 43702 584367 43754 584373
rect 43702 584309 43754 584315
rect 43510 581407 43562 581413
rect 43510 581349 43562 581355
rect 43414 579853 43466 579859
rect 43414 579795 43466 579801
rect 43714 579360 43742 584309
rect 43798 584293 43850 584299
rect 43798 584235 43850 584241
rect 43522 579332 43742 579360
rect 43522 577195 43550 579332
rect 43810 579212 43838 584235
rect 43618 579184 43838 579212
rect 43510 577189 43562 577195
rect 43510 577131 43562 577137
rect 43618 573495 43646 579184
rect 43606 573489 43658 573495
rect 43606 573431 43658 573437
rect 41782 558393 41834 558399
rect 41780 558358 41782 558367
rect 43222 558393 43274 558399
rect 41834 558358 41836 558367
rect 43222 558335 43274 558341
rect 41780 558293 41836 558302
rect 41780 557914 41836 557923
rect 41780 557849 41782 557858
rect 41834 557849 41836 557858
rect 43606 557875 43658 557881
rect 41782 557817 41834 557823
rect 43606 557817 43658 557823
rect 42260 555398 42316 555407
rect 42260 555333 42316 555342
rect 41588 554658 41644 554667
rect 41588 554593 41644 554602
rect 34388 554066 34444 554075
rect 34388 554001 34444 554010
rect 23060 547554 23116 547563
rect 23060 547489 23116 547498
rect 23074 547119 23102 547489
rect 23060 547110 23116 547119
rect 23060 547045 23116 547054
rect 34402 541495 34430 554001
rect 41602 553219 41630 554593
rect 41684 554066 41740 554075
rect 41684 554001 41740 554010
rect 41590 553213 41642 553219
rect 41590 553155 41642 553161
rect 34484 552142 34540 552151
rect 34484 552077 34540 552086
rect 34498 541643 34526 552077
rect 41492 551698 41548 551707
rect 41492 551633 41548 551642
rect 41396 549182 41452 549191
rect 41396 549117 41452 549126
rect 34484 541634 34540 541643
rect 34484 541569 34540 541578
rect 34388 541486 34444 541495
rect 34388 541421 34444 541430
rect 41410 541379 41438 549117
rect 41398 541373 41450 541379
rect 41398 541315 41450 541321
rect 41506 541305 41534 551633
rect 41588 550218 41644 550227
rect 41588 550153 41590 550162
rect 41642 550153 41644 550162
rect 41590 550121 41642 550127
rect 41698 541347 41726 554001
rect 42164 553326 42220 553335
rect 42164 553261 42220 553270
rect 41780 552882 41836 552891
rect 41780 552817 41836 552826
rect 41684 541338 41740 541347
rect 41494 541299 41546 541305
rect 41684 541273 41740 541282
rect 41494 541241 41546 541247
rect 41794 541009 41822 552817
rect 41972 551328 42028 551337
rect 41972 551263 42028 551272
rect 41876 550958 41932 550967
rect 41876 550893 41932 550902
rect 41890 550481 41918 550893
rect 41878 550475 41930 550481
rect 41878 550417 41930 550423
rect 41876 548886 41932 548895
rect 41876 548821 41878 548830
rect 41930 548821 41932 548830
rect 41878 548789 41930 548795
rect 41876 547406 41932 547415
rect 41876 547341 41878 547350
rect 41930 547341 41932 547350
rect 41878 547309 41930 547315
rect 41986 541051 42014 551263
rect 42178 549908 42206 553261
rect 42082 549880 42206 549908
rect 42082 541823 42110 549880
rect 42164 549774 42220 549783
rect 42164 549709 42220 549718
rect 42070 541817 42122 541823
rect 42070 541759 42122 541765
rect 42178 541051 42206 549709
rect 42274 542859 42302 555333
rect 42838 553213 42890 553219
rect 42838 553155 42890 553161
rect 42742 550179 42794 550185
rect 42742 550121 42794 550127
rect 42262 542853 42314 542859
rect 42262 542795 42314 542801
rect 42754 541643 42782 550121
rect 42850 550094 42878 553155
rect 43126 550475 43178 550481
rect 43126 550417 43178 550423
rect 42850 550066 42974 550094
rect 42838 548847 42890 548853
rect 42838 548789 42890 548795
rect 42740 541634 42796 541643
rect 42740 541569 42796 541578
rect 42742 541521 42794 541527
rect 42742 541463 42794 541469
rect 41972 541042 42028 541051
rect 41782 541003 41834 541009
rect 41972 540977 42028 540986
rect 42164 541042 42220 541051
rect 42164 540977 42220 540986
rect 41782 540945 41834 540951
rect 41782 540781 41834 540787
rect 41782 540723 41834 540729
rect 41794 540245 41822 540723
rect 42070 538931 42122 538937
rect 42070 538873 42122 538879
rect 42082 538424 42110 538873
rect 42754 538345 42782 541463
rect 42166 538339 42218 538345
rect 42166 538281 42218 538287
rect 42742 538339 42794 538345
rect 42742 538281 42794 538287
rect 42178 537758 42206 538281
rect 42070 537081 42122 537087
rect 42070 537023 42122 537029
rect 42082 536574 42110 537023
rect 42850 535829 42878 548789
rect 42946 538937 42974 550066
rect 43138 543248 43166 550417
rect 43138 543220 43262 543248
rect 43030 542853 43082 542859
rect 43234 542804 43262 543220
rect 43030 542795 43082 542801
rect 42934 538931 42986 538937
rect 42934 538873 42986 538879
rect 42934 538783 42986 538789
rect 42934 538725 42986 538731
rect 42070 535823 42122 535829
rect 42070 535765 42122 535771
rect 42838 535823 42890 535829
rect 42838 535765 42890 535771
rect 42082 535390 42110 535765
rect 42836 535714 42892 535723
rect 42836 535649 42892 535658
rect 42164 535122 42220 535131
rect 42164 535057 42220 535066
rect 42178 534724 42206 535057
rect 42166 534491 42218 534497
rect 42166 534433 42218 534439
rect 42178 534058 42206 534433
rect 42166 533973 42218 533979
rect 42166 533915 42218 533921
rect 42178 533776 42206 533915
rect 42082 533748 42206 533776
rect 42082 533540 42110 533748
rect 42850 531537 42878 535649
rect 42946 534497 42974 538725
rect 42934 534491 42986 534497
rect 42934 534433 42986 534439
rect 42166 531531 42218 531537
rect 42166 531473 42218 531479
rect 42838 531531 42890 531537
rect 42838 531473 42890 531479
rect 42178 531024 42206 531473
rect 42836 531422 42892 531431
rect 42836 531357 42892 531366
rect 41972 530682 42028 530691
rect 41972 530617 42028 530626
rect 41986 530401 42014 530617
rect 42070 530199 42122 530205
rect 42070 530141 42122 530147
rect 42082 529766 42110 530141
rect 41780 529646 41836 529655
rect 41780 529581 41836 529590
rect 41794 529205 41822 529581
rect 42178 527245 42206 527365
rect 42166 527239 42218 527245
rect 42166 527181 42218 527187
rect 42850 527097 42878 531357
rect 43042 527245 43070 542795
rect 43138 542776 43262 542804
rect 43138 541916 43166 542776
rect 43138 541888 43358 541916
rect 43126 541817 43178 541823
rect 43126 541759 43178 541765
rect 43138 533979 43166 541759
rect 43222 541373 43274 541379
rect 43222 541315 43274 541321
rect 43234 538789 43262 541315
rect 43222 538783 43274 538789
rect 43222 538725 43274 538731
rect 43330 537087 43358 541888
rect 43414 541299 43466 541305
rect 43414 541241 43466 541247
rect 43318 537081 43370 537087
rect 43318 537023 43370 537029
rect 43126 533973 43178 533979
rect 43126 533915 43178 533921
rect 43426 533776 43454 541241
rect 43138 533748 43454 533776
rect 43138 530205 43166 533748
rect 43126 530199 43178 530205
rect 43126 530141 43178 530147
rect 43618 529934 43646 557817
rect 43234 529906 43646 529934
rect 43030 527239 43082 527245
rect 43030 527181 43082 527187
rect 42070 527091 42122 527097
rect 42070 527033 42122 527039
rect 42838 527091 42890 527097
rect 42838 527033 42890 527039
rect 42082 526732 42110 527033
rect 41780 526538 41836 526547
rect 41780 526473 41836 526482
rect 41794 526066 41822 526473
rect 41782 432297 41834 432303
rect 41780 432262 41782 432271
rect 41834 432262 41836 432271
rect 41780 432197 41836 432206
rect 41782 431779 41834 431785
rect 41780 431744 41782 431753
rect 41834 431744 41836 431753
rect 41780 431679 41836 431688
rect 41590 431409 41642 431415
rect 41588 431374 41590 431383
rect 41642 431374 41644 431383
rect 41588 431309 41644 431318
rect 43234 430823 43262 529906
rect 41782 430817 41834 430823
rect 41780 430782 41782 430791
rect 43222 430817 43274 430823
rect 41834 430782 41836 430791
rect 43222 430759 43274 430765
rect 41780 430717 41836 430726
rect 41780 430264 41836 430273
rect 41780 430199 41782 430208
rect 41834 430199 41836 430208
rect 43318 430225 43370 430231
rect 41782 430167 41834 430173
rect 43318 430167 43370 430173
rect 40724 429894 40780 429903
rect 40724 429829 40780 429838
rect 40738 429015 40766 429829
rect 40724 429006 40780 429015
rect 40724 428941 40780 428950
rect 28820 419978 28876 419987
rect 28820 419913 28876 419922
rect 28834 419543 28862 419913
rect 28820 419534 28876 419543
rect 28820 419469 28876 419478
rect 40738 417577 40766 428941
rect 41588 428562 41644 428571
rect 41588 428497 41590 428506
rect 41642 428497 41644 428506
rect 43222 428523 43274 428529
rect 41590 428465 41642 428471
rect 43222 428465 43274 428471
rect 41876 425232 41932 425241
rect 41876 425167 41932 425176
rect 41780 423308 41836 423317
rect 41780 423243 41836 423252
rect 41588 421606 41644 421615
rect 41588 421541 41644 421550
rect 41602 421129 41630 421541
rect 41590 421123 41642 421129
rect 41590 421065 41642 421071
rect 41588 421014 41644 421023
rect 41588 420949 41590 420958
rect 41642 420949 41644 420958
rect 41590 420917 41642 420923
rect 41794 420537 41822 423243
rect 41782 420531 41834 420537
rect 41782 420473 41834 420479
rect 41780 419830 41836 419839
rect 41780 419765 41782 419774
rect 41834 419765 41836 419774
rect 41782 419733 41834 419739
rect 40726 417571 40778 417577
rect 40726 417513 40778 417519
rect 41890 413433 41918 425167
rect 41972 422790 42028 422799
rect 41972 422725 42028 422734
rect 41986 420759 42014 422725
rect 43030 421123 43082 421129
rect 43030 421065 43082 421071
rect 42934 420975 42986 420981
rect 42934 420917 42986 420923
rect 41974 420753 42026 420759
rect 41974 420695 42026 420701
rect 42838 420531 42890 420537
rect 42838 420473 42890 420479
rect 41878 413427 41930 413433
rect 41878 413369 41930 413375
rect 41878 413205 41930 413211
rect 41878 413147 41930 413153
rect 41890 412624 41918 413147
rect 41972 411246 42028 411255
rect 41972 411181 42028 411190
rect 41986 410805 42014 411181
rect 42070 410541 42122 410547
rect 42070 410483 42122 410489
rect 42082 410182 42110 410483
rect 42850 409511 42878 420473
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42838 409505 42890 409511
rect 42838 409447 42890 409453
rect 42178 408965 42206 409447
rect 42946 408253 42974 420917
rect 42166 408247 42218 408253
rect 42166 408189 42218 408195
rect 42934 408247 42986 408253
rect 42934 408189 42986 408195
rect 42178 407769 42206 408189
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 43042 406921 43070 421065
rect 43126 420753 43178 420759
rect 43126 420695 43178 420701
rect 43138 407513 43166 420695
rect 43126 407507 43178 407513
rect 43126 407449 43178 407455
rect 42166 406915 42218 406921
rect 42166 406857 42218 406863
rect 43030 406915 43082 406921
rect 43030 406857 43082 406863
rect 42178 406482 42206 406857
rect 41780 406066 41836 406075
rect 41780 406001 41836 406010
rect 41794 405929 41822 406001
rect 41780 403846 41836 403855
rect 41780 403781 41836 403790
rect 41794 403448 41822 403781
rect 41780 403106 41836 403115
rect 41780 403041 41836 403050
rect 41794 402782 41822 403041
rect 41780 402514 41836 402523
rect 41780 402449 41836 402458
rect 41794 402157 41822 402449
rect 41780 401922 41836 401931
rect 41780 401857 41836 401866
rect 41794 401598 41822 401857
rect 41780 399998 41836 400007
rect 41780 399933 41836 399942
rect 41794 399748 41822 399933
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41876 398962 41932 398971
rect 41876 398897 41932 398906
rect 41890 398490 41918 398897
rect 41876 390962 41932 390971
rect 41876 390897 41932 390906
rect 41890 389351 41918 390897
rect 41876 389342 41932 389351
rect 41876 389277 41932 389286
rect 41782 389081 41834 389087
rect 41780 389046 41782 389055
rect 41834 389046 41836 389055
rect 41780 388981 41836 388990
rect 41590 388785 41642 388791
rect 41588 388750 41590 388759
rect 41642 388750 41644 388759
rect 41588 388685 41644 388694
rect 41782 388045 41834 388051
rect 41780 388010 41782 388019
rect 41834 388010 41836 388019
rect 41780 387945 41836 387954
rect 41782 387601 41834 387607
rect 41780 387566 41782 387575
rect 41834 387566 41836 387575
rect 41780 387501 41836 387510
rect 41780 387048 41836 387057
rect 41780 386983 41782 386992
rect 41834 386983 41836 386992
rect 41782 386951 41834 386957
rect 41890 386095 41918 389277
rect 41876 386086 41932 386095
rect 41876 386021 41932 386030
rect 43234 385239 43262 428465
rect 43330 387607 43358 430167
rect 44278 417571 44330 417577
rect 44278 417513 44330 417519
rect 43318 387601 43370 387607
rect 43318 387543 43370 387549
rect 43510 387009 43562 387015
rect 43510 386951 43562 386957
rect 41590 385233 41642 385239
rect 34484 385198 34540 385207
rect 34484 385133 34540 385142
rect 41588 385198 41590 385207
rect 43222 385233 43274 385239
rect 41642 385198 41644 385207
rect 43222 385175 43274 385181
rect 41588 385133 41644 385142
rect 34498 381613 34526 385133
rect 41876 382016 41932 382025
rect 41876 381951 41932 381960
rect 34486 381607 34538 381613
rect 34486 381549 34538 381555
rect 41780 380166 41836 380175
rect 41780 380101 41782 380110
rect 41834 380101 41836 380110
rect 41782 380069 41834 380075
rect 41780 379574 41836 379583
rect 41780 379509 41836 379518
rect 41588 378834 41644 378843
rect 41588 378769 41644 378778
rect 41602 378505 41630 378769
rect 41590 378499 41642 378505
rect 41590 378441 41642 378447
rect 41588 378390 41644 378399
rect 41794 378357 41822 379509
rect 41588 378325 41644 378334
rect 41782 378351 41834 378357
rect 41602 378283 41630 378325
rect 41782 378293 41834 378299
rect 41590 378277 41642 378283
rect 41590 378219 41642 378225
rect 41780 378094 41836 378103
rect 41780 378029 41836 378038
rect 41794 377617 41822 378029
rect 41782 377611 41834 377617
rect 41782 377553 41834 377559
rect 40244 377354 40300 377363
rect 40244 377289 40300 377298
rect 28820 376762 28876 376771
rect 28820 376697 28876 376706
rect 28834 376327 28862 376697
rect 40258 376581 40286 377289
rect 41780 376614 41836 376623
rect 40246 376575 40298 376581
rect 41780 376549 41782 376558
rect 40246 376517 40298 376523
rect 41834 376549 41836 376558
rect 41782 376517 41834 376523
rect 28820 376318 28876 376327
rect 28820 376253 28876 376262
rect 41890 370217 41918 381951
rect 43318 381607 43370 381613
rect 43318 381549 43370 381555
rect 42838 380127 42890 380133
rect 42838 380069 42890 380075
rect 42742 378351 42794 378357
rect 42742 378293 42794 378299
rect 41878 370211 41930 370217
rect 41878 370153 41930 370159
rect 41878 369989 41930 369995
rect 41878 369931 41930 369937
rect 41890 369445 41918 369931
rect 41972 368178 42028 368187
rect 41972 368113 42028 368122
rect 41986 367632 42014 368113
rect 42070 367399 42122 367405
rect 42070 367341 42122 367347
rect 42082 366966 42110 367341
rect 42070 366289 42122 366295
rect 42070 366231 42122 366237
rect 42082 365782 42110 366231
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42178 364569 42206 364973
rect 42754 364445 42782 378293
rect 42850 366295 42878 380069
rect 43126 378499 43178 378505
rect 43126 378441 43178 378447
rect 43030 378277 43082 378283
rect 43030 378219 43082 378225
rect 42934 377611 42986 377617
rect 42934 377553 42986 377559
rect 42838 366289 42890 366295
rect 42838 366231 42890 366237
rect 42946 365037 42974 377553
rect 42934 365031 42986 365037
rect 42934 364973 42986 364979
rect 42070 364439 42122 364445
rect 42070 364381 42122 364387
rect 42742 364439 42794 364445
rect 42742 364381 42794 364387
rect 42082 363932 42110 364381
rect 43042 363705 43070 378219
rect 42166 363699 42218 363705
rect 42166 363641 42218 363647
rect 43030 363699 43082 363705
rect 43030 363641 43082 363647
rect 42178 363266 42206 363641
rect 41780 362850 41836 362859
rect 41780 362785 41836 362794
rect 41794 362748 41822 362785
rect 43138 360671 43166 378441
rect 42166 360665 42218 360671
rect 42166 360607 42218 360613
rect 43126 360665 43178 360671
rect 43126 360607 43178 360613
rect 42178 360232 42206 360607
rect 41780 359890 41836 359899
rect 41780 359825 41836 359834
rect 41794 359601 41822 359825
rect 41780 359446 41836 359455
rect 41780 359381 41836 359390
rect 41794 358974 41822 359381
rect 41780 358706 41836 358715
rect 41780 358641 41836 358650
rect 41794 358382 41822 358641
rect 41780 356930 41836 356939
rect 41780 356865 41836 356874
rect 41794 356565 41822 356865
rect 41780 356486 41836 356495
rect 41780 356421 41836 356430
rect 41794 355940 41822 356421
rect 41780 355598 41836 355607
rect 41780 355533 41836 355542
rect 41794 355274 41822 355533
rect 41782 345939 41834 345945
rect 41780 345904 41782 345913
rect 41834 345904 41836 345913
rect 41780 345839 41836 345848
rect 41590 345569 41642 345575
rect 41588 345534 41590 345543
rect 41642 345534 41644 345543
rect 41588 345469 41644 345478
rect 41782 344829 41834 344835
rect 41780 344794 41782 344803
rect 41834 344794 41836 344803
rect 41780 344729 41836 344738
rect 41782 344385 41834 344391
rect 41780 344350 41782 344359
rect 41834 344350 41836 344359
rect 41780 344285 41836 344294
rect 41780 343906 41836 343915
rect 41780 343841 41782 343850
rect 41834 343841 41836 343850
rect 43222 343867 43274 343873
rect 41782 343809 41834 343815
rect 43222 343809 43274 343815
rect 41782 343349 41834 343355
rect 41780 343314 41782 343323
rect 41834 343314 41836 343323
rect 41780 343249 41836 343258
rect 41782 342387 41834 342393
rect 41780 342352 41782 342361
rect 41834 342352 41836 342361
rect 41780 342287 41836 342296
rect 41590 342017 41642 342023
rect 41588 341982 41590 341991
rect 41642 341982 41644 341991
rect 41588 341917 41644 341926
rect 41876 338874 41932 338883
rect 41876 338809 41932 338818
rect 41780 336950 41836 336959
rect 41780 336885 41836 336894
rect 41588 336210 41644 336219
rect 41588 336145 41644 336154
rect 41602 335289 41630 336145
rect 41590 335283 41642 335289
rect 41590 335225 41642 335231
rect 41588 335174 41644 335183
rect 41588 335109 41644 335118
rect 41602 334697 41630 335109
rect 41794 334993 41822 336885
rect 41782 334987 41834 334993
rect 41782 334929 41834 334935
rect 41780 334878 41836 334887
rect 41780 334813 41836 334822
rect 41590 334691 41642 334697
rect 41590 334633 41642 334639
rect 41794 334549 41822 334813
rect 41782 334543 41834 334549
rect 41782 334485 41834 334491
rect 28820 333546 28876 333555
rect 28820 333481 28876 333490
rect 28834 333111 28862 333481
rect 41780 333398 41836 333407
rect 41780 333333 41782 333342
rect 41834 333333 41836 333342
rect 41782 333301 41834 333307
rect 28820 333102 28876 333111
rect 28820 333037 28876 333046
rect 41890 327075 41918 338809
rect 42452 335766 42508 335775
rect 42508 335724 42590 335752
rect 42452 335701 42508 335710
rect 42562 328334 42590 335724
rect 43126 335283 43178 335289
rect 43126 335225 43178 335231
rect 42934 334987 42986 334993
rect 42934 334929 42986 334935
rect 42838 334543 42890 334549
rect 42838 334485 42890 334491
rect 42466 328306 42590 328334
rect 41878 327069 41930 327075
rect 41878 327011 41930 327017
rect 41878 326773 41930 326779
rect 41878 326715 41930 326721
rect 41890 326266 41918 326715
rect 42466 326557 42494 328306
rect 42454 326551 42506 326557
rect 42454 326493 42506 326499
rect 41780 324962 41836 324971
rect 41780 324897 41836 324906
rect 41794 324416 41822 324897
rect 42166 324183 42218 324189
rect 42166 324125 42218 324131
rect 42178 323750 42206 324125
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42178 322566 42206 323089
rect 42850 321821 42878 334485
rect 42946 323153 42974 334929
rect 43030 334691 43082 334697
rect 43030 334633 43082 334639
rect 43042 326705 43070 334633
rect 43030 326699 43082 326705
rect 43030 326641 43082 326647
rect 43030 326551 43082 326557
rect 43030 326493 43082 326499
rect 42934 323147 42986 323153
rect 42934 323089 42986 323095
rect 42934 322999 42986 323005
rect 42934 322941 42986 322947
rect 42070 321815 42122 321821
rect 42070 321757 42122 321763
rect 42838 321815 42890 321821
rect 42838 321757 42890 321763
rect 42082 321382 42110 321757
rect 42166 321075 42218 321081
rect 42166 321017 42218 321023
rect 42178 320716 42206 321017
rect 42946 320637 42974 322941
rect 42166 320631 42218 320637
rect 42166 320573 42218 320579
rect 42934 320631 42986 320637
rect 42934 320573 42986 320579
rect 42178 320081 42206 320573
rect 41780 319782 41836 319791
rect 41780 319717 41836 319726
rect 41794 319532 41822 319717
rect 43042 317529 43070 326493
rect 43138 321081 43166 335225
rect 43126 321075 43178 321081
rect 43126 321017 43178 321023
rect 42166 317523 42218 317529
rect 42166 317465 42218 317471
rect 43030 317523 43082 317529
rect 43030 317465 43082 317471
rect 42178 317045 42206 317465
rect 41780 316822 41836 316831
rect 41780 316757 41836 316766
rect 41794 316424 41822 316757
rect 41780 316082 41836 316091
rect 41780 316017 41836 316026
rect 41794 315758 41822 316017
rect 41780 315490 41836 315499
rect 41780 315425 41836 315434
rect 41794 315205 41822 315425
rect 41876 313714 41932 313723
rect 41876 313649 41932 313658
rect 41890 313390 41918 313649
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312724 41822 313205
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 41782 302723 41834 302729
rect 41780 302688 41782 302697
rect 41834 302688 41836 302697
rect 41780 302623 41836 302632
rect 41590 302353 41642 302359
rect 41588 302318 41590 302327
rect 41642 302318 41644 302327
rect 41588 302253 41644 302262
rect 41782 301613 41834 301619
rect 41780 301578 41782 301587
rect 41834 301578 41836 301587
rect 41780 301513 41836 301522
rect 43234 301249 43262 343809
rect 43330 342023 43358 381549
rect 43522 344391 43550 386951
rect 44182 385233 44234 385239
rect 44182 385175 44234 385181
rect 43510 344385 43562 344391
rect 43510 344327 43562 344333
rect 43414 343349 43466 343355
rect 43414 343291 43466 343297
rect 43318 342017 43370 342023
rect 43318 341959 43370 341965
rect 43318 326699 43370 326705
rect 43318 326641 43370 326647
rect 43330 323005 43358 326641
rect 43318 322999 43370 323005
rect 43318 322941 43370 322947
rect 43426 318417 43454 343291
rect 43510 342387 43562 342393
rect 43510 342329 43562 342335
rect 43414 318411 43466 318417
rect 43414 318353 43466 318359
rect 43522 318288 43550 342329
rect 43330 318260 43550 318288
rect 41782 301243 41834 301249
rect 41780 301208 41782 301217
rect 43222 301243 43274 301249
rect 41834 301208 41836 301217
rect 43222 301185 43274 301191
rect 41780 301143 41836 301152
rect 41780 300690 41836 300699
rect 41780 300625 41782 300634
rect 41834 300625 41836 300634
rect 41782 300593 41834 300599
rect 41782 300133 41834 300139
rect 41780 300098 41782 300107
rect 41834 300098 41836 300107
rect 41780 300033 41836 300042
rect 41782 299689 41834 299695
rect 41780 299654 41782 299663
rect 41834 299654 41836 299663
rect 41780 299589 41836 299598
rect 41590 299393 41642 299399
rect 41588 299358 41590 299367
rect 43222 299393 43274 299399
rect 41642 299358 41644 299367
rect 43222 299335 43274 299341
rect 41588 299293 41644 299302
rect 41782 298653 41834 298659
rect 41780 298618 41782 298627
rect 41834 298618 41836 298627
rect 41780 298553 41836 298562
rect 43234 296654 43262 299335
rect 43330 298659 43358 318260
rect 43414 318189 43466 318195
rect 43414 318131 43466 318137
rect 43426 299695 43454 318131
rect 43606 300651 43658 300657
rect 43606 300593 43658 300599
rect 43510 300133 43562 300139
rect 43510 300075 43562 300081
rect 43414 299689 43466 299695
rect 43414 299631 43466 299637
rect 43318 298653 43370 298659
rect 43318 298595 43370 298601
rect 43522 296654 43550 300075
rect 43234 296626 43358 296654
rect 41972 295658 42028 295667
rect 41972 295593 42028 295602
rect 41780 293734 41836 293743
rect 41780 293669 41836 293678
rect 41588 292994 41644 293003
rect 41588 292929 41644 292938
rect 41602 291629 41630 292929
rect 41590 291623 41642 291629
rect 41590 291565 41642 291571
rect 41588 291514 41644 291523
rect 41588 291449 41644 291458
rect 41602 291185 41630 291449
rect 41590 291179 41642 291185
rect 41590 291121 41642 291127
rect 41794 290963 41822 293669
rect 41876 292624 41932 292633
rect 41876 292559 41932 292568
rect 41890 292369 41918 292559
rect 41878 292363 41930 292369
rect 41878 292305 41930 292311
rect 41876 292254 41932 292263
rect 41876 292189 41932 292198
rect 41890 291111 41918 292189
rect 41878 291105 41930 291111
rect 41878 291047 41930 291053
rect 41782 290957 41834 290963
rect 41782 290899 41834 290905
rect 28820 290478 28876 290487
rect 28820 290413 28876 290422
rect 28834 289895 28862 290413
rect 41780 290182 41836 290191
rect 41780 290117 41782 290126
rect 41834 290117 41836 290126
rect 41782 290085 41834 290091
rect 28820 289886 28876 289895
rect 28820 289821 28876 289830
rect 41986 283859 42014 295593
rect 43126 292363 43178 292369
rect 43126 292305 43178 292311
rect 43030 291623 43082 291629
rect 43030 291565 43082 291571
rect 42742 291179 42794 291185
rect 42742 291121 42794 291127
rect 41974 283853 42026 283859
rect 41974 283795 42026 283801
rect 41974 283557 42026 283563
rect 41974 283499 42026 283505
rect 41986 283050 42014 283499
rect 41780 281746 41836 281755
rect 41780 281681 41836 281690
rect 41794 281200 41822 281681
rect 42166 281115 42218 281121
rect 42166 281057 42218 281063
rect 42178 280534 42206 281057
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42754 278605 42782 291121
rect 42934 291105 42986 291111
rect 42934 291047 42986 291053
rect 42838 290957 42890 290963
rect 42838 290899 42890 290905
rect 42850 279937 42878 290899
rect 42838 279931 42890 279937
rect 42838 279873 42890 279879
rect 42166 278599 42218 278605
rect 42166 278541 42218 278547
rect 42742 278599 42794 278605
rect 42742 278541 42794 278547
rect 42178 278166 42206 278541
rect 42166 277859 42218 277865
rect 42166 277801 42218 277807
rect 42178 277500 42206 277801
rect 42946 277421 42974 291047
rect 43042 277865 43070 291565
rect 43030 277859 43082 277865
rect 43030 277801 43082 277807
rect 42070 277415 42122 277421
rect 42070 277357 42122 277363
rect 42934 277415 42986 277421
rect 42934 277357 42986 277363
rect 42082 276908 42110 277357
rect 41780 276566 41836 276575
rect 41780 276501 41836 276510
rect 41794 276316 41822 276501
rect 43138 274313 43166 292305
rect 42166 274307 42218 274313
rect 42166 274249 42218 274255
rect 43126 274307 43178 274313
rect 43126 274249 43178 274255
rect 42178 273845 42206 274249
rect 41780 273606 41836 273615
rect 41780 273541 41836 273550
rect 41794 273208 41822 273541
rect 41780 272866 41836 272875
rect 41780 272801 41836 272810
rect 41794 272542 41822 272801
rect 41780 272422 41836 272431
rect 41780 272357 41836 272366
rect 41794 272024 41822 272357
rect 41780 270498 41836 270507
rect 41780 270433 41836 270442
rect 41794 270174 41822 270433
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41780 269166 41836 269175
rect 41780 269101 41836 269110
rect 41794 268877 41822 269101
rect 41590 259729 41642 259735
rect 41588 259694 41590 259703
rect 41642 259694 41644 259703
rect 41588 259629 41644 259638
rect 43222 259211 43274 259217
rect 43222 259153 43274 259159
rect 41782 258989 41834 258995
rect 41780 258954 41782 258963
rect 41834 258954 41836 258963
rect 41780 258889 41836 258898
rect 41782 258397 41834 258403
rect 41780 258362 41782 258371
rect 41834 258362 41836 258371
rect 41780 258297 41836 258306
rect 41782 258027 41834 258033
rect 41780 257992 41782 258001
rect 41834 257992 41836 258001
rect 41780 257927 41836 257936
rect 41780 257474 41836 257483
rect 41780 257409 41782 257418
rect 41834 257409 41836 257418
rect 41782 257377 41834 257383
rect 43234 256923 43262 259153
rect 41782 256917 41834 256923
rect 41780 256882 41782 256891
rect 43222 256917 43274 256923
rect 41834 256882 41836 256891
rect 43222 256859 43274 256865
rect 41780 256817 41836 256826
rect 41782 256547 41834 256553
rect 41780 256512 41782 256521
rect 41834 256512 41836 256521
rect 41780 256447 41836 256456
rect 41780 255994 41836 256003
rect 41780 255929 41782 255938
rect 41834 255929 41836 255938
rect 41782 255897 41834 255903
rect 41782 255437 41834 255443
rect 41780 255402 41782 255411
rect 41834 255402 41836 255411
rect 41780 255337 41836 255346
rect 41876 252442 41932 252451
rect 41876 252377 41932 252386
rect 41780 250518 41836 250527
rect 41780 250453 41836 250462
rect 41588 249778 41644 249787
rect 41588 249713 41644 249722
rect 41602 249301 41630 249713
rect 41590 249295 41642 249301
rect 41590 249237 41642 249243
rect 41588 249186 41644 249195
rect 41588 249121 41644 249130
rect 41602 248413 41630 249121
rect 41590 248407 41642 248413
rect 41590 248349 41642 248355
rect 41588 248298 41644 248307
rect 41588 248233 41644 248242
rect 41602 248117 41630 248233
rect 41590 248111 41642 248117
rect 41590 248053 41642 248059
rect 41794 247969 41822 250453
rect 41782 247963 41834 247969
rect 41782 247905 41834 247911
rect 41590 247741 41642 247747
rect 41588 247706 41590 247715
rect 41642 247706 41644 247715
rect 41588 247641 41644 247650
rect 41588 247262 41644 247271
rect 41588 247197 41644 247206
rect 41602 244861 41630 247197
rect 41684 246670 41740 246679
rect 41684 246605 41740 246614
rect 41590 244855 41642 244861
rect 41590 244797 41642 244803
rect 41698 243381 41726 246605
rect 41686 243375 41738 243381
rect 41686 243317 41738 243323
rect 41890 240643 41918 252377
rect 43126 249295 43178 249301
rect 43126 249237 43178 249243
rect 41972 249038 42028 249047
rect 41972 248973 42028 248982
rect 41986 247895 42014 248973
rect 42838 248407 42890 248413
rect 42838 248349 42890 248355
rect 42742 247963 42794 247969
rect 42742 247905 42794 247911
rect 41974 247889 42026 247895
rect 41974 247831 42026 247837
rect 41878 240637 41930 240643
rect 41878 240579 41930 240585
rect 41878 240415 41930 240421
rect 41878 240357 41930 240363
rect 41890 239834 41918 240357
rect 41780 238382 41836 238391
rect 41780 238317 41836 238326
rect 41794 237984 41822 238317
rect 42754 236721 42782 247905
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42742 236715 42794 236721
rect 42742 236657 42794 236663
rect 42178 236165 42206 236657
rect 42850 236592 42878 248349
rect 42934 248111 42986 248117
rect 42934 248053 42986 248059
rect 42754 236564 42878 236592
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42166 234865 42218 234871
rect 42166 234807 42218 234813
rect 42178 234325 42206 234807
rect 42070 234051 42122 234057
rect 42070 233993 42122 233999
rect 42082 233692 42110 233993
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 42754 231097 42782 236564
rect 42838 236493 42890 236499
rect 42838 236435 42890 236441
rect 42850 234871 42878 236435
rect 42946 235463 42974 248053
rect 43030 247889 43082 247895
rect 43030 247831 43082 247837
rect 42934 235457 42986 235463
rect 42934 235399 42986 235405
rect 42838 234865 42890 234871
rect 42838 234807 42890 234813
rect 43042 234057 43070 247831
rect 43138 236499 43166 249237
rect 43126 236493 43178 236499
rect 43126 236435 43178 236441
rect 43030 234051 43082 234057
rect 43030 233993 43082 233999
rect 42070 231091 42122 231097
rect 42070 231033 42122 231039
rect 42742 231091 42794 231097
rect 42742 231033 42794 231039
rect 42082 230658 42110 231033
rect 41780 230390 41836 230399
rect 41780 230325 41836 230334
rect 41794 229992 41822 230325
rect 41780 229798 41836 229807
rect 41780 229733 41836 229742
rect 41794 229357 41822 229733
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 41876 227430 41932 227439
rect 41876 227365 41932 227374
rect 41890 226958 41918 227365
rect 41780 226838 41836 226847
rect 41780 226773 41836 226782
rect 41794 226321 41822 226773
rect 41972 226246 42028 226255
rect 41972 226181 42028 226190
rect 41986 225700 42014 226181
rect 41590 216513 41642 216519
rect 41588 216478 41590 216487
rect 41642 216478 41644 216487
rect 41588 216413 41644 216422
rect 41782 215773 41834 215779
rect 41780 215738 41782 215747
rect 41834 215738 41836 215747
rect 41780 215673 41836 215682
rect 41782 215255 41834 215261
rect 41780 215220 41782 215229
rect 41834 215220 41836 215229
rect 41780 215155 41836 215164
rect 41590 215033 41642 215039
rect 41588 214998 41590 215007
rect 41642 214998 41644 215007
rect 41588 214933 41644 214942
rect 41782 214293 41834 214299
rect 41780 214258 41782 214267
rect 41834 214258 41836 214267
rect 41780 214193 41836 214202
rect 41782 213701 41834 213707
rect 41780 213666 41782 213675
rect 41834 213666 41836 213675
rect 41780 213601 41836 213610
rect 43234 213337 43262 256859
rect 43330 255443 43358 296626
rect 43426 296626 43550 296654
rect 43426 256553 43454 296626
rect 43618 258033 43646 300593
rect 44194 278499 44222 385175
rect 44290 293849 44318 417513
rect 44386 302581 44414 599849
rect 44482 558959 44510 945799
rect 44468 558950 44524 558959
rect 44468 558885 44524 558894
rect 44470 547367 44522 547373
rect 44470 547309 44522 547315
rect 44374 302575 44426 302581
rect 44374 302517 44426 302523
rect 44278 293843 44330 293849
rect 44278 293785 44330 293791
rect 44180 278490 44236 278499
rect 44180 278425 44236 278434
rect 43606 258027 43658 258033
rect 43606 257969 43658 257975
rect 43510 257435 43562 257441
rect 43510 257377 43562 257383
rect 43414 256547 43466 256553
rect 43414 256489 43466 256495
rect 43414 255955 43466 255961
rect 43414 255897 43466 255903
rect 43426 255443 43454 255897
rect 43318 255437 43370 255443
rect 43318 255379 43370 255385
rect 43414 255437 43466 255443
rect 43414 255379 43466 255385
rect 41782 213331 41834 213337
rect 41780 213296 41782 213305
rect 43222 213331 43274 213337
rect 41834 213296 41836 213305
rect 43222 213273 43274 213279
rect 41780 213231 41836 213240
rect 41590 212961 41642 212967
rect 41588 212926 41590 212935
rect 41642 212926 41644 212935
rect 41588 212861 41644 212870
rect 43426 212227 43454 255379
rect 43522 215039 43550 257377
rect 44482 249153 44510 547309
rect 44470 249147 44522 249153
rect 44470 249089 44522 249095
rect 43510 215033 43562 215039
rect 43510 214975 43562 214981
rect 44578 212967 44606 987535
rect 44674 213707 44702 987609
rect 44854 987519 44906 987525
rect 44854 987461 44906 987467
rect 44758 987445 44810 987451
rect 44758 987387 44810 987393
rect 44770 255443 44798 987387
rect 44866 259217 44894 987461
rect 44950 987075 45002 987081
rect 44950 987017 45002 987023
rect 44962 299399 44990 987017
rect 45058 943643 45086 989237
rect 45142 987149 45194 987155
rect 45142 987091 45194 987097
rect 45046 943637 45098 943643
rect 45046 943579 45098 943585
rect 45046 932167 45098 932173
rect 45046 932109 45098 932115
rect 44950 299393 45002 299399
rect 44950 299335 45002 299341
rect 44950 285185 45002 285191
rect 44950 285127 45002 285133
rect 44854 259211 44906 259217
rect 44854 259153 44906 259159
rect 44758 255437 44810 255443
rect 44758 255379 44810 255385
rect 44854 242709 44906 242715
rect 44854 242651 44906 242657
rect 44758 242635 44810 242641
rect 44758 242577 44810 242583
rect 44662 213701 44714 213707
rect 44662 213643 44714 213649
rect 44566 212961 44618 212967
rect 44566 212903 44618 212909
rect 41782 212221 41834 212227
rect 41780 212186 41782 212195
rect 43414 212221 43466 212227
rect 41834 212186 41836 212195
rect 43414 212163 43466 212169
rect 41780 212121 41836 212130
rect 41972 209226 42028 209235
rect 41972 209161 42028 209170
rect 41986 207374 42014 209161
rect 41986 207346 42110 207374
rect 41588 207154 41644 207163
rect 41588 207089 41644 207098
rect 41602 205197 41630 207089
rect 41780 206784 41836 206793
rect 41780 206719 41836 206728
rect 41794 205937 41822 206719
rect 41876 206266 41932 206275
rect 41876 206201 41878 206210
rect 41930 206201 41932 206210
rect 41878 206169 41930 206175
rect 41782 205931 41834 205937
rect 41782 205873 41834 205879
rect 41780 205822 41836 205831
rect 41780 205757 41836 205766
rect 41590 205191 41642 205197
rect 41590 205133 41642 205139
rect 41588 205082 41644 205091
rect 41588 205017 41644 205026
rect 41602 204901 41630 205017
rect 41686 204969 41738 204975
rect 41684 204934 41686 204943
rect 41738 204934 41740 204943
rect 41590 204895 41642 204901
rect 41684 204869 41740 204878
rect 41590 204837 41642 204843
rect 41794 204605 41822 205757
rect 41782 204599 41834 204605
rect 41782 204541 41834 204547
rect 41782 204377 41834 204383
rect 41780 204342 41782 204351
rect 41834 204342 41836 204351
rect 41780 204277 41836 204286
rect 41782 203785 41834 203791
rect 41780 203750 41782 203759
rect 41834 203750 41836 203759
rect 41780 203685 41836 203694
rect 42082 197427 42110 207346
rect 42742 206227 42794 206233
rect 42742 206169 42794 206175
rect 42070 197421 42122 197427
rect 42070 197363 42122 197369
rect 42070 197199 42122 197205
rect 42070 197141 42122 197147
rect 42082 196618 42110 197141
rect 42754 196909 42782 206169
rect 43126 205931 43178 205937
rect 43126 205873 43178 205879
rect 42934 205191 42986 205197
rect 42934 205133 42986 205139
rect 42838 204895 42890 204901
rect 42838 204837 42890 204843
rect 42742 196903 42794 196909
rect 42742 196845 42794 196851
rect 41780 195166 41836 195175
rect 41780 195101 41836 195110
rect 41794 194805 41822 195101
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42850 192247 42878 204837
rect 42946 193505 42974 205133
rect 43030 204599 43082 204605
rect 43030 204541 43082 204547
rect 42934 193499 42986 193505
rect 42934 193441 42986 193447
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42838 192241 42890 192247
rect 42838 192183 42890 192189
rect 42178 191769 42206 192183
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42082 191142 42110 191443
rect 43042 191063 43070 204541
rect 43138 191507 43166 205873
rect 44770 204383 44798 242577
rect 44758 204377 44810 204383
rect 44758 204319 44810 204325
rect 44866 203791 44894 242651
rect 44962 215779 44990 285127
rect 45058 246267 45086 932109
rect 45154 300139 45182 987091
rect 45238 986779 45290 986785
rect 45238 986721 45290 986727
rect 45250 342393 45278 986721
rect 45334 986705 45386 986711
rect 45334 986647 45386 986653
rect 45346 343355 45374 986647
rect 62038 986483 62090 986489
rect 62038 986425 62090 986431
rect 61942 983671 61994 983677
rect 61942 983613 61994 983619
rect 61846 983597 61898 983603
rect 61846 983539 61898 983545
rect 60982 983079 61034 983085
rect 60982 983021 61034 983027
rect 57622 982931 57674 982937
rect 57622 982873 57674 982879
rect 48982 982857 49034 982863
rect 48982 982799 49034 982805
rect 48994 976407 49022 982799
rect 55414 979231 55466 979237
rect 55414 979173 55466 979179
rect 52054 977751 52106 977757
rect 52054 977693 52106 977699
rect 48898 976379 49022 976407
rect 48898 972059 48926 976379
rect 51958 974939 52010 974945
rect 51958 974881 52010 974887
rect 51862 973533 51914 973539
rect 51862 973475 51914 973481
rect 45622 972053 45674 972059
rect 45622 971995 45674 972001
rect 48886 972053 48938 972059
rect 48886 971995 48938 972001
rect 45526 967761 45578 967767
rect 45526 967703 45578 967709
rect 45430 806441 45482 806447
rect 45430 806383 45482 806389
rect 45334 343349 45386 343355
rect 45334 343291 45386 343297
rect 45238 342387 45290 342393
rect 45238 342329 45290 342335
rect 45238 311085 45290 311091
rect 45238 311027 45290 311033
rect 45142 300133 45194 300139
rect 45142 300075 45194 300081
rect 45142 296729 45194 296735
rect 45142 296671 45194 296677
rect 45046 246261 45098 246267
rect 45046 246203 45098 246209
rect 45046 242857 45098 242863
rect 45046 242799 45098 242805
rect 44950 215773 45002 215779
rect 44950 215715 45002 215721
rect 45058 204975 45086 242799
rect 45154 216519 45182 296671
rect 45142 216513 45194 216519
rect 45142 216455 45194 216461
rect 45250 215261 45278 311027
rect 45442 246489 45470 806383
rect 45538 784617 45566 967703
rect 45526 784611 45578 784617
rect 45526 784553 45578 784559
rect 45526 763299 45578 763305
rect 45526 763241 45578 763247
rect 45430 246483 45482 246489
rect 45430 246425 45482 246431
rect 45538 246341 45566 763241
rect 45634 741401 45662 971995
rect 48982 969241 49034 969247
rect 48982 969183 49034 969189
rect 46678 968501 46730 968507
rect 46678 968443 46730 968449
rect 46690 966139 46718 968443
rect 46678 966133 46730 966139
rect 46678 966075 46730 966081
rect 46006 965023 46058 965029
rect 46006 964965 46058 964971
rect 45718 964801 45770 964807
rect 45718 964743 45770 964749
rect 45730 784321 45758 964743
rect 45910 959103 45962 959109
rect 45910 959045 45962 959051
rect 45718 784315 45770 784321
rect 45718 784257 45770 784263
rect 45716 772958 45772 772967
rect 45716 772893 45772 772902
rect 45622 741395 45674 741401
rect 45622 741337 45674 741343
rect 45622 720231 45674 720237
rect 45622 720173 45674 720179
rect 45634 246415 45662 720173
rect 45730 316123 45758 772893
rect 45814 757453 45866 757459
rect 45814 757395 45866 757401
rect 45718 316117 45770 316123
rect 45718 316059 45770 316065
rect 45826 305319 45854 757395
rect 45922 685975 45950 959045
rect 46018 694707 46046 964965
rect 48994 964881 49022 969183
rect 50326 969167 50378 969173
rect 50326 969109 50378 969115
rect 48982 964875 49034 964881
rect 48982 964817 49034 964823
rect 47542 961989 47594 961995
rect 47542 961931 47594 961937
rect 47446 951925 47498 951931
rect 47446 951867 47498 951873
rect 46006 694701 46058 694707
rect 46006 694643 46058 694649
rect 45910 685969 45962 685975
rect 45910 685911 45962 685917
rect 45910 676941 45962 676947
rect 45910 676883 45962 676889
rect 45814 305313 45866 305319
rect 45814 305255 45866 305261
rect 45922 246637 45950 676883
rect 46006 633947 46058 633953
rect 46006 633889 46058 633895
rect 45910 246631 45962 246637
rect 45910 246573 45962 246579
rect 46018 246563 46046 633889
rect 47458 607651 47486 951867
rect 47554 943865 47582 961931
rect 50338 959109 50366 969109
rect 51874 967767 51902 973475
rect 51970 968507 51998 974881
rect 52066 970653 52094 977693
rect 52054 970647 52106 970653
rect 52054 970589 52106 970595
rect 51958 968501 52010 968507
rect 51958 968443 52010 968449
rect 51862 967761 51914 967767
rect 51862 967703 51914 967709
rect 55426 965029 55454 979173
rect 57634 976444 57662 982873
rect 58198 979305 58250 979311
rect 58198 979247 58250 979253
rect 57538 976416 57662 976444
rect 56278 973607 56330 973613
rect 56278 973549 56330 973555
rect 56086 973459 56138 973465
rect 56086 973401 56138 973407
rect 55414 965023 55466 965029
rect 55414 964965 55466 964971
rect 51862 964949 51914 964955
rect 51862 964891 51914 964897
rect 50326 959103 50378 959109
rect 50326 959045 50378 959051
rect 51874 956316 51902 964891
rect 56098 964881 56126 973401
rect 56290 964955 56318 973549
rect 57538 969247 57566 976416
rect 58210 973613 58238 979247
rect 60994 979237 61022 983021
rect 60982 979231 61034 979237
rect 60982 979173 61034 979179
rect 58870 976493 58922 976499
rect 58870 976435 58922 976441
rect 58198 973607 58250 973613
rect 58198 973549 58250 973555
rect 57526 969241 57578 969247
rect 57526 969183 57578 969189
rect 58882 969173 58910 976435
rect 58966 976419 59018 976425
rect 58966 976361 59018 976367
rect 58978 973539 59006 976361
rect 59540 976014 59596 976023
rect 59540 975949 59596 975958
rect 58966 973533 59018 973539
rect 58966 973475 59018 973481
rect 59554 970727 59582 975949
rect 59542 970721 59594 970727
rect 59542 970663 59594 970669
rect 58870 969167 58922 969173
rect 58870 969109 58922 969115
rect 56278 964949 56330 964955
rect 56278 964891 56330 964897
rect 52438 964875 52490 964881
rect 52438 964817 52490 964823
rect 56086 964875 56138 964881
rect 56086 964817 56138 964823
rect 51778 956288 51902 956316
rect 48982 953331 49034 953337
rect 48982 953273 49034 953279
rect 48994 945863 49022 953273
rect 51778 951931 51806 956288
rect 52450 953337 52478 964817
rect 59540 962990 59596 962999
rect 59540 962925 59596 962934
rect 59554 961995 59582 962925
rect 59542 961989 59594 961995
rect 59542 961931 59594 961937
rect 52438 953331 52490 953337
rect 52438 953273 52490 953279
rect 51766 951925 51818 951931
rect 51766 951867 51818 951873
rect 59540 949966 59596 949975
rect 59540 949901 59596 949910
rect 59554 947565 59582 949901
rect 59542 947559 59594 947565
rect 59542 947501 59594 947507
rect 48982 945857 49034 945863
rect 48982 945799 49034 945805
rect 47542 943859 47594 943865
rect 47542 943801 47594 943807
rect 59542 938901 59594 938907
rect 59542 938843 59594 938849
rect 59554 936951 59582 938843
rect 59540 936942 59596 936951
rect 59540 936877 59596 936886
rect 58580 923770 58636 923779
rect 58580 923705 58636 923714
rect 58594 921665 58622 923705
rect 58582 921659 58634 921665
rect 58582 921601 58634 921607
rect 59540 910746 59596 910755
rect 59540 910681 59596 910690
rect 59554 910121 59582 910681
rect 50422 910115 50474 910121
rect 50422 910057 50474 910063
rect 59542 910115 59594 910121
rect 59542 910057 59594 910063
rect 47638 895759 47690 895765
rect 47638 895701 47690 895707
rect 47542 869859 47594 869865
rect 47542 869801 47594 869807
rect 47554 757533 47582 869801
rect 47650 819323 47678 895701
rect 47638 819317 47690 819323
rect 47638 819259 47690 819265
rect 50434 818065 50462 910057
rect 59540 897870 59596 897879
rect 59540 897805 59596 897814
rect 59554 895765 59582 897805
rect 59542 895759 59594 895765
rect 59542 895701 59594 895707
rect 58004 884846 58060 884855
rect 58004 884781 58060 884790
rect 58018 884221 58046 884781
rect 53398 884215 53450 884221
rect 53398 884157 53450 884163
rect 58006 884215 58058 884221
rect 58006 884157 58058 884163
rect 53206 858315 53258 858321
rect 53206 858257 53258 858263
rect 50518 832415 50570 832421
rect 50518 832357 50570 832363
rect 50422 818059 50474 818065
rect 50422 818001 50474 818007
rect 50326 817985 50378 817991
rect 50326 817927 50378 817933
rect 47638 806515 47690 806521
rect 47638 806457 47690 806463
rect 47542 757527 47594 757533
rect 47542 757469 47594 757475
rect 47650 731855 47678 806457
rect 47830 792085 47882 792091
rect 47830 792027 47882 792033
rect 47734 751755 47786 751761
rect 47734 751697 47786 751703
rect 47638 731849 47690 731855
rect 47638 731791 47690 731797
rect 47542 714311 47594 714317
rect 47542 714253 47594 714259
rect 47554 627885 47582 714253
rect 47638 699881 47690 699887
rect 47638 699823 47690 699829
rect 47650 645423 47678 699823
rect 47746 688639 47774 751697
rect 47842 732891 47870 792027
rect 47926 740211 47978 740217
rect 47926 740153 47978 740159
rect 47830 732885 47882 732891
rect 47830 732827 47882 732833
rect 47938 689527 47966 740153
rect 50338 714391 50366 817927
rect 50530 775367 50558 832357
rect 50518 775361 50570 775367
rect 50518 775303 50570 775309
rect 53218 774849 53246 858257
rect 53302 843885 53354 843891
rect 53302 843827 53354 843833
rect 53314 776107 53342 843827
rect 53410 818583 53438 884157
rect 59540 871674 59596 871683
rect 59540 871609 59596 871618
rect 59554 869865 59582 871609
rect 59542 869859 59594 869865
rect 59542 869801 59594 869807
rect 58388 858650 58444 858659
rect 58388 858585 58444 858594
rect 58402 858321 58430 858585
rect 58390 858315 58442 858321
rect 58390 858257 58442 858263
rect 59540 845626 59596 845635
rect 59540 845561 59596 845570
rect 59554 843891 59582 845561
rect 59542 843885 59594 843891
rect 59542 843827 59594 843833
rect 59540 832602 59596 832611
rect 59540 832537 59596 832546
rect 59554 832421 59582 832537
rect 59542 832415 59594 832421
rect 59542 832357 59594 832363
rect 59540 819430 59596 819439
rect 59540 819365 59596 819374
rect 53398 818577 53450 818583
rect 53398 818519 53450 818525
rect 59554 817991 59582 819365
rect 59542 817985 59594 817991
rect 59542 817927 59594 817933
rect 59540 806554 59596 806563
rect 59540 806489 59542 806498
rect 59594 806489 59596 806498
rect 59542 806457 59594 806463
rect 59540 793530 59596 793539
rect 59540 793465 59596 793474
rect 59554 792091 59582 793465
rect 59542 792085 59594 792091
rect 59542 792027 59594 792033
rect 59540 780506 59596 780515
rect 59540 780441 59596 780450
rect 59554 777661 59582 780441
rect 53398 777655 53450 777661
rect 53398 777597 53450 777603
rect 59542 777655 59594 777661
rect 59542 777597 59594 777603
rect 53302 776101 53354 776107
rect 53302 776043 53354 776049
rect 53206 774843 53258 774849
rect 53206 774785 53258 774791
rect 53206 766111 53258 766117
rect 53206 766053 53258 766059
rect 50518 725855 50570 725861
rect 50518 725797 50570 725803
rect 50326 714385 50378 714391
rect 50326 714327 50378 714333
rect 47926 689521 47978 689527
rect 47926 689463 47978 689469
rect 50530 688935 50558 725797
rect 50518 688929 50570 688935
rect 50518 688871 50570 688877
rect 47734 688633 47786 688639
rect 47734 688575 47786 688581
rect 50422 688411 50474 688417
rect 50422 688353 50474 688359
rect 50326 662437 50378 662443
rect 50326 662379 50378 662385
rect 47638 645417 47690 645423
rect 47638 645359 47690 645365
rect 47734 636537 47786 636543
rect 47734 636479 47786 636485
rect 47542 627879 47594 627885
rect 47542 627821 47594 627827
rect 47542 622107 47594 622113
rect 47542 622049 47594 622055
rect 47444 607642 47500 607651
rect 47444 607577 47500 607586
rect 47554 602799 47582 622049
rect 47638 610637 47690 610643
rect 47638 610579 47690 610585
rect 47542 602793 47594 602799
rect 47542 602735 47594 602741
rect 47542 596207 47594 596213
rect 47542 596149 47594 596155
rect 47446 590731 47498 590737
rect 47446 590673 47498 590679
rect 47458 246711 47486 590673
rect 47554 285117 47582 596149
rect 47650 541527 47678 610579
rect 47746 603095 47774 636479
rect 47734 603089 47786 603095
rect 47734 603031 47786 603037
rect 50338 584743 50366 662379
rect 50434 646311 50462 688353
rect 53218 671101 53246 766053
rect 53410 732151 53438 777597
rect 59540 767482 59596 767491
rect 59540 767417 59596 767426
rect 59554 766117 59582 767417
rect 59542 766111 59594 766117
rect 59542 766053 59594 766059
rect 59540 754310 59596 754319
rect 59540 754245 59596 754254
rect 59554 751761 59582 754245
rect 59542 751755 59594 751761
rect 59542 751697 59594 751703
rect 58580 741286 58636 741295
rect 58580 741221 58636 741230
rect 58594 740217 58622 741221
rect 58582 740211 58634 740217
rect 58582 740153 58634 740159
rect 53398 732145 53450 732151
rect 53398 732087 53450 732093
rect 59156 728262 59212 728271
rect 59156 728197 59212 728206
rect 59170 725861 59198 728197
rect 59158 725855 59210 725861
rect 59158 725797 59210 725803
rect 59540 715386 59596 715395
rect 59540 715321 59596 715330
rect 59554 714317 59582 715321
rect 59542 714311 59594 714317
rect 59542 714253 59594 714259
rect 59540 702214 59596 702223
rect 59540 702149 59596 702158
rect 59554 699887 59582 702149
rect 59542 699881 59594 699887
rect 59542 699823 59594 699829
rect 59540 689190 59596 689199
rect 59540 689125 59596 689134
rect 59554 688417 59582 689125
rect 59542 688411 59594 688417
rect 59542 688353 59594 688359
rect 59060 676166 59116 676175
rect 59060 676101 59116 676110
rect 59074 673987 59102 676101
rect 53302 673981 53354 673987
rect 53302 673923 53354 673929
rect 59062 673981 59114 673987
rect 59062 673923 59114 673929
rect 53206 671095 53258 671101
rect 53206 671037 53258 671043
rect 53206 648081 53258 648087
rect 53206 648023 53258 648029
rect 50422 646305 50474 646311
rect 50422 646247 50474 646253
rect 53218 602207 53246 648023
rect 53314 645793 53342 673923
rect 58100 663142 58156 663151
rect 58100 663077 58156 663086
rect 58114 662443 58142 663077
rect 58102 662437 58154 662443
rect 58102 662379 58154 662385
rect 59540 650118 59596 650127
rect 59540 650053 59596 650062
rect 59554 648087 59582 650053
rect 59542 648081 59594 648087
rect 59542 648023 59594 648029
rect 53302 645787 53354 645793
rect 53302 645729 53354 645735
rect 59540 637094 59596 637103
rect 59540 637029 59596 637038
rect 59554 636543 59582 637029
rect 59542 636537 59594 636543
rect 59542 636479 59594 636485
rect 59540 624070 59596 624079
rect 59540 624005 59596 624014
rect 59554 622113 59582 624005
rect 59542 622107 59594 622113
rect 59542 622049 59594 622055
rect 59252 611046 59308 611055
rect 59252 610981 59308 610990
rect 59266 610643 59294 610981
rect 59254 610637 59306 610643
rect 59254 610579 59306 610585
rect 53206 602201 53258 602207
rect 53206 602143 53258 602149
rect 59348 598022 59404 598031
rect 59348 597957 59404 597966
rect 59362 596213 59390 597957
rect 53206 596207 53258 596213
rect 53206 596149 53258 596155
rect 59350 596207 59402 596213
rect 59350 596149 59402 596155
rect 50326 584737 50378 584743
rect 50326 584679 50378 584685
rect 50422 584737 50474 584743
rect 50422 584679 50474 584685
rect 50434 559879 50462 584679
rect 50422 559873 50474 559879
rect 50422 559815 50474 559821
rect 53218 558843 53246 596149
rect 59540 584850 59596 584859
rect 59540 584785 59596 584794
rect 59554 584743 59582 584785
rect 59542 584737 59594 584743
rect 59542 584679 59594 584685
rect 59540 571826 59596 571835
rect 59540 571761 59596 571770
rect 59554 570313 59582 571761
rect 59542 570307 59594 570313
rect 59542 570249 59594 570255
rect 53206 558837 53258 558843
rect 53206 558779 53258 558785
rect 59540 558802 59596 558811
rect 50326 558763 50378 558769
rect 59540 558737 59542 558746
rect 50326 558705 50378 558711
rect 59594 558737 59596 558746
rect 59542 558705 59594 558711
rect 47638 541521 47690 541527
rect 47638 541463 47690 541469
rect 47638 532863 47690 532869
rect 47638 532805 47690 532811
rect 47650 432303 47678 532805
rect 47830 518433 47882 518439
rect 47830 518375 47882 518381
rect 47734 504077 47786 504083
rect 47734 504019 47786 504025
rect 47638 432297 47690 432303
rect 47638 432239 47690 432245
rect 47638 419791 47690 419797
rect 47638 419733 47690 419739
rect 47542 285111 47594 285117
rect 47542 285053 47594 285059
rect 47650 249375 47678 419733
rect 47746 367405 47774 504019
rect 47842 431785 47870 518375
rect 48022 478177 48074 478183
rect 48022 478119 48074 478125
rect 47926 440733 47978 440739
rect 47926 440675 47978 440681
rect 47830 431779 47882 431785
rect 47830 431721 47882 431727
rect 47830 376575 47882 376581
rect 47830 376517 47882 376523
rect 47734 367399 47786 367405
rect 47734 367341 47786 367347
rect 47734 348529 47786 348535
rect 47734 348471 47786 348477
rect 47746 258403 47774 348471
rect 47734 258397 47786 258403
rect 47734 258339 47786 258345
rect 47638 249369 47690 249375
rect 47638 249311 47690 249317
rect 47842 249301 47870 376517
rect 47938 344835 47966 440675
rect 48034 389087 48062 478119
rect 50338 410547 50366 558705
rect 59540 545926 59596 545935
rect 59540 545861 59596 545870
rect 59554 544413 59582 545861
rect 53302 544407 53354 544413
rect 53302 544349 53354 544355
rect 59542 544407 59594 544413
rect 59542 544349 59594 544355
rect 50422 492533 50474 492539
rect 50422 492475 50474 492481
rect 50326 410541 50378 410547
rect 50326 410483 50378 410489
rect 50326 400403 50378 400409
rect 50326 400345 50378 400351
rect 48022 389081 48074 389087
rect 48022 389023 48074 389029
rect 48022 362959 48074 362965
rect 48022 362901 48074 362907
rect 47926 344829 47978 344835
rect 47926 344771 47978 344777
rect 47926 333359 47978 333365
rect 47926 333301 47978 333307
rect 47830 249295 47882 249301
rect 47830 249237 47882 249243
rect 47938 249227 47966 333301
rect 48034 302359 48062 362901
rect 49270 316117 49322 316123
rect 49270 316059 49322 316065
rect 49282 305245 49310 316059
rect 49270 305239 49322 305245
rect 49270 305181 49322 305187
rect 48022 302353 48074 302359
rect 48022 302295 48074 302301
rect 48022 290143 48074 290149
rect 48022 290085 48074 290091
rect 48034 249449 48062 290085
rect 50338 281121 50366 400345
rect 50434 388051 50462 492475
rect 53206 452203 53258 452209
rect 53206 452145 53258 452151
rect 50614 414759 50666 414765
rect 50614 414701 50666 414707
rect 50422 388045 50474 388051
rect 50422 387987 50474 387993
rect 50518 374429 50570 374435
rect 50518 374371 50570 374377
rect 50422 337059 50474 337065
rect 50422 337001 50474 337007
rect 50326 281115 50378 281121
rect 50326 281057 50378 281063
rect 50434 259735 50462 337001
rect 50530 302729 50558 374371
rect 50626 345575 50654 414701
rect 50614 345569 50666 345575
rect 50614 345511 50666 345517
rect 53218 324189 53246 452145
rect 53314 431415 53342 544349
rect 59540 532902 59596 532911
rect 59540 532837 59542 532846
rect 59594 532837 59596 532846
rect 59542 532805 59594 532811
rect 59540 519730 59596 519739
rect 59540 519665 59596 519674
rect 59554 518439 59582 519665
rect 59542 518433 59594 518439
rect 59542 518375 59594 518381
rect 59540 506706 59596 506715
rect 59540 506641 59596 506650
rect 59554 504083 59582 506641
rect 59542 504077 59594 504083
rect 59542 504019 59594 504025
rect 59540 493682 59596 493691
rect 59540 493617 59596 493626
rect 59554 492539 59582 493617
rect 59542 492533 59594 492539
rect 59542 492475 59594 492481
rect 59540 480658 59596 480667
rect 59540 480593 59596 480602
rect 59554 478183 59582 480593
rect 59542 478177 59594 478183
rect 59542 478119 59594 478125
rect 57812 467486 57868 467495
rect 57812 467421 57868 467430
rect 57826 466639 57854 467421
rect 53494 466633 53546 466639
rect 53494 466575 53546 466581
rect 57814 466633 57866 466639
rect 57814 466575 57866 466581
rect 53302 431409 53354 431415
rect 53302 431351 53354 431357
rect 53398 426303 53450 426309
rect 53398 426245 53450 426251
rect 53302 388859 53354 388865
rect 53302 388801 53354 388807
rect 53206 324183 53258 324189
rect 53206 324125 53258 324131
rect 53206 305239 53258 305245
rect 53206 305181 53258 305187
rect 50518 302723 50570 302729
rect 50518 302665 50570 302671
rect 53218 290963 53246 305181
rect 53314 301619 53342 388801
rect 53410 345945 53438 426245
rect 53506 388791 53534 466575
rect 59540 454610 59596 454619
rect 59540 454545 59596 454554
rect 59554 452209 59582 454545
rect 59542 452203 59594 452209
rect 59542 452145 59594 452151
rect 57812 441586 57868 441595
rect 57812 441521 57868 441530
rect 57826 440739 57854 441521
rect 57814 440733 57866 440739
rect 57814 440675 57866 440681
rect 59540 428562 59596 428571
rect 59540 428497 59596 428506
rect 59554 426309 59582 428497
rect 59542 426303 59594 426309
rect 59542 426245 59594 426251
rect 59540 415390 59596 415399
rect 59540 415325 59596 415334
rect 59554 414765 59582 415325
rect 59542 414759 59594 414765
rect 59542 414701 59594 414707
rect 59540 402366 59596 402375
rect 59540 402301 59596 402310
rect 59554 400409 59582 402301
rect 59542 400403 59594 400409
rect 59542 400345 59594 400351
rect 59540 389342 59596 389351
rect 59540 389277 59596 389286
rect 59554 388865 59582 389277
rect 59542 388859 59594 388865
rect 59542 388801 59594 388807
rect 53494 388785 53546 388791
rect 53494 388727 53546 388733
rect 61858 381613 61886 983539
rect 61954 384467 61982 983613
rect 62050 938981 62078 986425
rect 62134 986409 62186 986415
rect 62134 986351 62186 986357
rect 62146 941793 62174 986351
rect 73474 983534 73502 989311
rect 89602 983534 89630 989977
rect 92962 989375 92990 1005591
rect 94102 1005575 94154 1005581
rect 109940 1005549 109996 1005558
rect 110516 1005614 110572 1005623
rect 110516 1005549 110518 1005558
rect 94102 1005517 94154 1005523
rect 110570 1005549 110572 1005558
rect 110518 1005517 110570 1005523
rect 94114 990041 94142 1005517
rect 102070 1005501 102122 1005507
rect 102068 1005466 102070 1005475
rect 102122 1005466 102124 1005475
rect 102068 1005401 102124 1005410
rect 107062 1005353 107114 1005359
rect 107060 1005318 107062 1005327
rect 124630 1005353 124682 1005359
rect 107114 1005318 107116 1005327
rect 124630 1005295 124682 1005301
rect 107060 1005253 107116 1005262
rect 98038 1005205 98090 1005211
rect 94964 1005170 95020 1005179
rect 94964 1005105 95020 1005114
rect 97172 1005170 97228 1005179
rect 97940 1005170 97996 1005179
rect 97228 1005128 97940 1005156
rect 97172 1005105 97228 1005114
rect 105430 1005205 105482 1005211
rect 98038 1005147 98090 1005153
rect 105428 1005170 105430 1005179
rect 108022 1005205 108074 1005211
rect 105482 1005170 105484 1005179
rect 97940 1005105 97996 1005114
rect 94978 1002254 95006 1005105
rect 97846 1002467 97898 1002473
rect 97846 1002409 97898 1002415
rect 95062 1002393 95114 1002399
rect 95062 1002335 95114 1002341
rect 94882 1002226 95006 1002254
rect 94102 990035 94154 990041
rect 94102 989977 94154 989983
rect 92950 989369 93002 989375
rect 92950 989311 93002 989317
rect 94882 983529 94910 1002226
rect 95074 999735 95102 1002335
rect 95062 999729 95114 999735
rect 95062 999671 95114 999677
rect 94964 995846 95020 995855
rect 94964 995781 94966 995790
rect 95018 995781 95020 995790
rect 94966 995749 95018 995755
rect 94964 995698 95020 995707
rect 94964 995633 95020 995642
rect 94978 995591 95006 995633
rect 94966 995585 95018 995591
rect 94966 995527 95018 995533
rect 97858 993815 97886 1002409
rect 98050 999439 98078 1005147
rect 105428 1005105 105484 1005114
rect 108020 1005170 108022 1005179
rect 108074 1005170 108076 1005179
rect 108020 1005105 108076 1005114
rect 103028 1002506 103084 1002515
rect 103028 1002441 103030 1002450
rect 103082 1002441 103084 1002450
rect 103030 1002409 103082 1002415
rect 101494 1002393 101546 1002399
rect 101492 1002358 101494 1002367
rect 101546 1002358 101548 1002367
rect 100534 1002319 100586 1002325
rect 101492 1002293 101548 1002302
rect 103604 1002358 103660 1002367
rect 103604 1002293 103606 1002302
rect 100534 1002261 100586 1002267
rect 103658 1002293 103660 1002302
rect 103606 1002261 103658 1002267
rect 100546 999513 100574 1002261
rect 100534 999507 100586 999513
rect 100534 999449 100586 999455
rect 98038 999433 98090 999439
rect 98038 999375 98090 999381
rect 106006 997953 106058 997959
rect 106004 997918 106006 997927
rect 106058 997918 106060 997927
rect 106004 997853 106060 997862
rect 108500 996290 108556 996299
rect 108500 996225 108502 996234
rect 108554 996225 108556 996234
rect 112438 996251 112490 996257
rect 108502 996193 108554 996199
rect 112438 996193 112490 996199
rect 100532 996142 100588 996151
rect 100532 996077 100588 996086
rect 103988 996142 104044 996151
rect 103988 996077 104044 996086
rect 104468 996142 104524 996151
rect 104468 996077 104524 996086
rect 108596 996142 108652 996151
rect 108596 996077 108652 996086
rect 109556 996142 109612 996151
rect 109556 996077 109612 996086
rect 100546 995887 100574 996077
rect 103604 995994 103660 996003
rect 103604 995929 103660 995938
rect 100534 995881 100586 995887
rect 100534 995823 100586 995829
rect 97846 993809 97898 993815
rect 97846 993751 97898 993757
rect 103618 993741 103646 995929
rect 104002 994079 104030 996077
rect 103988 994070 104044 994079
rect 103988 994005 104044 994014
rect 104482 993783 104510 996077
rect 104468 993774 104524 993783
rect 103606 993735 103658 993741
rect 104468 993709 104524 993718
rect 103606 993677 103658 993683
rect 105814 990701 105866 990707
rect 105814 990643 105866 990649
rect 105826 983534 105854 990643
rect 108610 989301 108638 996077
rect 109570 990707 109598 996077
rect 112340 995846 112396 995855
rect 112340 995781 112396 995790
rect 110324 993922 110380 993931
rect 110324 993857 110380 993866
rect 109558 990701 109610 990707
rect 109558 990643 109610 990649
rect 110338 989449 110366 993857
rect 110326 989443 110378 989449
rect 110326 989385 110378 989391
rect 108598 989295 108650 989301
rect 108598 989237 108650 989243
rect 112354 986489 112382 995781
rect 112342 986483 112394 986489
rect 112342 986425 112394 986431
rect 112450 986415 112478 996193
rect 115222 996177 115274 996183
rect 115222 996119 115274 996125
rect 115234 996003 115262 996119
rect 124642 996035 124670 1005295
rect 126646 1005205 126698 1005211
rect 126646 1005147 126698 1005153
rect 126658 996109 126686 1005147
rect 143830 1004835 143882 1004841
rect 143830 1004777 143882 1004783
rect 143734 999433 143786 999439
rect 143734 999375 143786 999381
rect 126646 996103 126698 996109
rect 126646 996045 126698 996051
rect 124630 996029 124682 996035
rect 115220 995994 115276 996003
rect 124630 995971 124682 995977
rect 115220 995929 115276 995938
rect 133652 995846 133708 995855
rect 133440 995804 133652 995832
rect 137972 995846 138028 995855
rect 137760 995804 137972 995832
rect 133652 995781 133708 995790
rect 142656 995813 143006 995832
rect 143746 995813 143774 999375
rect 142656 995807 143018 995813
rect 142656 995804 142966 995807
rect 137972 995781 138028 995790
rect 142966 995749 143018 995755
rect 143734 995807 143786 995813
rect 143734 995749 143786 995755
rect 143842 995739 143870 1004777
rect 143926 1002319 143978 1002325
rect 143926 1002261 143978 1002267
rect 141046 995733 141098 995739
rect 137396 995698 137452 995707
rect 137136 995656 137396 995684
rect 138960 995665 139358 995684
rect 140784 995681 141046 995684
rect 140784 995675 141098 995681
rect 143830 995733 143882 995739
rect 143830 995675 143882 995681
rect 138960 995659 139370 995665
rect 138960 995656 139318 995659
rect 137396 995633 137452 995642
rect 140784 995656 141086 995675
rect 143938 995665 143966 1002261
rect 143926 995659 143978 995665
rect 139318 995601 139370 995607
rect 143926 995601 143978 995607
rect 136724 995550 136780 995559
rect 128482 993741 128510 995522
rect 129120 995508 129374 995536
rect 129346 993889 129374 995508
rect 129334 993883 129386 993889
rect 129334 993825 129386 993831
rect 129730 993783 129758 995522
rect 131616 995508 131870 995536
rect 132144 995508 132446 995536
rect 131842 993815 131870 995508
rect 132418 995411 132446 995508
rect 132404 995402 132460 995411
rect 132404 995337 132460 995346
rect 132802 994227 132830 995522
rect 135936 995508 136190 995536
rect 136464 995508 136724 995536
rect 132788 994218 132844 994227
rect 132788 994153 132844 994162
rect 136162 993931 136190 995508
rect 140160 995508 140414 995536
rect 136724 995485 136780 995494
rect 140386 995147 140414 995508
rect 140374 995141 140426 995147
rect 140374 995083 140426 995089
rect 136148 993922 136204 993931
rect 136148 993857 136204 993866
rect 131830 993809 131882 993815
rect 129716 993774 129772 993783
rect 128470 993735 128522 993741
rect 131830 993751 131882 993757
rect 129716 993709 129772 993718
rect 128470 993677 128522 993683
rect 138262 989739 138314 989745
rect 138262 989681 138314 989687
rect 122038 989443 122090 989449
rect 122038 989385 122090 989391
rect 112438 986409 112490 986415
rect 112438 986351 112490 986357
rect 122050 983534 122078 989385
rect 138274 983534 138302 989681
rect 146626 986563 146654 1007917
rect 158516 1005614 158572 1005623
rect 158516 1005549 158518 1005558
rect 158570 1005549 158572 1005558
rect 172918 1005575 172970 1005581
rect 158518 1005517 158570 1005523
rect 172918 1005517 172970 1005523
rect 151126 1005501 151178 1005507
rect 161398 1005501 161450 1005507
rect 151126 1005443 151178 1005449
rect 161396 1005466 161398 1005475
rect 161450 1005466 161452 1005475
rect 146902 996325 146954 996331
rect 146902 996267 146954 996273
rect 146806 996029 146858 996035
rect 146708 995994 146764 996003
rect 146806 995971 146858 995977
rect 146708 995929 146710 995938
rect 146762 995929 146764 995938
rect 146710 995897 146762 995903
rect 146710 995807 146762 995813
rect 146710 995749 146762 995755
rect 146722 995411 146750 995749
rect 146818 995707 146846 995971
rect 146804 995698 146860 995707
rect 146804 995633 146860 995642
rect 146708 995402 146764 995411
rect 146708 995337 146764 995346
rect 146914 993889 146942 996267
rect 149686 996251 149738 996257
rect 149686 996193 149738 996199
rect 149698 994227 149726 996193
rect 149684 994218 149740 994227
rect 149684 994153 149740 994162
rect 146902 993883 146954 993889
rect 146902 993825 146954 993831
rect 151138 989745 151166 1005443
rect 152662 1005427 152714 1005433
rect 161396 1005401 161452 1005410
rect 161876 1005466 161932 1005475
rect 161876 1005401 161878 1005410
rect 152662 1005369 152714 1005375
rect 161930 1005401 161932 1005410
rect 161878 1005369 161930 1005375
rect 151988 996142 152044 996151
rect 151988 996077 152044 996086
rect 152372 996142 152428 996151
rect 152372 996077 152428 996086
rect 152002 995961 152030 996077
rect 152386 996035 152414 996077
rect 152374 996029 152426 996035
rect 152374 995971 152426 995977
rect 151990 995955 152042 995961
rect 151990 995897 152042 995903
rect 151126 989739 151178 989745
rect 151126 989681 151178 989687
rect 152674 989227 152702 1005369
rect 159478 1005353 159530 1005359
rect 159476 1005318 159478 1005327
rect 172822 1005353 172874 1005359
rect 159530 1005318 159532 1005327
rect 159476 1005253 159532 1005262
rect 161492 1005318 161548 1005327
rect 172822 1005295 172874 1005301
rect 161492 1005253 161494 1005262
rect 161546 1005253 161548 1005262
rect 169942 1005279 169994 1005285
rect 161494 1005221 161546 1005227
rect 169942 1005221 169994 1005227
rect 160918 1005205 160970 1005211
rect 160916 1005170 160918 1005179
rect 166964 1005205 167016 1005211
rect 160970 1005170 160972 1005179
rect 160916 1005105 160972 1005114
rect 166962 1005153 166964 1005179
rect 167016 1005153 167018 1005179
rect 166962 1005105 167018 1005153
rect 156980 1004874 157036 1004883
rect 156980 1004809 156982 1004818
rect 157034 1004809 157036 1004818
rect 156982 1004777 157034 1004783
rect 153044 1002358 153100 1002367
rect 153044 1002293 153046 1002302
rect 153098 1002293 153100 1002302
rect 153046 1002261 153098 1002267
rect 154966 999433 155018 999439
rect 154964 999398 154966 999407
rect 155018 999398 155020 999407
rect 154964 999333 155020 999342
rect 154390 996325 154442 996331
rect 153428 996290 153484 996299
rect 153428 996225 153430 996234
rect 153482 996225 153484 996234
rect 154388 996290 154390 996299
rect 154442 996290 154444 996299
rect 154388 996225 154444 996234
rect 159956 996290 160012 996299
rect 159956 996225 159958 996234
rect 153430 996193 153482 996199
rect 160010 996225 160012 996234
rect 159958 996193 160010 996199
rect 166978 996183 167006 1005105
rect 166966 996177 167018 996183
rect 154004 996142 154060 996151
rect 154004 996077 154060 996086
rect 156500 996142 156556 996151
rect 156500 996077 156556 996086
rect 157364 996142 157420 996151
rect 157364 996077 157420 996086
rect 158900 996142 158956 996151
rect 166966 996119 167018 996125
rect 158900 996077 158902 996086
rect 154018 995813 154046 996077
rect 156212 995994 156268 996003
rect 156212 995929 156268 995938
rect 154006 995807 154058 995813
rect 154006 995749 154058 995755
rect 156226 993815 156254 995929
rect 156214 993809 156266 993815
rect 156214 993751 156266 993757
rect 156514 993741 156542 996077
rect 157378 993783 157406 996077
rect 158954 996077 158956 996086
rect 164278 996103 164330 996109
rect 158902 996045 158954 996051
rect 164278 996045 164330 996051
rect 158914 995887 158942 996045
rect 159668 995994 159724 996003
rect 159668 995929 159670 995938
rect 159722 995929 159724 995938
rect 164182 995955 164234 995961
rect 159670 995897 159722 995903
rect 164182 995897 164234 995903
rect 158902 995881 158954 995887
rect 158902 995823 158954 995829
rect 157364 993774 157420 993783
rect 156502 993735 156554 993741
rect 157364 993709 157420 993718
rect 156502 993677 156554 993683
rect 152662 989221 152714 989227
rect 152662 989163 152714 989169
rect 154486 989221 154538 989227
rect 154486 989163 154538 989169
rect 146614 986557 146666 986563
rect 146614 986499 146666 986505
rect 154498 983534 154526 989163
rect 164194 986637 164222 995897
rect 164182 986631 164234 986637
rect 164182 986573 164234 986579
rect 164290 983751 164318 996045
rect 164278 983745 164330 983751
rect 164278 983687 164330 983693
rect 169954 983548 169982 1005221
rect 172834 996109 172862 1005295
rect 172822 996103 172874 996109
rect 172822 996045 172874 996051
rect 172930 996035 172958 1005517
rect 197206 1005501 197258 1005507
rect 207382 1005501 207434 1005507
rect 197206 1005443 197258 1005449
rect 207380 1005466 207382 1005475
rect 207434 1005466 207436 1005475
rect 195190 1000839 195242 1000845
rect 195190 1000781 195242 1000787
rect 195094 999433 195146 999439
rect 195094 999375 195146 999381
rect 172918 996029 172970 996035
rect 172918 995971 172970 995977
rect 185108 995846 185164 995855
rect 184848 995804 185108 995832
rect 188544 995813 188894 995832
rect 189168 995813 189470 995832
rect 188544 995807 188906 995813
rect 188544 995804 188854 995807
rect 185108 995781 185164 995790
rect 189168 995807 189482 995813
rect 189168 995804 189430 995807
rect 188854 995749 188906 995755
rect 189430 995749 189482 995755
rect 195106 995739 195134 999375
rect 194422 995733 194474 995739
rect 184340 995698 184396 995707
rect 184176 995656 184340 995684
rect 190580 995698 190636 995707
rect 190368 995656 190580 995684
rect 184340 995633 184396 995642
rect 192192 995665 192542 995684
rect 194064 995681 194422 995684
rect 194064 995675 194474 995681
rect 195094 995733 195146 995739
rect 195094 995675 195146 995681
rect 192192 995659 192554 995665
rect 192192 995656 192502 995659
rect 190580 995633 190636 995642
rect 194064 995656 194462 995675
rect 195202 995665 195230 1000781
rect 195190 995659 195242 995665
rect 192502 995601 192554 995607
rect 195190 995601 195242 995607
rect 183284 995550 183340 995559
rect 179842 993815 179870 995522
rect 180514 993889 180542 995522
rect 181152 995508 181406 995536
rect 183024 995508 183284 995536
rect 180502 993883 180554 993889
rect 180502 993825 180554 993831
rect 179830 993809 179882 993815
rect 179830 993751 179882 993757
rect 181378 993741 181406 995508
rect 188084 995550 188140 995559
rect 183552 995517 183806 995536
rect 183552 995511 183818 995517
rect 183552 995508 183766 995511
rect 183284 995485 183340 995494
rect 183766 995453 183818 995459
rect 187330 995263 187358 995522
rect 187872 995508 188084 995536
rect 188084 995485 188140 995494
rect 187316 995254 187372 995263
rect 187316 995189 187372 995198
rect 186934 995067 186986 995073
rect 186934 995009 186986 995015
rect 181366 993735 181418 993741
rect 181366 993677 181418 993683
rect 94870 983523 94922 983529
rect 169954 983520 170736 983548
rect 186946 983534 186974 995009
rect 191554 993783 191582 995522
rect 197218 995115 197246 1005443
rect 207380 1005401 207436 1005410
rect 210838 1005353 210890 1005359
rect 210836 1005318 210838 1005327
rect 227350 1005353 227402 1005359
rect 210890 1005318 210892 1005327
rect 201622 1005279 201674 1005285
rect 210836 1005253 210892 1005262
rect 212852 1005318 212908 1005327
rect 227350 1005295 227402 1005301
rect 212852 1005253 212854 1005262
rect 201622 1005221 201674 1005227
rect 212906 1005253 212908 1005262
rect 212854 1005221 212906 1005227
rect 201526 996251 201578 996257
rect 201526 996193 201578 996199
rect 198644 995994 198700 996003
rect 198644 995929 198700 995938
rect 198742 995955 198794 995961
rect 197204 995106 197260 995115
rect 197204 995041 197260 995050
rect 191540 993774 191596 993783
rect 191540 993709 191596 993718
rect 198658 986859 198686 995929
rect 198742 995897 198794 995903
rect 198754 993889 198782 995897
rect 201538 995411 201566 996193
rect 201524 995402 201580 995411
rect 201524 995337 201580 995346
rect 198742 993883 198794 993889
rect 198742 993825 198794 993831
rect 201634 988857 201662 1005221
rect 209878 1005205 209930 1005211
rect 209876 1005170 209878 1005179
rect 225430 1005205 225482 1005211
rect 209930 1005170 209932 1005179
rect 225430 1005147 225482 1005153
rect 209876 1005105 209932 1005114
rect 208436 1000878 208492 1000887
rect 208436 1000813 208438 1000822
rect 208490 1000813 208492 1000822
rect 208438 1000781 208490 1000787
rect 206326 999433 206378 999439
rect 206324 999398 206326 999407
rect 206378 999398 206380 999407
rect 206324 999333 206380 999342
rect 204884 996290 204940 996299
rect 204884 996225 204886 996234
rect 204938 996225 204940 996234
rect 204886 996193 204938 996199
rect 211414 996177 211466 996183
rect 202292 996142 202348 996151
rect 202292 996077 202348 996086
rect 202868 996142 202924 996151
rect 202868 996077 202924 996086
rect 203924 996142 203980 996151
rect 203924 996077 203980 996086
rect 205268 996142 205324 996151
rect 205268 996077 205324 996086
rect 205940 996142 205996 996151
rect 205940 996077 205996 996086
rect 207860 996142 207916 996151
rect 207860 996077 207916 996086
rect 210836 996142 210892 996151
rect 210836 996077 210838 996086
rect 202306 995813 202334 996077
rect 202294 995807 202346 995813
rect 202294 995749 202346 995755
rect 202882 995559 202910 996077
rect 203938 995887 203966 996077
rect 203926 995881 203978 995887
rect 203926 995823 203978 995829
rect 202868 995550 202924 995559
rect 205282 995517 205310 996077
rect 205954 995961 205982 996077
rect 205942 995955 205994 995961
rect 205942 995897 205994 995903
rect 202868 995485 202924 995494
rect 205270 995511 205322 995517
rect 205270 995453 205322 995459
rect 207874 993815 207902 996077
rect 210890 996077 210892 996086
rect 211412 996142 211414 996151
rect 216022 996177 216074 996183
rect 211466 996142 211468 996151
rect 211412 996077 211468 996086
rect 212756 996142 212812 996151
rect 216022 996119 216074 996125
rect 219092 996142 219148 996151
rect 212756 996077 212758 996086
rect 210838 996045 210890 996051
rect 212810 996077 212812 996086
rect 212758 996045 212810 996051
rect 216034 996003 216062 996119
rect 216118 996103 216170 996109
rect 219092 996077 219148 996086
rect 216118 996045 216170 996051
rect 210164 995994 210220 996003
rect 210164 995929 210220 995938
rect 216020 995994 216076 996003
rect 216020 995929 216076 995938
rect 210178 995887 210206 995929
rect 210166 995881 210218 995887
rect 210166 995823 210218 995829
rect 213142 995881 213194 995887
rect 213142 995823 213194 995829
rect 209108 995550 209164 995559
rect 209108 995485 209164 995494
rect 207862 993809 207914 993815
rect 207862 993751 207914 993757
rect 209122 993741 209150 995485
rect 209110 993735 209162 993741
rect 209110 993677 209162 993683
rect 201622 988851 201674 988857
rect 201622 988793 201674 988799
rect 203158 988851 203210 988857
rect 203158 988793 203210 988799
rect 198646 986853 198698 986859
rect 198646 986795 198698 986801
rect 203170 983534 203198 988793
rect 213154 986933 213182 995823
rect 216130 989523 216158 996045
rect 216598 995955 216650 995961
rect 216598 995897 216650 995903
rect 216118 989517 216170 989523
rect 216118 989459 216170 989465
rect 216610 987007 216638 995897
rect 216598 987001 216650 987007
rect 216598 986943 216650 986949
rect 213142 986927 213194 986933
rect 213142 986869 213194 986875
rect 219106 983548 219134 996077
rect 225442 995961 225470 1005147
rect 227362 996109 227390 1005295
rect 246934 1002467 246986 1002473
rect 246934 1002409 246986 1002415
rect 246550 1002393 246602 1002399
rect 246550 1002335 246602 1002341
rect 246562 999532 246590 1002335
rect 246838 1002319 246890 1002325
rect 246838 1002261 246890 1002267
rect 246466 999504 246590 999532
rect 246646 999581 246698 999587
rect 246646 999523 246698 999529
rect 227350 996103 227402 996109
rect 227350 996045 227402 996051
rect 225430 995955 225482 995961
rect 225430 995897 225482 995903
rect 246466 995887 246494 999504
rect 246550 999433 246602 999439
rect 246550 999375 246602 999381
rect 246454 995881 246506 995887
rect 240212 995846 240268 995855
rect 239952 995804 240212 995832
rect 241844 995846 241900 995855
rect 240576 995813 240926 995832
rect 240576 995807 240938 995813
rect 240576 995804 240886 995807
rect 240212 995781 240268 995790
rect 241776 995804 241844 995832
rect 245424 995813 245726 995832
rect 246454 995823 246506 995829
rect 246562 995813 246590 999375
rect 245424 995807 245738 995813
rect 245424 995804 245686 995807
rect 241844 995781 241900 995790
rect 240886 995749 240938 995755
rect 245686 995749 245738 995755
rect 246550 995807 246602 995813
rect 246550 995749 246602 995755
rect 246658 995739 246686 999523
rect 246742 996547 246794 996553
rect 246742 996489 246794 996495
rect 243958 995733 244010 995739
rect 232148 995698 232204 995707
rect 231936 995656 232148 995684
rect 235584 995665 235838 995684
rect 243600 995681 243958 995684
rect 243600 995675 244010 995681
rect 246646 995733 246698 995739
rect 246646 995675 246698 995681
rect 235584 995659 235850 995665
rect 235584 995656 235798 995659
rect 232148 995633 232204 995642
rect 243600 995656 243998 995675
rect 246754 995665 246782 996489
rect 246742 995659 246794 995665
rect 235798 995601 235850 995607
rect 246742 995601 246794 995607
rect 236470 995585 236522 995591
rect 235220 995550 235276 995559
rect 231264 995508 231518 995536
rect 231490 994079 231518 995508
rect 231476 994070 231532 994079
rect 231476 994005 231532 994014
rect 232546 993741 232574 995522
rect 234370 994227 234398 995522
rect 234960 995508 235220 995536
rect 236256 995533 236470 995536
rect 236256 995527 236522 995533
rect 236256 995508 236510 995527
rect 235220 995485 235276 995494
rect 238690 994375 238718 995522
rect 239280 995517 239582 995536
rect 239280 995511 239594 995517
rect 239280 995508 239542 995511
rect 242976 995508 243230 995536
rect 246850 995517 246878 1002261
rect 246946 996003 246974 1002409
rect 247030 999507 247082 999513
rect 247030 999449 247082 999455
rect 246932 995994 246988 996003
rect 246932 995929 246988 995938
rect 247042 995559 247070 999449
rect 247028 995550 247084 995559
rect 239542 995453 239594 995459
rect 238676 994366 238732 994375
rect 238676 994301 238732 994310
rect 234356 994218 234412 994227
rect 234356 994153 234412 994162
rect 243202 993931 243230 995508
rect 246838 995511 246890 995517
rect 247028 995485 247084 995494
rect 246838 995453 246890 995459
rect 243188 993922 243244 993931
rect 243188 993857 243244 993866
rect 232534 993735 232586 993741
rect 232534 993677 232586 993683
rect 235606 989517 235658 989523
rect 235606 989459 235658 989465
rect 219106 983520 219408 983548
rect 235618 983534 235646 989459
rect 250498 989301 250526 1016205
rect 353410 1007991 353438 1016205
rect 351284 1007982 351340 1007991
rect 351284 1007917 351340 1007926
rect 353396 1007982 353452 1007991
rect 353396 1007917 353452 1007926
rect 261332 1006502 261388 1006511
rect 261332 1006437 261334 1006446
rect 261386 1006437 261388 1006446
rect 276598 1006463 276650 1006469
rect 261334 1006405 261386 1006411
rect 276598 1006405 276650 1006411
rect 262292 1005910 262348 1005919
rect 262292 1005845 262294 1005854
rect 262346 1005845 262348 1005854
rect 276502 1005871 276554 1005877
rect 262294 1005813 262346 1005819
rect 276502 1005813 276554 1005819
rect 255284 1002506 255340 1002515
rect 255284 1002441 255286 1002450
rect 255338 1002441 255340 1002450
rect 255286 1002409 255338 1002415
rect 253654 1002393 253706 1002399
rect 253652 1002358 253654 1002367
rect 253706 1002358 253708 1002367
rect 253652 1002293 253708 1002302
rect 254228 1002358 254284 1002367
rect 254228 1002293 254230 1002302
rect 254282 1002293 254284 1002302
rect 254230 1002261 254282 1002267
rect 259798 999581 259850 999587
rect 256628 999546 256684 999555
rect 256628 999481 256630 999490
rect 256682 999481 256684 999490
rect 259796 999546 259798 999555
rect 259850 999546 259852 999555
rect 259796 999481 259852 999490
rect 256630 999449 256682 999455
rect 257782 999433 257834 999439
rect 257780 999398 257782 999407
rect 257834 999398 257836 999407
rect 257780 999333 257836 999342
rect 256244 996586 256300 996595
rect 256244 996521 256246 996530
rect 256298 996521 256300 996530
rect 256246 996489 256298 996495
rect 276514 996183 276542 1005813
rect 262774 996177 262826 996183
rect 252308 996142 252364 996151
rect 252692 996142 252748 996151
rect 252364 996100 252692 996128
rect 252308 996077 252364 996086
rect 252692 996077 252748 996086
rect 254804 996142 254860 996151
rect 254804 996077 254860 996086
rect 258740 996142 258796 996151
rect 258740 996077 258796 996086
rect 260372 996142 260428 996151
rect 260372 996077 260428 996086
rect 262772 996142 262774 996151
rect 276502 996177 276554 996183
rect 262826 996142 262828 996151
rect 262772 996077 262828 996086
rect 263732 996142 263788 996151
rect 263732 996077 263734 996086
rect 254818 995591 254846 996077
rect 254806 995585 254858 995591
rect 254806 995527 254858 995533
rect 258754 994227 258782 996077
rect 258740 994218 258796 994227
rect 258740 994153 258796 994162
rect 251828 993774 251884 993783
rect 260386 993741 260414 996077
rect 263786 996077 263788 996086
rect 270740 996142 270796 996151
rect 276502 996119 276554 996125
rect 270740 996077 270796 996086
rect 263734 996045 263786 996051
rect 262486 996029 262538 996035
rect 261524 995994 261580 996003
rect 261524 995929 261526 995938
rect 261578 995929 261580 995938
rect 262484 995994 262486 996003
rect 268054 996029 268106 996035
rect 262538 995994 262540 996003
rect 267860 995994 267916 996003
rect 262484 995929 262540 995938
rect 265174 995955 265226 995961
rect 261526 995897 261578 995903
rect 268054 995971 268106 995977
rect 267860 995929 267916 995938
rect 265174 995897 265226 995903
rect 251828 993709 251884 993718
rect 260374 993735 260426 993741
rect 250486 989295 250538 989301
rect 250486 989237 250538 989243
rect 251842 983534 251870 993709
rect 260374 993677 260426 993683
rect 265186 989375 265214 995897
rect 265174 989369 265226 989375
rect 265174 989311 265226 989317
rect 267874 983548 267902 995929
rect 267956 995846 268012 995855
rect 267956 995781 268012 995790
rect 267970 989523 267998 995781
rect 267958 989517 268010 989523
rect 267958 989459 268010 989465
rect 268066 987229 268094 995971
rect 270754 989449 270782 996077
rect 276610 996035 276638 1006405
rect 316438 1005353 316490 1005359
rect 313844 1005318 313900 1005327
rect 313844 1005253 313846 1005262
rect 313898 1005253 313900 1005262
rect 316436 1005318 316438 1005327
rect 331222 1005353 331274 1005359
rect 316490 1005318 316492 1005327
rect 331222 1005295 331274 1005301
rect 316436 1005253 316492 1005262
rect 329686 1005279 329738 1005285
rect 313846 1005221 313898 1005227
rect 329686 1005221 329738 1005227
rect 298486 1005205 298538 1005211
rect 308278 1005205 308330 1005211
rect 298486 1005147 298538 1005153
rect 308276 1005170 308278 1005179
rect 312886 1005205 312938 1005211
rect 308330 1005170 308332 1005179
rect 298238 1000173 298290 1000179
rect 298238 1000115 298290 1000121
rect 298142 999581 298194 999587
rect 298058 999529 298142 999532
rect 298058 999523 298194 999529
rect 298058 999504 298182 999523
rect 276598 996029 276650 996035
rect 276598 995971 276650 995977
rect 286772 995846 286828 995855
rect 286560 995804 286772 995832
rect 291764 995846 291820 995855
rect 291504 995804 291764 995832
rect 286772 995781 286828 995790
rect 292176 995813 292574 995832
rect 297072 995813 297374 995832
rect 292176 995807 292586 995813
rect 292176 995804 292534 995807
rect 291764 995781 291820 995790
rect 297072 995807 297386 995813
rect 297072 995804 297334 995807
rect 292534 995749 292586 995755
rect 297334 995749 297386 995755
rect 298058 995739 298086 999504
rect 298142 999433 298194 999439
rect 298142 999375 298194 999381
rect 298154 995813 298182 999375
rect 298250 995887 298278 1000115
rect 298334 999507 298386 999513
rect 298334 999449 298386 999455
rect 298238 995881 298290 995887
rect 298238 995823 298290 995829
rect 298142 995807 298194 995813
rect 298142 995749 298194 995755
rect 295414 995733 295466 995739
rect 293588 995698 293644 995707
rect 290352 995665 290654 995684
rect 290352 995659 290666 995665
rect 290352 995656 290614 995659
rect 293376 995656 293588 995684
rect 295200 995681 295414 995684
rect 295200 995675 295466 995681
rect 298046 995733 298098 995739
rect 298046 995675 298098 995681
rect 295200 995656 295454 995675
rect 293588 995633 293644 995642
rect 290614 995601 290666 995607
rect 298346 995591 298374 999449
rect 298498 996003 298526 1005147
rect 308276 1005105 308332 1005114
rect 312884 1005170 312886 1005179
rect 312938 1005170 312940 1005179
rect 312884 1005105 312940 1005114
rect 299542 1002689 299594 1002695
rect 306742 1002689 306794 1002695
rect 299542 1002631 299594 1002637
rect 306740 1002654 306742 1002663
rect 306794 1002654 306796 1002663
rect 299446 996547 299498 996553
rect 299446 996489 299498 996495
rect 298484 995994 298540 996003
rect 298484 995929 298540 995938
rect 299458 995665 299486 996489
rect 299554 995855 299582 1002631
rect 299734 1002615 299786 1002621
rect 306740 1002589 306796 1002598
rect 307316 1002654 307372 1002663
rect 307316 1002589 307318 1002598
rect 299734 1002557 299786 1002563
rect 307370 1002589 307372 1002598
rect 307318 1002557 307370 1002563
rect 299638 1002467 299690 1002473
rect 299638 1002409 299690 1002415
rect 299650 1000179 299678 1002409
rect 299638 1000173 299690 1000179
rect 299638 1000115 299690 1000121
rect 299540 995846 299596 995855
rect 299540 995781 299596 995790
rect 299746 995707 299774 1002557
rect 300118 1002541 300170 1002547
rect 307894 1002541 307946 1002547
rect 300118 1002483 300170 1002489
rect 305300 1002506 305356 1002515
rect 300022 1002393 300074 1002399
rect 300022 1002335 300074 1002341
rect 299830 1002319 299882 1002325
rect 299830 1002261 299882 1002267
rect 299842 999513 299870 1002261
rect 299830 999507 299882 999513
rect 299830 999449 299882 999455
rect 299732 995698 299788 995707
rect 299446 995659 299498 995665
rect 299732 995633 299788 995642
rect 299446 995601 299498 995607
rect 291190 995585 291242 995591
rect 284372 995550 284428 995559
rect 282850 994079 282878 995522
rect 283522 994227 283550 995522
rect 284160 995508 284372 995536
rect 284372 995485 284428 995494
rect 286018 994523 286046 995522
rect 287184 995508 287486 995536
rect 287856 995517 287966 995536
rect 290880 995533 291190 995536
rect 290880 995527 291242 995533
rect 298334 995585 298386 995591
rect 298334 995527 298386 995533
rect 287856 995511 287978 995517
rect 287856 995508 287926 995511
rect 287458 995411 287486 995508
rect 290880 995508 291230 995527
rect 287926 995453 287978 995459
rect 287444 995402 287500 995411
rect 287444 995337 287500 995346
rect 286004 994514 286060 994523
rect 286004 994449 286060 994458
rect 283508 994218 283564 994227
rect 283508 994153 283564 994162
rect 282836 994070 282892 994079
rect 282836 994005 282892 994014
rect 294562 993783 294590 995522
rect 300034 995517 300062 1002335
rect 300022 995511 300074 995517
rect 300022 995453 300074 995459
rect 300130 995411 300158 1002483
rect 305300 1002441 305302 1002450
rect 305354 1002441 305356 1002450
rect 307892 1002506 307894 1002515
rect 307946 1002506 307948 1002515
rect 307892 1002441 307948 1002450
rect 305302 1002409 305354 1002415
rect 306358 1002393 306410 1002399
rect 305780 1002358 305836 1002367
rect 305780 1002293 305782 1002302
rect 305834 1002293 305836 1002302
rect 306356 1002358 306358 1002367
rect 306410 1002358 306412 1002367
rect 306356 1002293 306412 1002302
rect 305782 1002261 305834 1002267
rect 311446 999581 311498 999587
rect 311444 999546 311446 999555
rect 311498 999546 311500 999555
rect 311444 999481 311500 999490
rect 309334 999433 309386 999439
rect 309332 999398 309334 999407
rect 309386 999398 309388 999407
rect 309332 999333 309388 999342
rect 309812 996586 309868 996595
rect 309812 996521 309814 996530
rect 309866 996521 309868 996530
rect 309814 996489 309866 996495
rect 314230 996177 314282 996183
rect 304436 996142 304492 996151
rect 304916 996142 304972 996151
rect 304492 996100 304916 996128
rect 304436 996077 304492 996086
rect 304916 996077 304972 996086
rect 305300 996142 305356 996151
rect 305300 996077 305356 996086
rect 310868 996142 310924 996151
rect 314228 996142 314230 996151
rect 321622 996177 321674 996183
rect 314282 996142 314284 996151
rect 310868 996077 310924 996086
rect 313846 996103 313898 996109
rect 304820 995994 304876 996003
rect 304820 995929 304876 995938
rect 303380 995846 303436 995855
rect 303380 995781 303436 995790
rect 300116 995402 300172 995411
rect 300116 995337 300172 995346
rect 303394 994523 303422 995781
rect 303380 994514 303436 994523
rect 303380 994449 303436 994458
rect 304834 994227 304862 995929
rect 304820 994218 304876 994227
rect 304820 994153 304876 994162
rect 294548 993774 294604 993783
rect 294548 993709 294604 993718
rect 300502 989517 300554 989523
rect 300502 989459 300554 989465
rect 270742 989443 270794 989449
rect 270742 989385 270794 989391
rect 284278 989443 284330 989449
rect 284278 989385 284330 989391
rect 268054 987223 268106 987229
rect 268054 987165 268106 987171
rect 267874 983520 268080 983548
rect 284290 983534 284318 989385
rect 300514 983534 300542 989459
rect 305314 989449 305342 996077
rect 310882 994079 310910 996077
rect 314228 996077 314284 996086
rect 319604 996142 319660 996151
rect 321622 996119 321674 996125
rect 319604 996077 319660 996086
rect 313846 996045 313898 996051
rect 313078 996029 313130 996035
rect 313076 995994 313078 996003
rect 313858 996003 313886 996045
rect 317206 996029 317258 996035
rect 313130 995994 313132 996003
rect 313076 995929 313132 995938
rect 313844 995994 313900 996003
rect 317206 995971 317258 995977
rect 313844 995929 313900 995938
rect 310868 994070 310924 994079
rect 310868 994005 310924 994014
rect 316724 993922 316780 993931
rect 316724 993857 316780 993866
rect 305302 989443 305354 989449
rect 305302 989385 305354 989391
rect 316738 983534 316766 993857
rect 317218 987303 317246 995971
rect 319618 989523 319646 996077
rect 319700 995994 319756 996003
rect 319700 995929 319756 995938
rect 319714 989597 319742 995929
rect 319702 989591 319754 989597
rect 319702 989533 319754 989539
rect 319606 989517 319658 989523
rect 319606 989459 319658 989465
rect 321634 987377 321662 996119
rect 329698 987821 329726 1005221
rect 329782 1005205 329834 1005211
rect 329782 1005147 329834 1005153
rect 329686 987815 329738 987821
rect 329686 987757 329738 987763
rect 329794 987747 329822 1005147
rect 331234 992631 331262 1005295
rect 331222 992625 331274 992631
rect 331222 992567 331274 992573
rect 332566 992625 332618 992631
rect 332566 992567 332618 992573
rect 329782 987741 329834 987747
rect 329782 987683 329834 987689
rect 321622 987371 321674 987377
rect 321622 987313 321674 987319
rect 317206 987297 317258 987303
rect 317206 987239 317258 987245
rect 332578 983548 332606 992567
rect 351298 989523 351326 1007917
rect 356374 1006093 356426 1006099
rect 356372 1006058 356374 1006067
rect 371638 1006093 371690 1006099
rect 356426 1006058 356428 1006067
rect 356372 1005993 356428 1006002
rect 357908 1006058 357964 1006067
rect 558166 1006093 558218 1006099
rect 371638 1006035 371690 1006041
rect 558164 1006058 558166 1006067
rect 574678 1006093 574730 1006099
rect 558218 1006058 558220 1006067
rect 357908 1005993 357910 1006002
rect 357962 1005993 357964 1006002
rect 357910 1005961 357962 1005967
rect 358774 1005945 358826 1005951
rect 358772 1005910 358774 1005919
rect 358826 1005910 358828 1005919
rect 358772 1005845 358828 1005854
rect 359348 1005910 359404 1005919
rect 359348 1005845 359350 1005854
rect 359402 1005845 359404 1005854
rect 359350 1005813 359402 1005819
rect 361844 1005762 361900 1005771
rect 361844 1005697 361846 1005706
rect 361898 1005697 361900 1005706
rect 361846 1005665 361898 1005671
rect 358294 1005649 358346 1005655
rect 356756 1005614 356812 1005623
rect 356756 1005549 356758 1005558
rect 356810 1005549 356812 1005558
rect 357140 1005614 357196 1005623
rect 357140 1005549 357196 1005558
rect 358292 1005614 358294 1005623
rect 358346 1005614 358348 1005623
rect 358292 1005549 358348 1005558
rect 371542 1005575 371594 1005581
rect 356758 1005517 356810 1005523
rect 357154 1005507 357182 1005549
rect 371542 1005517 371594 1005523
rect 357142 1005501 357194 1005507
rect 357142 1005443 357194 1005449
rect 361268 1005466 361324 1005475
rect 361268 1005401 361270 1005410
rect 361322 1005401 361324 1005410
rect 361270 1005369 361322 1005375
rect 360886 1005353 360938 1005359
rect 360884 1005318 360886 1005327
rect 360938 1005318 360940 1005327
rect 360884 1005253 360940 1005262
rect 362324 1005318 362380 1005327
rect 362324 1005253 362326 1005262
rect 362378 1005253 362380 1005262
rect 362326 1005221 362378 1005227
rect 362806 1005205 362858 1005211
rect 362804 1005170 362806 1005179
rect 362858 1005170 362860 1005179
rect 362804 1005105 362860 1005114
rect 371554 1004989 371582 1005517
rect 371542 1004983 371594 1004989
rect 371542 1004925 371594 1004931
rect 371650 1004915 371678 1006035
rect 377302 1006019 377354 1006025
rect 574678 1006035 574730 1006041
rect 558164 1005993 558220 1006002
rect 377302 1005961 377354 1005967
rect 372022 1005501 372074 1005507
rect 372022 1005443 372074 1005449
rect 372034 1005063 372062 1005443
rect 374998 1005427 375050 1005433
rect 374998 1005369 375050 1005375
rect 374518 1005353 374570 1005359
rect 374518 1005295 374570 1005301
rect 374422 1005205 374474 1005211
rect 374422 1005147 374474 1005153
rect 372022 1005057 372074 1005063
rect 372022 1004999 372074 1005005
rect 371638 1004909 371690 1004915
rect 371638 1004851 371690 1004857
rect 374434 1000993 374462 1005147
rect 374422 1000987 374474 1000993
rect 374422 1000929 374474 1000935
rect 359732 1000878 359788 1000887
rect 359732 1000813 359734 1000822
rect 359786 1000813 359788 1000822
rect 359734 1000781 359786 1000787
rect 374422 996177 374474 996183
rect 363860 996142 363916 996151
rect 363860 996077 363916 996086
rect 366260 996142 366316 996151
rect 366260 996077 366316 996086
rect 366740 996142 366796 996151
rect 366740 996077 366742 996086
rect 360020 995698 360076 995707
rect 360020 995633 360076 995642
rect 362900 995698 362956 995707
rect 362900 995633 362956 995642
rect 363476 995698 363532 995707
rect 363476 995633 363532 995642
rect 360034 993741 360062 995633
rect 360022 993735 360074 993741
rect 360022 993677 360074 993683
rect 362914 993223 362942 995633
rect 362902 993217 362954 993223
rect 362902 993159 362954 993165
rect 349174 989517 349226 989523
rect 349174 989459 349226 989465
rect 351286 989517 351338 989523
rect 351286 989459 351338 989465
rect 332578 983520 332976 983548
rect 349186 983534 349214 989459
rect 362914 987451 362942 993159
rect 363490 987599 363518 995633
rect 363874 993149 363902 996077
rect 366274 996035 366302 996077
rect 366794 996077 366796 996086
rect 371540 996142 371596 996151
rect 374422 996119 374474 996125
rect 371540 996077 371596 996086
rect 371638 996103 371690 996109
rect 366742 996045 366794 996051
rect 366262 996029 366314 996035
rect 366262 995971 366314 995977
rect 364436 995698 364492 995707
rect 364436 995633 364492 995642
rect 363862 993143 363914 993149
rect 363862 993085 363914 993091
rect 363478 987593 363530 987599
rect 363478 987535 363530 987541
rect 363874 987525 363902 993085
rect 364450 987673 364478 995633
rect 371554 989671 371582 996077
rect 371638 996045 371690 996051
rect 371650 989745 371678 996045
rect 371734 996029 371786 996035
rect 374434 996003 374462 996119
rect 371734 995971 371786 995977
rect 374420 995994 374476 996003
rect 371638 989739 371690 989745
rect 371638 989681 371690 989687
rect 371542 989665 371594 989671
rect 371542 989607 371594 989613
rect 371746 989597 371774 995971
rect 374420 995929 374476 995938
rect 374530 993931 374558 1005295
rect 374614 1005279 374666 1005285
rect 374614 1005221 374666 1005227
rect 374516 993922 374572 993931
rect 374516 993857 374572 993866
rect 374626 993783 374654 1005221
rect 375010 1000919 375038 1005369
rect 374998 1000913 375050 1000919
rect 374998 1000855 375050 1000861
rect 377314 997145 377342 1005961
rect 378838 1005945 378890 1005951
rect 425686 1005945 425738 1005951
rect 378838 1005887 378890 1005893
rect 425684 1005910 425686 1005919
rect 471670 1005945 471722 1005951
rect 425738 1005910 425740 1005919
rect 377302 997139 377354 997145
rect 377302 997081 377354 997087
rect 378850 996553 378878 1005887
rect 380086 1005871 380138 1005877
rect 425684 1005845 425740 1005854
rect 429716 1005910 429772 1005919
rect 471670 1005887 471722 1005893
rect 551636 1005910 551692 1005919
rect 429716 1005845 429718 1005854
rect 380086 1005813 380138 1005819
rect 429770 1005845 429772 1005854
rect 466486 1005871 466538 1005877
rect 429718 1005813 429770 1005819
rect 466486 1005813 466538 1005819
rect 379990 1005649 380042 1005655
rect 379990 1005591 380042 1005597
rect 380002 1002254 380030 1005591
rect 380098 1005156 380126 1005813
rect 428278 1005797 428330 1005803
rect 428276 1005762 428278 1005771
rect 460822 1005797 460874 1005803
rect 428330 1005762 428332 1005771
rect 383638 1005723 383690 1005729
rect 428276 1005697 428332 1005706
rect 428660 1005762 428716 1005771
rect 460822 1005739 460874 1005745
rect 428660 1005697 428662 1005706
rect 383638 1005665 383690 1005671
rect 428714 1005697 428716 1005706
rect 428662 1005665 428714 1005671
rect 380098 1005128 380318 1005156
rect 380182 1005057 380234 1005063
rect 380182 1004999 380234 1005005
rect 380002 1002226 380126 1002254
rect 380098 996572 380126 1002226
rect 380194 999513 380222 1004999
rect 380182 999507 380234 999513
rect 380182 999449 380234 999455
rect 380290 999439 380318 1005128
rect 380374 1004983 380426 1004989
rect 380374 1004925 380426 1004931
rect 380278 999433 380330 999439
rect 380278 999375 380330 999381
rect 378838 996547 378890 996553
rect 380098 996544 380222 996572
rect 378838 996489 378890 996495
rect 380194 995707 380222 996544
rect 380180 995698 380236 995707
rect 380180 995633 380236 995642
rect 380386 995517 380414 1004925
rect 380470 1004909 380522 1004915
rect 380470 1004851 380522 1004857
rect 380374 995511 380426 995517
rect 380374 995453 380426 995459
rect 380482 995443 380510 1004851
rect 383446 1000987 383498 1000993
rect 383446 1000929 383498 1000935
rect 383350 1000913 383402 1000919
rect 383350 1000855 383402 1000861
rect 382870 999507 382922 999513
rect 382870 999449 382922 999455
rect 382678 997139 382730 997145
rect 382678 997081 382730 997087
rect 382690 996035 382718 997081
rect 382774 996547 382826 996553
rect 382774 996489 382826 996495
rect 382678 996029 382730 996035
rect 382678 995971 382730 995977
rect 382786 995855 382814 996489
rect 382772 995846 382828 995855
rect 382772 995781 382828 995790
rect 382882 995591 382910 999449
rect 382966 999433 383018 999439
rect 382966 999375 383018 999381
rect 382978 995961 383006 999375
rect 382966 995955 383018 995961
rect 382966 995897 383018 995903
rect 383362 995665 383390 1000855
rect 383458 995887 383486 1000929
rect 383542 1000839 383594 1000845
rect 383542 1000781 383594 1000787
rect 383446 995881 383498 995887
rect 383446 995823 383498 995829
rect 383554 995739 383582 1000781
rect 383650 995813 383678 1005665
rect 426742 1005649 426794 1005655
rect 425300 1005614 425356 1005623
rect 425300 1005549 425302 1005558
rect 425354 1005549 425356 1005558
rect 426740 1005614 426742 1005623
rect 426794 1005614 426796 1005623
rect 426740 1005549 426796 1005558
rect 425302 1005517 425354 1005523
rect 423766 1005501 423818 1005507
rect 423764 1005466 423766 1005475
rect 423818 1005466 423820 1005475
rect 423764 1005401 423820 1005410
rect 424724 1005466 424780 1005475
rect 424724 1005401 424726 1005410
rect 424778 1005401 424780 1005410
rect 424726 1005369 424778 1005375
rect 424150 1005353 424202 1005359
rect 424148 1005318 424150 1005327
rect 424202 1005318 424204 1005327
rect 424148 1005253 424204 1005262
rect 426164 1005318 426220 1005327
rect 426164 1005253 426166 1005262
rect 426218 1005253 426220 1005262
rect 426166 1005221 426218 1005227
rect 417524 1005170 417580 1005179
rect 417524 1005105 417580 1005114
rect 420788 1005170 420844 1005179
rect 421556 1005170 421612 1005179
rect 420844 1005128 421556 1005156
rect 420788 1005105 420844 1005114
rect 421556 1005105 421612 1005114
rect 399922 999433 399974 999439
rect 399922 999375 399974 999381
rect 399934 999219 399962 999375
rect 399874 999191 399962 999219
rect 388820 995846 388876 995855
rect 384418 995813 384672 995832
rect 383638 995807 383690 995813
rect 383638 995749 383690 995755
rect 384406 995807 384672 995813
rect 384458 995804 384672 995807
rect 385968 995813 386078 995832
rect 388066 995813 388368 995832
rect 385968 995807 386090 995813
rect 385968 995804 386038 995807
rect 384406 995749 384458 995755
rect 386038 995749 386090 995755
rect 388054 995807 388368 995813
rect 388106 995804 388368 995807
rect 388876 995804 388992 995832
rect 393058 995813 393312 995832
rect 393046 995807 393312 995813
rect 388820 995781 388876 995790
rect 388054 995749 388106 995755
rect 393098 995804 393312 995807
rect 396336 995813 396638 995832
rect 399874 995813 399902 999191
rect 396336 995807 396650 995813
rect 396336 995804 396598 995807
rect 393046 995749 393098 995755
rect 396598 995749 396650 995755
rect 399862 995807 399914 995813
rect 399862 995749 399914 995755
rect 383542 995733 383594 995739
rect 383542 995675 383594 995681
rect 384982 995733 385034 995739
rect 394868 995698 394924 995707
rect 385034 995681 385296 995684
rect 384982 995675 385296 995681
rect 383350 995659 383402 995665
rect 384994 995656 385296 995675
rect 387490 995665 387792 995684
rect 387478 995659 387792 995665
rect 383350 995601 383402 995607
rect 387530 995656 387792 995659
rect 394924 995656 395184 995684
rect 394868 995633 394924 995642
rect 387478 995601 387530 995607
rect 382870 995585 382922 995591
rect 382870 995527 382922 995533
rect 389398 995585 389450 995591
rect 389450 995533 389664 995536
rect 389398 995527 389664 995533
rect 389410 995508 389664 995527
rect 380470 995437 380522 995443
rect 380470 995379 380522 995385
rect 392098 993931 392126 995522
rect 392386 995517 392688 995536
rect 392374 995511 392688 995517
rect 392426 995508 392688 995511
rect 393730 995508 393984 995536
rect 392374 995453 392426 995459
rect 393730 995443 393758 995508
rect 393718 995437 393770 995443
rect 393718 995379 393770 995385
rect 392084 993922 392140 993931
rect 392084 993857 392140 993866
rect 396994 993783 397022 995522
rect 373940 993774 373996 993783
rect 373940 993709 373996 993718
rect 374612 993774 374668 993783
rect 374612 993709 374668 993718
rect 396980 993774 397036 993783
rect 398818 993741 398846 995522
rect 396980 993709 397036 993718
rect 398806 993735 398858 993741
rect 373954 990707 373982 993709
rect 398806 993677 398858 993683
rect 373942 990701 373994 990707
rect 373942 990643 373994 990649
rect 381622 990701 381674 990707
rect 381622 990643 381674 990649
rect 365398 989591 365450 989597
rect 365398 989533 365450 989539
rect 371734 989591 371786 989597
rect 371734 989533 371786 989539
rect 364438 987667 364490 987673
rect 364438 987609 364490 987615
rect 363862 987519 363914 987525
rect 363862 987461 363914 987467
rect 362902 987445 362954 987451
rect 362902 987387 362954 987393
rect 365410 983534 365438 989533
rect 381634 983534 381662 990643
rect 397846 989739 397898 989745
rect 397846 989681 397898 989687
rect 397858 983534 397886 989681
rect 414070 989665 414122 989671
rect 414070 989607 414122 989613
rect 414082 983534 414110 989607
rect 417538 987451 417566 1005105
rect 430196 1001026 430252 1001035
rect 430196 1000961 430198 1000970
rect 430250 1000961 430252 1000970
rect 430198 1000929 430250 1000935
rect 429238 1000913 429290 1000919
rect 427124 1000878 427180 1000887
rect 427124 1000813 427126 1000822
rect 427178 1000813 427180 1000822
rect 429236 1000878 429238 1000887
rect 429290 1000878 429292 1000887
rect 429236 1000813 429292 1000822
rect 427126 1000781 427178 1000787
rect 460834 999439 460862 1005739
rect 446518 999433 446570 999439
rect 446518 999375 446570 999381
rect 460822 999433 460874 999439
rect 460822 999375 460874 999381
rect 432790 996177 432842 996183
rect 430196 996142 430252 996151
rect 430196 996077 430252 996086
rect 431252 996142 431308 996151
rect 431252 996077 431308 996086
rect 432788 996142 432790 996151
rect 440662 996177 440714 996183
rect 432842 996142 432844 996151
rect 432788 996077 432844 996086
rect 433556 996142 433612 996151
rect 433556 996077 433612 996086
rect 434132 996142 434188 996151
rect 437972 996142 438028 996151
rect 434132 996077 434134 996086
rect 427412 995698 427468 995707
rect 427412 995633 427468 995642
rect 427426 993741 427454 995633
rect 427414 993735 427466 993741
rect 427414 993677 427466 993683
rect 430210 993001 430238 996077
rect 430868 995550 430924 995559
rect 430868 995485 430924 995494
rect 430882 993223 430910 995485
rect 430870 993217 430922 993223
rect 430870 993159 430922 993165
rect 431266 993075 431294 996077
rect 433570 996035 433598 996077
rect 434186 996077 434188 996086
rect 437782 996103 437834 996109
rect 434134 996045 434186 996051
rect 440662 996119 440714 996125
rect 437972 996077 438028 996086
rect 437782 996045 437834 996051
rect 433558 996029 433610 996035
rect 433558 995971 433610 995977
rect 431828 995550 431884 995559
rect 431828 995485 431884 995494
rect 431842 993149 431870 995485
rect 431830 993143 431882 993149
rect 431830 993085 431882 993091
rect 434902 993143 434954 993149
rect 434902 993085 434954 993091
rect 431254 993069 431306 993075
rect 431254 993011 431306 993017
rect 430198 992995 430250 993001
rect 430198 992937 430250 992943
rect 417526 987445 417578 987451
rect 417526 987387 417578 987393
rect 430210 987081 430238 992937
rect 430294 989591 430346 989597
rect 430294 989533 430346 989539
rect 430198 987075 430250 987081
rect 430198 987017 430250 987023
rect 430306 983534 430334 989533
rect 431266 987155 431294 993011
rect 434914 993001 434942 993085
rect 434902 992995 434954 993001
rect 434902 992937 434954 992943
rect 437794 989745 437822 996045
rect 437878 996029 437930 996035
rect 437878 995971 437930 995977
rect 437782 989739 437834 989745
rect 437782 989681 437834 989687
rect 437890 989597 437918 995971
rect 437986 989671 438014 996077
rect 440674 996003 440702 996119
rect 440660 995994 440716 996003
rect 440660 995929 440716 995938
rect 437974 989665 438026 989671
rect 437974 989607 438026 989613
rect 437878 989591 437930 989597
rect 437878 989533 437930 989539
rect 431254 987149 431306 987155
rect 431254 987091 431306 987097
rect 446530 983534 446558 999375
rect 466498 998052 466526 1005813
rect 469270 1005723 469322 1005729
rect 469270 1005665 469322 1005671
rect 469282 999513 469310 1005665
rect 469270 999507 469322 999513
rect 469270 999449 469322 999455
rect 469366 999433 469418 999439
rect 469366 999375 469418 999381
rect 466498 998024 466622 998052
rect 466594 993783 466622 998024
rect 469378 995443 469406 999375
rect 469366 995437 469418 995443
rect 469366 995379 469418 995385
rect 471682 993931 471710 1005887
rect 551636 1005845 551638 1005854
rect 551690 1005845 551692 1005854
rect 571606 1005871 571658 1005877
rect 551638 1005813 551690 1005819
rect 571606 1005813 571658 1005819
rect 502294 1005797 502346 1005803
rect 501716 1005762 501772 1005771
rect 501716 1005697 501718 1005706
rect 501770 1005697 501772 1005706
rect 502292 1005762 502294 1005771
rect 518518 1005797 518570 1005803
rect 502346 1005762 502348 1005771
rect 553654 1005797 553706 1005803
rect 518518 1005739 518570 1005745
rect 553652 1005762 553654 1005771
rect 571318 1005797 571370 1005803
rect 553706 1005762 553708 1005771
rect 502292 1005697 502348 1005706
rect 501718 1005665 501770 1005671
rect 472054 1005649 472106 1005655
rect 472054 1005591 472106 1005597
rect 502676 1005614 502732 1005623
rect 471862 1005575 471914 1005581
rect 471862 1005517 471914 1005523
rect 471766 1005501 471818 1005507
rect 471766 1005443 471818 1005449
rect 471778 995961 471806 1005443
rect 471874 996003 471902 1005517
rect 471958 1005353 472010 1005359
rect 471958 1005295 472010 1005301
rect 471860 995994 471916 996003
rect 471766 995955 471818 995961
rect 471860 995929 471916 995938
rect 471766 995897 471818 995903
rect 471970 995559 471998 1005295
rect 472066 995591 472094 1005591
rect 502676 1005549 502678 1005558
rect 502730 1005549 502732 1005558
rect 502678 1005517 502730 1005523
rect 500758 1005501 500810 1005507
rect 500756 1005466 500758 1005475
rect 509686 1005501 509738 1005507
rect 500810 1005466 500812 1005475
rect 472150 1005427 472202 1005433
rect 500756 1005401 500812 1005410
rect 503732 1005466 503788 1005475
rect 509686 1005443 509738 1005449
rect 518422 1005501 518474 1005507
rect 518422 1005443 518474 1005449
rect 503732 1005401 503734 1005410
rect 472150 1005369 472202 1005375
rect 503786 1005401 503788 1005410
rect 503734 1005369 503786 1005375
rect 472162 995855 472190 1005369
rect 505270 1005353 505322 1005359
rect 503252 1005318 503308 1005327
rect 472246 1005279 472298 1005285
rect 503252 1005253 503254 1005262
rect 472246 1005221 472298 1005227
rect 503306 1005253 503308 1005262
rect 505268 1005318 505270 1005327
rect 505322 1005318 505324 1005327
rect 505268 1005253 505324 1005262
rect 503254 1005221 503306 1005227
rect 472258 995887 472286 1005221
rect 501142 1005205 501194 1005211
rect 501140 1005170 501142 1005179
rect 506710 1005205 506762 1005211
rect 501194 1005170 501196 1005179
rect 501140 1005105 501196 1005114
rect 506708 1005170 506710 1005179
rect 506762 1005170 506764 1005179
rect 506708 1005105 506764 1005114
rect 505652 1002358 505708 1002367
rect 505652 1002293 505654 1002302
rect 505706 1002293 505708 1002302
rect 505654 1002261 505706 1002267
rect 509698 1002251 509726 1005443
rect 509782 1005131 509834 1005137
rect 509782 1005073 509834 1005079
rect 509686 1002245 509738 1002251
rect 509686 1002187 509738 1002193
rect 472642 1000993 472766 1001012
rect 472630 1000987 472766 1000993
rect 472682 1000984 472766 1000987
rect 472630 1000929 472682 1000935
rect 472534 1000913 472586 1000919
rect 472534 1000855 472586 1000861
rect 472438 999507 472490 999513
rect 472438 999449 472490 999455
rect 472246 995881 472298 995887
rect 472148 995846 472204 995855
rect 472246 995823 472298 995829
rect 472148 995781 472204 995790
rect 472054 995585 472106 995591
rect 471956 995550 472012 995559
rect 472054 995527 472106 995533
rect 472450 995517 472478 999449
rect 472546 995739 472574 1000855
rect 472630 1000839 472682 1000845
rect 472630 1000781 472682 1000787
rect 472642 995813 472670 1000781
rect 472630 995807 472682 995813
rect 472630 995749 472682 995755
rect 472534 995733 472586 995739
rect 472534 995675 472586 995681
rect 472738 995665 472766 1000984
rect 507188 1000878 507244 1000887
rect 507188 1000813 507190 1000822
rect 507242 1000813 507244 1000822
rect 507190 1000781 507242 1000787
rect 506228 1000730 506284 1000739
rect 506228 1000665 506230 1000674
rect 506282 1000665 506284 1000674
rect 506230 1000633 506282 1000639
rect 504212 999546 504268 999555
rect 504212 999481 504214 999490
rect 504266 999481 504268 999490
rect 504214 999449 504266 999455
rect 509794 999439 509822 1005073
rect 515830 1002245 515882 1002251
rect 515830 1002187 515882 1002193
rect 509782 999433 509834 999439
rect 509782 999375 509834 999381
rect 509782 996177 509834 996183
rect 499124 996142 499180 996151
rect 499124 996077 499180 996086
rect 509780 996142 509782 996151
rect 510742 996177 510794 996183
rect 509834 996142 509836 996151
rect 509780 996077 509836 996086
rect 510740 996142 510742 996151
rect 515734 996177 515786 996183
rect 510794 996142 510796 996151
rect 510740 996077 510796 996086
rect 511124 996142 511180 996151
rect 515540 996142 515596 996151
rect 511124 996077 511180 996086
rect 512662 996103 512714 996109
rect 499138 995855 499166 996077
rect 511138 996035 511166 996077
rect 515734 996119 515786 996125
rect 515540 996077 515596 996086
rect 512662 996045 512714 996051
rect 511126 996029 511178 996035
rect 507860 995994 507916 996003
rect 507860 995929 507916 995938
rect 508436 995994 508492 996003
rect 512674 996003 512702 996045
rect 511126 995971 511178 995977
rect 512660 995994 512716 996003
rect 508436 995929 508492 995938
rect 512660 995929 512716 995938
rect 478388 995846 478444 995855
rect 474082 995813 474336 995832
rect 477730 995813 477984 995832
rect 474070 995807 474336 995813
rect 474122 995804 474336 995807
rect 477718 995807 477984 995813
rect 474070 995749 474122 995755
rect 477770 995804 477984 995807
rect 482036 995846 482092 995855
rect 478444 995804 478656 995832
rect 478388 995781 478444 995790
rect 495284 995846 495340 995855
rect 482092 995804 482352 995832
rect 482722 995813 482976 995832
rect 482710 995807 482976 995813
rect 482036 995781 482092 995790
rect 477718 995749 477770 995755
rect 482762 995804 482976 995807
rect 495284 995781 495340 995790
rect 499124 995846 499180 995855
rect 499124 995781 499180 995790
rect 482710 995749 482762 995755
rect 473302 995733 473354 995739
rect 473354 995681 473664 995684
rect 473302 995675 473664 995681
rect 472726 995659 472778 995665
rect 473314 995656 473664 995675
rect 474658 995665 474960 995684
rect 474646 995659 474960 995665
rect 472726 995601 472778 995607
rect 474698 995656 474960 995659
rect 474646 995601 474698 995607
rect 476950 995585 477002 995591
rect 476386 995517 476784 995536
rect 480982 995585 481034 995591
rect 477002 995533 477360 995536
rect 476950 995527 477360 995533
rect 481364 995550 481420 995559
rect 481034 995533 481104 995536
rect 480982 995527 481104 995533
rect 471956 995485 472012 995494
rect 472438 995511 472490 995517
rect 472438 995453 472490 995459
rect 476374 995511 476784 995517
rect 476426 995508 476784 995511
rect 476962 995508 477360 995527
rect 480994 995508 481104 995527
rect 485588 995550 485644 995559
rect 481420 995508 481680 995536
rect 481364 995485 481420 995494
rect 476374 995453 476426 995459
rect 484162 993931 484190 995522
rect 485376 995508 485588 995536
rect 491828 995550 491884 995559
rect 485588 995485 485644 995494
rect 471668 993922 471724 993931
rect 471668 993857 471724 993866
rect 484148 993922 484204 993931
rect 484148 993857 484204 993866
rect 485986 993783 486014 995522
rect 466580 993774 466636 993783
rect 466580 993709 466636 993718
rect 485972 993774 486028 993783
rect 487810 993741 487838 995522
rect 491828 995485 491884 995494
rect 485972 993709 486028 993718
rect 487798 993735 487850 993741
rect 487798 993677 487850 993683
rect 462742 989739 462794 989745
rect 462742 989681 462794 989687
rect 462754 983534 462782 989681
rect 491842 989671 491870 995485
rect 478966 989665 479018 989671
rect 478966 989607 479018 989613
rect 491830 989665 491882 989671
rect 491830 989607 491882 989613
rect 478978 983534 479006 989607
rect 495190 989591 495242 989597
rect 495190 989533 495242 989539
rect 495202 983534 495230 989533
rect 495298 987081 495326 995781
rect 504404 995550 504460 995559
rect 504404 995485 504460 995494
rect 507284 995550 507340 995559
rect 507284 995485 507340 995494
rect 504418 993741 504446 995485
rect 504406 993735 504458 993741
rect 504406 993677 504458 993683
rect 507298 993001 507326 995485
rect 507874 993149 507902 995929
rect 507862 993143 507914 993149
rect 507862 993085 507914 993091
rect 507286 992995 507338 993001
rect 507286 992937 507338 992943
rect 495286 987075 495338 987081
rect 495286 987017 495338 987023
rect 507298 986785 507326 992937
rect 508450 992927 508478 995929
rect 508820 995550 508876 995559
rect 508820 995485 508876 995494
rect 508834 993075 508862 995485
rect 508822 993069 508874 993075
rect 508822 993011 508874 993017
rect 508438 992921 508490 992927
rect 508438 992863 508490 992869
rect 507286 986779 507338 986785
rect 507286 986721 507338 986727
rect 508450 986711 508478 992863
rect 515554 989671 515582 996077
rect 515638 996029 515690 996035
rect 515638 995971 515690 995977
rect 515650 989745 515678 995971
rect 515638 989739 515690 989745
rect 515638 989681 515690 989687
rect 511414 989665 511466 989671
rect 511414 989607 511466 989613
rect 515542 989665 515594 989671
rect 515542 989607 515594 989613
rect 508438 986705 508490 986711
rect 508438 986647 508490 986653
rect 511426 983534 511454 989607
rect 515746 989597 515774 996119
rect 515842 994037 515870 1002187
rect 517860 1000878 517916 1000887
rect 517860 1000813 517862 1000822
rect 517914 1000813 517916 1000822
rect 517862 1000781 517914 1000787
rect 518084 1000730 518140 1000739
rect 518084 1000665 518086 1000674
rect 518138 1000665 518140 1000674
rect 518086 1000633 518138 1000639
rect 518086 999507 518138 999513
rect 518086 999449 518138 999455
rect 517750 999433 517802 999439
rect 518098 999407 518126 999449
rect 517750 999375 517802 999381
rect 518084 999398 518140 999407
rect 517762 994185 517790 999375
rect 518084 999333 518140 999342
rect 518434 995411 518462 1005443
rect 518530 995559 518558 1005739
rect 523990 1005723 524042 1005729
rect 553652 1005697 553708 1005706
rect 554612 1005762 554668 1005771
rect 571318 1005739 571370 1005745
rect 554612 1005697 554614 1005706
rect 523990 1005665 524042 1005671
rect 554666 1005697 554668 1005706
rect 554614 1005665 554666 1005671
rect 520534 1005427 520586 1005433
rect 520534 1005369 520586 1005375
rect 520342 1005353 520394 1005359
rect 520342 1005295 520394 1005301
rect 520354 1002769 520382 1005295
rect 520342 1002763 520394 1002769
rect 520342 1002705 520394 1002711
rect 520546 999703 520574 1005369
rect 521302 1005279 521354 1005285
rect 521302 1005221 521354 1005227
rect 520532 999694 520588 999703
rect 520532 999629 520588 999638
rect 521314 999555 521342 1005221
rect 521494 1005131 521546 1005137
rect 521494 1005073 521546 1005079
rect 521398 1002319 521450 1002325
rect 521398 1002261 521450 1002267
rect 521300 999546 521356 999555
rect 521300 999481 521356 999490
rect 521410 995855 521438 1002261
rect 521506 996003 521534 1005073
rect 521590 1002763 521642 1002769
rect 521590 1002705 521642 1002711
rect 521492 995994 521548 996003
rect 521492 995929 521548 995938
rect 521396 995846 521452 995855
rect 521396 995781 521452 995790
rect 521602 995707 521630 1002705
rect 524002 1002254 524030 1005665
rect 554038 1005649 554090 1005655
rect 554036 1005614 554038 1005623
rect 554090 1005614 554092 1005623
rect 554036 1005549 554092 1005558
rect 555190 1005501 555242 1005507
rect 555188 1005466 555190 1005475
rect 555242 1005466 555244 1005475
rect 555188 1005401 555244 1005410
rect 552598 1005353 552650 1005359
rect 552212 1005318 552268 1005327
rect 552212 1005253 552214 1005262
rect 552266 1005253 552268 1005262
rect 552596 1005318 552598 1005327
rect 561526 1005353 561578 1005359
rect 552650 1005318 552652 1005327
rect 561526 1005295 561578 1005301
rect 552596 1005253 552652 1005262
rect 561046 1005279 561098 1005285
rect 552214 1005221 552266 1005227
rect 561046 1005221 561098 1005227
rect 552982 1005205 553034 1005211
rect 552980 1005170 552982 1005179
rect 553034 1005170 553036 1005179
rect 552980 1005105 553036 1005114
rect 561058 1002399 561086 1005221
rect 561046 1002393 561098 1002399
rect 558548 1002358 558604 1002367
rect 561046 1002335 561098 1002341
rect 561538 1002344 561566 1005295
rect 564310 1005131 564362 1005137
rect 564310 1005073 564362 1005079
rect 561538 1002316 561662 1002344
rect 558548 1002293 558550 1002302
rect 558602 1002293 558604 1002302
rect 558550 1002261 558602 1002267
rect 523810 1002226 524030 1002254
rect 523604 999694 523660 999703
rect 523604 999629 523660 999638
rect 521588 995698 521644 995707
rect 521588 995633 521644 995642
rect 523618 995591 523646 999629
rect 523700 999546 523756 999555
rect 523700 999481 523756 999490
rect 523714 995961 523742 999481
rect 523702 995955 523754 995961
rect 523702 995897 523754 995903
rect 523810 995665 523838 1002226
rect 523892 1000878 523948 1000887
rect 523892 1000813 523948 1000822
rect 523906 995887 523934 1000813
rect 523988 1000730 524044 1000739
rect 523988 1000665 524044 1000674
rect 523894 995881 523946 995887
rect 523894 995823 523946 995829
rect 524002 995739 524030 1000665
rect 540310 999581 540362 999587
rect 540310 999523 540362 999529
rect 524084 999398 524140 999407
rect 524084 999333 524140 999342
rect 524098 995813 524126 999333
rect 527924 995846 527980 995855
rect 525346 995813 525744 995832
rect 526114 995813 526368 995832
rect 524086 995807 524138 995813
rect 524086 995749 524138 995755
rect 525334 995807 525744 995813
rect 525386 995804 525744 995807
rect 526102 995807 526368 995813
rect 525334 995749 525386 995755
rect 526154 995804 526368 995807
rect 537236 995846 537292 995855
rect 527980 995804 528192 995832
rect 529090 995813 529392 995832
rect 529078 995807 529392 995813
rect 527924 995781 527980 995790
rect 526102 995749 526154 995755
rect 529130 995804 529392 995807
rect 536784 995813 537182 995832
rect 536784 995807 537194 995813
rect 536784 995804 537142 995807
rect 529078 995749 529130 995755
rect 537292 995804 537408 995832
rect 540322 995813 540350 999523
rect 561634 999513 561662 1002316
rect 561622 999507 561674 999513
rect 561622 999449 561674 999455
rect 564322 999439 564350 1005073
rect 564406 1002393 564458 1002399
rect 564406 1002335 564458 1002341
rect 564310 999433 564362 999439
rect 564310 999375 564362 999381
rect 564418 999384 564446 1002335
rect 567382 1002319 567434 1002325
rect 567382 1002261 567434 1002267
rect 564418 999356 564542 999384
rect 564514 998181 564542 999356
rect 564502 998175 564554 998181
rect 564502 998117 564554 998123
rect 567394 997737 567422 1002261
rect 567382 997731 567434 997737
rect 567382 997673 567434 997679
rect 555574 997657 555626 997663
rect 555572 997622 555574 997631
rect 555626 997622 555628 997631
rect 555572 997557 555628 997566
rect 557590 997509 557642 997515
rect 557588 997474 557590 997483
rect 557642 997474 557644 997483
rect 557588 997409 557644 997418
rect 555956 996142 556012 996151
rect 555956 996077 556012 996086
rect 559124 996142 559180 996151
rect 559124 996077 559180 996086
rect 561140 996142 561196 996151
rect 561140 996077 561142 996086
rect 540310 995807 540362 995813
rect 537236 995781 537292 995790
rect 537142 995749 537194 995755
rect 540310 995749 540362 995755
rect 523990 995733 524042 995739
rect 523990 995675 524042 995681
rect 524758 995733 524810 995739
rect 532244 995698 532300 995707
rect 524810 995681 525072 995684
rect 524758 995675 525072 995681
rect 523798 995659 523850 995665
rect 524770 995656 525072 995675
rect 529762 995665 530064 995684
rect 529750 995659 530064 995665
rect 523798 995601 523850 995607
rect 529802 995656 530064 995659
rect 532300 995656 532512 995684
rect 532244 995633 532300 995642
rect 529750 995601 529802 995607
rect 523606 995585 523658 995591
rect 518516 995550 518572 995559
rect 523606 995527 523658 995533
rect 528406 995585 528458 995591
rect 533396 995550 533452 995559
rect 528458 995533 528768 995536
rect 528406 995527 528768 995533
rect 528418 995508 528768 995527
rect 532834 995508 533088 995536
rect 518516 995485 518572 995494
rect 518420 995402 518476 995411
rect 518420 995337 518476 995346
rect 532834 994185 532862 995508
rect 533452 995508 533712 995536
rect 533396 995485 533452 995494
rect 517750 994179 517802 994185
rect 517750 994121 517802 994127
rect 532822 994179 532874 994185
rect 532822 994121 532874 994127
rect 534370 994037 534398 995522
rect 535330 995508 535584 995536
rect 538978 995508 539232 995536
rect 535330 995411 535358 995508
rect 535316 995402 535372 995411
rect 535316 995337 535372 995346
rect 515830 994031 515882 994037
rect 515830 993973 515882 993979
rect 534358 994031 534410 994037
rect 534358 993973 534410 993979
rect 538978 993741 539006 995508
rect 555970 993741 555998 996077
rect 538966 993735 539018 993741
rect 538966 993677 539018 993683
rect 555958 993735 556010 993741
rect 555958 993677 556010 993683
rect 559138 993149 559166 996077
rect 561194 996077 561196 996086
rect 561908 996142 561964 996151
rect 561908 996077 561910 996086
rect 561142 996045 561194 996051
rect 561962 996077 561964 996086
rect 569876 996142 569932 996151
rect 569876 996077 569932 996086
rect 569974 996103 570026 996109
rect 561910 996045 561962 996051
rect 560180 995994 560236 996003
rect 560180 995929 560236 995938
rect 569780 995994 569836 996003
rect 569780 995929 569836 995938
rect 559126 993143 559178 993149
rect 559126 993085 559178 993091
rect 560194 993075 560222 995929
rect 567188 995846 567244 995855
rect 567188 995781 567244 995790
rect 565844 995698 565900 995707
rect 565844 995633 565900 995642
rect 561620 995254 561676 995263
rect 561620 995189 561676 995198
rect 561634 993815 561662 995189
rect 561622 993809 561674 993815
rect 561622 993751 561674 993757
rect 560182 993069 560234 993075
rect 560182 993011 560234 993017
rect 527638 989739 527690 989745
rect 527638 989681 527690 989687
rect 515734 989591 515786 989597
rect 515734 989533 515786 989539
rect 527650 983534 527678 989681
rect 543766 989665 543818 989671
rect 543766 989607 543818 989613
rect 543778 983534 543806 989607
rect 560086 989591 560138 989597
rect 560086 989533 560138 989539
rect 560098 983534 560126 989533
rect 565462 985077 565514 985083
rect 565462 985019 565514 985025
rect 565474 983603 565502 985019
rect 565858 985009 565886 995633
rect 566036 995550 566092 995559
rect 566036 995485 566092 995494
rect 566050 985083 566078 995485
rect 567202 989597 567230 995781
rect 567380 995402 567436 995411
rect 567380 995337 567436 995346
rect 567394 994079 567422 995337
rect 567380 994070 567436 994079
rect 567380 994005 567436 994014
rect 569794 989819 569822 995929
rect 569782 989813 569834 989819
rect 569782 989755 569834 989761
rect 569890 989745 569918 996077
rect 569974 996045 570026 996051
rect 569878 989739 569930 989745
rect 569878 989681 569930 989687
rect 569986 989671 570014 996045
rect 571330 993963 571358 1005739
rect 571318 993957 571370 993963
rect 571318 993899 571370 993905
rect 569974 989665 570026 989671
rect 569974 989607 570026 989613
rect 567190 989591 567242 989597
rect 567190 989533 567242 989539
rect 571618 986711 571646 1005813
rect 573046 1005723 573098 1005729
rect 573046 1005665 573098 1005671
rect 572950 1005649 573002 1005655
rect 572950 1005591 573002 1005597
rect 571990 1005501 572042 1005507
rect 571990 1005443 572042 1005449
rect 572002 997589 572030 1005443
rect 572854 999581 572906 999587
rect 572854 999523 572906 999529
rect 571990 997583 572042 997589
rect 571990 997525 572042 997531
rect 572866 996553 572894 999523
rect 572854 996547 572906 996553
rect 572854 996489 572906 996495
rect 572962 993783 572990 1005591
rect 573058 994375 573086 1005665
rect 573142 999359 573194 999365
rect 573142 999301 573194 999307
rect 573154 994523 573182 999301
rect 573238 998175 573290 998181
rect 573238 998117 573290 998123
rect 573140 994514 573196 994523
rect 573140 994449 573196 994458
rect 573044 994366 573100 994375
rect 573044 994301 573100 994310
rect 573250 994227 573278 998117
rect 573236 994218 573292 994227
rect 573236 994153 573292 994162
rect 574690 993931 574718 1006035
rect 590710 999729 590762 999735
rect 590710 999671 590762 999677
rect 625558 999729 625610 999735
rect 625558 999671 625610 999677
rect 590614 999581 590666 999587
rect 590614 999523 590666 999529
rect 574870 999507 574922 999513
rect 574870 999449 574922 999455
rect 590518 999507 590570 999513
rect 590518 999449 590570 999455
rect 574882 997441 574910 999449
rect 590530 997737 590558 999449
rect 590518 997731 590570 997737
rect 590518 997673 590570 997679
rect 590626 997515 590654 999523
rect 590614 997509 590666 997515
rect 590614 997451 590666 997457
rect 590722 997441 590750 999671
rect 609046 999655 609098 999661
rect 609046 999597 609098 999603
rect 609058 997589 609086 999597
rect 609046 997583 609098 997589
rect 609046 997525 609098 997531
rect 574870 997435 574922 997441
rect 574870 997377 574922 997383
rect 590710 997435 590762 997441
rect 590710 997377 590762 997383
rect 576310 996547 576362 996553
rect 576310 996489 576362 996495
rect 574676 993922 574732 993931
rect 574676 993857 574732 993866
rect 572948 993774 573004 993783
rect 572948 993709 573004 993718
rect 571606 986705 571658 986711
rect 571606 986647 571658 986653
rect 566038 985077 566090 985083
rect 566038 985019 566090 985025
rect 565846 985003 565898 985009
rect 565846 984945 565898 984951
rect 566326 985003 566378 985009
rect 566326 984945 566378 984951
rect 566338 983677 566366 984945
rect 566326 983671 566378 983677
rect 566326 983613 566378 983619
rect 565462 983597 565514 983603
rect 565462 983539 565514 983545
rect 576322 983534 576350 996489
rect 625570 995961 625598 999671
rect 625846 999655 625898 999661
rect 625846 999597 625898 999603
rect 625750 999581 625802 999587
rect 625750 999523 625802 999529
rect 625654 999507 625706 999513
rect 625654 999449 625706 999455
rect 625558 995955 625610 995961
rect 625558 995897 625610 995903
rect 625666 995887 625694 999449
rect 625654 995881 625706 995887
rect 625654 995823 625706 995829
rect 625762 995739 625790 999523
rect 625858 997756 625886 999597
rect 625858 997728 625982 997756
rect 625846 997657 625898 997663
rect 625846 997599 625898 997605
rect 625858 995813 625886 997599
rect 625846 995807 625898 995813
rect 625846 995749 625898 995755
rect 625750 995733 625802 995739
rect 625750 995675 625802 995681
rect 625954 995665 625982 997728
rect 627106 995813 627504 995832
rect 627874 995813 628176 995832
rect 634594 995813 634896 995832
rect 627094 995807 627504 995813
rect 627146 995804 627504 995807
rect 627862 995807 628176 995813
rect 627094 995749 627146 995755
rect 627914 995804 628176 995807
rect 634582 995807 634896 995813
rect 627862 995749 627914 995755
rect 634634 995804 634896 995807
rect 634582 995749 634634 995755
rect 626518 995733 626570 995739
rect 626570 995681 626880 995684
rect 626518 995675 626880 995681
rect 625942 995659 625994 995665
rect 626530 995656 626880 995675
rect 630178 995665 630576 995684
rect 630166 995659 630576 995665
rect 625942 995601 625994 995607
rect 630218 995656 630576 995659
rect 630166 995601 630218 995607
rect 629986 994079 630014 995522
rect 630946 995508 631200 995536
rect 630946 994375 630974 995508
rect 631810 994523 631838 995522
rect 631796 994514 631852 994523
rect 631796 994449 631852 994458
rect 630932 994366 630988 994375
rect 630932 994301 630988 994310
rect 629972 994070 630028 994079
rect 629972 994005 630028 994014
rect 634306 993815 634334 995522
rect 635266 995508 635520 995536
rect 635266 993963 635294 995508
rect 636130 994227 636158 995522
rect 636116 994218 636172 994227
rect 636116 994153 636172 994162
rect 635254 993957 635306 993963
rect 635254 993899 635306 993905
rect 634294 993809 634346 993815
rect 637378 993783 637406 995522
rect 638530 993783 638558 995522
rect 639202 993931 639230 995522
rect 639188 993922 639244 993931
rect 639188 993857 639244 993866
rect 634294 993751 634346 993757
rect 637364 993774 637420 993783
rect 637364 993709 637420 993718
rect 638516 993774 638572 993783
rect 641026 993741 641054 995522
rect 641108 993774 641164 993783
rect 638516 993709 638572 993718
rect 641014 993735 641066 993741
rect 641108 993709 641164 993718
rect 641014 993677 641066 993683
rect 592438 989813 592490 989819
rect 592438 989755 592490 989761
rect 592450 983534 592478 989755
rect 608758 989739 608810 989745
rect 608758 989681 608810 989687
rect 608770 983534 608798 989681
rect 624982 989665 625034 989671
rect 624982 989607 625034 989613
rect 624994 983534 625022 989607
rect 641122 983534 641150 993709
rect 660886 989591 660938 989597
rect 660886 989533 660938 989539
rect 649558 989517 649610 989523
rect 649558 989459 649610 989465
rect 649462 987445 649514 987451
rect 649462 987387 649514 987393
rect 649366 987075 649418 987081
rect 649366 987017 649418 987023
rect 94870 983465 94922 983471
rect 65110 983449 65162 983455
rect 65110 983391 65162 983397
rect 63382 983375 63434 983381
rect 63382 983317 63434 983323
rect 63190 983301 63242 983307
rect 63190 983243 63242 983249
rect 62902 983227 62954 983233
rect 62902 983169 62954 983175
rect 62914 974945 62942 983169
rect 63094 983153 63146 983159
rect 63094 983095 63146 983101
rect 63106 977757 63134 983095
rect 63202 979311 63230 983243
rect 63286 983005 63338 983011
rect 63286 982947 63338 982953
rect 63190 979305 63242 979311
rect 63190 979247 63242 979253
rect 63094 977751 63146 977757
rect 63094 977693 63146 977699
rect 63298 976499 63326 982947
rect 63286 976493 63338 976499
rect 63286 976435 63338 976441
rect 62902 974939 62954 974945
rect 62902 974881 62954 974887
rect 63394 973539 63422 983317
rect 65122 976425 65150 983391
rect 65110 976419 65162 976425
rect 65110 976361 65162 976367
rect 63382 973533 63434 973539
rect 63382 973475 63434 973481
rect 62134 941787 62186 941793
rect 62134 941729 62186 941735
rect 62038 938975 62090 938981
rect 62038 938917 62090 938923
rect 62038 823757 62090 823763
rect 62038 823699 62090 823705
rect 61940 384458 61996 384467
rect 61940 384393 61996 384402
rect 61846 381607 61898 381613
rect 61846 381549 61898 381555
rect 59444 376318 59500 376327
rect 59444 376253 59500 376262
rect 59458 374435 59486 376253
rect 59446 374429 59498 374435
rect 59446 374371 59498 374377
rect 58388 363294 58444 363303
rect 58388 363229 58444 363238
rect 58402 362965 58430 363229
rect 58390 362959 58442 362965
rect 58390 362901 58442 362907
rect 59540 350270 59596 350279
rect 59540 350205 59596 350214
rect 59554 348535 59582 350205
rect 59542 348529 59594 348535
rect 59542 348471 59594 348477
rect 53398 345939 53450 345945
rect 53398 345881 53450 345887
rect 59540 337246 59596 337255
rect 59540 337181 59596 337190
rect 59554 337065 59582 337181
rect 59542 337059 59594 337065
rect 59542 337001 59594 337007
rect 59540 324222 59596 324231
rect 59540 324157 59596 324166
rect 59554 322635 59582 324157
rect 53398 322629 53450 322635
rect 53398 322571 53450 322577
rect 59542 322629 59594 322635
rect 59542 322571 59594 322577
rect 53302 301613 53354 301619
rect 53302 301555 53354 301561
rect 53206 290957 53258 290963
rect 53206 290899 53258 290905
rect 50422 259729 50474 259735
rect 50422 259671 50474 259677
rect 53410 258995 53438 322571
rect 58580 311198 58636 311207
rect 58580 311133 58636 311142
rect 58594 311091 58622 311133
rect 58582 311085 58634 311091
rect 58582 311027 58634 311033
rect 58966 305239 59018 305245
rect 58966 305181 59018 305187
rect 53686 302575 53738 302581
rect 53686 302517 53738 302523
rect 53698 301175 53726 302517
rect 53686 301169 53738 301175
rect 53686 301111 53738 301117
rect 55318 301169 55370 301175
rect 55318 301111 55370 301117
rect 55330 293849 55358 301111
rect 55318 293843 55370 293849
rect 55318 293785 55370 293791
rect 57526 290957 57578 290963
rect 57526 290899 57578 290905
rect 57538 285265 57566 290899
rect 57526 285259 57578 285265
rect 57526 285201 57578 285207
rect 58978 278605 59006 305181
rect 59540 298026 59596 298035
rect 59540 297961 59596 297970
rect 59554 296735 59582 297961
rect 59542 296729 59594 296735
rect 59542 296671 59594 296677
rect 60310 293843 60362 293849
rect 60310 293785 60362 293791
rect 59542 285185 59594 285191
rect 59540 285150 59542 285159
rect 59594 285150 59596 285159
rect 59540 285085 59596 285094
rect 60322 278679 60350 293785
rect 60406 293769 60458 293775
rect 60406 293711 60458 293717
rect 60418 287948 60446 293711
rect 60418 287920 60638 287948
rect 60406 285111 60458 285117
rect 60406 285053 60458 285059
rect 60418 282176 60446 285053
rect 60418 282148 60542 282176
rect 60310 278673 60362 278679
rect 60310 278615 60362 278621
rect 58966 278599 59018 278605
rect 58966 278541 59018 278547
rect 60514 278531 60542 282148
rect 60502 278525 60554 278531
rect 60502 278467 60554 278473
rect 60610 278457 60638 287920
rect 60598 278451 60650 278457
rect 60598 278393 60650 278399
rect 62050 278351 62078 823699
rect 62228 389194 62284 389203
rect 62228 389129 62284 389138
rect 62036 278342 62092 278351
rect 62036 278277 62092 278286
rect 62242 278203 62270 389129
rect 63286 285259 63338 285265
rect 63286 285201 63338 285207
rect 63298 282324 63326 285201
rect 63298 282296 63422 282324
rect 62228 278194 62284 278203
rect 62228 278129 62284 278138
rect 63394 278055 63422 282296
rect 320950 278081 321002 278087
rect 63380 278046 63436 278055
rect 422518 278081 422570 278087
rect 320950 278023 321002 278029
rect 63380 277981 63436 277990
rect 317878 278007 317930 278013
rect 317878 277949 317930 277955
rect 65890 269323 65918 277870
rect 67042 269471 67070 277870
rect 68194 270761 68222 277870
rect 69442 272283 69470 277870
rect 69428 272274 69484 272283
rect 69428 272209 69484 272218
rect 68182 270755 68234 270761
rect 68182 270697 68234 270703
rect 69046 270755 69098 270761
rect 69046 270697 69098 270703
rect 67028 269462 67084 269471
rect 67028 269397 67084 269406
rect 65876 269314 65932 269323
rect 65876 269249 65932 269258
rect 53398 258989 53450 258995
rect 53398 258931 53450 258937
rect 48022 249443 48074 249449
rect 48022 249385 48074 249391
rect 47926 249221 47978 249227
rect 47926 249163 47978 249169
rect 69058 246785 69086 270697
rect 70594 269619 70622 277870
rect 71746 272135 71774 277870
rect 72994 272167 73022 277870
rect 72982 272161 73034 272167
rect 71732 272126 71788 272135
rect 72982 272103 73034 272109
rect 71732 272061 71788 272070
rect 70580 269610 70636 269619
rect 70580 269545 70636 269554
rect 74050 269355 74078 277870
rect 75298 271205 75326 277870
rect 75286 271199 75338 271205
rect 75286 271141 75338 271147
rect 76450 269503 76478 277870
rect 77494 271199 77546 271205
rect 77494 271141 77546 271147
rect 76438 269497 76490 269503
rect 76438 269439 76490 269445
rect 74038 269349 74090 269355
rect 74038 269291 74090 269297
rect 77506 246859 77534 271141
rect 77698 269281 77726 277870
rect 78850 269429 78878 277870
rect 80098 273499 80126 277870
rect 80086 273493 80138 273499
rect 80086 273435 80138 273441
rect 81250 272315 81278 277870
rect 81238 272309 81290 272315
rect 81238 272251 81290 272257
rect 82402 272241 82430 277870
rect 82390 272235 82442 272241
rect 82390 272177 82442 272183
rect 83554 269577 83582 277870
rect 84802 273573 84830 277870
rect 84790 273567 84842 273573
rect 84790 273509 84842 273515
rect 85954 269651 85982 277870
rect 87106 272389 87134 277870
rect 87094 272383 87146 272389
rect 87094 272325 87146 272331
rect 88354 269725 88382 277870
rect 89506 271945 89534 277870
rect 90658 272463 90686 277870
rect 90646 272457 90698 272463
rect 90646 272399 90698 272405
rect 89494 271939 89546 271945
rect 89494 271881 89546 271887
rect 91810 269799 91838 277870
rect 93058 272537 93086 277870
rect 93046 272531 93098 272537
rect 93046 272473 93098 272479
rect 94210 271797 94238 277870
rect 95458 272685 95486 277870
rect 95446 272679 95498 272685
rect 95446 272621 95498 272627
rect 94198 271791 94250 271797
rect 94198 271733 94250 271739
rect 96610 269873 96638 277870
rect 97762 272019 97790 277870
rect 97750 272013 97802 272019
rect 97750 271955 97802 271961
rect 98914 269947 98942 277870
rect 100162 272611 100190 277870
rect 100150 272605 100202 272611
rect 100150 272547 100202 272553
rect 101314 272093 101342 277870
rect 102562 272759 102590 277870
rect 102550 272753 102602 272759
rect 102550 272695 102602 272701
rect 101302 272087 101354 272093
rect 101302 272029 101354 272035
rect 103714 270095 103742 277870
rect 104866 271723 104894 277870
rect 104854 271717 104906 271723
rect 104854 271659 104906 271665
rect 103702 270089 103754 270095
rect 103702 270031 103754 270037
rect 106018 270021 106046 277870
rect 107170 272833 107198 277870
rect 107158 272827 107210 272833
rect 107158 272769 107210 272775
rect 108418 271649 108446 277870
rect 109570 272907 109598 277870
rect 109558 272901 109610 272907
rect 109558 272843 109610 272849
rect 108406 271643 108458 271649
rect 108406 271585 108458 271591
rect 110818 270169 110846 277870
rect 111970 271871 111998 277870
rect 113218 273055 113246 277870
rect 113206 273049 113258 273055
rect 113206 272991 113258 272997
rect 111958 271865 112010 271871
rect 111958 271807 112010 271813
rect 114274 270243 114302 277870
rect 115522 270761 115550 277870
rect 116674 273129 116702 277870
rect 116662 273123 116714 273129
rect 116662 273065 116714 273071
rect 115510 270755 115562 270761
rect 115510 270697 115562 270703
rect 117922 270317 117950 277870
rect 119074 273351 119102 277870
rect 119062 273345 119114 273351
rect 119062 273287 119114 273293
rect 120226 272981 120254 277870
rect 120886 273345 120938 273351
rect 120886 273287 120938 273293
rect 120214 272975 120266 272981
rect 120214 272917 120266 272923
rect 118006 270755 118058 270761
rect 118006 270697 118058 270703
rect 117910 270311 117962 270317
rect 117910 270253 117962 270259
rect 114262 270237 114314 270243
rect 114262 270179 114314 270185
rect 110806 270163 110858 270169
rect 110806 270105 110858 270111
rect 106006 270015 106058 270021
rect 106006 269957 106058 269963
rect 98902 269941 98954 269947
rect 98902 269883 98954 269889
rect 96598 269867 96650 269873
rect 96598 269809 96650 269815
rect 91798 269793 91850 269799
rect 91798 269735 91850 269741
rect 88342 269719 88394 269725
rect 88342 269661 88394 269667
rect 85942 269645 85994 269651
rect 85942 269587 85994 269593
rect 83542 269571 83594 269577
rect 83542 269513 83594 269519
rect 78838 269423 78890 269429
rect 78838 269365 78890 269371
rect 77686 269275 77738 269281
rect 77686 269217 77738 269223
rect 118018 247007 118046 270697
rect 120898 249523 120926 273287
rect 121378 270391 121406 277870
rect 122530 270761 122558 277870
rect 123778 273203 123806 277870
rect 123766 273197 123818 273203
rect 123766 273139 123818 273145
rect 122518 270755 122570 270761
rect 122518 270697 122570 270703
rect 123766 270755 123818 270761
rect 123766 270697 123818 270703
rect 121366 270385 121418 270391
rect 121366 270327 121418 270333
rect 120886 249517 120938 249523
rect 120886 249459 120938 249465
rect 118006 247001 118058 247007
rect 118006 246943 118058 246949
rect 123778 246933 123806 270697
rect 124930 270465 124958 277870
rect 126178 271575 126206 277870
rect 127330 273277 127358 277870
rect 127318 273271 127370 273277
rect 127318 273213 127370 273219
rect 126166 271569 126218 271575
rect 126166 271511 126218 271517
rect 124918 270459 124970 270465
rect 124918 270401 124970 270407
rect 128578 269767 128606 277870
rect 129634 271501 129662 277870
rect 129622 271495 129674 271501
rect 129622 271437 129674 271443
rect 130882 269915 130910 277870
rect 132034 273351 132062 277870
rect 132022 273345 132074 273351
rect 132022 273287 132074 273293
rect 133282 271427 133310 277870
rect 133270 271421 133322 271427
rect 133270 271363 133322 271369
rect 134434 270539 134462 277870
rect 134422 270533 134474 270539
rect 134422 270475 134474 270481
rect 130868 269906 130924 269915
rect 130868 269841 130924 269850
rect 128564 269758 128620 269767
rect 128564 269693 128620 269702
rect 135682 269207 135710 277870
rect 136834 271279 136862 277870
rect 136822 271273 136874 271279
rect 136822 271215 136874 271221
rect 137890 270613 137918 277870
rect 139138 273425 139166 277870
rect 139126 273419 139178 273425
rect 139126 273361 139178 273367
rect 140290 271131 140318 277870
rect 140278 271125 140330 271131
rect 140278 271067 140330 271073
rect 137878 270607 137930 270613
rect 137878 270549 137930 270555
rect 135670 269201 135722 269207
rect 135670 269143 135722 269149
rect 141538 269133 141566 277870
rect 142390 273567 142442 273573
rect 142390 273509 142442 273515
rect 141526 269127 141578 269133
rect 141526 269069 141578 269075
rect 142402 262473 142430 273509
rect 142486 273493 142538 273499
rect 142486 273435 142538 273441
rect 142390 262467 142442 262473
rect 142390 262409 142442 262415
rect 123766 246927 123818 246933
rect 123766 246869 123818 246875
rect 77494 246853 77546 246859
rect 77494 246795 77546 246801
rect 69046 246779 69098 246785
rect 69046 246721 69098 246727
rect 47446 246705 47498 246711
rect 47446 246647 47498 246653
rect 46006 246557 46058 246563
rect 46006 246499 46058 246505
rect 45622 246409 45674 246415
rect 45622 246351 45674 246357
rect 45526 246335 45578 246341
rect 45526 246277 45578 246283
rect 45334 242783 45386 242789
rect 45334 242725 45386 242731
rect 45238 215255 45290 215261
rect 45238 215197 45290 215203
rect 45346 214299 45374 242725
rect 45334 214293 45386 214299
rect 45334 214235 45386 214241
rect 45046 204969 45098 204975
rect 45046 204911 45098 204917
rect 44854 203785 44906 203791
rect 44854 203727 44906 203733
rect 43222 196903 43274 196909
rect 43222 196845 43274 196851
rect 43126 191501 43178 191507
rect 43126 191443 43178 191449
rect 42166 191057 42218 191063
rect 42166 190999 42218 191005
rect 43030 191057 43082 191063
rect 43030 190999 43082 191005
rect 42178 190476 42206 190999
rect 41780 190134 41836 190143
rect 41780 190069 41836 190078
rect 41794 189929 41822 190069
rect 43234 187881 43262 196845
rect 42166 187875 42218 187881
rect 42166 187817 42218 187823
rect 43222 187875 43274 187881
rect 43222 187817 43274 187823
rect 42178 187442 42206 187817
rect 41780 187174 41836 187183
rect 41780 187109 41836 187118
rect 41794 186776 41822 187109
rect 41780 186730 41836 186739
rect 41780 186665 41836 186674
rect 41794 186184 41822 186665
rect 41780 185842 41836 185851
rect 41780 185777 41836 185786
rect 41794 185592 41822 185777
rect 41780 184066 41836 184075
rect 41780 184001 41836 184010
rect 41794 183742 41822 184001
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183121 41822 183557
rect 41780 183030 41836 183039
rect 41780 182965 41836 182974
rect 41794 182484 41822 182965
rect 142508 178280 142536 273435
rect 142582 271939 142634 271945
rect 142582 271881 142634 271887
rect 142594 178428 142622 271881
rect 142690 270687 142718 277870
rect 142774 271791 142826 271797
rect 142774 271733 142826 271739
rect 142678 270681 142730 270687
rect 142678 270623 142730 270629
rect 142678 262467 142730 262473
rect 142678 262409 142730 262415
rect 142690 180130 142718 262409
rect 142786 182128 142814 271733
rect 143062 271569 143114 271575
rect 143062 271511 143114 271517
rect 142966 271495 143018 271501
rect 142966 271437 143018 271443
rect 142870 271421 142922 271427
rect 142870 271363 142922 271369
rect 142882 187012 142910 271363
rect 142978 187308 143006 271437
rect 143074 187456 143102 271511
rect 143158 271273 143210 271279
rect 143158 271215 143210 271221
rect 143170 190101 143198 271215
rect 143254 271125 143306 271131
rect 143254 271067 143306 271073
rect 143158 190095 143210 190101
rect 143158 190037 143210 190043
rect 143266 190027 143294 271067
rect 143938 270761 143966 277870
rect 143926 270755 143978 270761
rect 143926 270697 143978 270703
rect 144994 269059 145022 277870
rect 146242 273499 146270 277870
rect 146230 273493 146282 273499
rect 146230 273435 146282 273441
rect 147394 270761 147422 277870
rect 145366 270755 145418 270761
rect 145366 270697 145418 270703
rect 147382 270755 147434 270761
rect 147382 270697 147434 270703
rect 144982 269053 145034 269059
rect 144982 268995 145034 269001
rect 143254 190021 143306 190027
rect 143254 189963 143306 189969
rect 145378 189953 145406 270697
rect 148642 268985 148670 277870
rect 149794 273573 149822 277870
rect 149782 273567 149834 273573
rect 149782 273509 149834 273515
rect 151042 270761 151070 277870
rect 151126 272013 151178 272019
rect 151126 271955 151178 271961
rect 149686 270755 149738 270761
rect 149686 270697 149738 270703
rect 151030 270755 151082 270761
rect 151030 270697 151082 270703
rect 148630 268979 148682 268985
rect 148630 268921 148682 268927
rect 145558 249517 145610 249523
rect 145558 249459 145610 249465
rect 145462 246853 145514 246859
rect 145462 246795 145514 246801
rect 145366 189947 145418 189953
rect 145366 189889 145418 189895
rect 143074 187428 143390 187456
rect 142978 187280 143294 187308
rect 143158 187209 143210 187215
rect 143158 187151 143210 187157
rect 143170 187012 143198 187151
rect 143266 187067 143294 187280
rect 143362 187141 143390 187428
rect 143350 187135 143402 187141
rect 143350 187077 143402 187083
rect 142882 186984 143198 187012
rect 143254 187061 143306 187067
rect 143254 187003 143306 187009
rect 142786 182100 143102 182128
rect 143074 181443 143102 182100
rect 143062 181437 143114 181443
rect 143062 181379 143114 181385
rect 142690 180102 143102 180130
rect 143074 178557 143102 180102
rect 143062 178551 143114 178557
rect 143062 178493 143114 178499
rect 142594 178409 143102 178428
rect 142594 178403 143114 178409
rect 142594 178400 143062 178403
rect 143062 178345 143114 178351
rect 143158 178329 143210 178335
rect 142508 178277 143158 178280
rect 142508 178271 143210 178277
rect 142508 178252 143198 178271
rect 145474 175671 145502 246795
rect 145570 184255 145598 249459
rect 145654 247001 145706 247007
rect 145654 246943 145706 246949
rect 145666 184329 145694 246943
rect 145750 246779 145802 246785
rect 145750 246721 145802 246727
rect 145762 201571 145790 246721
rect 149396 244598 149452 244607
rect 149396 244533 149452 244542
rect 148244 242082 148300 242091
rect 148244 242017 148300 242026
rect 146900 229946 146956 229955
rect 146900 229881 146956 229890
rect 145750 201565 145802 201571
rect 145750 201507 145802 201513
rect 146914 188843 146942 229881
rect 146996 228170 147052 228179
rect 146996 228105 147052 228114
rect 146902 188837 146954 188843
rect 146902 188779 146954 188785
rect 145654 184323 145706 184329
rect 145654 184265 145706 184271
rect 145558 184249 145610 184255
rect 145558 184191 145610 184197
rect 145462 175665 145514 175671
rect 145462 175607 145514 175613
rect 146900 165566 146956 165575
rect 146900 165501 146956 165510
rect 146914 123871 146942 165501
rect 147010 164497 147038 228105
rect 148148 222694 148204 222703
rect 148148 222629 148204 222638
rect 148052 221510 148108 221519
rect 148052 221445 148108 221454
rect 147380 217810 147436 217819
rect 147380 217745 147436 217754
rect 147394 216889 147422 217745
rect 147382 216883 147434 216889
rect 147382 216825 147434 216831
rect 147284 216626 147340 216635
rect 147284 216561 147340 216570
rect 147298 216297 147326 216561
rect 147286 216291 147338 216297
rect 147286 216233 147338 216239
rect 147380 214850 147436 214859
rect 147380 214785 147436 214794
rect 147394 213337 147422 214785
rect 147382 213331 147434 213337
rect 147382 213273 147434 213279
rect 147092 212926 147148 212935
rect 147092 212861 147148 212870
rect 147106 212523 147134 212861
rect 147094 212517 147146 212523
rect 147094 212459 147146 212465
rect 147380 211742 147436 211751
rect 147380 211677 147436 211686
rect 147394 210377 147422 211677
rect 147382 210371 147434 210377
rect 147382 210313 147434 210319
rect 147284 209226 147340 209235
rect 147284 209161 147340 209170
rect 147298 207491 147326 209161
rect 147286 207485 147338 207491
rect 147286 207427 147338 207433
rect 147956 201678 148012 201687
rect 147956 201613 148012 201622
rect 147860 198422 147916 198431
rect 147860 198357 147916 198366
rect 147764 192206 147820 192215
rect 147764 192141 147820 192150
rect 147572 191022 147628 191031
rect 147572 190957 147628 190966
rect 147586 190249 147614 190957
rect 147574 190243 147626 190249
rect 147574 190185 147626 190191
rect 147476 189838 147532 189847
rect 147476 189773 147532 189782
rect 147286 188837 147338 188843
rect 147286 188779 147338 188785
rect 147188 177702 147244 177711
rect 147188 177637 147244 177646
rect 147202 176781 147230 177637
rect 147190 176775 147242 176781
rect 147190 176717 147242 176723
rect 147188 176518 147244 176527
rect 147188 176453 147244 176462
rect 147092 175186 147148 175195
rect 147092 175121 147148 175130
rect 146998 164491 147050 164497
rect 146998 164433 147050 164439
rect 146996 164382 147052 164391
rect 146996 164317 147052 164326
rect 146902 123865 146954 123871
rect 146902 123807 146954 123813
rect 147010 123797 147038 164317
rect 147106 129569 147134 175121
rect 147202 132455 147230 176453
rect 147298 170417 147326 188779
rect 147380 178886 147436 178895
rect 147380 178821 147382 178830
rect 147434 178821 147436 178830
rect 147382 178789 147434 178795
rect 147380 174002 147436 174011
rect 147380 173937 147436 173946
rect 147286 170411 147338 170417
rect 147286 170353 147338 170359
rect 147284 170302 147340 170311
rect 147284 170237 147340 170246
rect 147190 132449 147242 132455
rect 147190 132391 147242 132397
rect 147094 129563 147146 129569
rect 147094 129505 147146 129511
rect 147092 129158 147148 129167
rect 147092 129093 147148 129102
rect 146998 123791 147050 123797
rect 146998 123733 147050 123739
rect 146996 120574 147052 120583
rect 146996 120509 147052 120518
rect 146900 111990 146956 111999
rect 146900 111925 146956 111934
rect 146914 92125 146942 111925
rect 147010 97897 147038 120509
rect 147106 103595 147134 129093
rect 147298 126683 147326 170237
rect 147394 129495 147422 173937
rect 147490 141039 147518 189773
rect 147668 187470 147724 187479
rect 147668 187405 147724 187414
rect 147572 183770 147628 183779
rect 147572 183705 147628 183714
rect 147478 141033 147530 141039
rect 147478 140975 147530 140981
rect 147586 135341 147614 183705
rect 147682 141428 147710 187405
rect 147778 143796 147806 192141
rect 147874 143999 147902 198357
rect 147970 146663 147998 201613
rect 148066 158429 148094 221445
rect 148162 161241 148190 222629
rect 148258 172785 148286 242017
rect 149410 241975 149438 244533
rect 149398 241969 149450 241975
rect 149398 241911 149450 241917
rect 148724 240898 148780 240907
rect 148724 240833 148780 240842
rect 148532 238530 148588 238539
rect 148532 238465 148588 238474
rect 148340 236754 148396 236763
rect 148340 236689 148396 236698
rect 148246 172779 148298 172785
rect 148246 172721 148298 172727
rect 148246 170411 148298 170417
rect 148246 170353 148298 170359
rect 148258 163757 148286 170353
rect 148354 169825 148382 236689
rect 148436 233646 148492 233655
rect 148436 233581 148492 233590
rect 148342 169819 148394 169825
rect 148342 169761 148394 169767
rect 148450 167013 148478 233581
rect 148546 169899 148574 238465
rect 148628 231130 148684 231139
rect 148628 231065 148684 231074
rect 148534 169893 148586 169899
rect 148534 169835 148586 169841
rect 148438 167007 148490 167013
rect 148438 166949 148490 166955
rect 148642 164127 148670 231065
rect 148738 172711 148766 240833
rect 149396 239714 149452 239723
rect 149396 239649 149452 239658
rect 149410 239089 149438 239649
rect 149398 239083 149450 239089
rect 149398 239025 149450 239031
rect 149012 236014 149068 236023
rect 149012 235949 149068 235958
rect 148820 226394 148876 226403
rect 148820 226329 148876 226338
rect 148726 172705 148778 172711
rect 148726 172647 148778 172653
rect 148630 164121 148682 164127
rect 148630 164063 148682 164069
rect 148246 163751 148298 163757
rect 148246 163693 148298 163699
rect 148150 161235 148202 161241
rect 148150 161177 148202 161183
rect 148834 161167 148862 226329
rect 148916 219734 148972 219743
rect 148916 219669 148972 219678
rect 148930 198611 148958 219669
rect 148918 198605 148970 198611
rect 148918 198547 148970 198553
rect 148918 198457 148970 198463
rect 148918 198399 148970 198405
rect 148930 189879 148958 198399
rect 148918 189873 148970 189879
rect 148918 189815 148970 189821
rect 148916 184510 148972 184519
rect 148916 184445 148972 184454
rect 148930 178483 148958 184445
rect 148918 178477 148970 178483
rect 148918 178419 148970 178425
rect 148916 172818 148972 172827
rect 148916 172753 148972 172762
rect 148930 169548 148958 172753
rect 149026 169751 149054 235949
rect 149396 234830 149452 234839
rect 149396 234765 149452 234774
rect 149410 234427 149438 234765
rect 149398 234421 149450 234427
rect 149398 234363 149450 234369
rect 149204 232314 149260 232323
rect 149204 232249 149260 232258
rect 149108 225210 149164 225219
rect 149108 225145 149164 225154
rect 149014 169745 149066 169751
rect 149014 169687 149066 169693
rect 148930 169520 149054 169548
rect 148916 168082 148972 168091
rect 148916 168017 148972 168026
rect 148822 161161 148874 161167
rect 148822 161103 148874 161109
rect 148340 159498 148396 159507
rect 148340 159433 148396 159442
rect 148054 158423 148106 158429
rect 148054 158365 148106 158371
rect 148244 156982 148300 156991
rect 148244 156917 148300 156926
rect 148052 148546 148108 148555
rect 148052 148481 148108 148490
rect 148066 148069 148094 148481
rect 148054 148063 148106 148069
rect 148054 148005 148106 148011
rect 148052 147362 148108 147371
rect 148052 147297 148108 147306
rect 148066 147033 148094 147297
rect 148054 147027 148106 147033
rect 148054 146969 148106 146975
rect 147958 146657 148010 146663
rect 147958 146599 148010 146605
rect 147956 146178 148012 146187
rect 147956 146113 148012 146122
rect 147970 145849 147998 146113
rect 147958 145843 148010 145849
rect 147958 145785 148010 145791
rect 147956 144402 148012 144411
rect 147956 144337 147958 144346
rect 148010 144337 148012 144346
rect 147958 144305 148010 144311
rect 147862 143993 147914 143999
rect 147862 143935 147914 143941
rect 147778 143768 147998 143796
rect 147860 143662 147916 143671
rect 147860 143597 147916 143606
rect 147874 142593 147902 143597
rect 147862 142587 147914 142593
rect 147862 142529 147914 142535
rect 147860 142478 147916 142487
rect 147860 142413 147916 142422
rect 147874 141557 147902 142413
rect 147862 141551 147914 141557
rect 147862 141493 147914 141499
rect 147682 141400 147902 141428
rect 147668 141294 147724 141303
rect 147668 141229 147670 141238
rect 147722 141229 147724 141238
rect 147670 141197 147722 141203
rect 147874 138227 147902 141400
rect 147970 141113 147998 143768
rect 147958 141107 148010 141113
rect 147958 141049 148010 141055
rect 147956 138778 148012 138787
rect 147956 138713 148012 138722
rect 147862 138221 147914 138227
rect 147862 138163 147914 138169
rect 147574 135335 147626 135341
rect 147574 135277 147626 135283
rect 147860 135078 147916 135087
rect 147860 135013 147916 135022
rect 147668 133894 147724 133903
rect 147668 133829 147724 133838
rect 147572 130934 147628 130943
rect 147572 130869 147628 130878
rect 147382 129489 147434 129495
rect 147382 129431 147434 129437
rect 147286 126677 147338 126683
rect 147188 126642 147244 126651
rect 147286 126619 147338 126625
rect 147188 126577 147244 126586
rect 147094 103589 147146 103595
rect 147094 103531 147146 103537
rect 147202 100783 147230 126577
rect 147284 125458 147340 125467
rect 147284 125393 147340 125402
rect 147190 100777 147242 100783
rect 147190 100719 147242 100725
rect 147298 100709 147326 125393
rect 147380 124274 147436 124283
rect 147380 124209 147436 124218
rect 147286 100703 147338 100709
rect 147286 100645 147338 100651
rect 147394 100635 147422 124209
rect 147476 122498 147532 122507
rect 147476 122433 147532 122442
rect 147382 100629 147434 100635
rect 147382 100571 147434 100577
rect 146998 97891 147050 97897
rect 146998 97833 147050 97839
rect 147490 97823 147518 122433
rect 147586 103669 147614 130869
rect 147682 106555 147710 133829
rect 147764 130342 147820 130351
rect 147764 130277 147820 130286
rect 147670 106549 147722 106555
rect 147670 106491 147722 106497
rect 147574 103663 147626 103669
rect 147574 103605 147626 103611
rect 147668 103554 147724 103563
rect 147778 103521 147806 130277
rect 147874 106407 147902 135013
rect 147970 109441 147998 138713
rect 148052 137594 148108 137603
rect 148052 137529 148108 137538
rect 147958 109435 148010 109441
rect 147958 109377 148010 109383
rect 148066 106481 148094 137529
rect 148148 132710 148204 132719
rect 148148 132645 148204 132654
rect 148054 106475 148106 106481
rect 148054 106417 148106 106423
rect 147862 106401 147914 106407
rect 147862 106343 147914 106349
rect 147956 106070 148012 106079
rect 147956 106005 148012 106014
rect 147668 103489 147724 103498
rect 147766 103515 147818 103521
rect 147478 97817 147530 97823
rect 147478 97759 147530 97765
rect 147572 94970 147628 94979
rect 147572 94905 147628 94914
rect 146902 92119 146954 92125
rect 146902 92061 146954 92067
rect 147586 80507 147614 94905
rect 147682 86353 147710 103489
rect 147766 103457 147818 103463
rect 147970 89239 147998 106005
rect 148052 104738 148108 104747
rect 148052 104673 148108 104682
rect 147958 89233 148010 89239
rect 147958 89175 148010 89181
rect 148066 86427 148094 104673
rect 148162 103447 148190 132645
rect 148258 112327 148286 156917
rect 148354 115213 148382 159433
rect 148820 157722 148876 157731
rect 148820 157657 148876 157666
rect 148436 155798 148492 155807
rect 148436 155733 148492 155742
rect 148342 115207 148394 115213
rect 148342 115149 148394 115155
rect 148246 112321 148298 112327
rect 148246 112263 148298 112269
rect 148450 112179 148478 155733
rect 148628 154614 148684 154623
rect 148628 154549 148684 154558
rect 148532 150914 148588 150923
rect 148532 150849 148588 150858
rect 148438 112173 148490 112179
rect 148438 112115 148490 112121
rect 148340 109474 148396 109483
rect 148340 109409 148396 109418
rect 148150 103441 148202 103447
rect 148150 103383 148202 103389
rect 148244 99854 148300 99863
rect 148244 99789 148300 99798
rect 148148 98670 148204 98679
rect 148148 98605 148204 98614
rect 148054 86421 148106 86427
rect 148054 86363 148106 86369
rect 147670 86347 147722 86353
rect 147670 86289 147722 86295
rect 148162 83319 148190 98605
rect 148258 83541 148286 99789
rect 148354 89091 148382 109409
rect 148546 109293 148574 150849
rect 148642 112253 148670 154549
rect 148724 152098 148780 152107
rect 148724 152033 148780 152042
rect 148630 112247 148682 112253
rect 148630 112189 148682 112195
rect 148738 109367 148766 152033
rect 148834 115139 148862 157657
rect 148930 126609 148958 168017
rect 149026 163905 149054 169520
rect 149014 163899 149066 163905
rect 149014 163841 149066 163847
rect 149012 161866 149068 161875
rect 149012 161801 149068 161810
rect 148918 126603 148970 126609
rect 148918 126545 148970 126551
rect 149026 120837 149054 161801
rect 149122 161093 149150 225145
rect 149218 166939 149246 232249
rect 149396 227430 149452 227439
rect 149396 227365 149452 227374
rect 149300 206414 149356 206423
rect 149300 206349 149356 206358
rect 149314 204531 149342 206349
rect 149302 204525 149354 204531
rect 149302 204467 149354 204473
rect 149300 199606 149356 199615
rect 149300 199541 149356 199550
rect 149314 198833 149342 199541
rect 149302 198827 149354 198833
rect 149302 198769 149354 198775
rect 149302 195941 149354 195947
rect 149300 195906 149302 195915
rect 149354 195906 149356 195915
rect 149300 195841 149356 195850
rect 149410 194856 149438 227365
rect 149492 223878 149548 223887
rect 149492 223813 149548 223822
rect 149506 216014 149534 223813
rect 149588 218994 149644 219003
rect 149588 218929 149590 218938
rect 149642 218929 149644 218938
rect 149590 218897 149642 218903
rect 149506 215986 149630 216014
rect 149492 214110 149548 214119
rect 149492 214045 149548 214054
rect 149506 213189 149534 214045
rect 149494 213183 149546 213189
rect 149494 213125 149546 213131
rect 149492 210410 149548 210419
rect 149492 210345 149548 210354
rect 149506 210303 149534 210345
rect 149494 210297 149546 210303
rect 149494 210239 149546 210245
rect 149492 208042 149548 208051
rect 149492 207977 149548 207986
rect 149506 207417 149534 207977
rect 149494 207411 149546 207417
rect 149494 207353 149546 207359
rect 149492 205674 149548 205683
rect 149492 205609 149548 205618
rect 149506 204605 149534 205609
rect 149494 204599 149546 204605
rect 149494 204541 149546 204547
rect 149492 203306 149548 203315
rect 149492 203241 149548 203250
rect 149506 201645 149534 203241
rect 149494 201639 149546 201645
rect 149494 201581 149546 201587
rect 149492 200790 149548 200799
rect 149492 200725 149548 200734
rect 149506 198759 149534 200725
rect 149494 198753 149546 198759
rect 149494 198695 149546 198701
rect 149494 198605 149546 198611
rect 149494 198547 149546 198553
rect 149314 194828 149438 194856
rect 149206 166933 149258 166939
rect 149206 166875 149258 166881
rect 149204 166306 149260 166315
rect 149204 166241 149260 166250
rect 149110 161087 149162 161093
rect 149110 161029 149162 161035
rect 149108 160682 149164 160691
rect 149108 160617 149164 160626
rect 149122 120985 149150 160617
rect 149218 150215 149246 166241
rect 149314 164053 149342 194828
rect 149396 194722 149452 194731
rect 149396 194657 149398 194666
rect 149450 194657 149452 194666
rect 149398 194625 149450 194631
rect 149396 193094 149452 193103
rect 149396 193029 149398 193038
rect 149450 193029 149452 193038
rect 149398 192997 149450 193003
rect 149396 188062 149452 188071
rect 149396 187997 149452 188006
rect 149410 187289 149438 187997
rect 149398 187283 149450 187289
rect 149398 187225 149450 187231
rect 149396 186286 149452 186295
rect 149396 186221 149452 186230
rect 149410 184403 149438 186221
rect 149398 184397 149450 184403
rect 149398 184339 149450 184345
rect 149396 182586 149452 182595
rect 149396 182521 149452 182530
rect 149410 181517 149438 182521
rect 149398 181511 149450 181517
rect 149398 181453 149450 181459
rect 149396 179626 149452 179635
rect 149396 179561 149398 179570
rect 149450 179561 149452 179570
rect 149398 179529 149450 179535
rect 149396 171042 149452 171051
rect 149396 170977 149452 170986
rect 149410 169973 149438 170977
rect 149398 169967 149450 169973
rect 149398 169909 149450 169915
rect 149396 169118 149452 169127
rect 149396 169053 149452 169062
rect 149410 167087 149438 169053
rect 149398 167081 149450 167087
rect 149398 167023 149450 167029
rect 149302 164047 149354 164053
rect 149302 163989 149354 163995
rect 149302 163899 149354 163905
rect 149302 163841 149354 163847
rect 149206 150209 149258 150215
rect 149206 150151 149258 150157
rect 149206 140959 149258 140965
rect 149206 140901 149258 140907
rect 149218 139971 149246 140901
rect 149204 139962 149260 139971
rect 149204 139897 149260 139906
rect 149204 135818 149260 135827
rect 149204 135753 149260 135762
rect 149218 123372 149246 135753
rect 149314 129421 149342 163841
rect 149396 163198 149452 163207
rect 149396 163133 149452 163142
rect 149302 129415 149354 129421
rect 149302 129357 149354 129363
rect 149300 127974 149356 127983
rect 149300 127909 149356 127918
rect 149314 123520 149342 127909
rect 149410 125444 149438 163133
rect 149506 158355 149534 198547
rect 149602 161019 149630 215986
rect 149698 204624 149726 270697
rect 149698 204596 149822 204624
rect 149684 204490 149740 204499
rect 149684 204425 149740 204434
rect 149698 201719 149726 204425
rect 149686 201713 149738 201719
rect 149686 201655 149738 201661
rect 149794 201516 149822 204596
rect 149698 201488 149822 201516
rect 149698 198463 149726 201488
rect 149686 198457 149738 198463
rect 149686 198399 149738 198405
rect 149684 197090 149740 197099
rect 149684 197025 149740 197034
rect 149698 195873 149726 197025
rect 149686 195867 149738 195873
rect 149686 195809 149738 195815
rect 149684 181402 149740 181411
rect 151138 181369 151166 271955
rect 152194 268911 152222 277870
rect 152566 270755 152618 270761
rect 152566 270697 152618 270703
rect 152182 268905 152234 268911
rect 152182 268847 152234 268853
rect 151510 216883 151562 216889
rect 151510 216825 151562 216831
rect 151222 216291 151274 216297
rect 151222 216233 151274 216239
rect 149684 181337 149740 181346
rect 151126 181363 151178 181369
rect 149698 178631 149726 181337
rect 151126 181305 151178 181311
rect 149686 178625 149738 178631
rect 149686 178567 149738 178573
rect 149686 178477 149738 178483
rect 149686 178419 149738 178425
rect 149590 161013 149642 161019
rect 149590 160955 149642 160961
rect 149494 158349 149546 158355
rect 149494 158291 149546 158297
rect 149698 155534 149726 178419
rect 151126 176775 151178 176781
rect 151126 176717 151178 176723
rect 149506 155506 149726 155534
rect 149506 135267 149534 155506
rect 149686 150209 149738 150215
rect 149686 150151 149738 150157
rect 149588 149878 149644 149887
rect 149588 149813 149644 149822
rect 149494 135261 149546 135267
rect 149494 135203 149546 135209
rect 149410 125416 149534 125444
rect 149506 123723 149534 125416
rect 149494 123717 149546 123723
rect 149494 123659 149546 123665
rect 149314 123492 149534 123520
rect 149218 123344 149438 123372
rect 149300 121758 149356 121767
rect 149300 121693 149356 121702
rect 149110 120979 149162 120985
rect 149110 120921 149162 120927
rect 149014 120831 149066 120837
rect 149014 120773 149066 120779
rect 149204 119390 149260 119399
rect 149204 119325 149260 119334
rect 148916 118206 148972 118215
rect 148916 118141 148972 118150
rect 148822 115133 148874 115139
rect 148822 115075 148874 115081
rect 148820 110954 148876 110963
rect 148820 110889 148876 110898
rect 148726 109361 148778 109367
rect 148726 109303 148778 109309
rect 148534 109287 148586 109293
rect 148534 109229 148586 109235
rect 148436 108438 148492 108447
rect 148436 108373 148492 108382
rect 148450 89165 148478 108373
rect 148628 107254 148684 107263
rect 148628 107189 148684 107198
rect 148532 102370 148588 102379
rect 148532 102305 148588 102314
rect 148438 89159 148490 89165
rect 148438 89101 148490 89107
rect 148342 89085 148394 89091
rect 148342 89027 148394 89033
rect 148546 86279 148574 102305
rect 148642 89017 148670 107189
rect 148724 97486 148780 97495
rect 148724 97421 148780 97430
rect 148630 89011 148682 89017
rect 148630 88953 148682 88959
rect 148534 86273 148586 86279
rect 148534 86215 148586 86221
rect 148340 85350 148396 85359
rect 148340 85285 148396 85294
rect 148246 83535 148298 83541
rect 148246 83477 148298 83483
rect 148150 83313 148202 83319
rect 148150 83255 148202 83261
rect 147574 80501 147626 80507
rect 147574 80443 147626 80449
rect 148354 74809 148382 85285
rect 148532 84166 148588 84175
rect 148532 84101 148588 84110
rect 148436 81650 148492 81659
rect 148436 81585 148492 81594
rect 148342 74803 148394 74809
rect 148342 74745 148394 74751
rect 148450 71997 148478 81585
rect 148546 74735 148574 84101
rect 148738 83467 148766 97421
rect 148834 92051 148862 110889
rect 148930 95011 148958 118141
rect 149108 116874 149164 116883
rect 149108 116809 149164 116818
rect 149012 114506 149068 114515
rect 149012 114441 149068 114450
rect 148918 95005 148970 95011
rect 148918 94947 148970 94953
rect 148916 92602 148972 92611
rect 148916 92537 148972 92546
rect 148822 92045 148874 92051
rect 148822 91987 148874 91993
rect 148820 86534 148876 86543
rect 148820 86469 148876 86478
rect 148726 83461 148778 83467
rect 148726 83403 148778 83409
rect 148724 80466 148780 80475
rect 148724 80401 148780 80410
rect 148628 77950 148684 77959
rect 148628 77885 148684 77894
rect 148534 74729 148586 74735
rect 148534 74671 148586 74677
rect 148438 71991 148490 71997
rect 148438 71933 148490 71939
rect 148642 69111 148670 77885
rect 148738 71923 148766 80401
rect 148834 74883 148862 86469
rect 148930 80433 148958 92537
rect 149026 91903 149054 114441
rect 149122 94863 149150 116809
rect 149218 94937 149246 119325
rect 149314 97749 149342 121693
rect 149410 106333 149438 123344
rect 149506 120708 149534 123492
rect 149602 120911 149630 149813
rect 149698 123649 149726 150151
rect 151138 132381 151166 176717
rect 151234 155321 151262 216233
rect 151414 213331 151466 213337
rect 151414 213273 151466 213279
rect 151318 210371 151370 210377
rect 151318 210313 151370 210319
rect 151222 155315 151274 155321
rect 151222 155257 151274 155263
rect 151330 152657 151358 210313
rect 151426 155469 151454 213273
rect 151522 158281 151550 216825
rect 151702 212517 151754 212523
rect 151702 212459 151754 212465
rect 151606 207485 151658 207491
rect 151606 207427 151658 207433
rect 151510 158275 151562 158281
rect 151510 158217 151562 158223
rect 151414 155463 151466 155469
rect 151414 155405 151466 155411
rect 151318 152651 151370 152657
rect 151318 152593 151370 152599
rect 151618 152583 151646 207427
rect 151714 155395 151742 212459
rect 152578 192987 152606 270697
rect 153346 268837 153374 277870
rect 154006 271717 154058 271723
rect 154006 271659 154058 271665
rect 153334 268831 153386 268837
rect 153334 268773 153386 268779
rect 152566 192981 152618 192987
rect 152566 192923 152618 192929
rect 151798 190243 151850 190249
rect 151798 190185 151850 190191
rect 151702 155389 151754 155395
rect 151702 155331 151754 155337
rect 151606 152577 151658 152583
rect 151606 152519 151658 152525
rect 151702 148063 151754 148069
rect 151702 148005 151754 148011
rect 151222 147027 151274 147033
rect 151222 146969 151274 146975
rect 151126 132375 151178 132381
rect 151126 132317 151178 132323
rect 149686 123643 149738 123649
rect 149686 123585 149738 123591
rect 149590 120905 149642 120911
rect 149590 120847 149642 120853
rect 149506 120680 149726 120708
rect 149588 115690 149644 115699
rect 149588 115625 149644 115634
rect 149492 113174 149548 113183
rect 149492 113109 149548 113118
rect 149398 106327 149450 106333
rect 149398 106269 149450 106275
rect 149506 106204 149534 113109
rect 149410 106176 149534 106204
rect 149302 97743 149354 97749
rect 149302 97685 149354 97691
rect 149206 94931 149258 94937
rect 149206 94873 149258 94879
rect 149110 94857 149162 94863
rect 149110 94799 149162 94805
rect 149204 93786 149260 93795
rect 149204 93721 149260 93730
rect 149014 91897 149066 91903
rect 149014 91839 149066 91845
rect 149012 91418 149068 91427
rect 149012 91353 149068 91362
rect 148918 80427 148970 80433
rect 148918 80369 148970 80375
rect 149026 77769 149054 91353
rect 149108 90234 149164 90243
rect 149108 90169 149164 90178
rect 149014 77763 149066 77769
rect 149014 77705 149066 77711
rect 149122 77695 149150 90169
rect 149218 80655 149246 93721
rect 149410 91977 149438 106176
rect 149492 95710 149548 95719
rect 149492 95645 149548 95654
rect 149398 91971 149450 91977
rect 149398 91913 149450 91919
rect 149300 89050 149356 89059
rect 149300 88985 149356 88994
rect 149206 80649 149258 80655
rect 149206 80591 149258 80597
rect 149110 77689 149162 77695
rect 149110 77631 149162 77637
rect 149314 77547 149342 88985
rect 149396 87274 149452 87283
rect 149396 87209 149452 87218
rect 149410 77621 149438 87209
rect 149506 80581 149534 95645
rect 149602 94789 149630 115625
rect 149698 101024 149726 120680
rect 151234 118025 151262 146969
rect 151606 145843 151658 145849
rect 151606 145785 151658 145791
rect 151318 144363 151370 144369
rect 151318 144305 151370 144311
rect 151330 118099 151358 144305
rect 151510 141551 151562 141557
rect 151510 141493 151562 141499
rect 151414 141255 151466 141261
rect 151414 141197 151466 141203
rect 151318 118093 151370 118099
rect 151318 118035 151370 118041
rect 151222 118019 151274 118025
rect 151222 117961 151274 117967
rect 151426 115065 151454 141197
rect 151414 115059 151466 115065
rect 151414 115001 151466 115007
rect 151522 114991 151550 141493
rect 151618 117951 151646 145785
rect 151714 120763 151742 148005
rect 151810 140891 151838 190185
rect 154018 181295 154046 271659
rect 154498 270761 154526 277870
rect 155650 271797 155678 277870
rect 156898 272019 156926 277870
rect 158064 277856 158366 277884
rect 156886 272013 156938 272019
rect 156886 271955 156938 271961
rect 155638 271791 155690 271797
rect 155638 271733 155690 271739
rect 156886 271643 156938 271649
rect 156886 271585 156938 271591
rect 154486 270755 154538 270761
rect 154486 270697 154538 270703
rect 155446 270755 155498 270761
rect 155446 270697 155498 270703
rect 154102 193055 154154 193061
rect 154102 192997 154154 193003
rect 154006 181289 154058 181295
rect 154006 181231 154058 181237
rect 151894 142587 151946 142593
rect 151894 142529 151946 142535
rect 151798 140885 151850 140891
rect 151798 140827 151850 140833
rect 151702 120757 151754 120763
rect 151702 120699 151754 120705
rect 151606 117945 151658 117951
rect 151606 117887 151658 117893
rect 151906 117877 151934 142529
rect 154114 140817 154142 192997
rect 155458 192913 155486 270697
rect 155446 192907 155498 192913
rect 155446 192849 155498 192855
rect 156898 184181 156926 271585
rect 157078 247741 157130 247747
rect 157078 247683 157130 247689
rect 156982 244855 157034 244861
rect 156982 244797 157034 244803
rect 156886 184175 156938 184181
rect 156886 184117 156938 184123
rect 156886 179587 156938 179593
rect 156886 179529 156938 179535
rect 154198 178847 154250 178853
rect 154198 178789 154250 178795
rect 154102 140811 154154 140817
rect 154102 140753 154154 140759
rect 154210 132307 154238 178789
rect 154198 132301 154250 132307
rect 154198 132243 154250 132249
rect 156898 132233 156926 179529
rect 156994 175597 157022 244797
rect 157090 221773 157118 247683
rect 157078 221767 157130 221773
rect 157078 221709 157130 221715
rect 157078 194683 157130 194689
rect 157078 194625 157130 194631
rect 156982 175591 157034 175597
rect 156982 175533 157034 175539
rect 157090 143925 157118 194625
rect 158338 192839 158366 277856
rect 159298 268689 159326 277870
rect 159766 272087 159818 272093
rect 159766 272029 159818 272035
rect 159286 268683 159338 268689
rect 159286 268625 159338 268631
rect 158326 192833 158378 192839
rect 158326 192775 158378 192781
rect 159778 181221 159806 272029
rect 160450 268763 160478 277870
rect 161602 271649 161630 277870
rect 162646 271865 162698 271871
rect 162646 271807 162698 271813
rect 161590 271643 161642 271649
rect 161590 271585 161642 271591
rect 160438 268757 160490 268763
rect 160438 268699 160490 268705
rect 159862 234421 159914 234427
rect 159862 234363 159914 234369
rect 159766 181215 159818 181221
rect 159766 181157 159818 181163
rect 159874 166865 159902 234363
rect 159958 198827 160010 198833
rect 159958 198769 160010 198775
rect 159862 166859 159914 166865
rect 159862 166801 159914 166807
rect 159970 146811 159998 198769
rect 162658 184107 162686 271807
rect 162754 271797 162782 277870
rect 164002 272093 164030 277870
rect 163990 272087 164042 272093
rect 163990 272029 164042 272035
rect 162742 271791 162794 271797
rect 162742 271733 162794 271739
rect 164086 271643 164138 271649
rect 164086 271585 164138 271591
rect 162742 195941 162794 195947
rect 162742 195883 162794 195889
rect 162646 184101 162698 184107
rect 162646 184043 162698 184049
rect 162646 178625 162698 178631
rect 162646 178567 162698 178573
rect 159958 146805 160010 146811
rect 159958 146747 160010 146753
rect 157078 143919 157130 143925
rect 157078 143861 157130 143867
rect 162658 135193 162686 178567
rect 162754 143851 162782 195883
rect 164098 192765 164126 271585
rect 165154 270761 165182 277870
rect 165142 270755 165194 270761
rect 165142 270697 165194 270703
rect 166402 268615 166430 277870
rect 166966 270755 167018 270761
rect 166966 270697 167018 270703
rect 166390 268609 166442 268615
rect 166390 268551 166442 268557
rect 165526 218955 165578 218961
rect 165526 218897 165578 218903
rect 164086 192759 164138 192765
rect 164086 192701 164138 192707
rect 165538 158207 165566 218897
rect 166978 195799 167006 270697
rect 167554 268541 167582 277870
rect 168706 271945 168734 277870
rect 169858 272112 169886 277870
rect 169762 272084 169886 272112
rect 168694 271939 168746 271945
rect 168694 271881 168746 271887
rect 169762 271427 169790 272084
rect 169846 271939 169898 271945
rect 169846 271881 169898 271887
rect 169750 271421 169802 271427
rect 169750 271363 169802 271369
rect 167542 268535 167594 268541
rect 167542 268477 167594 268483
rect 168502 246927 168554 246933
rect 168502 246869 168554 246875
rect 168406 241969 168458 241975
rect 168406 241911 168458 241917
rect 166966 195793 167018 195799
rect 166966 195735 167018 195741
rect 165622 187283 165674 187289
rect 165622 187225 165674 187231
rect 165526 158201 165578 158207
rect 165526 158143 165578 158149
rect 162742 143845 162794 143851
rect 162742 143787 162794 143793
rect 165634 138153 165662 187225
rect 168418 172637 168446 241911
rect 168514 186993 168542 246869
rect 168598 204599 168650 204605
rect 168598 204541 168650 204547
rect 168502 186987 168554 186993
rect 168502 186929 168554 186935
rect 168406 172631 168458 172637
rect 168406 172573 168458 172579
rect 168610 149771 168638 204541
rect 169858 195725 169886 271881
rect 171010 271871 171038 277870
rect 172272 277856 172766 277884
rect 170998 271865 171050 271871
rect 170998 271807 171050 271813
rect 171286 195867 171338 195873
rect 171286 195809 171338 195815
rect 169846 195719 169898 195725
rect 169846 195661 169898 195667
rect 168694 184397 168746 184403
rect 168694 184339 168746 184345
rect 168598 149765 168650 149771
rect 168598 149707 168650 149713
rect 165622 138147 165674 138153
rect 165622 138089 165674 138095
rect 168706 138079 168734 184339
rect 171298 143777 171326 195809
rect 172738 195651 172766 277856
rect 173410 268467 173438 277870
rect 173398 268461 173450 268467
rect 173398 268403 173450 268409
rect 174658 268393 174686 277870
rect 175810 271131 175838 277870
rect 176962 271205 176990 277870
rect 178114 271723 178142 277870
rect 179362 271945 179390 277870
rect 179350 271939 179402 271945
rect 179350 271881 179402 271887
rect 178102 271717 178154 271723
rect 178102 271659 178154 271665
rect 176950 271199 177002 271205
rect 176950 271141 177002 271147
rect 175798 271125 175850 271131
rect 175798 271067 175850 271073
rect 178486 271125 178538 271131
rect 178486 271067 178538 271073
rect 177046 269793 177098 269799
rect 177046 269735 177098 269741
rect 174646 268387 174698 268393
rect 174646 268329 174698 268335
rect 177058 268319 177086 269735
rect 177046 268313 177098 268319
rect 177046 268255 177098 268261
rect 174166 239083 174218 239089
rect 174166 239025 174218 239031
rect 172726 195645 172778 195651
rect 172726 195587 172778 195593
rect 171382 181511 171434 181517
rect 171382 181453 171434 181459
rect 171286 143771 171338 143777
rect 171286 143713 171338 143719
rect 168694 138073 168746 138079
rect 168694 138015 168746 138021
rect 162646 135187 162698 135193
rect 162646 135129 162698 135135
rect 171394 135119 171422 181453
rect 174178 169677 174206 239025
rect 177046 207411 177098 207417
rect 177046 207353 177098 207359
rect 174262 204525 174314 204531
rect 174262 204467 174314 204473
rect 174166 169671 174218 169677
rect 174166 169613 174218 169619
rect 174274 149697 174302 204467
rect 174262 149691 174314 149697
rect 174262 149633 174314 149639
rect 177058 149549 177086 207353
rect 177142 198753 177194 198759
rect 177142 198695 177194 198701
rect 177046 149543 177098 149549
rect 177046 149485 177098 149491
rect 177154 146737 177182 198695
rect 178498 198611 178526 271067
rect 180514 268245 180542 277870
rect 181366 271939 181418 271945
rect 181366 271881 181418 271887
rect 180502 268239 180554 268245
rect 180502 268181 180554 268187
rect 179926 210297 179978 210303
rect 179926 210239 179978 210245
rect 178486 198605 178538 198611
rect 178486 198547 178538 198553
rect 179938 152509 179966 210239
rect 180022 201713 180074 201719
rect 180022 201655 180074 201661
rect 179926 152503 179978 152509
rect 179926 152445 179978 152451
rect 180034 149623 180062 201655
rect 181378 198685 181406 271881
rect 181762 271501 181790 277870
rect 182914 271945 182942 277870
rect 182902 271939 182954 271945
rect 182902 271881 182954 271887
rect 181750 271495 181802 271501
rect 181750 271437 181802 271443
rect 184162 268171 184190 277870
rect 184246 271939 184298 271945
rect 184246 271881 184298 271887
rect 184150 268165 184202 268171
rect 184150 268107 184202 268113
rect 182806 213183 182858 213189
rect 182806 213125 182858 213131
rect 181366 198679 181418 198685
rect 181366 198621 181418 198627
rect 180118 169967 180170 169973
rect 180118 169909 180170 169915
rect 180022 149617 180074 149623
rect 180022 149559 180074 149565
rect 177142 146731 177194 146737
rect 177142 146673 177194 146679
rect 171382 135113 171434 135119
rect 171382 135055 171434 135061
rect 156886 132227 156938 132233
rect 156886 132169 156938 132175
rect 180130 129347 180158 169909
rect 182818 154951 182846 213125
rect 182902 201639 182954 201645
rect 182902 201581 182954 201587
rect 182806 154945 182858 154951
rect 182806 154887 182858 154893
rect 182914 146885 182942 201581
rect 184258 197691 184286 271881
rect 185218 271353 185246 277870
rect 186370 271649 186398 277870
rect 185398 271643 185450 271649
rect 185398 271585 185450 271591
rect 186358 271643 186410 271649
rect 186358 271585 186410 271591
rect 185206 271347 185258 271353
rect 185206 271289 185258 271295
rect 185302 242857 185354 242863
rect 185302 242799 185354 242805
rect 184342 221767 184394 221773
rect 184342 221709 184394 221715
rect 184354 219595 184382 221709
rect 185314 221075 185342 242799
rect 185300 221066 185356 221075
rect 185300 221001 185356 221010
rect 184340 219586 184396 219595
rect 184340 219521 184396 219530
rect 184342 201565 184394 201571
rect 184342 201507 184394 201513
rect 184354 199763 184382 201507
rect 184340 199754 184396 199763
rect 184340 199689 184396 199698
rect 184342 198679 184394 198685
rect 184342 198621 184394 198627
rect 184244 197682 184300 197691
rect 184244 197617 184300 197626
rect 184354 196803 184382 198621
rect 184438 198605 184490 198611
rect 184438 198547 184490 198553
rect 184340 196794 184396 196803
rect 184340 196729 184396 196738
rect 184450 196063 184478 198547
rect 185410 198283 185438 271585
rect 187618 271057 187646 277870
rect 188770 271131 188798 277870
rect 189730 277856 190032 277884
rect 188758 271125 188810 271131
rect 188758 271067 188810 271073
rect 187606 271051 187658 271057
rect 187606 270993 187658 270999
rect 189730 266395 189758 277856
rect 191170 271871 191198 277870
rect 191158 271865 191210 271871
rect 191158 271807 191210 271813
rect 192322 271575 192350 277870
rect 193076 272274 193132 272283
rect 193076 272209 193132 272218
rect 192982 271791 193034 271797
rect 192982 271733 193034 271739
rect 192310 271569 192362 271575
rect 192310 271511 192362 271517
rect 192596 269462 192652 269471
rect 192596 269397 192652 269406
rect 192404 269314 192460 269323
rect 192404 269249 192460 269258
rect 187222 266389 187274 266395
rect 187222 266331 187274 266337
rect 189718 266389 189770 266395
rect 189718 266331 189770 266337
rect 186838 249443 186890 249449
rect 186838 249385 186890 249391
rect 186742 249369 186794 249375
rect 186742 249311 186794 249317
rect 186454 249147 186506 249153
rect 186454 249089 186506 249095
rect 186166 246631 186218 246637
rect 186166 246573 186218 246579
rect 186070 246483 186122 246489
rect 186070 246425 186122 246431
rect 185878 246261 185930 246267
rect 185878 246203 185930 246209
rect 185590 243375 185642 243381
rect 185590 243317 185642 243323
rect 185494 242709 185546 242715
rect 185494 242651 185546 242657
rect 185506 220335 185534 242651
rect 185492 220326 185548 220335
rect 185492 220261 185548 220270
rect 185602 218855 185630 243317
rect 185782 242635 185834 242641
rect 185782 242577 185834 242583
rect 185686 224727 185738 224733
rect 185686 224669 185738 224675
rect 185588 218846 185644 218855
rect 185588 218781 185644 218790
rect 185396 198274 185452 198283
rect 185396 198209 185452 198218
rect 184436 196054 184492 196063
rect 184436 195989 184492 195998
rect 184534 195793 184586 195799
rect 184534 195735 184586 195741
rect 184438 195719 184490 195725
rect 184438 195661 184490 195667
rect 184342 195645 184394 195651
rect 184342 195587 184394 195593
rect 184354 195323 184382 195587
rect 184340 195314 184396 195323
rect 184340 195249 184396 195258
rect 184450 194435 184478 195661
rect 184436 194426 184492 194435
rect 184436 194361 184492 194370
rect 184546 193843 184574 195735
rect 184532 193834 184588 193843
rect 184532 193769 184588 193778
rect 184630 192981 184682 192987
rect 184436 192946 184492 192955
rect 184630 192923 184682 192929
rect 184436 192881 184492 192890
rect 184534 192907 184586 192913
rect 184342 192833 184394 192839
rect 184342 192775 184394 192781
rect 184354 192363 184382 192775
rect 184450 192765 184478 192881
rect 184534 192849 184586 192855
rect 184438 192759 184490 192765
rect 184438 192701 184490 192707
rect 184340 192354 184396 192363
rect 184340 192289 184396 192298
rect 184546 191475 184574 192849
rect 184532 191466 184588 191475
rect 184532 191401 184588 191410
rect 184642 190735 184670 192923
rect 184628 190726 184684 190735
rect 184628 190661 184684 190670
rect 184630 190095 184682 190101
rect 184630 190037 184682 190043
rect 184534 190021 184586 190027
rect 184340 189986 184396 189995
rect 184534 189963 184586 189969
rect 184340 189921 184396 189930
rect 184438 189947 184490 189953
rect 184354 189879 184382 189921
rect 184438 189889 184490 189895
rect 184342 189873 184394 189879
rect 184342 189815 184394 189821
rect 184450 189255 184478 189889
rect 184436 189246 184492 189255
rect 184436 189181 184492 189190
rect 184546 188515 184574 189963
rect 184532 188506 184588 188515
rect 184532 188441 184588 188450
rect 184642 187627 184670 190037
rect 184628 187618 184684 187627
rect 184628 187553 184684 187562
rect 184438 187209 184490 187215
rect 184438 187151 184490 187157
rect 184342 187061 184394 187067
rect 184342 187003 184394 187009
rect 184354 186147 184382 187003
rect 184450 186887 184478 187151
rect 184630 187135 184682 187141
rect 184630 187077 184682 187083
rect 184534 186987 184586 186993
rect 184534 186929 184586 186935
rect 184436 186878 184492 186887
rect 184436 186813 184492 186822
rect 184340 186138 184396 186147
rect 184340 186073 184396 186082
rect 184546 184667 184574 186929
rect 184642 185407 184670 187077
rect 184628 185398 184684 185407
rect 184628 185333 184684 185342
rect 184532 184658 184588 184667
rect 184532 184593 184588 184602
rect 184534 184323 184586 184329
rect 184534 184265 184586 184271
rect 184342 184249 184394 184255
rect 184342 184191 184394 184197
rect 184354 183927 184382 184191
rect 184438 184101 184490 184107
rect 184438 184043 184490 184049
rect 184340 183918 184396 183927
rect 184340 183853 184396 183862
rect 184450 182447 184478 184043
rect 184546 183187 184574 184265
rect 184630 184175 184682 184181
rect 184630 184117 184682 184123
rect 184532 183178 184588 183187
rect 184532 183113 184588 183122
rect 184436 182438 184492 182447
rect 184436 182373 184492 182382
rect 184642 181559 184670 184117
rect 184628 181550 184684 181559
rect 184628 181485 184684 181494
rect 184630 181437 184682 181443
rect 184630 181379 184682 181385
rect 184534 181363 184586 181369
rect 184534 181305 184586 181311
rect 184342 181289 184394 181295
rect 184342 181231 184394 181237
rect 184354 180819 184382 181231
rect 184438 181215 184490 181221
rect 184438 181157 184490 181163
rect 184340 180810 184396 180819
rect 184340 180745 184396 180754
rect 184450 180079 184478 181157
rect 184436 180070 184492 180079
rect 184436 180005 184492 180014
rect 184546 179339 184574 181305
rect 184532 179330 184588 179339
rect 184532 179265 184588 179274
rect 184642 178599 184670 181379
rect 184628 178590 184684 178599
rect 184438 178551 184490 178557
rect 184628 178525 184684 178534
rect 184438 178493 184490 178499
rect 184342 178403 184394 178409
rect 184342 178345 184394 178351
rect 184354 177711 184382 178345
rect 184340 177702 184396 177711
rect 184340 177637 184396 177646
rect 184450 177119 184478 178493
rect 184534 178477 184586 178483
rect 184534 178419 184586 178425
rect 184436 177110 184492 177119
rect 184436 177045 184492 177054
rect 184546 176231 184574 178419
rect 184532 176222 184588 176231
rect 184532 176157 184588 176166
rect 184342 175665 184394 175671
rect 184340 175630 184342 175639
rect 184394 175630 184396 175639
rect 184340 175565 184396 175574
rect 184438 175591 184490 175597
rect 184438 175533 184490 175539
rect 184450 174011 184478 175533
rect 184436 174002 184492 174011
rect 184436 173937 184492 173946
rect 184438 172779 184490 172785
rect 184438 172721 184490 172727
rect 184342 172631 184394 172637
rect 184342 172573 184394 172579
rect 184354 172531 184382 172573
rect 184340 172522 184396 172531
rect 184340 172457 184396 172466
rect 184450 170903 184478 172721
rect 184534 172705 184586 172711
rect 184534 172647 184586 172653
rect 184436 170894 184492 170903
rect 184436 170829 184492 170838
rect 184546 170311 184574 172647
rect 184532 170302 184588 170311
rect 184532 170237 184588 170246
rect 184438 169893 184490 169899
rect 184438 169835 184490 169841
rect 184342 169671 184394 169677
rect 184342 169613 184394 169619
rect 184354 169423 184382 169613
rect 184340 169414 184396 169423
rect 184340 169349 184396 169358
rect 184450 168683 184478 169835
rect 184534 169819 184586 169825
rect 184534 169761 184586 169767
rect 184436 168674 184492 168683
rect 184436 168609 184492 168618
rect 184546 167943 184574 169761
rect 184630 169745 184682 169751
rect 184630 169687 184682 169693
rect 184532 167934 184588 167943
rect 184532 167869 184588 167878
rect 184642 167203 184670 169687
rect 184628 167194 184684 167203
rect 184628 167129 184684 167138
rect 182998 167081 183050 167087
rect 182998 167023 183050 167029
rect 182902 146879 182954 146885
rect 182902 146821 182954 146827
rect 180118 129341 180170 129347
rect 180118 129283 180170 129289
rect 183010 126535 183038 167023
rect 184438 167007 184490 167013
rect 184438 166949 184490 166955
rect 184342 166859 184394 166865
rect 184342 166801 184394 166807
rect 184354 166463 184382 166801
rect 184340 166454 184396 166463
rect 184340 166389 184396 166398
rect 184450 165723 184478 166949
rect 184534 166933 184586 166939
rect 184534 166875 184586 166881
rect 184436 165714 184492 165723
rect 184436 165649 184492 165658
rect 184546 164835 184574 166875
rect 184532 164826 184588 164835
rect 184532 164761 184588 164770
rect 184342 164121 184394 164127
rect 184340 164086 184342 164095
rect 184394 164086 184396 164095
rect 184340 164021 184396 164030
rect 184534 164047 184586 164053
rect 184534 163989 184586 163995
rect 184438 163973 184490 163979
rect 184438 163915 184490 163921
rect 184342 163899 184394 163905
rect 184342 163841 184394 163847
rect 184354 163355 184382 163841
rect 184340 163346 184396 163355
rect 184340 163281 184396 163290
rect 184450 162615 184478 163915
rect 184436 162606 184492 162615
rect 184436 162541 184492 162550
rect 184546 161875 184574 163989
rect 184532 161866 184588 161875
rect 184532 161801 184588 161810
rect 184630 161235 184682 161241
rect 184630 161177 184682 161183
rect 184342 161161 184394 161167
rect 184342 161103 184394 161109
rect 184354 160987 184382 161103
rect 184438 161087 184490 161093
rect 184438 161029 184490 161035
rect 184340 160978 184396 160987
rect 184340 160913 184396 160922
rect 184450 160395 184478 161029
rect 184534 161013 184586 161019
rect 184534 160955 184586 160961
rect 184436 160386 184492 160395
rect 184436 160321 184492 160330
rect 184546 159507 184574 160955
rect 184532 159498 184588 159507
rect 184532 159433 184588 159442
rect 184642 158915 184670 161177
rect 184628 158906 184684 158915
rect 184628 158841 184684 158850
rect 184438 158423 184490 158429
rect 184438 158365 184490 158371
rect 184342 158201 184394 158207
rect 184342 158143 184394 158149
rect 184354 156547 184382 158143
rect 184450 158027 184478 158365
rect 184534 158349 184586 158355
rect 184534 158291 184586 158297
rect 184436 158018 184492 158027
rect 184436 157953 184492 157962
rect 184546 157435 184574 158291
rect 184630 158275 184682 158281
rect 184630 158217 184682 158223
rect 184532 157426 184588 157435
rect 184532 157361 184588 157370
rect 184340 156538 184396 156547
rect 184340 156473 184396 156482
rect 184642 155659 184670 158217
rect 184628 155650 184684 155659
rect 184628 155585 184684 155594
rect 184438 155463 184490 155469
rect 184438 155405 184490 155411
rect 184342 155315 184394 155321
rect 184342 155257 184394 155263
rect 184354 155067 184382 155257
rect 184340 155058 184396 155067
rect 184340 154993 184396 155002
rect 184450 154179 184478 155405
rect 184534 155389 184586 155395
rect 184534 155331 184586 155337
rect 184436 154170 184492 154179
rect 184436 154105 184492 154114
rect 184546 152699 184574 155331
rect 184726 154945 184778 154951
rect 184726 154887 184778 154893
rect 184738 153587 184766 154887
rect 184724 153578 184780 153587
rect 184724 153513 184780 153522
rect 184532 152690 184588 152699
rect 184342 152651 184394 152657
rect 184532 152625 184588 152634
rect 184342 152593 184394 152599
rect 184354 151959 184382 152593
rect 184438 152577 184490 152583
rect 184438 152519 184490 152525
rect 184340 151950 184396 151959
rect 184340 151885 184396 151894
rect 184450 150479 184478 152519
rect 184534 152503 184586 152509
rect 184534 152445 184586 152451
rect 184546 151219 184574 152445
rect 184532 151210 184588 151219
rect 184532 151145 184588 151154
rect 184436 150470 184492 150479
rect 184436 150405 184492 150414
rect 184438 149765 184490 149771
rect 184438 149707 184490 149713
rect 184628 149730 184684 149739
rect 184342 149691 184394 149697
rect 184342 149633 184394 149639
rect 184354 148999 184382 149633
rect 184340 148990 184396 148999
rect 184340 148925 184396 148934
rect 184450 148111 184478 149707
rect 184628 149665 184684 149674
rect 184534 149617 184586 149623
rect 184534 149559 184586 149565
rect 184436 148102 184492 148111
rect 184436 148037 184492 148046
rect 184546 147371 184574 149559
rect 184642 149549 184670 149665
rect 184630 149543 184682 149549
rect 184630 149485 184682 149491
rect 184532 147362 184588 147371
rect 184532 147297 184588 147306
rect 184438 146805 184490 146811
rect 184438 146747 184490 146753
rect 184342 146657 184394 146663
rect 184342 146599 184394 146605
rect 184354 145891 184382 146599
rect 184340 145882 184396 145891
rect 184340 145817 184396 145826
rect 184450 144411 184478 146747
rect 184534 146731 184586 146737
rect 184534 146673 184586 146679
rect 184546 145151 184574 146673
rect 184532 145142 184588 145151
rect 184532 145077 184588 145086
rect 184436 144402 184492 144411
rect 184436 144337 184492 144346
rect 184438 143993 184490 143999
rect 184438 143935 184490 143941
rect 184342 143771 184394 143777
rect 184342 143713 184394 143719
rect 184354 142783 184382 143713
rect 184450 143671 184478 143935
rect 184630 143919 184682 143925
rect 184630 143861 184682 143867
rect 184534 143845 184586 143851
rect 184534 143787 184586 143793
rect 184436 143662 184492 143671
rect 184436 143597 184492 143606
rect 184340 142774 184396 142783
rect 184340 142709 184396 142718
rect 184546 142191 184574 143787
rect 184532 142182 184588 142191
rect 184532 142117 184588 142126
rect 184642 141303 184670 143861
rect 184628 141294 184684 141303
rect 184628 141229 184684 141238
rect 184534 141107 184586 141113
rect 184534 141049 184586 141055
rect 184438 140885 184490 140891
rect 184438 140827 184490 140833
rect 184342 140811 184394 140817
rect 184342 140753 184394 140759
rect 184354 140563 184382 140753
rect 184340 140554 184396 140563
rect 184340 140489 184396 140498
rect 184450 138935 184478 140827
rect 184546 139823 184574 141049
rect 184630 141033 184682 141039
rect 184630 140975 184682 140981
rect 184532 139814 184588 139823
rect 184532 139749 184588 139758
rect 184436 138926 184492 138935
rect 184436 138861 184492 138870
rect 184642 138343 184670 140975
rect 185698 140965 185726 224669
rect 185794 173271 185822 242577
rect 185890 201391 185918 246203
rect 185974 242783 186026 242789
rect 185974 242725 186026 242731
rect 185876 201382 185932 201391
rect 185876 201317 185932 201326
rect 185986 195854 186014 242725
rect 186082 202871 186110 246425
rect 186178 207311 186206 246573
rect 186358 246409 186410 246415
rect 186358 246351 186410 246357
rect 186262 246335 186314 246341
rect 186262 246277 186314 246283
rect 186164 207302 186220 207311
rect 186164 207237 186220 207246
rect 186274 204351 186302 246277
rect 186370 205239 186398 246351
rect 186466 212047 186494 249089
rect 186646 246705 186698 246711
rect 186646 246647 186698 246653
rect 186550 246557 186602 246563
rect 186550 246499 186602 246505
rect 186452 212038 186508 212047
rect 186452 211973 186508 211982
rect 186562 209087 186590 246499
rect 186658 210567 186686 246647
rect 186754 213527 186782 249311
rect 186850 218115 186878 249385
rect 186934 249295 186986 249301
rect 186934 249237 186986 249243
rect 186836 218106 186892 218115
rect 186836 218041 186892 218050
rect 186946 215007 186974 249237
rect 187030 249221 187082 249227
rect 187030 249163 187082 249169
rect 187042 216487 187070 249163
rect 187124 243414 187180 243423
rect 187124 243349 187180 243358
rect 187138 224733 187166 243349
rect 187126 224727 187178 224733
rect 187126 224669 187178 224675
rect 187028 216478 187084 216487
rect 187028 216413 187084 216422
rect 186932 214998 186988 215007
rect 186932 214933 186988 214942
rect 186740 213518 186796 213527
rect 186740 213453 186796 213462
rect 186644 210558 186700 210567
rect 186644 210493 186700 210502
rect 186548 209078 186604 209087
rect 186548 209013 186604 209022
rect 186356 205230 186412 205239
rect 186356 205165 186412 205174
rect 186260 204342 186316 204351
rect 186260 204277 186316 204286
rect 186068 202862 186124 202871
rect 186068 202797 186124 202806
rect 187234 199171 187262 266331
rect 192418 263810 192446 269249
rect 192610 263824 192638 269397
rect 192994 268097 193022 271733
rect 192982 268091 193034 268097
rect 192982 268033 193034 268039
rect 193090 263824 193118 272209
rect 193174 271643 193226 271649
rect 193174 271585 193226 271591
rect 193186 268023 193214 271585
rect 193474 271279 193502 277870
rect 194722 272167 194750 277870
rect 194422 272161 194474 272167
rect 194228 272126 194284 272135
rect 194422 272103 194474 272109
rect 194710 272161 194762 272167
rect 194710 272103 194762 272109
rect 194228 272061 194284 272070
rect 193462 271273 193514 271279
rect 193462 271215 193514 271221
rect 193748 269610 193804 269619
rect 193748 269545 193804 269554
rect 193174 268017 193226 268023
rect 193174 267959 193226 267965
rect 192610 263796 192864 263824
rect 193090 263796 193344 263824
rect 193762 263810 193790 269545
rect 194242 263810 194270 272061
rect 194434 263824 194462 272103
rect 195874 271797 195902 277870
rect 196822 272309 196874 272315
rect 196822 272251 196874 272257
rect 195862 271791 195914 271797
rect 195862 271733 195914 271739
rect 195670 269497 195722 269503
rect 195670 269439 195722 269445
rect 194998 269349 195050 269355
rect 194998 269291 195050 269297
rect 195010 263824 195038 269291
rect 194434 263796 194736 263824
rect 195010 263796 195264 263824
rect 195682 263810 195710 269439
rect 196630 269423 196682 269429
rect 196630 269365 196682 269371
rect 196150 269275 196202 269281
rect 196150 269217 196202 269223
rect 196162 263810 196190 269217
rect 196642 263810 196670 269365
rect 196834 263824 196862 272251
rect 197122 269281 197150 277870
rect 197398 272235 197450 272241
rect 197398 272177 197450 272183
rect 197110 269275 197162 269281
rect 197110 269217 197162 269223
rect 197410 263824 197438 272177
rect 198274 270983 198302 277870
rect 199030 272383 199082 272389
rect 199030 272325 199082 272331
rect 198646 271421 198698 271427
rect 198646 271363 198698 271369
rect 198262 270977 198314 270983
rect 198262 270919 198314 270925
rect 198658 269651 198686 271363
rect 198550 269645 198602 269651
rect 198550 269587 198602 269593
rect 198646 269645 198698 269651
rect 198646 269587 198698 269593
rect 198070 269571 198122 269577
rect 198070 269513 198122 269519
rect 196834 263796 197088 263824
rect 197410 263796 197664 263824
rect 198082 263810 198110 269513
rect 198562 263810 198590 269587
rect 199042 263810 199070 272325
rect 199522 271427 199550 277870
rect 199702 272457 199754 272463
rect 199702 272399 199754 272405
rect 199510 271421 199562 271427
rect 199510 271363 199562 271369
rect 199222 269719 199274 269725
rect 199222 269661 199274 269667
rect 199234 263824 199262 269661
rect 199714 263824 199742 272399
rect 200578 269355 200606 277870
rect 201142 272679 201194 272685
rect 201142 272621 201194 272627
rect 200950 272531 201002 272537
rect 200950 272473 201002 272479
rect 200566 269349 200618 269355
rect 200566 269291 200618 269297
rect 200470 268313 200522 268319
rect 200470 268255 200522 268261
rect 199234 263796 199488 263824
rect 199714 263796 199968 263824
rect 200482 263810 200510 268255
rect 200962 263810 200990 272473
rect 201154 263824 201182 272621
rect 201826 271649 201854 277870
rect 202870 272605 202922 272611
rect 202870 272547 202922 272553
rect 201814 271643 201866 271649
rect 201814 271585 201866 271591
rect 202294 269941 202346 269947
rect 202294 269883 202346 269889
rect 201622 269867 201674 269873
rect 201622 269809 201674 269815
rect 201634 263824 201662 269809
rect 201154 263796 201408 263824
rect 201634 263796 201888 263824
rect 202306 263810 202334 269883
rect 202882 263810 202910 272547
rect 202978 269429 203006 277870
rect 203350 272753 203402 272759
rect 203350 272695 203402 272701
rect 202966 269423 203018 269429
rect 202966 269365 203018 269371
rect 203362 263810 203390 272695
rect 204022 271199 204074 271205
rect 204022 271141 204074 271147
rect 203542 270089 203594 270095
rect 203542 270031 203594 270037
rect 203554 263824 203582 270031
rect 204034 269799 204062 271141
rect 204022 269793 204074 269799
rect 204022 269735 204074 269741
rect 204130 269503 204158 277870
rect 205270 272901 205322 272907
rect 205270 272843 205322 272849
rect 204694 272827 204746 272833
rect 204694 272769 204746 272775
rect 204214 270015 204266 270021
rect 204214 269957 204266 269963
rect 204118 269497 204170 269503
rect 204118 269439 204170 269445
rect 204226 263824 204254 269957
rect 203554 263796 203808 263824
rect 204226 263796 204288 263824
rect 204706 263810 204734 272769
rect 205282 263810 205310 272843
rect 205378 271205 205406 277870
rect 205942 273049 205994 273055
rect 205942 272991 205994 272997
rect 205366 271199 205418 271205
rect 205366 271141 205418 271147
rect 205846 271051 205898 271057
rect 205846 270993 205898 270999
rect 205750 270163 205802 270169
rect 205750 270105 205802 270111
rect 205366 268313 205418 268319
rect 205366 268255 205418 268261
rect 205378 268171 205406 268255
rect 205474 268245 205694 268264
rect 205462 268239 205706 268245
rect 205514 268236 205654 268239
rect 205462 268181 205514 268187
rect 205654 268181 205706 268187
rect 205366 268165 205418 268171
rect 205366 268107 205418 268113
rect 205762 263810 205790 270105
rect 205858 269725 205886 270993
rect 205846 269719 205898 269725
rect 205846 269661 205898 269667
rect 205954 263824 205982 272991
rect 206422 270237 206474 270243
rect 206422 270179 206474 270185
rect 206434 263824 206462 270179
rect 206530 269577 206558 277870
rect 207670 273567 207722 273573
rect 207670 273509 207722 273515
rect 207286 273419 207338 273425
rect 207286 273361 207338 273367
rect 206998 273345 207050 273351
rect 206998 273287 207050 273293
rect 206518 269571 206570 269577
rect 206518 269513 206570 269519
rect 207010 267991 207038 273287
rect 207094 273123 207146 273129
rect 207094 273065 207146 273071
rect 206996 267982 207052 267991
rect 206996 267917 207052 267926
rect 205954 263796 206208 263824
rect 206434 263796 206688 263824
rect 207106 263810 207134 273065
rect 207298 268097 207326 273361
rect 207478 271939 207530 271945
rect 207478 271881 207530 271887
rect 207382 271717 207434 271723
rect 207382 271659 207434 271665
rect 207394 270169 207422 271659
rect 207382 270163 207434 270169
rect 207382 270105 207434 270111
rect 207490 269947 207518 271881
rect 207682 270317 207710 273509
rect 207778 272389 207806 277870
rect 207958 272975 208010 272981
rect 207958 272917 208010 272923
rect 207766 272383 207818 272389
rect 207766 272325 207818 272331
rect 207862 272087 207914 272093
rect 207862 272029 207914 272035
rect 207766 272013 207818 272019
rect 207766 271955 207818 271961
rect 207574 270311 207626 270317
rect 207574 270253 207626 270259
rect 207670 270311 207722 270317
rect 207670 270253 207722 270259
rect 207478 269941 207530 269947
rect 207478 269883 207530 269889
rect 207286 268091 207338 268097
rect 207286 268033 207338 268039
rect 207586 263810 207614 270253
rect 207778 267875 207806 271955
rect 207874 267949 207902 272029
rect 207862 267943 207914 267949
rect 207862 267885 207914 267891
rect 207766 267869 207818 267875
rect 207766 267811 207818 267817
rect 207970 263824 207998 272917
rect 208834 272537 208862 277870
rect 209974 273271 210026 273277
rect 209974 273213 210026 273219
rect 209014 273197 209066 273203
rect 209014 273139 209066 273145
rect 208822 272531 208874 272537
rect 208822 272473 208874 272479
rect 208342 270385 208394 270391
rect 208342 270327 208394 270333
rect 208354 263824 208382 270327
rect 207970 263796 208128 263824
rect 208354 263796 208608 263824
rect 209026 263810 209054 273139
rect 209494 270459 209546 270465
rect 209494 270401 209546 270407
rect 209506 263810 209534 270401
rect 209986 263810 210014 273213
rect 210082 272315 210110 277870
rect 210166 273493 210218 273499
rect 210166 273435 210218 273441
rect 210070 272309 210122 272315
rect 210070 272251 210122 272257
rect 210178 270243 210206 273435
rect 211234 271945 211262 277870
rect 212482 272611 212510 277870
rect 213634 272833 213662 277870
rect 214882 272907 214910 277870
rect 214870 272901 214922 272907
rect 214870 272843 214922 272849
rect 213622 272827 213674 272833
rect 213622 272769 213674 272775
rect 215938 272759 215966 277870
rect 217186 273129 217214 277870
rect 217174 273123 217226 273129
rect 217174 273065 217226 273071
rect 218338 273055 218366 277870
rect 219586 273277 219614 277870
rect 219574 273271 219626 273277
rect 219574 273213 219626 273219
rect 218326 273049 218378 273055
rect 218326 272991 218378 272997
rect 220738 272981 220766 277870
rect 220726 272975 220778 272981
rect 220726 272917 220778 272923
rect 215926 272753 215978 272759
rect 215926 272695 215978 272701
rect 212470 272605 212522 272611
rect 212470 272547 212522 272553
rect 211222 271939 211274 271945
rect 211222 271881 211274 271887
rect 221590 271791 221642 271797
rect 221590 271733 221642 271739
rect 210454 271495 210506 271501
rect 210454 271437 210506 271443
rect 210358 271347 210410 271353
rect 210358 271289 210410 271295
rect 210262 271125 210314 271131
rect 210262 271067 210314 271073
rect 210166 270237 210218 270243
rect 210166 270179 210218 270185
rect 210274 269873 210302 271067
rect 210370 270021 210398 271289
rect 210466 270095 210494 271437
rect 221494 271421 221546 271427
rect 221494 271363 221546 271369
rect 214294 270681 214346 270687
rect 214294 270623 214346 270629
rect 212662 270607 212714 270613
rect 212662 270549 212714 270555
rect 211894 270533 211946 270539
rect 211894 270475 211946 270481
rect 210454 270089 210506 270095
rect 210454 270031 210506 270037
rect 210358 270015 210410 270021
rect 210358 269957 210410 269963
rect 210740 269906 210796 269915
rect 210262 269867 210314 269873
rect 210740 269841 210796 269850
rect 210262 269809 210314 269815
rect 210260 269758 210316 269767
rect 210260 269693 210316 269702
rect 210274 263824 210302 269693
rect 210754 263824 210782 269841
rect 211412 267982 211468 267991
rect 211412 267917 211468 267926
rect 210274 263796 210528 263824
rect 210754 263796 211008 263824
rect 211426 263810 211454 267917
rect 211906 263810 211934 270475
rect 212374 269201 212426 269207
rect 212374 269143 212426 269149
rect 212386 263810 212414 269143
rect 212674 263824 212702 270549
rect 213814 269127 213866 269133
rect 213814 269069 213866 269075
rect 213334 268091 213386 268097
rect 213334 268033 213386 268039
rect 212674 263796 212928 263824
rect 213346 263810 213374 268033
rect 213826 263810 213854 269069
rect 214306 263810 214334 270623
rect 216214 270311 216266 270317
rect 216214 270253 216266 270259
rect 214966 270237 215018 270243
rect 214966 270179 215018 270185
rect 214486 269053 214538 269059
rect 214486 268995 214538 269001
rect 214498 263824 214526 268995
rect 214978 263824 215006 270179
rect 215734 268979 215786 268985
rect 215734 268921 215786 268927
rect 214498 263796 214752 263824
rect 214978 263796 215232 263824
rect 215746 263810 215774 268921
rect 216226 263810 216254 270253
rect 221206 269645 221258 269651
rect 221206 269587 221258 269593
rect 216694 268905 216746 268911
rect 216694 268847 216746 268853
rect 216706 263810 216734 268847
rect 216886 268831 216938 268837
rect 216886 268773 216938 268779
rect 216898 263824 216926 268773
rect 218902 268757 218954 268763
rect 218902 268699 218954 268705
rect 218614 268683 218666 268689
rect 218614 268625 218666 268631
rect 217366 268017 217418 268023
rect 217366 267959 217418 267965
rect 217378 263824 217406 267959
rect 218134 267869 218186 267875
rect 218134 267811 218186 267817
rect 216898 263796 217152 263824
rect 217378 263796 217632 263824
rect 218146 263810 218174 267811
rect 218626 263810 218654 268625
rect 218914 263824 218942 268699
rect 220534 268609 220586 268615
rect 220534 268551 220586 268557
rect 219286 268165 219338 268171
rect 219286 268107 219338 268113
rect 219298 263824 219326 268107
rect 219958 267943 220010 267949
rect 219958 267885 220010 267891
rect 218914 263796 219072 263824
rect 219298 263796 219552 263824
rect 219970 263810 219998 267885
rect 220546 263810 220574 268551
rect 221014 268535 221066 268541
rect 221014 268477 221066 268483
rect 221026 263810 221054 268477
rect 221218 263824 221246 269587
rect 221506 268097 221534 271363
rect 221494 268091 221546 268097
rect 221494 268033 221546 268039
rect 221602 268023 221630 271733
rect 221686 271273 221738 271279
rect 221686 271215 221738 271221
rect 221590 268017 221642 268023
rect 221590 267959 221642 267965
rect 221698 267875 221726 271215
rect 221890 271057 221918 277870
rect 221974 271569 222026 271575
rect 221974 271511 222026 271517
rect 221878 271051 221930 271057
rect 221878 270993 221930 270999
rect 221782 269941 221834 269947
rect 221782 269883 221834 269889
rect 221686 267869 221738 267875
rect 221686 267811 221738 267817
rect 221794 263824 221822 269883
rect 221986 267949 222014 271511
rect 223138 270983 223166 277870
rect 223126 270977 223178 270983
rect 223126 270919 223178 270925
rect 224194 270909 224222 277870
rect 224566 272161 224618 272167
rect 224566 272103 224618 272109
rect 224278 271643 224330 271649
rect 224278 271585 224330 271591
rect 224182 270903 224234 270909
rect 224182 270845 224234 270851
rect 223606 270163 223658 270169
rect 223606 270105 223658 270111
rect 223414 269793 223466 269799
rect 223414 269735 223466 269741
rect 222358 268461 222410 268467
rect 222358 268403 222410 268409
rect 221974 267943 222026 267949
rect 221974 267885 222026 267891
rect 221218 263796 221472 263824
rect 221794 263796 221952 263824
rect 222370 263810 222398 268403
rect 222838 268387 222890 268393
rect 222838 268329 222890 268335
rect 222850 263810 222878 268329
rect 223426 263810 223454 269735
rect 223618 263824 223646 270105
rect 224290 268245 224318 271585
rect 224086 268239 224138 268245
rect 224086 268181 224138 268187
rect 224278 268239 224330 268245
rect 224278 268181 224330 268187
rect 224098 263824 224126 268181
rect 224578 268171 224606 272103
rect 225442 270835 225470 277870
rect 225430 270829 225482 270835
rect 225430 270771 225482 270777
rect 226594 270761 226622 277870
rect 227842 272167 227870 277870
rect 228994 272241 229022 277870
rect 228982 272235 229034 272241
rect 228982 272177 229034 272183
rect 227830 272161 227882 272167
rect 227830 272103 227882 272109
rect 230242 272093 230270 277870
rect 230230 272087 230282 272093
rect 230230 272029 230282 272035
rect 231394 272019 231422 277870
rect 232546 272463 232574 277870
rect 233698 272685 233726 277870
rect 233686 272679 233738 272685
rect 233686 272621 233738 272627
rect 234358 272531 234410 272537
rect 234358 272473 234410 272479
rect 232534 272457 232586 272463
rect 232534 272399 232586 272405
rect 233878 272383 233930 272389
rect 233878 272325 233930 272331
rect 231382 272013 231434 272019
rect 231382 271955 231434 271961
rect 227158 271865 227210 271871
rect 227158 271807 227210 271813
rect 226582 270755 226634 270761
rect 226582 270697 226634 270703
rect 224758 270089 224810 270095
rect 224758 270031 224810 270037
rect 224566 268165 224618 268171
rect 224566 268107 224618 268113
rect 223618 263796 223872 263824
rect 224098 263796 224352 263824
rect 224770 263810 224798 270031
rect 225526 270015 225578 270021
rect 225526 269957 225578 269963
rect 225238 268313 225290 268319
rect 225238 268255 225290 268261
rect 225250 263810 225278 268255
rect 225538 263824 225566 269957
rect 226678 269867 226730 269873
rect 226678 269809 226730 269815
rect 226006 269719 226058 269725
rect 226006 269661 226058 269667
rect 226018 263824 226046 269661
rect 225538 263796 225792 263824
rect 226018 263796 226272 263824
rect 226690 263810 226718 269809
rect 227170 263810 227198 271807
rect 232630 271199 232682 271205
rect 232630 271141 232682 271147
rect 230038 270681 230090 270687
rect 230038 270623 230090 270629
rect 229558 269275 229610 269281
rect 229558 269217 229610 269223
rect 228406 268165 228458 268171
rect 228406 268107 228458 268113
rect 227638 267943 227690 267949
rect 227638 267885 227690 267891
rect 227650 263810 227678 267885
rect 227830 267869 227882 267875
rect 227830 267811 227882 267817
rect 227842 263824 227870 267811
rect 228418 263824 228446 268107
rect 229078 268017 229130 268023
rect 229078 267959 229130 267965
rect 227842 263796 228096 263824
rect 228418 263796 228672 263824
rect 229090 263810 229118 267959
rect 229570 263810 229598 269217
rect 230050 263810 230078 270623
rect 232150 269497 232202 269503
rect 232150 269439 232202 269445
rect 231958 269423 232010 269429
rect 231958 269365 232010 269371
rect 230998 269349 231050 269355
rect 230998 269291 231050 269297
rect 230422 268091 230474 268097
rect 230422 268033 230474 268039
rect 230434 264120 230462 268033
rect 230434 264092 230510 264120
rect 230482 263810 230510 264092
rect 231010 263810 231038 269291
rect 231478 268239 231530 268245
rect 231478 268181 231530 268187
rect 231490 263810 231518 268181
rect 231970 263810 231998 269365
rect 232162 263824 232190 269439
rect 232642 263824 232670 271141
rect 233398 269571 233450 269577
rect 233398 269513 233450 269519
rect 232162 263796 232416 263824
rect 232642 263796 232896 263824
rect 233410 263810 233438 269513
rect 233890 263810 233918 272325
rect 234370 263810 234398 272473
rect 234946 272315 234974 277870
rect 235702 272605 235754 272611
rect 235702 272547 235754 272553
rect 234550 272309 234602 272315
rect 234550 272251 234602 272257
rect 234934 272309 234986 272315
rect 234934 272251 234986 272257
rect 234562 263824 234590 272251
rect 235030 271939 235082 271945
rect 235030 271881 235082 271887
rect 235042 263824 235070 271881
rect 234562 263796 234816 263824
rect 235042 263796 235296 263824
rect 235714 263810 235742 272547
rect 236098 272389 236126 277870
rect 236470 272901 236522 272907
rect 236470 272843 236522 272849
rect 236278 272827 236330 272833
rect 236278 272769 236330 272775
rect 236086 272383 236138 272389
rect 236086 272325 236138 272331
rect 236290 263810 236318 272769
rect 236482 263824 236510 272843
rect 236950 272753 237002 272759
rect 236950 272695 237002 272701
rect 236962 263824 236990 272695
rect 237250 271353 237278 277870
rect 237622 273123 237674 273129
rect 237622 273065 237674 273071
rect 237238 271347 237290 271353
rect 237238 271289 237290 271295
rect 236482 263796 236736 263824
rect 236962 263796 237216 263824
rect 237634 263810 237662 273065
rect 238102 273049 238154 273055
rect 238102 272991 238154 272997
rect 238114 263810 238142 272991
rect 238498 271279 238526 277870
rect 238678 273271 238730 273277
rect 238678 273213 238730 273219
rect 238486 271273 238538 271279
rect 238486 271215 238538 271221
rect 238690 263810 238718 273213
rect 239158 272975 239210 272981
rect 239158 272917 239210 272923
rect 239170 263824 239198 272917
rect 239554 271205 239582 277870
rect 239542 271199 239594 271205
rect 239542 271141 239594 271147
rect 240802 271131 240830 277870
rect 240790 271125 240842 271131
rect 240790 271067 240842 271073
rect 241954 271057 241982 277870
rect 242422 272235 242474 272241
rect 242422 272177 242474 272183
rect 242134 272161 242186 272167
rect 242134 272103 242186 272109
rect 239350 271051 239402 271057
rect 239350 270993 239402 270999
rect 241942 271051 241994 271057
rect 241942 270993 241994 270999
rect 239136 263796 239198 263824
rect 239362 263824 239390 270993
rect 240022 270977 240074 270983
rect 240022 270919 240074 270925
rect 239362 263796 239616 263824
rect 240034 263810 240062 270919
rect 240502 270903 240554 270909
rect 240502 270845 240554 270851
rect 240514 263810 240542 270845
rect 241078 270829 241130 270835
rect 241078 270771 241130 270777
rect 241090 263810 241118 270771
rect 241270 270755 241322 270761
rect 241270 270697 241322 270703
rect 241282 263824 241310 270697
rect 242146 263824 242174 272103
rect 241282 263796 241536 263824
rect 242016 263796 242174 263824
rect 242434 263810 242462 272177
rect 242902 272087 242954 272093
rect 242902 272029 242954 272035
rect 242914 263810 242942 272029
rect 243094 272013 243146 272019
rect 243094 271955 243146 271961
rect 243106 263824 243134 271955
rect 243202 270983 243230 277870
rect 244054 272679 244106 272685
rect 244054 272621 244106 272627
rect 243670 272457 243722 272463
rect 243670 272399 243722 272405
rect 243190 270977 243242 270983
rect 243190 270919 243242 270925
rect 243682 263824 243710 272399
rect 244066 263824 244094 272621
rect 244354 270909 244382 277870
rect 245302 272383 245354 272389
rect 245302 272325 245354 272331
rect 244822 272309 244874 272315
rect 244822 272251 244874 272257
rect 244342 270903 244394 270909
rect 244342 270845 244394 270851
rect 243106 263796 243360 263824
rect 243682 263796 243936 263824
rect 244066 263796 244368 263824
rect 244834 263810 244862 272251
rect 245314 263810 245342 272325
rect 245494 271347 245546 271353
rect 245494 271289 245546 271295
rect 245506 263824 245534 271289
rect 245602 270835 245630 277870
rect 246070 271273 246122 271279
rect 246070 271215 246122 271221
rect 245590 270829 245642 270835
rect 245590 270771 245642 270777
rect 246082 263824 246110 271215
rect 246454 271199 246506 271205
rect 246454 271141 246506 271147
rect 246466 263824 246494 271141
rect 246754 270761 246782 277870
rect 247222 271125 247274 271131
rect 247222 271067 247274 271073
rect 246742 270755 246794 270761
rect 246742 270697 246794 270703
rect 245506 263796 245760 263824
rect 246082 263796 246336 263824
rect 246466 263796 246768 263824
rect 247234 263810 247262 271067
rect 247702 271051 247754 271057
rect 247702 270993 247754 270999
rect 247714 263810 247742 270993
rect 247906 268393 247934 277870
rect 247990 270977 248042 270983
rect 247990 270919 248042 270925
rect 247894 268387 247946 268393
rect 247894 268329 247946 268335
rect 248002 263824 248030 270919
rect 248662 270903 248714 270909
rect 248662 270845 248714 270851
rect 248002 263796 248160 263824
rect 248674 263810 248702 270845
rect 249058 269651 249086 277870
rect 250320 277856 250526 277884
rect 249142 270829 249194 270835
rect 249142 270771 249194 270777
rect 250498 270780 250526 277856
rect 249046 269645 249098 269651
rect 249046 269587 249098 269593
rect 249154 263810 249182 270771
rect 249622 270755 249674 270761
rect 250498 270752 250718 270780
rect 249622 270697 249674 270703
rect 249634 263810 249662 270697
rect 250294 269645 250346 269651
rect 250294 269587 250346 269593
rect 249814 268387 249866 268393
rect 249814 268329 249866 268335
rect 249826 263824 249854 268329
rect 250306 263824 250334 269587
rect 250690 263824 250718 270752
rect 251458 263824 251486 277870
rect 252322 277856 252624 277884
rect 252322 263824 252350 277856
rect 253366 269571 253418 269577
rect 253366 269513 253418 269519
rect 253174 268535 253226 268541
rect 253174 268477 253226 268483
rect 252694 268387 252746 268393
rect 252694 268329 252746 268335
rect 252706 263824 252734 268329
rect 253186 263824 253214 268477
rect 249826 263796 250080 263824
rect 250306 263796 250560 263824
rect 250690 263796 250992 263824
rect 251458 263796 251568 263824
rect 252048 263796 252350 263824
rect 252480 263796 252734 263824
rect 252960 263796 253214 263824
rect 253378 263810 253406 269513
rect 253858 268393 253886 277870
rect 253942 270311 253994 270317
rect 253942 270253 253994 270259
rect 253846 268387 253898 268393
rect 253846 268329 253898 268335
rect 253954 263810 253982 270253
rect 255010 268541 255038 277870
rect 255286 270237 255338 270243
rect 255286 270179 255338 270185
rect 254998 268535 255050 268541
rect 254998 268477 255050 268483
rect 254614 268239 254666 268245
rect 254614 268181 254666 268187
rect 254626 263824 254654 268181
rect 255094 267943 255146 267949
rect 255094 267885 255146 267891
rect 255106 263824 255134 267885
rect 254400 263796 254654 263824
rect 254880 263796 255134 263824
rect 255298 263810 255326 270179
rect 255766 269719 255818 269725
rect 255766 269661 255818 269667
rect 255778 263810 255806 269661
rect 256162 269577 256190 277870
rect 257314 270317 257342 277870
rect 257302 270311 257354 270317
rect 257302 270253 257354 270259
rect 256150 269571 256202 269577
rect 256150 269513 256202 269519
rect 256246 269497 256298 269503
rect 256246 269439 256298 269445
rect 256258 263810 256286 269439
rect 258166 269349 258218 269355
rect 258166 269291 258218 269297
rect 257014 268831 257066 268837
rect 257014 268773 257066 268779
rect 257026 263824 257054 268773
rect 257686 268757 257738 268763
rect 257686 268699 257738 268705
rect 257494 268313 257546 268319
rect 257494 268255 257546 268261
rect 257506 263824 257534 268255
rect 256800 263796 257054 263824
rect 257280 263796 257534 263824
rect 257698 263810 257726 268699
rect 258178 263810 258206 269291
rect 258562 268245 258590 277870
rect 258646 269867 258698 269873
rect 258646 269809 258698 269815
rect 258550 268239 258602 268245
rect 258550 268181 258602 268187
rect 258658 263810 258686 269809
rect 259414 268535 259466 268541
rect 259414 268477 259466 268483
rect 259426 263824 259454 268477
rect 259714 267949 259742 277870
rect 260962 270243 260990 277870
rect 262006 270681 262058 270687
rect 262006 270623 262058 270629
rect 260950 270237 261002 270243
rect 260950 270179 261002 270185
rect 260086 269275 260138 269281
rect 260086 269217 260138 269223
rect 259894 269127 259946 269133
rect 259894 269069 259946 269075
rect 259702 267943 259754 267949
rect 259702 267885 259754 267891
rect 259906 263824 259934 269069
rect 259200 263796 259454 263824
rect 259680 263796 259934 263824
rect 260098 263810 260126 269217
rect 260566 269201 260618 269207
rect 260566 269143 260618 269149
rect 260578 263810 260606 269143
rect 261814 269053 261866 269059
rect 261814 268995 261866 269001
rect 261238 268387 261290 268393
rect 261238 268329 261290 268335
rect 261250 263824 261278 268329
rect 261826 263824 261854 268995
rect 261024 263796 261278 263824
rect 261600 263796 261854 263824
rect 262018 263810 262046 270623
rect 262114 269725 262142 277870
rect 262966 270607 263018 270613
rect 262966 270549 263018 270555
rect 262486 270459 262538 270465
rect 262486 270401 262538 270407
rect 262102 269719 262154 269725
rect 262102 269661 262154 269667
rect 262498 263810 262526 270401
rect 262978 263810 263006 270549
rect 263266 269503 263294 277870
rect 263254 269497 263306 269503
rect 263254 269439 263306 269445
rect 264118 268905 264170 268911
rect 264118 268847 264170 268853
rect 263638 268239 263690 268245
rect 263638 268181 263690 268187
rect 263650 263824 263678 268181
rect 264130 263824 264158 268847
rect 264418 268837 264446 277870
rect 264886 270311 264938 270317
rect 264886 270253 264938 270259
rect 264694 270163 264746 270169
rect 264694 270105 264746 270111
rect 264406 268831 264458 268837
rect 264406 268773 264458 268779
rect 264706 263824 264734 270105
rect 263424 263796 263678 263824
rect 263904 263796 264158 263824
rect 264432 263796 264734 263824
rect 264898 263810 264926 270253
rect 265366 270089 265418 270095
rect 265366 270031 265418 270037
rect 265378 263810 265406 270031
rect 265570 268319 265598 277870
rect 266038 270237 266090 270243
rect 266038 270179 266090 270185
rect 265558 268313 265610 268319
rect 265558 268255 265610 268261
rect 266050 263824 266078 270179
rect 266518 270015 266570 270021
rect 266518 269957 266570 269963
rect 266530 263824 266558 269957
rect 266818 268763 266846 277870
rect 267286 269719 267338 269725
rect 267286 269661 267338 269667
rect 267094 269571 267146 269577
rect 267094 269513 267146 269519
rect 266806 268757 266858 268763
rect 266806 268699 266858 268705
rect 267106 263824 267134 269513
rect 265824 263796 266078 263824
rect 266304 263796 266558 263824
rect 266832 263796 267134 263824
rect 267298 263810 267326 269661
rect 267766 269497 267818 269503
rect 267766 269439 267818 269445
rect 267778 263824 267806 269439
rect 267970 269355 267998 277870
rect 269218 269873 269246 277870
rect 270262 272531 270314 272537
rect 270262 272473 270314 272479
rect 269878 270311 269930 270317
rect 269878 270253 269930 270259
rect 269890 270169 269918 270253
rect 269878 270163 269930 270169
rect 269878 270105 269930 270111
rect 269494 269941 269546 269947
rect 269494 269883 269546 269889
rect 269206 269867 269258 269873
rect 269206 269809 269258 269815
rect 268438 269793 268490 269799
rect 268438 269735 268490 269741
rect 267958 269349 268010 269355
rect 267958 269291 268010 269297
rect 268450 263824 268478 269735
rect 269206 269645 269258 269651
rect 269206 269587 269258 269593
rect 268630 269423 268682 269429
rect 268630 269365 268682 269371
rect 267744 263796 267806 263824
rect 268224 263796 268478 263824
rect 268642 263810 268670 269365
rect 269218 263810 269246 269587
rect 269506 269577 269534 269883
rect 269494 269571 269546 269577
rect 269494 269513 269546 269519
rect 269686 269571 269738 269577
rect 269686 269513 269738 269519
rect 269698 263810 269726 269513
rect 270274 263824 270302 272473
rect 270370 268541 270398 277870
rect 271030 272753 271082 272759
rect 271030 272695 271082 272701
rect 270550 271939 270602 271945
rect 270550 271881 270602 271887
rect 270358 268535 270410 268541
rect 270358 268477 270410 268483
rect 270144 263796 270302 263824
rect 270562 263676 270590 271881
rect 271042 263810 271070 272695
rect 271522 269133 271550 277870
rect 271798 272457 271850 272463
rect 271798 272399 271850 272405
rect 271510 269127 271562 269133
rect 271510 269069 271562 269075
rect 271810 263824 271838 272399
rect 272278 271865 272330 271871
rect 272278 271807 272330 271813
rect 272290 263824 272318 271807
rect 272674 269281 272702 277870
rect 273922 276494 273950 277870
rect 273826 276466 273950 276494
rect 272758 272383 272810 272389
rect 272758 272325 272810 272331
rect 272662 269275 272714 269281
rect 272662 269217 272714 269223
rect 272770 263824 272798 272325
rect 273430 272309 273482 272315
rect 273430 272251 273482 272257
rect 272950 272013 273002 272019
rect 272950 271955 273002 271961
rect 271536 263796 271838 263824
rect 272064 263796 272318 263824
rect 272544 263796 272798 263824
rect 272962 263810 272990 271955
rect 273442 263810 273470 272251
rect 273826 269207 273854 276466
rect 273910 272087 273962 272093
rect 273910 272029 273962 272035
rect 273814 269201 273866 269207
rect 273814 269143 273866 269149
rect 273922 263810 273950 272029
rect 274678 269349 274730 269355
rect 274678 269291 274730 269297
rect 274690 263824 274718 269291
rect 275074 268393 275102 277870
rect 276322 276494 276350 277870
rect 276226 276466 276350 276494
rect 275350 273493 275402 273499
rect 275350 273435 275402 273441
rect 275158 272235 275210 272241
rect 275158 272177 275210 272183
rect 275062 268387 275114 268393
rect 275062 268329 275114 268335
rect 275170 263824 275198 272177
rect 274464 263796 274718 263824
rect 274944 263796 275198 263824
rect 275362 263810 275390 273435
rect 276226 269059 276254 276466
rect 276310 273419 276362 273425
rect 276310 273361 276362 273367
rect 276214 269053 276266 269059
rect 276214 268995 276266 269001
rect 275830 268683 275882 268689
rect 275830 268625 275882 268631
rect 275842 263810 275870 268625
rect 276322 263810 276350 273361
rect 277078 272161 277130 272167
rect 277078 272103 277130 272109
rect 277090 263824 277118 272103
rect 277474 270465 277502 277870
rect 277750 273567 277802 273573
rect 277750 273509 277802 273515
rect 277462 270459 277514 270465
rect 277462 270401 277514 270407
rect 277558 268905 277610 268911
rect 277558 268847 277610 268853
rect 277570 263824 277598 268847
rect 276864 263796 277118 263824
rect 277344 263796 277598 263824
rect 277762 263810 277790 273509
rect 278230 273345 278282 273351
rect 278230 273287 278282 273293
rect 278242 263810 278270 273287
rect 278722 270317 278750 277870
rect 279670 273197 279722 273203
rect 279670 273139 279722 273145
rect 279286 273049 279338 273055
rect 279286 272991 279338 272997
rect 278710 270311 278762 270317
rect 278710 270253 278762 270259
rect 278902 268979 278954 268985
rect 278902 268921 278954 268927
rect 278914 263824 278942 268921
rect 279298 263824 279326 272991
rect 278688 263796 278942 263824
rect 279168 263796 279326 263824
rect 279682 263810 279710 273139
rect 279778 270391 279806 277870
rect 280630 273123 280682 273129
rect 280630 273065 280682 273071
rect 279766 270385 279818 270391
rect 279766 270327 279818 270333
rect 280150 269053 280202 269059
rect 280150 268995 280202 269001
rect 280162 263810 280190 268995
rect 280642 263810 280670 273065
rect 281026 268245 281054 277870
rect 281302 273271 281354 273277
rect 281302 273213 281354 273219
rect 281014 268239 281066 268245
rect 281014 268181 281066 268187
rect 281314 263824 281342 273213
rect 281782 269201 281834 269207
rect 281782 269143 281834 269149
rect 281794 263824 281822 269143
rect 282178 268837 282206 277870
rect 283330 270095 283358 277870
rect 283702 270681 283754 270687
rect 283702 270623 283754 270629
rect 283318 270089 283370 270095
rect 283318 270031 283370 270037
rect 282550 269127 282602 269133
rect 282550 269069 282602 269075
rect 282166 268831 282218 268837
rect 282166 268773 282218 268779
rect 282070 268757 282122 268763
rect 282070 268699 282122 268705
rect 281088 263796 281342 263824
rect 281568 263796 281822 263824
rect 282082 263810 282110 268699
rect 282562 263810 282590 269069
rect 283030 268831 283082 268837
rect 283030 268773 283082 268779
rect 283042 263810 283070 268773
rect 283714 263824 283742 270623
rect 284182 270607 284234 270613
rect 284182 270549 284234 270555
rect 284194 263824 284222 270549
rect 284578 270169 284606 277870
rect 284950 272901 285002 272907
rect 284950 272843 285002 272849
rect 284566 270163 284618 270169
rect 284566 270105 284618 270111
rect 284470 267351 284522 267357
rect 284470 267293 284522 267299
rect 283488 263796 283742 263824
rect 283968 263796 284222 263824
rect 284482 263810 284510 267293
rect 284962 263810 284990 272843
rect 285622 270533 285674 270539
rect 285622 270475 285674 270481
rect 285634 263824 285662 270475
rect 285730 270021 285758 277870
rect 286294 270459 286346 270465
rect 286294 270401 286346 270407
rect 285718 270015 285770 270021
rect 285718 269957 285770 269963
rect 286102 267425 286154 267431
rect 286102 267367 286154 267373
rect 286114 263824 286142 267367
rect 285408 263796 285662 263824
rect 285888 263796 286142 263824
rect 286306 263810 286334 270401
rect 286774 270385 286826 270391
rect 286774 270327 286826 270333
rect 286786 263810 286814 270327
rect 286882 270243 286910 277870
rect 287926 272827 287978 272833
rect 287926 272769 287978 272775
rect 286870 270237 286922 270243
rect 286870 270179 286922 270185
rect 287350 267203 287402 267209
rect 287350 267145 287402 267151
rect 287362 263810 287390 267145
rect 287938 263824 287966 272769
rect 288034 269873 288062 277870
rect 288502 272975 288554 272981
rect 288502 272917 288554 272923
rect 288022 269867 288074 269873
rect 288022 269809 288074 269815
rect 288514 263824 288542 272917
rect 289174 270237 289226 270243
rect 289174 270179 289226 270185
rect 288694 267277 288746 267283
rect 288694 267219 288746 267225
rect 287808 263796 287966 263824
rect 288288 263796 288542 263824
rect 288706 263810 288734 267219
rect 289186 263810 289214 270179
rect 289282 269947 289310 277870
rect 289942 270163 289994 270169
rect 289942 270105 289994 270111
rect 289270 269941 289322 269947
rect 289270 269883 289322 269889
rect 289954 263824 289982 270105
rect 290434 269725 290462 277870
rect 290614 270311 290666 270317
rect 290614 270253 290666 270259
rect 290422 269719 290474 269725
rect 290422 269661 290474 269667
rect 290422 267055 290474 267061
rect 290422 266997 290474 267003
rect 290434 263824 290462 266997
rect 289728 263796 289982 263824
rect 290208 263796 290462 263824
rect 290626 263810 290654 270253
rect 291094 270089 291146 270095
rect 291094 270031 291146 270037
rect 291106 263810 291134 270031
rect 291682 269503 291710 277870
rect 292726 272679 292778 272685
rect 292726 272621 292778 272627
rect 292246 269941 292298 269947
rect 292246 269883 292298 269889
rect 291670 269497 291722 269503
rect 291670 269439 291722 269445
rect 291574 267129 291626 267135
rect 291574 267071 291626 267077
rect 291586 263810 291614 267071
rect 292258 263824 292286 269883
rect 292738 263824 292766 272621
rect 292834 269799 292862 277870
rect 293014 276231 293066 276237
rect 293014 276173 293066 276179
rect 292822 269793 292874 269799
rect 292822 269735 292874 269741
rect 292032 263796 292286 263824
rect 292608 263796 292766 263824
rect 293026 263810 293054 276173
rect 293974 270015 294026 270021
rect 293974 269957 294026 269963
rect 293494 269867 293546 269873
rect 293494 269809 293546 269815
rect 293506 263810 293534 269809
rect 293986 263810 294014 269957
rect 294082 269429 294110 277870
rect 294646 276157 294698 276163
rect 294646 276099 294698 276105
rect 294070 269423 294122 269429
rect 294070 269365 294122 269371
rect 294658 263824 294686 276099
rect 295138 269651 295166 277870
rect 295894 276083 295946 276089
rect 295894 276025 295946 276031
rect 295414 272605 295466 272611
rect 295414 272547 295466 272553
rect 295126 269645 295178 269651
rect 295126 269587 295178 269593
rect 295222 267869 295274 267875
rect 295222 267811 295274 267817
rect 295234 263824 295262 267811
rect 294432 263796 294686 263824
rect 295008 263796 295262 263824
rect 295426 263810 295454 272547
rect 295906 263810 295934 276025
rect 296386 269577 296414 277870
rect 297334 276009 297386 276015
rect 297334 275951 297386 275957
rect 296470 269793 296522 269799
rect 296470 269735 296522 269741
rect 296374 269571 296426 269577
rect 296374 269513 296426 269519
rect 296482 263824 296510 269735
rect 297046 269719 297098 269725
rect 297046 269661 297098 269667
rect 297058 263824 297086 269661
rect 296352 263796 296510 263824
rect 296832 263796 297086 263824
rect 297346 263810 297374 275951
rect 297538 272537 297566 277870
rect 297526 272531 297578 272537
rect 297526 272473 297578 272479
rect 298294 272531 298346 272537
rect 298294 272473 298346 272479
rect 297814 266981 297866 266987
rect 297814 266923 297866 266929
rect 297826 263810 297854 266923
rect 298306 263810 298334 272473
rect 298690 271945 298718 277870
rect 298966 275935 299018 275941
rect 298966 275877 299018 275883
rect 298678 271939 298730 271945
rect 298678 271881 298730 271887
rect 298978 263824 299006 275877
rect 299938 272759 299966 277870
rect 300214 275861 300266 275867
rect 300214 275803 300266 275809
rect 299926 272753 299978 272759
rect 299926 272695 299978 272701
rect 299446 271939 299498 271945
rect 299446 271881 299498 271887
rect 299458 268763 299486 271881
rect 299638 269645 299690 269651
rect 299638 269587 299690 269593
rect 299446 268757 299498 268763
rect 299446 268699 299498 268705
rect 299446 266833 299498 266839
rect 299446 266775 299498 266781
rect 299458 263824 299486 266775
rect 298752 263796 299006 263824
rect 299232 263796 299486 263824
rect 299650 263810 299678 269587
rect 300226 263810 300254 275803
rect 301090 272463 301118 277870
rect 301750 275787 301802 275793
rect 301750 275729 301802 275735
rect 301078 272457 301130 272463
rect 301078 272399 301130 272405
rect 301366 272457 301418 272463
rect 301366 272399 301418 272405
rect 300694 266907 300746 266913
rect 300694 266849 300746 266855
rect 300706 263810 300734 266849
rect 301378 263824 301406 272399
rect 301762 263824 301790 275729
rect 301846 272753 301898 272759
rect 301846 272695 301898 272701
rect 301858 267875 301886 272695
rect 302338 271871 302366 277870
rect 303286 275713 303338 275719
rect 303286 275655 303338 275661
rect 302326 271865 302378 271871
rect 302326 271807 302378 271813
rect 302614 269571 302666 269577
rect 302614 269513 302666 269519
rect 301846 267869 301898 267875
rect 301846 267811 301898 267817
rect 302038 266759 302090 266765
rect 302038 266701 302090 266707
rect 301152 263796 301406 263824
rect 301632 263796 301790 263824
rect 302050 263810 302078 266701
rect 302626 263810 302654 269513
rect 303298 263824 303326 275655
rect 303394 272389 303422 277870
rect 303766 275639 303818 275645
rect 303766 275581 303818 275587
rect 303382 272383 303434 272389
rect 303382 272325 303434 272331
rect 303778 263824 303806 275581
rect 304438 275565 304490 275571
rect 304438 275507 304490 275513
rect 303958 272383 304010 272389
rect 303958 272325 304010 272331
rect 303072 263796 303326 263824
rect 303552 263796 303806 263824
rect 303970 263810 303998 272325
rect 304450 263810 304478 275507
rect 304642 272019 304670 277870
rect 305014 275491 305066 275497
rect 305014 275433 305066 275439
rect 304630 272013 304682 272019
rect 304630 271955 304682 271961
rect 305026 263810 305054 275433
rect 305794 272315 305822 277870
rect 306358 275417 306410 275423
rect 306358 275359 306410 275365
rect 306166 275343 306218 275349
rect 306166 275285 306218 275291
rect 305782 272309 305834 272315
rect 305782 272251 305834 272257
rect 305686 269497 305738 269503
rect 305686 269439 305738 269445
rect 305698 263824 305726 269439
rect 306178 263824 306206 275285
rect 305472 263796 305726 263824
rect 305952 263796 306206 263824
rect 306370 263810 306398 275359
rect 306838 272309 306890 272315
rect 306838 272251 306890 272257
rect 306850 263810 306878 272251
rect 307042 272093 307070 277870
rect 308086 275269 308138 275275
rect 308086 275211 308138 275217
rect 307318 273937 307370 273943
rect 307318 273879 307370 273885
rect 307030 272087 307082 272093
rect 307030 272029 307082 272035
rect 307330 263810 307358 273879
rect 308098 263824 308126 275211
rect 308194 269355 308222 277870
rect 309442 272241 309470 277870
rect 310390 275195 310442 275201
rect 310390 275137 310442 275143
rect 309430 272235 309482 272241
rect 309430 272177 309482 272183
rect 309910 272235 309962 272241
rect 309910 272177 309962 272183
rect 308278 269423 308330 269429
rect 308278 269365 308330 269371
rect 308182 269349 308234 269355
rect 308182 269291 308234 269297
rect 307872 263796 308126 263824
rect 308290 263810 308318 269365
rect 308758 266685 308810 266691
rect 308758 266627 308810 266633
rect 308770 263810 308798 266627
rect 309238 266611 309290 266617
rect 309238 266553 309290 266559
rect 309250 263810 309278 266553
rect 309922 263824 309950 272177
rect 310402 263824 310430 275137
rect 310498 273499 310526 277870
rect 311638 274011 311690 274017
rect 311638 273953 311690 273959
rect 310486 273493 310538 273499
rect 310486 273435 310538 273441
rect 311158 268165 311210 268171
rect 311158 268107 311210 268113
rect 310678 266537 310730 266543
rect 310678 266479 310730 266485
rect 309696 263796 309950 263824
rect 310272 263796 310430 263824
rect 310690 263810 310718 266479
rect 311170 263810 311198 268107
rect 311650 263810 311678 273953
rect 311746 268689 311774 277870
rect 312790 273493 312842 273499
rect 312790 273435 312842 273441
rect 311734 268683 311786 268689
rect 311734 268625 311786 268631
rect 312310 266389 312362 266395
rect 312310 266331 312362 266337
rect 312322 263824 312350 266331
rect 312802 263824 312830 273435
rect 312898 273425 312926 277870
rect 313558 275047 313610 275053
rect 313558 274989 313610 274995
rect 312886 273419 312938 273425
rect 312886 273361 312938 273367
rect 313078 265427 313130 265433
rect 313078 265369 313130 265375
rect 312096 263796 312350 263824
rect 312672 263796 312830 263824
rect 313090 263810 313118 265369
rect 313570 263810 313598 274989
rect 313942 273419 313994 273425
rect 313942 273361 313994 273367
rect 313954 268837 313982 273361
rect 314146 272167 314174 277870
rect 314710 275121 314762 275127
rect 314710 275063 314762 275069
rect 314134 272161 314186 272167
rect 314134 272103 314186 272109
rect 313942 268831 313994 268837
rect 313942 268773 313994 268779
rect 314230 268091 314282 268097
rect 314230 268033 314282 268039
rect 314242 263824 314270 268033
rect 314722 263824 314750 275063
rect 315298 268911 315326 277870
rect 315958 274085 316010 274091
rect 315958 274027 316010 274033
rect 315478 272161 315530 272167
rect 315478 272103 315530 272109
rect 315286 268905 315338 268911
rect 315286 268847 315338 268853
rect 314902 265279 314954 265285
rect 314902 265221 314954 265227
rect 314016 263796 314270 263824
rect 314496 263796 314750 263824
rect 314914 263810 314942 265221
rect 315490 263810 315518 272103
rect 315970 263810 315998 274027
rect 316450 273573 316478 277870
rect 316630 277489 316682 277495
rect 316630 277431 316682 277437
rect 316438 273567 316490 273573
rect 316438 273509 316490 273515
rect 316642 263824 316670 277431
rect 317302 274159 317354 274165
rect 317302 274101 317354 274107
rect 317110 268239 317162 268245
rect 317110 268181 317162 268187
rect 317122 263824 317150 268181
rect 316416 263796 316670 263824
rect 316896 263796 317150 263824
rect 317314 263810 317342 274101
rect 317698 273351 317726 277870
rect 317686 273345 317738 273351
rect 317686 273287 317738 273293
rect 317890 263810 317918 277949
rect 319510 277933 319562 277939
rect 319510 277875 319562 277881
rect 318358 271125 318410 271131
rect 318358 271067 318410 271073
rect 318370 263810 318398 271067
rect 318754 268985 318782 277870
rect 318742 268979 318794 268985
rect 318742 268921 318794 268927
rect 319030 265353 319082 265359
rect 319030 265295 319082 265301
rect 319042 263824 319070 265295
rect 319522 263824 319550 277875
rect 320002 273055 320030 277870
rect 320182 274233 320234 274239
rect 320182 274175 320234 274181
rect 319990 273049 320042 273055
rect 319990 272991 320042 272997
rect 319702 268313 319754 268319
rect 319702 268255 319754 268261
rect 318816 263796 319070 263824
rect 319296 263796 319550 263824
rect 319714 263810 319742 268255
rect 320194 263810 320222 274175
rect 320962 263824 320990 278023
rect 415426 278013 415728 278032
rect 422570 278029 422832 278032
rect 422518 278023 422832 278029
rect 415414 278007 415728 278013
rect 415466 278004 415728 278007
rect 422530 278004 422832 278023
rect 415414 277949 415466 277955
rect 419062 277933 419114 277939
rect 321154 273203 321182 277870
rect 322102 277859 322154 277865
rect 322102 277801 322154 277807
rect 321622 274307 321674 274313
rect 321622 274249 321674 274255
rect 321142 273197 321194 273203
rect 321142 273139 321194 273145
rect 321430 271199 321482 271205
rect 321430 271141 321482 271147
rect 321442 263824 321470 271141
rect 320736 263796 320990 263824
rect 321216 263796 321470 263824
rect 321634 263810 321662 274249
rect 322114 263810 322142 277801
rect 322402 269059 322430 277870
rect 323554 273129 323582 277870
rect 323830 277785 323882 277791
rect 323830 277727 323882 277733
rect 323542 273123 323594 273129
rect 323542 273065 323594 273071
rect 322390 269053 322442 269059
rect 322390 268995 322442 269001
rect 322582 268387 322634 268393
rect 322582 268329 322634 268335
rect 322594 263810 322622 268329
rect 323350 265501 323402 265507
rect 323350 265443 323402 265449
rect 323362 263824 323390 265443
rect 323842 263824 323870 277727
rect 324802 273277 324830 277870
rect 325474 277856 325968 277884
rect 324982 277711 325034 277717
rect 324982 277653 325034 277659
rect 324790 273271 324842 273277
rect 324790 273213 324842 273219
rect 324022 271273 324074 271279
rect 324022 271215 324074 271221
rect 323136 263796 323390 263824
rect 323616 263796 323870 263824
rect 324034 263810 324062 271215
rect 324502 265575 324554 265581
rect 324502 265517 324554 265523
rect 324514 263810 324542 265517
rect 324994 263810 325022 277653
rect 325474 270780 325502 277856
rect 326422 277415 326474 277421
rect 326422 277357 326474 277363
rect 325942 274381 325994 274387
rect 325942 274323 325994 274329
rect 325378 270752 325502 270780
rect 325378 269207 325406 270752
rect 325366 269201 325418 269207
rect 325366 269143 325418 269149
rect 325750 268461 325802 268467
rect 325750 268403 325802 268409
rect 325762 263824 325790 268403
rect 325536 263796 325790 263824
rect 325954 263810 325982 274323
rect 326434 263810 326462 277357
rect 327106 271945 327134 277870
rect 328054 277637 328106 277643
rect 328054 277579 328106 277585
rect 327574 274455 327626 274461
rect 327574 274397 327626 274403
rect 327094 271939 327146 271945
rect 327094 271881 327146 271887
rect 326902 271347 326954 271353
rect 326902 271289 326954 271295
rect 326914 263810 326942 271289
rect 327586 263824 327614 274397
rect 328066 263824 328094 277579
rect 328258 269133 328286 277870
rect 329302 277341 329354 277347
rect 329302 277283 329354 277289
rect 328246 269127 328298 269133
rect 328246 269069 328298 269075
rect 328342 268535 328394 268541
rect 328342 268477 328394 268483
rect 327360 263796 327614 263824
rect 327840 263796 328094 263824
rect 328354 263810 328382 268477
rect 328822 265649 328874 265655
rect 328822 265591 328874 265597
rect 328834 263810 328862 265591
rect 329314 263810 329342 277283
rect 329506 273425 329534 277870
rect 330454 274529 330506 274535
rect 330454 274471 330506 274477
rect 329494 273419 329546 273425
rect 329494 273361 329546 273367
rect 329974 271421 330026 271427
rect 329974 271363 330026 271369
rect 329986 263824 330014 271363
rect 330466 263824 330494 274471
rect 330658 270687 330686 277870
rect 330742 277193 330794 277199
rect 330742 277135 330794 277141
rect 330646 270681 330698 270687
rect 330646 270623 330698 270629
rect 329760 263796 330014 263824
rect 330240 263796 330494 263824
rect 330754 263810 330782 277135
rect 331810 270613 331838 277870
rect 332374 277267 332426 277273
rect 332374 277209 332426 277215
rect 331798 270607 331850 270613
rect 331798 270549 331850 270555
rect 331222 268609 331274 268615
rect 331222 268551 331274 268557
rect 331234 263810 331262 268551
rect 331894 265723 331946 265729
rect 331894 265665 331946 265671
rect 331906 263824 331934 265665
rect 332386 263824 332414 277209
rect 332566 271495 332618 271501
rect 332566 271437 332618 271443
rect 331680 263796 331934 263824
rect 332160 263796 332414 263824
rect 332578 263810 332606 271437
rect 333058 267357 333086 277870
rect 333622 277119 333674 277125
rect 333622 277061 333674 277067
rect 333142 274603 333194 274609
rect 333142 274545 333194 274551
rect 333046 267351 333098 267357
rect 333046 267293 333098 267299
rect 333154 263810 333182 274545
rect 333634 263810 333662 277061
rect 334114 272907 334142 277870
rect 334102 272901 334154 272907
rect 334102 272843 334154 272849
rect 335362 270539 335390 277870
rect 336022 274677 336074 274683
rect 336022 274619 336074 274625
rect 335446 271569 335498 271575
rect 335446 271511 335498 271517
rect 335350 270533 335402 270539
rect 335350 270475 335402 270481
rect 334294 268683 334346 268689
rect 334294 268625 334346 268631
rect 334306 263824 334334 268625
rect 334966 268017 335018 268023
rect 334966 267959 335018 267965
rect 334774 265797 334826 265803
rect 334774 265739 334826 265745
rect 334786 263824 334814 265739
rect 334080 263796 334334 263824
rect 334560 263796 334814 263824
rect 334978 263810 335006 267959
rect 335458 263810 335486 271511
rect 336034 263810 336062 274619
rect 336514 267431 336542 277870
rect 336694 277045 336746 277051
rect 336694 276987 336746 276993
rect 336502 267425 336554 267431
rect 336502 267367 336554 267373
rect 336706 263824 336734 276987
rect 337762 270761 337790 277870
rect 338614 271643 338666 271649
rect 338614 271585 338666 271591
rect 337750 270755 337802 270761
rect 337750 270697 337802 270703
rect 336886 268757 336938 268763
rect 336886 268699 336938 268705
rect 336480 263796 336734 263824
rect 336898 263824 336926 268699
rect 337846 267943 337898 267949
rect 337846 267885 337898 267891
rect 337366 265871 337418 265877
rect 337366 265813 337418 265819
rect 336898 263796 336960 263824
rect 337378 263810 337406 265813
rect 337858 263810 337886 267885
rect 338626 263824 338654 271585
rect 338914 270391 338942 277870
rect 339094 274751 339146 274757
rect 339094 274693 339146 274699
rect 338902 270385 338954 270391
rect 338902 270327 338954 270333
rect 339106 263824 339134 274693
rect 339766 268905 339818 268911
rect 339766 268847 339818 268853
rect 339286 267869 339338 267875
rect 339286 267811 339338 267817
rect 338400 263796 338654 263824
rect 338880 263796 339134 263824
rect 339298 263810 339326 267811
rect 339778 263810 339806 268847
rect 340162 267209 340190 277870
rect 341314 272833 341342 277870
rect 341686 274825 341738 274831
rect 341686 274767 341738 274773
rect 341302 272827 341354 272833
rect 341302 272769 341354 272775
rect 341494 271717 341546 271723
rect 341494 271659 341546 271665
rect 340534 270829 340586 270835
rect 340534 270771 340586 270777
rect 340546 270317 340574 270771
rect 340534 270311 340586 270317
rect 340534 270253 340586 270259
rect 341014 268831 341066 268837
rect 341014 268773 341066 268779
rect 340150 267203 340202 267209
rect 340150 267145 340202 267151
rect 340246 265945 340298 265951
rect 340246 265887 340298 265893
rect 340258 263810 340286 265887
rect 341026 263824 341054 268773
rect 341506 263824 341534 271659
rect 340800 263796 341054 263824
rect 341280 263796 341534 263824
rect 341698 263810 341726 274767
rect 342166 273567 342218 273573
rect 342166 273509 342218 273515
rect 342178 263810 342206 273509
rect 342466 272981 342494 277870
rect 343330 277856 343632 277884
rect 342454 272975 342506 272981
rect 342454 272917 342506 272923
rect 342646 268979 342698 268985
rect 342646 268921 342698 268927
rect 342658 263810 342686 268921
rect 343330 267283 343358 277856
rect 344566 274899 344618 274905
rect 344566 274841 344618 274847
rect 344086 271791 344138 271797
rect 344086 271733 344138 271739
rect 343606 269053 343658 269059
rect 343606 268995 343658 269001
rect 343318 267277 343370 267283
rect 343318 267219 343370 267225
rect 343318 266019 343370 266025
rect 343318 265961 343370 265967
rect 343330 263824 343358 265961
rect 343104 263796 343358 263824
rect 343618 263810 343646 268995
rect 344098 263810 344126 271733
rect 344578 263810 344606 274841
rect 344866 270243 344894 277870
rect 345238 271865 345290 271871
rect 345238 271807 345290 271813
rect 344854 270237 344906 270243
rect 344854 270179 344906 270185
rect 345250 263824 345278 271807
rect 346018 270169 346046 277870
rect 346966 271939 347018 271945
rect 346966 271881 347018 271887
rect 346006 270163 346058 270169
rect 346006 270105 346058 270111
rect 345430 269201 345482 269207
rect 345430 269143 345482 269149
rect 345024 263796 345278 263824
rect 345442 263676 345470 269143
rect 346486 269127 346538 269133
rect 346486 269069 346538 269075
rect 346006 266093 346058 266099
rect 346006 266035 346058 266041
rect 346018 263810 346046 266035
rect 346498 263810 346526 269069
rect 346870 268017 346922 268023
rect 346870 267959 346922 267965
rect 346882 264915 346910 267959
rect 346870 264909 346922 264915
rect 346870 264851 346922 264857
rect 346978 263810 347006 271881
rect 347266 267061 347294 277870
rect 347638 274973 347690 274979
rect 347638 274915 347690 274921
rect 347254 267055 347306 267061
rect 347254 266997 347306 267003
rect 347650 263824 347678 274915
rect 348118 272087 348170 272093
rect 348118 272029 348170 272035
rect 348130 263824 348158 272029
rect 348418 270835 348446 277870
rect 348406 270829 348458 270835
rect 348406 270771 348458 270777
rect 348406 270681 348458 270687
rect 348406 270623 348458 270629
rect 347424 263796 347678 263824
rect 347904 263796 348158 263824
rect 348418 263810 348446 270623
rect 349462 270607 349514 270613
rect 349462 270549 349514 270555
rect 348886 266167 348938 266173
rect 348886 266109 348938 266115
rect 348898 263810 348926 266109
rect 349474 263824 349502 270549
rect 349570 270095 349598 277870
rect 350230 276453 350282 276459
rect 350230 276395 350282 276401
rect 350038 272013 350090 272019
rect 350038 271955 350090 271961
rect 349558 270089 349610 270095
rect 349558 270031 349610 270037
rect 350050 263824 350078 271955
rect 349344 263796 349502 263824
rect 349824 263796 350078 263824
rect 350242 263810 350270 276395
rect 350722 267135 350750 277870
rect 350998 273419 351050 273425
rect 350998 273361 351050 273367
rect 350710 267129 350762 267135
rect 350710 267071 350762 267077
rect 351010 263824 351038 273361
rect 351286 270459 351338 270465
rect 351286 270401 351338 270407
rect 350736 263796 351038 263824
rect 351298 263810 351326 270401
rect 351874 269947 351902 277870
rect 352630 273345 352682 273351
rect 352630 273287 352682 273293
rect 352438 270533 352490 270539
rect 352438 270475 352490 270481
rect 351862 269941 351914 269947
rect 351862 269883 351914 269889
rect 351958 266241 352010 266247
rect 351958 266183 352010 266189
rect 351970 263824 351998 266183
rect 352450 263824 352478 270475
rect 351744 263796 351998 263824
rect 352224 263796 352478 263824
rect 352642 263810 352670 273287
rect 353122 272685 353150 277870
rect 353398 276379 353450 276385
rect 353398 276321 353450 276327
rect 353110 272679 353162 272685
rect 353110 272621 353162 272627
rect 353410 263824 353438 276321
rect 354274 276237 354302 277870
rect 354262 276231 354314 276237
rect 354262 276173 354314 276179
rect 353686 273271 353738 273277
rect 353686 273213 353738 273219
rect 353136 263796 353438 263824
rect 353698 263810 353726 273213
rect 355030 270385 355082 270391
rect 355030 270327 355082 270333
rect 354070 270311 354122 270317
rect 354070 270253 354122 270259
rect 354082 264120 354110 270253
rect 354262 267869 354314 267875
rect 354262 267811 354314 267817
rect 354274 264989 354302 267811
rect 354838 266315 354890 266321
rect 354838 266257 354890 266263
rect 354262 264983 354314 264989
rect 354262 264925 354314 264931
rect 354082 264092 354158 264120
rect 354130 263810 354158 264092
rect 354850 263824 354878 266257
rect 354624 263796 354878 263824
rect 355042 263810 355070 270327
rect 355522 269873 355550 277870
rect 356182 276231 356234 276237
rect 356182 276173 356234 276179
rect 355798 273197 355850 273203
rect 355798 273139 355850 273145
rect 355510 269867 355562 269873
rect 355510 269809 355562 269815
rect 355810 263824 355838 273139
rect 356194 263824 356222 276173
rect 356674 270021 356702 277870
rect 357430 276305 357482 276311
rect 357430 276247 357482 276253
rect 356758 273123 356810 273129
rect 356758 273065 356810 273071
rect 356662 270015 356714 270021
rect 356662 269957 356714 269963
rect 356770 263824 356798 273065
rect 356950 270163 357002 270169
rect 356950 270105 357002 270111
rect 355536 263796 355838 263824
rect 355968 263796 356222 263824
rect 356544 263796 356798 263824
rect 356962 263810 356990 270105
rect 357442 263810 357470 276247
rect 357922 276163 357950 277870
rect 357910 276157 357962 276163
rect 357910 276099 357962 276105
rect 358978 272759 359006 277870
rect 359350 273049 359402 273055
rect 359350 272991 359402 272997
rect 358966 272753 359018 272759
rect 358966 272695 359018 272701
rect 358582 271051 358634 271057
rect 358582 270993 358634 270999
rect 357910 270237 357962 270243
rect 357910 270179 357962 270185
rect 357922 263810 357950 270179
rect 358594 263824 358622 270993
rect 359158 267795 359210 267801
rect 359158 267737 359210 267743
rect 359170 263824 359198 267737
rect 358368 263796 358622 263824
rect 358944 263796 359198 263824
rect 359362 263810 359390 272991
rect 360226 272611 360254 277870
rect 360310 276157 360362 276163
rect 360310 276099 360362 276105
rect 360214 272605 360266 272611
rect 360214 272547 360266 272553
rect 359830 270089 359882 270095
rect 359830 270031 359882 270037
rect 359842 263810 359870 270031
rect 359926 267869 359978 267875
rect 359926 267811 359978 267817
rect 359938 264841 359966 267811
rect 359926 264835 359978 264841
rect 359926 264777 359978 264783
rect 360322 263810 360350 276099
rect 361378 276089 361406 277870
rect 361366 276083 361418 276089
rect 361366 276025 361418 276031
rect 361270 272975 361322 272981
rect 361270 272917 361322 272923
rect 360982 270015 361034 270021
rect 360982 269957 361034 269963
rect 360994 263824 361022 269957
rect 360768 263796 361022 263824
rect 361282 263810 361310 272917
rect 362230 272901 362282 272907
rect 362230 272843 362282 272849
rect 361750 267721 361802 267727
rect 361750 267663 361802 267669
rect 361762 263810 361790 267663
rect 362242 263810 362270 272843
rect 362626 269799 362654 277870
rect 363382 276083 363434 276089
rect 363382 276025 363434 276031
rect 362806 269867 362858 269873
rect 362806 269809 362858 269815
rect 362614 269793 362666 269799
rect 362614 269735 362666 269741
rect 362818 263824 362846 269809
rect 363394 263824 363422 276025
rect 363574 269941 363626 269947
rect 363574 269883 363626 269889
rect 362688 263796 362846 263824
rect 363168 263796 363422 263824
rect 363586 263810 363614 269883
rect 363778 269725 363806 277870
rect 364930 276015 364958 277870
rect 364918 276009 364970 276015
rect 364918 275951 364970 275957
rect 365974 276009 366026 276015
rect 365974 275951 366026 275957
rect 364150 272827 364202 272833
rect 364150 272769 364202 272775
rect 363766 269719 363818 269725
rect 363766 269661 363818 269667
rect 364162 263810 364190 272769
rect 365302 272753 365354 272759
rect 365302 272695 365354 272701
rect 364630 267647 364682 267653
rect 364630 267589 364682 267595
rect 364642 263810 364670 267589
rect 365314 263824 365342 272695
rect 365686 269793 365738 269799
rect 365686 269735 365738 269741
rect 365698 263824 365726 269735
rect 365088 263796 365342 263824
rect 365568 263796 365726 263824
rect 365986 263810 366014 275951
rect 366082 266987 366110 277870
rect 367030 272679 367082 272685
rect 367030 272621 367082 272627
rect 366550 269719 366602 269725
rect 366550 269661 366602 269667
rect 366070 266981 366122 266987
rect 366070 266923 366122 266929
rect 366562 263810 366590 269661
rect 367042 263824 367070 272621
rect 367234 272537 367262 277870
rect 368482 275941 368510 277870
rect 369346 277856 369648 277884
rect 419114 277881 419376 277884
rect 419062 277875 419376 277881
rect 368948 276418 369004 276427
rect 368948 276353 369004 276362
rect 368470 275935 368522 275941
rect 368470 275877 368522 275883
rect 367894 272605 367946 272611
rect 367894 272547 367946 272553
rect 367222 272531 367274 272537
rect 367222 272473 367274 272479
rect 367126 269571 367178 269577
rect 367126 269513 367178 269519
rect 367138 269355 367166 269513
rect 367126 269349 367178 269355
rect 367126 269291 367178 269297
rect 367702 267573 367754 267579
rect 367702 267515 367754 267521
rect 367714 263824 367742 267515
rect 367008 263796 367070 263824
rect 367488 263796 367742 263824
rect 367906 263810 367934 272547
rect 368372 268870 368428 268879
rect 368372 268805 368428 268814
rect 368386 263810 368414 268805
rect 368962 263810 368990 276353
rect 369346 266839 369374 277856
rect 370100 271978 370156 271987
rect 370100 271913 370156 271922
rect 369622 269645 369674 269651
rect 369622 269587 369674 269593
rect 369334 266833 369386 266839
rect 369334 266775 369386 266781
rect 369634 263824 369662 269587
rect 370114 263824 370142 271913
rect 370882 269577 370910 277870
rect 372034 275867 372062 277870
rect 372502 275935 372554 275941
rect 372502 275877 372554 275883
rect 372022 275861 372074 275867
rect 372022 275803 372074 275809
rect 371252 273606 371308 273615
rect 371252 273541 371308 273550
rect 370870 269571 370922 269577
rect 370870 269513 370922 269519
rect 370292 269314 370348 269323
rect 370292 269249 370348 269258
rect 369408 263796 369662 263824
rect 369888 263796 370142 263824
rect 370306 263810 370334 269249
rect 370774 267499 370826 267505
rect 370774 267441 370826 267447
rect 370786 263810 370814 267441
rect 371266 263810 371294 273541
rect 372022 267425 372074 267431
rect 372022 267367 372074 267373
rect 372034 263824 372062 267367
rect 372514 263824 372542 275877
rect 372692 269018 372748 269027
rect 372692 268953 372748 268962
rect 371808 263796 372062 263824
rect 372288 263796 372542 263824
rect 372706 263810 372734 268953
rect 373174 267351 373226 267357
rect 373174 267293 373226 267299
rect 373186 263810 373214 267293
rect 373282 266913 373310 277870
rect 374134 272531 374186 272537
rect 374134 272473 374186 272479
rect 373846 267277 373898 267283
rect 373846 267219 373898 267225
rect 373270 266907 373322 266913
rect 373270 266849 373322 266855
rect 373858 263824 373886 267219
rect 373632 263796 373886 263824
rect 374146 263676 374174 272473
rect 374338 272463 374366 277870
rect 375094 275861 375146 275867
rect 375094 275803 375146 275809
rect 374326 272457 374378 272463
rect 374326 272399 374378 272405
rect 374614 267203 374666 267209
rect 374614 267145 374666 267151
rect 374626 263810 374654 267145
rect 375106 263810 375134 275803
rect 375586 275793 375614 277870
rect 375574 275787 375626 275793
rect 375574 275729 375626 275735
rect 376054 273049 376106 273055
rect 376054 272991 376106 272997
rect 375574 272753 375626 272759
rect 375574 272695 375626 272701
rect 375586 272611 375614 272695
rect 375574 272605 375626 272611
rect 375574 272547 375626 272553
rect 376066 271057 376094 272991
rect 376054 271051 376106 271057
rect 376054 270993 376106 270999
rect 375572 269166 375628 269175
rect 375572 269101 375628 269110
rect 375586 263810 375614 269101
rect 376246 266981 376298 266987
rect 376246 266923 376298 266929
rect 376258 263824 376286 266923
rect 376738 266765 376766 277870
rect 377012 273458 377068 273467
rect 377012 273393 377068 273402
rect 376822 267055 376874 267061
rect 376822 266997 376874 267003
rect 376726 266759 376778 266765
rect 376726 266701 376778 266707
rect 376834 263824 376862 266997
rect 376032 263796 376286 263824
rect 376608 263796 376862 263824
rect 377026 263810 377054 273393
rect 377986 269355 378014 277870
rect 379138 275719 379166 277870
rect 379126 275713 379178 275719
rect 379126 275655 379178 275661
rect 380386 275645 380414 277870
rect 380566 275787 380618 275793
rect 380566 275729 380618 275735
rect 380374 275639 380426 275645
rect 380374 275581 380426 275587
rect 378262 273863 378314 273869
rect 378262 273805 378314 273811
rect 377974 269349 378026 269355
rect 377974 269291 378026 269297
rect 377494 267129 377546 267135
rect 377494 267071 377546 267077
rect 377506 263810 377534 267071
rect 378274 263824 378302 273805
rect 379892 273310 379948 273319
rect 379892 273245 379948 273254
rect 378644 270646 378700 270655
rect 378644 270581 378700 270590
rect 378658 263824 378686 270581
rect 379126 269423 379178 269429
rect 379126 269365 379178 269371
rect 379138 263824 379166 269365
rect 379414 266907 379466 266913
rect 379414 266849 379466 266855
rect 378000 263796 378302 263824
rect 378432 263796 378686 263824
rect 378912 263796 379166 263824
rect 379426 263810 379454 266849
rect 379906 263810 379934 273245
rect 380578 263824 380606 275729
rect 381046 275713 381098 275719
rect 381046 275655 381098 275661
rect 381058 263824 381086 275655
rect 381538 272389 381566 277870
rect 381812 276270 381868 276279
rect 381812 276205 381868 276214
rect 381526 272383 381578 272389
rect 381526 272325 381578 272331
rect 381236 270498 381292 270507
rect 381236 270433 381292 270442
rect 380352 263796 380606 263824
rect 380832 263796 381086 263824
rect 381250 263810 381278 270433
rect 381826 263810 381854 276205
rect 382594 275571 382622 277870
rect 383636 276122 383692 276131
rect 383636 276057 383692 276066
rect 383446 275639 383498 275645
rect 383446 275581 383498 275587
rect 382582 275565 382634 275571
rect 382582 275507 382634 275513
rect 382966 272383 383018 272389
rect 382966 272325 383018 272331
rect 382294 266833 382346 266839
rect 382294 266775 382346 266781
rect 382306 263810 382334 266775
rect 382978 263824 383006 272325
rect 383458 263824 383486 275581
rect 382752 263796 383006 263824
rect 383232 263796 383486 263824
rect 383650 263810 383678 276057
rect 383842 275497 383870 277870
rect 384884 275974 384940 275983
rect 384884 275909 384940 275918
rect 383830 275491 383882 275497
rect 383830 275433 383882 275439
rect 384118 269275 384170 269281
rect 384118 269217 384170 269223
rect 384130 263810 384158 269217
rect 384898 263824 384926 275909
rect 384994 269577 385022 277870
rect 386242 275349 386270 277870
rect 386518 275565 386570 275571
rect 386518 275507 386570 275513
rect 386230 275343 386282 275349
rect 386230 275285 386282 275291
rect 386326 275343 386378 275349
rect 386326 275285 386378 275291
rect 385556 273162 385612 273171
rect 385556 273097 385612 273106
rect 384982 269571 385034 269577
rect 384982 269513 385034 269519
rect 385366 266759 385418 266765
rect 385366 266701 385418 266707
rect 385378 263824 385406 266701
rect 384672 263796 384926 263824
rect 385152 263796 385406 263824
rect 385570 263810 385598 273097
rect 386338 263824 386366 275285
rect 386064 263796 386366 263824
rect 386530 263810 386558 275507
rect 387394 275423 387422 277870
rect 387764 275826 387820 275835
rect 387764 275761 387820 275770
rect 387382 275417 387434 275423
rect 387382 275359 387434 275365
rect 387284 270350 387340 270359
rect 387284 270285 387340 270294
rect 387298 263824 387326 270285
rect 387778 263824 387806 275761
rect 388642 272315 388670 277870
rect 389698 273943 389726 277870
rect 390836 275678 390892 275687
rect 390836 275613 390892 275622
rect 390358 275343 390410 275349
rect 390358 275285 390410 275291
rect 389686 273937 389738 273943
rect 389686 273879 389738 273885
rect 388918 273789 388970 273795
rect 388918 273731 388970 273737
rect 388630 272309 388682 272315
rect 388630 272251 388682 272257
rect 388726 272309 388778 272315
rect 388726 272251 388778 272257
rect 387956 266798 388012 266807
rect 387956 266733 388012 266742
rect 387072 263796 387326 263824
rect 387552 263796 387806 263824
rect 387970 263810 387998 266733
rect 388738 263824 388766 272251
rect 388464 263796 388766 263824
rect 388930 263810 388958 273731
rect 390164 270202 390220 270211
rect 390164 270137 390220 270146
rect 389684 266946 389740 266955
rect 389684 266881 389740 266890
rect 389698 263824 389726 266881
rect 390178 263824 390206 270137
rect 389472 263796 389726 263824
rect 389952 263796 390206 263824
rect 390370 263810 390398 275285
rect 390850 263810 390878 275613
rect 390946 275275 390974 277870
rect 391988 275530 392044 275539
rect 391988 275465 392044 275474
rect 390934 275269 390986 275275
rect 390934 275211 390986 275217
rect 391508 273014 391564 273023
rect 391508 272949 391564 272958
rect 391522 263824 391550 272949
rect 392002 263824 392030 275465
rect 392098 269355 392126 277870
rect 393236 275382 393292 275391
rect 393236 275317 393292 275326
rect 392758 269423 392810 269429
rect 392758 269365 392810 269371
rect 392086 269349 392138 269355
rect 392086 269291 392138 269297
rect 392278 266685 392330 266691
rect 392278 266627 392330 266633
rect 391296 263796 391550 263824
rect 391776 263796 392030 263824
rect 392290 263810 392318 266627
rect 392770 263810 392798 269365
rect 393250 263810 393278 275317
rect 393346 266617 393374 277870
rect 393910 276897 393962 276903
rect 393910 276839 393962 276845
rect 393334 266611 393386 266617
rect 393334 266553 393386 266559
rect 393922 263824 393950 276839
rect 394388 272866 394444 272875
rect 394388 272801 394444 272810
rect 394402 263824 394430 272801
rect 394498 266543 394526 277870
rect 395158 275269 395210 275275
rect 395158 275211 395210 275217
rect 394678 266611 394730 266617
rect 394678 266553 394730 266559
rect 394486 266537 394538 266543
rect 394486 266479 394538 266485
rect 393696 263796 393950 263824
rect 394176 263796 394430 263824
rect 394690 263810 394718 266553
rect 395170 263810 395198 275211
rect 395746 272241 395774 277870
rect 396790 276823 396842 276829
rect 396790 276765 396842 276771
rect 396308 275086 396364 275095
rect 396308 275021 396364 275030
rect 395734 272235 395786 272241
rect 395734 272177 395786 272183
rect 395636 270054 395692 270063
rect 395636 269989 395692 269998
rect 395650 263810 395678 269989
rect 396322 263824 396350 275021
rect 396802 263824 396830 276765
rect 396898 275201 396926 277870
rect 397556 275234 397612 275243
rect 396886 275195 396938 275201
rect 397556 275169 397612 275178
rect 396886 275137 396938 275143
rect 397078 272235 397130 272241
rect 397078 272177 397130 272183
rect 396096 263796 396350 263824
rect 396576 263796 396830 263824
rect 397090 263810 397118 272177
rect 397570 263810 397598 275169
rect 398050 266469 398078 277870
rect 398230 276749 398282 276755
rect 398230 276691 398282 276697
rect 398038 266463 398090 266469
rect 398038 266405 398090 266411
rect 398242 263824 398270 276691
rect 399094 275787 399146 275793
rect 399094 275729 399146 275735
rect 399106 273869 399134 275729
rect 399094 273863 399146 273869
rect 399094 273805 399146 273811
rect 398998 269349 399050 269355
rect 398998 269291 399050 269297
rect 399010 267854 399038 269291
rect 399202 268171 399230 277870
rect 399382 276601 399434 276607
rect 399382 276543 399434 276549
rect 399190 268165 399242 268171
rect 399190 268107 399242 268113
rect 398722 267826 399038 267854
rect 398722 263824 398750 267826
rect 398902 266537 398954 266543
rect 398902 266479 398954 266485
rect 398016 263796 398270 263824
rect 398496 263796 398750 263824
rect 398914 263810 398942 266479
rect 399394 263810 399422 276543
rect 400354 274017 400382 277870
rect 401110 276675 401162 276681
rect 401110 276617 401162 276623
rect 400342 274011 400394 274017
rect 400342 273953 400394 273959
rect 399956 272718 400012 272727
rect 399956 272653 400012 272662
rect 399970 263810 399998 272653
rect 400630 266463 400682 266469
rect 400630 266405 400682 266411
rect 400642 263824 400670 266405
rect 401122 263824 401150 276617
rect 401300 269906 401356 269915
rect 401300 269841 401356 269850
rect 400416 263796 400670 263824
rect 400896 263796 401150 263824
rect 401314 263810 401342 269841
rect 401602 266395 401630 277870
rect 402550 276527 402602 276533
rect 402550 276469 402602 276475
rect 401780 266650 401836 266659
rect 401780 266585 401836 266594
rect 401590 266389 401642 266395
rect 401590 266331 401642 266337
rect 401794 263810 401822 266585
rect 402562 263824 402590 276469
rect 402754 273499 402782 277870
rect 403702 273641 403754 273647
rect 403702 273583 403754 273589
rect 402742 273493 402794 273499
rect 402742 273435 402794 273441
rect 402838 273493 402890 273499
rect 402838 273435 402890 273441
rect 402850 269323 402878 273435
rect 403028 272570 403084 272579
rect 403028 272505 403084 272514
rect 402836 269314 402892 269323
rect 402836 269249 402892 269258
rect 403042 263824 403070 272505
rect 403222 266389 403274 266395
rect 403222 266331 403274 266337
rect 402336 263796 402590 263824
rect 402816 263796 403070 263824
rect 403234 263810 403262 266331
rect 403714 263810 403742 273583
rect 404002 265433 404030 277870
rect 404950 275195 405002 275201
rect 404950 275137 405002 275143
rect 404180 269758 404236 269767
rect 404180 269693 404236 269702
rect 403990 265427 404042 265433
rect 403990 265369 404042 265375
rect 404194 263810 404222 269693
rect 404962 263824 404990 275137
rect 405154 275053 405182 277870
rect 405430 276971 405482 276977
rect 405430 276913 405482 276919
rect 405142 275047 405194 275053
rect 405142 274989 405194 274995
rect 405442 263824 405470 276913
rect 406102 273715 406154 273721
rect 406102 273657 406154 273663
rect 405620 272422 405676 272431
rect 405620 272357 405676 272366
rect 404736 263796 404990 263824
rect 405216 263796 405470 263824
rect 405634 263810 405662 272357
rect 406114 263810 406142 273657
rect 406306 268097 406334 277870
rect 407458 275127 407486 277870
rect 408022 277563 408074 277569
rect 408022 277505 408074 277511
rect 407926 275343 407978 275349
rect 407926 275285 407978 275291
rect 407446 275121 407498 275127
rect 407446 275063 407498 275069
rect 407734 275121 407786 275127
rect 407734 275063 407786 275069
rect 407746 273721 407774 275063
rect 407938 273795 407966 275285
rect 407926 273789 407978 273795
rect 407926 273731 407978 273737
rect 407734 273715 407786 273721
rect 407734 273657 407786 273663
rect 407254 269275 407306 269281
rect 407254 269217 407306 269223
rect 406294 268091 406346 268097
rect 406294 268033 406346 268039
rect 406582 265427 406634 265433
rect 406582 265369 406634 265375
rect 406594 263810 406622 265369
rect 407266 263824 407294 269217
rect 407828 266354 407884 266363
rect 407828 266289 407884 266298
rect 407842 263824 407870 266289
rect 407040 263796 407294 263824
rect 407616 263796 407870 263824
rect 408034 263810 408062 277505
rect 408500 272274 408556 272283
rect 408500 272209 408556 272218
rect 408514 263810 408542 272209
rect 408706 265285 408734 277870
rect 409654 273715 409706 273721
rect 409654 273657 409706 273663
rect 409172 266502 409228 266511
rect 409172 266437 409228 266446
rect 408694 265279 408746 265285
rect 408694 265221 408746 265227
rect 409186 263824 409214 266437
rect 409666 263824 409694 273657
rect 409858 272167 409886 277870
rect 411106 274091 411134 277870
rect 412258 277495 412286 277870
rect 412246 277489 412298 277495
rect 412246 277431 412298 277437
rect 411094 274085 411146 274091
rect 411094 274027 411146 274033
rect 409846 272161 409898 272167
rect 409846 272103 409898 272109
rect 410902 272161 410954 272167
rect 410902 272103 410954 272109
rect 411764 272126 411820 272135
rect 409940 269610 409996 269619
rect 409940 269545 409996 269554
rect 408960 263796 409214 263824
rect 409440 263796 409694 263824
rect 409954 263810 409982 269545
rect 410420 269462 410476 269471
rect 410420 269397 410476 269406
rect 410434 263810 410462 269397
rect 410914 263810 410942 272103
rect 411764 272061 411820 272070
rect 411572 269314 411628 269323
rect 411572 269249 411628 269258
rect 411586 263824 411614 269249
rect 411360 263796 411614 263824
rect 411778 263824 411806 272061
rect 413410 268245 413438 277870
rect 414562 274165 414590 277870
rect 414550 274159 414602 274165
rect 414550 274101 414602 274107
rect 416962 271131 416990 277870
rect 416950 271125 417002 271131
rect 416950 271067 417002 271073
rect 413398 268239 413450 268245
rect 413398 268181 413450 268187
rect 418114 265359 418142 277870
rect 419074 277856 419376 277875
rect 420514 268319 420542 277870
rect 421666 274239 421694 277870
rect 421654 274233 421706 274239
rect 421654 274175 421706 274181
rect 424066 271205 424094 277870
rect 425218 274313 425246 277870
rect 426274 277865 426480 277884
rect 426262 277859 426480 277865
rect 426314 277856 426480 277859
rect 426262 277801 426314 277807
rect 425206 274307 425258 274313
rect 425206 274249 425258 274255
rect 424054 271199 424106 271205
rect 424054 271141 424106 271147
rect 427618 268393 427646 277870
rect 427606 268387 427658 268393
rect 427606 268329 427658 268335
rect 420502 268313 420554 268319
rect 420502 268255 420554 268261
rect 428866 265507 428894 277870
rect 429634 277856 429936 277884
rect 429634 277791 429662 277856
rect 429622 277785 429674 277791
rect 429622 277727 429674 277733
rect 431170 271279 431198 277870
rect 431158 271273 431210 271279
rect 431158 271215 431210 271221
rect 432322 265581 432350 277870
rect 433474 277717 433502 277870
rect 433462 277711 433514 277717
rect 433462 277653 433514 277659
rect 434722 268467 434750 277870
rect 435874 274387 435902 277870
rect 437026 277421 437054 277870
rect 437014 277415 437066 277421
rect 437014 277357 437066 277363
rect 435862 274381 435914 274387
rect 435862 274323 435914 274329
rect 438178 271353 438206 277870
rect 439426 274461 439454 277870
rect 440578 277643 440606 277870
rect 440566 277637 440618 277643
rect 440566 277579 440618 277585
rect 439414 274455 439466 274461
rect 439414 274397 439466 274403
rect 438166 271347 438218 271353
rect 438166 271289 438218 271295
rect 441826 268541 441854 277870
rect 441814 268535 441866 268541
rect 441814 268477 441866 268483
rect 434710 268461 434762 268467
rect 434710 268403 434762 268409
rect 442978 265655 443006 277870
rect 444226 277347 444254 277870
rect 444214 277341 444266 277347
rect 444214 277283 444266 277289
rect 445282 271427 445310 277870
rect 446530 274535 446558 277870
rect 447682 277199 447710 277870
rect 447670 277193 447722 277199
rect 447670 277135 447722 277141
rect 446518 274529 446570 274535
rect 446518 274471 446570 274477
rect 445270 271421 445322 271427
rect 445270 271363 445322 271369
rect 448834 268615 448862 277870
rect 448822 268609 448874 268615
rect 448822 268551 448874 268557
rect 450082 265729 450110 277870
rect 451234 277273 451262 277870
rect 451222 277267 451274 277273
rect 451222 277209 451274 277215
rect 452482 271501 452510 277870
rect 453538 274609 453566 277870
rect 454786 277125 454814 277870
rect 454774 277119 454826 277125
rect 454774 277061 454826 277067
rect 453526 274603 453578 274609
rect 453526 274545 453578 274551
rect 452470 271495 452522 271501
rect 452470 271437 452522 271443
rect 455938 268689 455966 277870
rect 455926 268683 455978 268689
rect 455926 268625 455978 268631
rect 457186 265803 457214 277870
rect 457174 265797 457226 265803
rect 457174 265739 457226 265745
rect 450070 265723 450122 265729
rect 450070 265665 450122 265671
rect 442966 265649 443018 265655
rect 442966 265591 443018 265597
rect 432310 265575 432362 265581
rect 432310 265517 432362 265523
rect 428854 265501 428906 265507
rect 428854 265443 428906 265449
rect 418102 265353 418154 265359
rect 418102 265295 418154 265301
rect 458338 264915 458366 277870
rect 459586 271575 459614 277870
rect 460642 274683 460670 277870
rect 461890 277051 461918 277870
rect 461878 277045 461930 277051
rect 461878 276987 461930 276993
rect 460630 274677 460682 274683
rect 460630 274619 460682 274625
rect 459574 271569 459626 271575
rect 459574 271511 459626 271517
rect 463042 268763 463070 277870
rect 463030 268757 463082 268763
rect 463030 268699 463082 268705
rect 464290 265877 464318 277870
rect 464278 265871 464330 265877
rect 464278 265813 464330 265819
rect 458326 264909 458378 264915
rect 458326 264851 458378 264857
rect 465442 264841 465470 277870
rect 466594 271649 466622 277870
rect 467842 274757 467870 277870
rect 467830 274751 467882 274757
rect 467830 274693 467882 274699
rect 466582 271643 466634 271649
rect 466582 271585 466634 271591
rect 468898 264989 468926 277870
rect 470146 268911 470174 277870
rect 470134 268905 470186 268911
rect 470134 268847 470186 268853
rect 471298 265951 471326 277870
rect 472546 268837 472574 277870
rect 473698 271723 473726 277870
rect 474946 274831 474974 277870
rect 474934 274825 474986 274831
rect 474934 274767 474986 274773
rect 476098 273573 476126 277870
rect 476086 273567 476138 273573
rect 476086 273509 476138 273515
rect 473686 271717 473738 271723
rect 473686 271659 473738 271665
rect 477250 268985 477278 277870
rect 477238 268979 477290 268985
rect 477238 268921 477290 268927
rect 472534 268831 472586 268837
rect 472534 268773 472586 268779
rect 478402 266025 478430 277870
rect 479650 269059 479678 277870
rect 480802 271797 480830 277870
rect 481954 274905 481982 277870
rect 481942 274899 481994 274905
rect 481942 274841 481994 274847
rect 480886 273715 480938 273721
rect 480886 273657 480938 273663
rect 480898 273573 480926 273657
rect 480886 273567 480938 273573
rect 480886 273509 480938 273515
rect 483202 271871 483230 277870
rect 483190 271865 483242 271871
rect 483190 271807 483242 271813
rect 480790 271791 480842 271797
rect 480790 271733 480842 271739
rect 484258 269207 484286 277870
rect 484246 269201 484298 269207
rect 484246 269143 484298 269149
rect 479638 269053 479690 269059
rect 479638 268995 479690 269001
rect 485506 266099 485534 277870
rect 486658 269133 486686 277870
rect 487906 271945 487934 277870
rect 489058 274979 489086 277870
rect 489046 274973 489098 274979
rect 489046 274915 489098 274921
rect 490306 272093 490334 277870
rect 490294 272087 490346 272093
rect 490294 272029 490346 272035
rect 487894 271939 487946 271945
rect 487894 271881 487946 271887
rect 491458 270687 491486 277870
rect 491446 270681 491498 270687
rect 491446 270623 491498 270629
rect 486646 269127 486698 269133
rect 486646 269069 486698 269075
rect 492610 266173 492638 277870
rect 493762 270613 493790 277870
rect 495010 272019 495038 277870
rect 496162 276459 496190 277870
rect 496150 276453 496202 276459
rect 496150 276395 496202 276401
rect 497410 273425 497438 277870
rect 497398 273419 497450 273425
rect 497398 273361 497450 273367
rect 494998 272013 495050 272019
rect 494998 271955 495050 271961
rect 493750 270607 493802 270613
rect 493750 270549 493802 270555
rect 498562 270465 498590 277870
rect 498550 270459 498602 270465
rect 498550 270401 498602 270407
rect 499714 266247 499742 277870
rect 500866 270539 500894 277870
rect 502018 273351 502046 277870
rect 503266 276385 503294 277870
rect 503254 276379 503306 276385
rect 503254 276321 503306 276327
rect 502006 273345 502058 273351
rect 502006 273287 502058 273293
rect 504418 273277 504446 277870
rect 504406 273271 504458 273277
rect 504406 273213 504458 273219
rect 500854 270533 500906 270539
rect 500854 270475 500906 270481
rect 505666 270317 505694 277870
rect 506530 277856 506832 277884
rect 505654 270311 505706 270317
rect 505654 270253 505706 270259
rect 506530 266321 506558 277856
rect 506806 273641 506858 273647
rect 506806 273583 506858 273589
rect 506818 273425 506846 273583
rect 506806 273419 506858 273425
rect 506806 273361 506858 273367
rect 507970 270391 507998 277870
rect 509122 273203 509150 277870
rect 510370 276237 510398 277870
rect 510358 276231 510410 276237
rect 510358 276173 510410 276179
rect 509110 273197 509162 273203
rect 509110 273139 509162 273145
rect 509206 273197 509258 273203
rect 509206 273139 509258 273145
rect 507958 270385 508010 270391
rect 507958 270327 508010 270333
rect 506518 266315 506570 266321
rect 506518 266257 506570 266263
rect 499702 266241 499754 266247
rect 499702 266183 499754 266189
rect 492598 266167 492650 266173
rect 492598 266109 492650 266115
rect 485494 266093 485546 266099
rect 485494 266035 485546 266041
rect 478390 266019 478442 266025
rect 478390 265961 478442 265967
rect 471286 265945 471338 265951
rect 471286 265887 471338 265893
rect 509218 265433 509246 273139
rect 511522 273129 511550 277870
rect 511510 273123 511562 273129
rect 511510 273065 511562 273071
rect 512770 270169 512798 277870
rect 513922 276311 513950 277870
rect 513910 276305 513962 276311
rect 513910 276247 513962 276253
rect 515074 270243 515102 277870
rect 516226 273055 516254 277870
rect 516214 273049 516266 273055
rect 516214 272991 516266 272997
rect 515062 270237 515114 270243
rect 515062 270179 515114 270185
rect 512758 270163 512810 270169
rect 512758 270105 512810 270111
rect 517378 267801 517406 277870
rect 518626 272981 518654 277870
rect 518614 272975 518666 272981
rect 518614 272917 518666 272923
rect 519778 270095 519806 277870
rect 521026 276163 521054 277870
rect 521014 276157 521066 276163
rect 521014 276099 521066 276105
rect 519766 270089 519818 270095
rect 519766 270031 519818 270037
rect 522178 270021 522206 277870
rect 523426 272907 523454 277870
rect 523414 272901 523466 272907
rect 523414 272843 523466 272849
rect 522166 270015 522218 270021
rect 522166 269957 522218 269963
rect 517366 267795 517418 267801
rect 517366 267737 517418 267743
rect 524482 267727 524510 277870
rect 525730 272833 525758 277870
rect 525718 272827 525770 272833
rect 525718 272769 525770 272775
rect 526882 269873 526910 277870
rect 528130 276089 528158 277870
rect 528118 276083 528170 276089
rect 528118 276025 528170 276031
rect 529282 269947 529310 277870
rect 530530 272759 530558 277870
rect 530518 272753 530570 272759
rect 530518 272695 530570 272701
rect 529270 269941 529322 269947
rect 529270 269883 529322 269889
rect 526870 269867 526922 269873
rect 526870 269809 526922 269815
rect 524470 267721 524522 267727
rect 524470 267663 524522 267669
rect 531586 267653 531614 277870
rect 532834 272611 532862 277870
rect 532822 272605 532874 272611
rect 532822 272547 532874 272553
rect 533986 269799 534014 277870
rect 535138 276015 535166 277870
rect 535126 276009 535178 276015
rect 535126 275951 535178 275957
rect 533974 269793 534026 269799
rect 533974 269735 534026 269741
rect 536386 269725 536414 277870
rect 537538 272685 537566 277870
rect 537526 272679 537578 272685
rect 537526 272621 537578 272627
rect 536374 269719 536426 269725
rect 536374 269661 536426 269667
rect 531574 267647 531626 267653
rect 531574 267589 531626 267595
rect 538786 267579 538814 277870
rect 539842 272537 539870 277870
rect 539830 272531 539882 272537
rect 539830 272473 539882 272479
rect 541090 268879 541118 277870
rect 542242 276427 542270 277870
rect 542228 276418 542284 276427
rect 542228 276353 542284 276362
rect 543490 269651 543518 277870
rect 544642 271987 544670 277870
rect 545890 273499 545918 277870
rect 546646 277563 546698 277569
rect 546646 277505 546698 277511
rect 546658 273499 546686 277505
rect 545878 273493 545930 273499
rect 545878 273435 545930 273441
rect 546646 273493 546698 273499
rect 546646 273435 546698 273441
rect 544628 271978 544684 271987
rect 544628 271913 544684 271922
rect 543478 269645 543530 269651
rect 543478 269587 543530 269593
rect 541076 268870 541132 268879
rect 541076 268805 541132 268814
rect 538774 267573 538826 267579
rect 538774 267515 538826 267521
rect 547042 267505 547070 277870
rect 548194 273615 548222 277870
rect 548180 273606 548236 273615
rect 548180 273541 548236 273550
rect 547030 267499 547082 267505
rect 547030 267441 547082 267447
rect 549346 267431 549374 277870
rect 550498 275941 550526 277870
rect 550486 275935 550538 275941
rect 550486 275877 550538 275883
rect 551746 269027 551774 277870
rect 551732 269018 551788 269027
rect 551732 268953 551788 268962
rect 549334 267425 549386 267431
rect 549334 267367 549386 267373
rect 552898 267357 552926 277870
rect 552886 267351 552938 267357
rect 552886 267293 552938 267299
rect 554146 267283 554174 277870
rect 555202 272463 555230 277870
rect 555190 272457 555242 272463
rect 555190 272399 555242 272405
rect 554134 267277 554186 267283
rect 554134 267219 554186 267225
rect 556450 267209 556478 277870
rect 557602 275867 557630 277870
rect 557590 275861 557642 275867
rect 557590 275803 557642 275809
rect 558850 269175 558878 277870
rect 558836 269166 558892 269175
rect 558836 269101 558892 269110
rect 556438 267203 556490 267209
rect 556438 267145 556490 267151
rect 560002 266987 560030 277870
rect 561250 267061 561278 277870
rect 562402 273467 562430 277870
rect 562388 273458 562444 273467
rect 562388 273393 562444 273402
rect 563554 267135 563582 277870
rect 564706 275793 564734 277870
rect 564694 275787 564746 275793
rect 564694 275729 564746 275735
rect 565858 270655 565886 277870
rect 565844 270646 565900 270655
rect 565844 270581 565900 270590
rect 567106 269577 567134 277870
rect 567094 269571 567146 269577
rect 567094 269513 567146 269519
rect 563542 267129 563594 267135
rect 563542 267071 563594 267077
rect 561238 267055 561290 267061
rect 561238 266997 561290 267003
rect 559990 266981 560042 266987
rect 559990 266923 560042 266929
rect 568258 266913 568286 277870
rect 569506 273319 569534 277870
rect 570658 275719 570686 277870
rect 570646 275713 570698 275719
rect 570646 275655 570698 275661
rect 571810 275645 571838 277870
rect 571798 275639 571850 275645
rect 571798 275581 571850 275587
rect 569492 273310 569548 273319
rect 569492 273245 569548 273254
rect 572962 270507 572990 277870
rect 574210 276279 574238 277870
rect 574196 276270 574252 276279
rect 574196 276205 574252 276214
rect 572948 270498 573004 270507
rect 572948 270433 573004 270442
rect 568246 266907 568298 266913
rect 568246 266849 568298 266855
rect 575362 266839 575390 277870
rect 576610 272389 576638 277870
rect 577762 275571 577790 277870
rect 578914 276131 578942 277870
rect 578900 276122 578956 276131
rect 578900 276057 578956 276066
rect 577750 275565 577802 275571
rect 577750 275507 577802 275513
rect 576598 272383 576650 272389
rect 576598 272325 576650 272331
rect 580066 269503 580094 277870
rect 581314 275983 581342 277870
rect 581300 275974 581356 275983
rect 581300 275909 581356 275918
rect 580054 269497 580106 269503
rect 580054 269439 580106 269445
rect 575350 266833 575402 266839
rect 575350 266775 575402 266781
rect 582466 266765 582494 277870
rect 583618 273171 583646 277870
rect 584866 275423 584894 277870
rect 586018 275497 586046 277870
rect 586006 275491 586058 275497
rect 586006 275433 586058 275439
rect 584854 275417 584906 275423
rect 584854 275359 584906 275365
rect 583604 273162 583660 273171
rect 583604 273097 583660 273106
rect 587170 270359 587198 277870
rect 588322 275835 588350 277870
rect 588308 275826 588364 275835
rect 588308 275761 588364 275770
rect 587156 270350 587212 270359
rect 587156 270285 587212 270294
rect 589570 266807 589598 277870
rect 590722 272315 590750 277870
rect 591970 275349 591998 277870
rect 591958 275343 592010 275349
rect 591958 275285 592010 275291
rect 590710 272309 590762 272315
rect 590710 272251 590762 272257
rect 593122 266955 593150 277870
rect 594370 270211 594398 277870
rect 595426 275275 595454 277870
rect 596674 275687 596702 277870
rect 596660 275678 596716 275687
rect 596660 275613 596716 275622
rect 595414 275269 595466 275275
rect 595414 275211 595466 275217
rect 597826 273023 597854 277870
rect 599074 275539 599102 277870
rect 599060 275530 599116 275539
rect 599060 275465 599116 275474
rect 597812 273014 597868 273023
rect 597812 272949 597868 272958
rect 594356 270202 594412 270211
rect 594356 270137 594412 270146
rect 593108 266946 593164 266955
rect 593108 266881 593164 266890
rect 589556 266798 589612 266807
rect 582454 266759 582506 266765
rect 589556 266733 589612 266742
rect 582454 266701 582506 266707
rect 600226 266691 600254 277870
rect 601378 269429 601406 277870
rect 602530 275391 602558 277870
rect 603682 276903 603710 277870
rect 603670 276897 603722 276903
rect 603670 276839 603722 276845
rect 602516 275382 602572 275391
rect 602516 275317 602572 275326
rect 604930 272875 604958 277870
rect 604916 272866 604972 272875
rect 604916 272801 604972 272810
rect 601366 269423 601418 269429
rect 601366 269365 601418 269371
rect 600214 266685 600266 266691
rect 600214 266627 600266 266633
rect 606082 266617 606110 277870
rect 607330 275201 607358 277870
rect 607318 275195 607370 275201
rect 607318 275137 607370 275143
rect 608482 270063 608510 277870
rect 609730 275095 609758 277870
rect 610786 276829 610814 277870
rect 610774 276823 610826 276829
rect 610774 276765 610826 276771
rect 609716 275086 609772 275095
rect 609716 275021 609772 275030
rect 612034 272241 612062 277870
rect 612982 276971 613034 276977
rect 612982 276913 613034 276919
rect 612994 273351 613022 276913
rect 613186 275243 613214 277870
rect 614434 276755 614462 277870
rect 614422 276749 614474 276755
rect 614422 276691 614474 276697
rect 613172 275234 613228 275243
rect 613172 275169 613228 275178
rect 612982 273345 613034 273351
rect 612982 273287 613034 273293
rect 612022 272235 612074 272241
rect 612022 272177 612074 272183
rect 608468 270054 608524 270063
rect 608468 269989 608524 269998
rect 615586 269355 615614 277870
rect 615574 269349 615626 269355
rect 615574 269291 615626 269297
rect 606070 266611 606122 266617
rect 606070 266553 606122 266559
rect 616738 266543 616766 277870
rect 617986 276607 618014 277870
rect 617974 276601 618026 276607
rect 617974 276543 618026 276549
rect 619042 272727 619070 277870
rect 619028 272718 619084 272727
rect 619028 272653 619084 272662
rect 616726 266537 616778 266543
rect 616726 266479 616778 266485
rect 620290 266469 620318 277870
rect 621442 276681 621470 277870
rect 621430 276675 621482 276681
rect 621430 276617 621482 276623
rect 622690 269915 622718 277870
rect 622676 269906 622732 269915
rect 622676 269841 622732 269850
rect 623842 266659 623870 277870
rect 625090 276533 625118 277870
rect 625078 276527 625130 276533
rect 625078 276469 625130 276475
rect 626146 272579 626174 277870
rect 626132 272570 626188 272579
rect 626132 272505 626188 272514
rect 623828 266650 623884 266659
rect 623828 266585 623884 266594
rect 620278 266463 620330 266469
rect 620278 266405 620330 266411
rect 627394 266395 627422 277870
rect 628546 273425 628574 277870
rect 628534 273419 628586 273425
rect 628534 273361 628586 273367
rect 629794 269767 629822 277870
rect 630946 275053 630974 277870
rect 630934 275047 630986 275053
rect 630934 274989 630986 274995
rect 632098 273351 632126 277870
rect 632086 273345 632138 273351
rect 632086 273287 632138 273293
rect 633346 272431 633374 277870
rect 634402 275127 634430 277870
rect 634390 275121 634442 275127
rect 634390 275063 634442 275069
rect 635650 273203 635678 277870
rect 635638 273197 635690 273203
rect 635638 273139 635690 273145
rect 633332 272422 633388 272431
rect 633332 272357 633388 272366
rect 629780 269758 629836 269767
rect 629780 269693 629836 269702
rect 636802 269281 636830 277870
rect 636790 269275 636842 269281
rect 636790 269217 636842 269223
rect 627382 266389 627434 266395
rect 638050 266363 638078 277870
rect 639202 273499 639230 277870
rect 639190 273493 639242 273499
rect 639190 273435 639242 273441
rect 640450 272283 640478 277870
rect 640436 272274 640492 272283
rect 640436 272209 640492 272218
rect 641602 266511 641630 277870
rect 642754 273573 642782 277870
rect 642742 273567 642794 273573
rect 642742 273509 642794 273515
rect 643906 269619 643934 277870
rect 643892 269610 643948 269619
rect 643892 269545 643948 269554
rect 645154 269471 645182 277870
rect 646306 272167 646334 277870
rect 646294 272161 646346 272167
rect 646294 272103 646346 272109
rect 645140 269462 645196 269471
rect 645140 269397 645196 269406
rect 647554 269323 647582 277870
rect 648706 272135 648734 277870
rect 648692 272126 648748 272135
rect 648692 272061 648748 272070
rect 647540 269314 647596 269323
rect 647540 269249 647596 269258
rect 641588 266502 641644 266511
rect 641588 266437 641644 266446
rect 627382 266331 627434 266337
rect 638036 266354 638092 266363
rect 638036 266289 638092 266298
rect 509206 265427 509258 265433
rect 509206 265369 509258 265375
rect 468886 264983 468938 264989
rect 468886 264925 468938 264931
rect 465430 264835 465482 264841
rect 465430 264777 465482 264783
rect 411778 263796 411840 263824
rect 270562 263648 270624 263676
rect 345442 263648 345504 263676
rect 374146 263648 374208 263676
rect 420404 262210 420460 262219
rect 420404 262145 420406 262154
rect 420458 262145 420460 262154
rect 606166 262171 606218 262177
rect 420406 262113 420458 262119
rect 606166 262113 606218 262119
rect 420404 259842 420460 259851
rect 420404 259777 420460 259786
rect 190004 259398 190060 259407
rect 190004 259333 190060 259342
rect 189908 251702 189964 251711
rect 189908 251637 189964 251646
rect 189922 224955 189950 251637
rect 190018 227545 190046 259333
rect 420418 259291 420446 259777
rect 420406 259285 420458 259291
rect 420406 259227 420458 259233
rect 603286 259285 603338 259291
rect 603286 259227 603338 259233
rect 420404 257030 420460 257039
rect 420404 256965 420460 256974
rect 420418 256405 420446 256965
rect 420406 256399 420458 256405
rect 420406 256341 420458 256347
rect 420404 255254 420460 255263
rect 420404 255189 420460 255198
rect 420418 253519 420446 255189
rect 420406 253513 420458 253519
rect 420406 253455 420458 253461
rect 420404 252886 420460 252895
rect 420404 252821 420460 252830
rect 420418 250633 420446 252821
rect 420406 250627 420458 250633
rect 420406 250569 420458 250575
rect 420308 250518 420364 250527
rect 420308 250453 420364 250462
rect 420322 247821 420350 250453
rect 420404 248150 420460 248159
rect 420404 248085 420460 248094
rect 420310 247815 420362 247821
rect 420310 247757 420362 247763
rect 420418 247747 420446 248085
rect 600406 247815 600458 247821
rect 600406 247757 600458 247763
rect 420406 247741 420458 247747
rect 420406 247683 420458 247689
rect 420404 245338 420460 245347
rect 420404 245273 420460 245282
rect 420418 244861 420446 245273
rect 420406 244855 420458 244861
rect 420406 244797 420458 244803
rect 420404 243562 420460 243571
rect 420404 243497 420460 243506
rect 420418 241975 420446 243497
rect 420406 241969 420458 241975
rect 420406 241911 420458 241917
rect 420404 241194 420460 241203
rect 420404 241129 420460 241138
rect 192418 233391 192446 239686
rect 192768 239672 192926 239700
rect 193152 239672 193406 239700
rect 192898 233613 192926 239672
rect 193378 236174 193406 239672
rect 193090 236146 193406 236174
rect 192886 233607 192938 233613
rect 192886 233549 192938 233555
rect 192406 233385 192458 233391
rect 192406 233327 192458 233333
rect 190006 227539 190058 227545
rect 190006 227481 190058 227487
rect 191542 227539 191594 227545
rect 191542 227481 191594 227487
rect 189910 224949 189962 224955
rect 189910 224891 189962 224897
rect 190774 224727 190826 224733
rect 190774 224669 190826 224675
rect 190786 221792 190814 224669
rect 190786 221764 190862 221792
rect 190834 221482 190862 221764
rect 191554 221482 191582 227481
rect 192310 224949 192362 224955
rect 192310 224891 192362 224897
rect 192322 221482 192350 224891
rect 193090 221792 193118 236146
rect 193474 233317 193502 239686
rect 193858 233391 193886 239686
rect 194242 233539 194270 239686
rect 194230 233533 194282 233539
rect 194230 233475 194282 233481
rect 194626 233465 194654 239686
rect 194976 239672 195230 239700
rect 195360 239672 195614 239700
rect 194614 233459 194666 233465
rect 194614 233401 194666 233407
rect 193750 233385 193802 233391
rect 193750 233327 193802 233333
rect 193846 233385 193898 233391
rect 193846 233327 193898 233333
rect 193462 233311 193514 233317
rect 193462 233253 193514 233259
rect 193042 221764 193118 221792
rect 193042 221482 193070 221764
rect 193762 221482 193790 233327
rect 195202 233317 195230 239672
rect 195586 233613 195614 239672
rect 195682 233687 195710 239686
rect 195670 233681 195722 233687
rect 195670 233623 195722 233629
rect 195286 233607 195338 233613
rect 195286 233549 195338 233555
rect 195574 233607 195626 233613
rect 195574 233549 195626 233555
rect 194614 233311 194666 233317
rect 194614 233253 194666 233259
rect 195190 233311 195242 233317
rect 195190 233253 195242 233259
rect 194626 221482 194654 233253
rect 195298 221792 195326 233549
rect 196162 233465 196190 239686
rect 196546 233761 196574 239686
rect 196930 233835 196958 239686
rect 197280 239672 197534 239700
rect 197664 239672 197918 239700
rect 197506 233983 197534 239672
rect 197494 233977 197546 233983
rect 197494 233919 197546 233925
rect 196918 233829 196970 233835
rect 196918 233771 196970 233777
rect 196534 233755 196586 233761
rect 196534 233697 196586 233703
rect 196054 233459 196106 233465
rect 196054 233401 196106 233407
rect 196150 233459 196202 233465
rect 196150 233401 196202 233407
rect 195298 221764 195374 221792
rect 195346 221482 195374 221764
rect 196066 221482 196094 233401
rect 196822 233385 196874 233391
rect 196822 233327 196874 233333
rect 196834 221482 196862 233327
rect 197890 233317 197918 239672
rect 197986 233391 198014 239686
rect 198370 234057 198398 239686
rect 198754 234131 198782 239686
rect 198742 234125 198794 234131
rect 198742 234067 198794 234073
rect 198358 234051 198410 234057
rect 198358 233993 198410 233999
rect 199138 233909 199166 239686
rect 199488 239672 199742 239700
rect 199968 239672 200222 239700
rect 199126 233903 199178 233909
rect 199126 233845 199178 233851
rect 198358 233533 198410 233539
rect 198358 233475 198410 233481
rect 197974 233385 198026 233391
rect 197974 233327 198026 233333
rect 197494 233311 197546 233317
rect 197494 233253 197546 233259
rect 197878 233311 197930 233317
rect 197878 233253 197930 233259
rect 197506 221792 197534 233253
rect 197506 221764 197582 221792
rect 197554 221482 197582 221764
rect 198370 221482 198398 233475
rect 199714 233465 199742 239672
rect 200194 234205 200222 239672
rect 200290 234279 200318 239686
rect 200278 234273 200330 234279
rect 200278 234215 200330 234221
rect 200182 234199 200234 234205
rect 200182 234141 200234 234147
rect 200566 233755 200618 233761
rect 200566 233697 200618 233703
rect 199798 233607 199850 233613
rect 199798 233549 199850 233555
rect 199126 233459 199178 233465
rect 199126 233401 199178 233407
rect 199702 233459 199754 233465
rect 199702 233401 199754 233407
rect 199138 221482 199166 233401
rect 199810 221792 199838 233549
rect 199810 221764 199886 221792
rect 199858 221482 199886 221764
rect 200578 221482 200606 233697
rect 200674 233539 200702 239686
rect 201058 233613 201086 239686
rect 201408 239672 201566 239700
rect 201792 239672 202046 239700
rect 202176 239672 202430 239700
rect 201538 233761 201566 239672
rect 202018 234501 202046 239672
rect 202006 234495 202058 234501
rect 202006 234437 202058 234443
rect 201526 233755 201578 233761
rect 201526 233697 201578 233703
rect 201334 233681 201386 233687
rect 201334 233623 201386 233629
rect 201046 233607 201098 233613
rect 201046 233549 201098 233555
rect 200662 233533 200714 233539
rect 200662 233475 200714 233481
rect 201346 221763 201374 233623
rect 202402 233317 202430 239672
rect 202498 233687 202526 239686
rect 202882 234575 202910 239686
rect 203266 234871 203294 239686
rect 203712 239672 203966 239700
rect 204096 239672 204254 239700
rect 203254 234865 203306 234871
rect 203254 234807 203306 234813
rect 202870 234569 202922 234575
rect 202870 234511 202922 234517
rect 202870 233829 202922 233835
rect 202870 233771 202922 233777
rect 202486 233681 202538 233687
rect 202486 233623 202538 233629
rect 202102 233311 202154 233317
rect 202102 233253 202154 233259
rect 202390 233311 202442 233317
rect 202390 233253 202442 233259
rect 202114 221792 202142 233253
rect 202114 221764 202190 221792
rect 201336 221713 201374 221763
rect 201336 221482 201364 221713
rect 202162 221482 202190 221764
rect 202882 221482 202910 233771
rect 203938 233391 203966 239672
rect 204226 233835 204254 239672
rect 204418 239672 204480 239700
rect 204418 234945 204446 239672
rect 204406 234939 204458 234945
rect 204406 234881 204458 234887
rect 204802 234649 204830 239686
rect 204790 234643 204842 234649
rect 204790 234585 204842 234591
rect 205186 233983 205214 239686
rect 204310 233977 204362 233983
rect 204310 233919 204362 233925
rect 205174 233977 205226 233983
rect 205174 233919 205226 233925
rect 204214 233829 204266 233835
rect 204214 233771 204266 233777
rect 203638 233385 203690 233391
rect 203638 233327 203690 233333
rect 203926 233385 203978 233391
rect 203926 233327 203978 233333
rect 203650 221482 203678 233327
rect 204322 221792 204350 233919
rect 205570 233909 205598 239686
rect 205920 239672 206174 239700
rect 206304 239672 206558 239700
rect 206688 239672 206942 239700
rect 206146 234427 206174 239672
rect 206530 234723 206558 239672
rect 206518 234717 206570 234723
rect 206518 234659 206570 234665
rect 206134 234421 206186 234427
rect 206134 234363 206186 234369
rect 206914 234057 206942 239672
rect 207010 234797 207038 239686
rect 206998 234791 207050 234797
rect 206998 234733 207050 234739
rect 207286 234643 207338 234649
rect 207286 234585 207338 234591
rect 207298 234224 207326 234585
rect 207382 234347 207434 234353
rect 207382 234289 207434 234295
rect 207394 234224 207422 234289
rect 207298 234196 207422 234224
rect 207490 234131 207518 239686
rect 207874 234649 207902 239686
rect 208224 239672 208478 239700
rect 208608 239672 208766 239700
rect 207862 234643 207914 234649
rect 207862 234585 207914 234591
rect 207382 234125 207434 234131
rect 207382 234067 207434 234073
rect 207478 234125 207530 234131
rect 207478 234067 207530 234073
rect 205942 234051 205994 234057
rect 205942 233993 205994 233999
rect 206902 234051 206954 234057
rect 206902 233993 206954 233999
rect 205078 233903 205130 233909
rect 205078 233845 205130 233851
rect 205558 233903 205610 233909
rect 205558 233845 205610 233851
rect 204322 221764 204398 221792
rect 204370 221482 204398 221764
rect 205090 221482 205118 233845
rect 205954 221496 205982 233993
rect 207286 233977 207338 233983
rect 207286 233919 207338 233925
rect 207298 233465 207326 233919
rect 206614 233459 206666 233465
rect 206614 233401 206666 233407
rect 207286 233459 207338 233465
rect 207286 233401 207338 233407
rect 205920 221468 205982 221496
rect 206626 221496 206654 233401
rect 206626 221468 206688 221496
rect 207394 221482 207422 234067
rect 208450 233539 208478 239672
rect 208738 233983 208766 239672
rect 208930 235093 208958 239686
rect 209314 235167 209342 239686
rect 209302 235161 209354 235167
rect 209302 235103 209354 235109
rect 208918 235087 208970 235093
rect 208918 235029 208970 235035
rect 209698 234205 209726 239686
rect 210082 235315 210110 239686
rect 210432 239672 210686 239700
rect 210816 239672 211070 239700
rect 210658 235907 210686 239672
rect 210646 235901 210698 235907
rect 210646 235843 210698 235849
rect 211042 235537 211070 239672
rect 211234 235981 211262 239686
rect 211222 235975 211274 235981
rect 211222 235917 211274 235923
rect 211618 235685 211646 239686
rect 212002 235759 212030 239686
rect 211990 235753 212042 235759
rect 211990 235695 212042 235701
rect 211606 235679 211658 235685
rect 211606 235621 211658 235627
rect 211030 235531 211082 235537
rect 211030 235473 211082 235479
rect 210070 235309 210122 235315
rect 210070 235251 210122 235257
rect 210358 234273 210410 234279
rect 210358 234215 210410 234221
rect 208822 234199 208874 234205
rect 208822 234141 208874 234147
rect 209686 234199 209738 234205
rect 209686 234141 209738 234147
rect 208726 233977 208778 233983
rect 208726 233919 208778 233925
rect 208150 233533 208202 233539
rect 208150 233475 208202 233481
rect 208438 233533 208490 233539
rect 208438 233475 208490 233481
rect 208162 221496 208190 233475
rect 208128 221468 208190 221496
rect 208834 221496 208862 234141
rect 209686 233607 209738 233613
rect 209686 233549 209738 233555
rect 208834 221468 208896 221496
rect 209698 221482 209726 233549
rect 210370 221792 210398 234215
rect 211894 233755 211946 233761
rect 211894 233697 211946 233703
rect 211126 233311 211178 233317
rect 211126 233253 211178 233259
rect 210370 221764 210446 221792
rect 210418 221482 210446 221764
rect 211138 221482 211166 233253
rect 211906 221482 211934 233697
rect 212386 226583 212414 239686
rect 212736 239672 212990 239700
rect 212962 235833 212990 239672
rect 213058 239672 213120 239700
rect 212950 235827 213002 235833
rect 212950 235769 213002 235775
rect 212566 233681 212618 233687
rect 212566 233623 212618 233629
rect 212374 226577 212426 226583
rect 212374 226519 212426 226525
rect 212578 221792 212606 233623
rect 213058 226879 213086 239672
rect 213442 235241 213470 239686
rect 213430 235235 213482 235241
rect 213430 235177 213482 235183
rect 213430 234495 213482 234501
rect 213430 234437 213482 234443
rect 213046 226873 213098 226879
rect 213046 226815 213098 226821
rect 212578 221764 212654 221792
rect 212626 221482 212654 221764
rect 213442 221749 213470 234437
rect 213826 226805 213854 239686
rect 214210 235611 214238 239686
rect 214198 235605 214250 235611
rect 214198 235547 214250 235553
rect 214198 233385 214250 233391
rect 214198 233327 214250 233333
rect 213814 226799 213866 226805
rect 213814 226741 213866 226747
rect 213442 221717 213490 221749
rect 213462 221482 213490 221717
rect 214210 221482 214238 233327
rect 214594 226731 214622 239686
rect 215040 239672 215294 239700
rect 215424 239672 215678 239700
rect 214870 234569 214922 234575
rect 214870 234511 214922 234517
rect 214582 226725 214634 226731
rect 214582 226667 214634 226673
rect 214882 221792 214910 234511
rect 215266 229025 215294 239672
rect 215542 233829 215594 233835
rect 215542 233771 215594 233777
rect 215254 229019 215306 229025
rect 215254 228961 215306 228967
rect 215554 224160 215582 233771
rect 215650 226139 215678 239672
rect 215746 226361 215774 239686
rect 216130 226657 216158 239686
rect 216528 239672 216734 239700
rect 216864 239672 217118 239700
rect 217248 239672 217502 239700
rect 217632 239672 217886 239700
rect 217968 239672 218270 239700
rect 216502 234865 216554 234871
rect 216502 234807 216554 234813
rect 216118 226651 216170 226657
rect 216118 226593 216170 226599
rect 215734 226355 215786 226361
rect 215734 226297 215786 226303
rect 215638 226133 215690 226139
rect 215638 226075 215690 226081
rect 215554 224132 215678 224160
rect 214882 221764 214958 221792
rect 214930 221482 214958 221764
rect 215650 221482 215678 224132
rect 216514 221482 216542 234807
rect 216706 229395 216734 239672
rect 216694 229389 216746 229395
rect 216694 229331 216746 229337
rect 217090 226287 217118 239672
rect 217174 233459 217226 233465
rect 217174 233401 217226 233407
rect 217078 226281 217130 226287
rect 217078 226223 217130 226229
rect 217186 221792 217214 233401
rect 217474 226435 217502 239672
rect 217858 234575 217886 239672
rect 217942 234939 217994 234945
rect 217942 234881 217994 234887
rect 217846 234569 217898 234575
rect 217846 234511 217898 234517
rect 217462 226429 217514 226435
rect 217462 226371 217514 226377
rect 217186 221764 217262 221792
rect 217234 221482 217262 221764
rect 217954 221482 217982 234881
rect 218242 232503 218270 239672
rect 218230 232497 218282 232503
rect 218230 232439 218282 232445
rect 218338 226213 218366 239686
rect 218710 233903 218762 233909
rect 218710 233845 218762 233851
rect 218326 226207 218378 226213
rect 218326 226149 218378 226155
rect 218722 221482 218750 233845
rect 218818 225917 218846 239686
rect 219168 239672 219422 239700
rect 219552 239672 219806 239700
rect 219936 239672 220190 239700
rect 220272 239672 220382 239700
rect 219394 235389 219422 239672
rect 219382 235383 219434 235389
rect 219382 235325 219434 235331
rect 219382 234347 219434 234353
rect 219382 234289 219434 234295
rect 218806 225911 218858 225917
rect 218806 225853 218858 225859
rect 219394 221792 219422 234289
rect 219778 232577 219806 239672
rect 219766 232571 219818 232577
rect 219766 232513 219818 232519
rect 220162 229617 220190 239672
rect 220246 234051 220298 234057
rect 220246 233993 220298 233999
rect 220150 229611 220202 229617
rect 220150 229553 220202 229559
rect 220258 221804 220286 233993
rect 220354 225843 220382 239672
rect 220642 235463 220670 239686
rect 220630 235457 220682 235463
rect 220630 235399 220682 235405
rect 220918 234421 220970 234427
rect 220918 234363 220970 234369
rect 220930 227534 220958 234363
rect 221026 232429 221054 239686
rect 221376 239672 221630 239700
rect 221014 232423 221066 232429
rect 221014 232365 221066 232371
rect 221602 229469 221630 239672
rect 221746 239404 221774 239686
rect 222144 239672 222398 239700
rect 221698 239376 221774 239404
rect 221590 229463 221642 229469
rect 221590 229405 221642 229411
rect 220930 227506 221054 227534
rect 220342 225837 220394 225843
rect 220342 225779 220394 225785
rect 219394 221764 219470 221792
rect 220258 221764 220296 221804
rect 219442 221482 219470 221764
rect 220268 221482 220296 221764
rect 221026 221482 221054 227506
rect 221698 226509 221726 239376
rect 222370 234871 222398 239672
rect 222358 234865 222410 234871
rect 222358 234807 222410 234813
rect 221782 234791 221834 234797
rect 221782 234733 221834 234739
rect 221686 226503 221738 226509
rect 221686 226445 221738 226451
rect 221794 221792 221822 234733
rect 222454 234717 222506 234723
rect 222454 234659 222506 234665
rect 221746 221764 221822 221792
rect 221746 221482 221774 221764
rect 222466 221482 222494 234659
rect 222562 232355 222590 239686
rect 222550 232349 222602 232355
rect 222550 232291 222602 232297
rect 222946 229543 222974 239686
rect 223222 233533 223274 233539
rect 223222 233475 223274 233481
rect 222934 229537 222986 229543
rect 222934 229479 222986 229485
rect 223234 221949 223262 233475
rect 223330 225695 223358 239686
rect 223680 239672 223934 239700
rect 224064 239672 224318 239700
rect 223906 234797 223934 239672
rect 223894 234791 223946 234797
rect 223894 234733 223946 234739
rect 223990 234125 224042 234131
rect 223990 234067 224042 234073
rect 223318 225689 223370 225695
rect 223318 225631 223370 225637
rect 223224 221905 223262 221949
rect 223224 221482 223252 221905
rect 224002 221792 224030 234067
rect 224290 232281 224318 239672
rect 224278 232275 224330 232281
rect 224278 232217 224330 232223
rect 224386 232207 224414 239686
rect 224784 239672 224990 239700
rect 224758 233977 224810 233983
rect 224758 233919 224810 233925
rect 224374 232201 224426 232207
rect 224374 232143 224426 232149
rect 224002 221764 224078 221792
rect 224050 221482 224078 221764
rect 224770 221482 224798 233919
rect 224962 225991 224990 239672
rect 225154 235019 225182 239686
rect 225142 235013 225194 235019
rect 225142 234955 225194 234961
rect 225538 234945 225566 239686
rect 225984 239672 226238 239700
rect 226368 239672 226622 239700
rect 225526 234939 225578 234945
rect 225526 234881 225578 234887
rect 225526 234643 225578 234649
rect 225526 234585 225578 234591
rect 224950 225985 225002 225991
rect 224950 225927 225002 225933
rect 225538 221482 225566 234585
rect 226210 229321 226238 239672
rect 226294 234199 226346 234205
rect 226294 234141 226346 234147
rect 226198 229315 226250 229321
rect 226198 229257 226250 229263
rect 226306 221792 226334 234141
rect 226594 227471 226622 239672
rect 226582 227465 226634 227471
rect 226582 227407 226634 227413
rect 226690 226065 226718 239686
rect 226966 235087 227018 235093
rect 226966 235029 227018 235035
rect 226678 226059 226730 226065
rect 226678 226001 226730 226007
rect 226258 221764 226334 221792
rect 226258 221482 226286 221764
rect 226978 221482 227006 235029
rect 227074 234723 227102 239686
rect 227062 234717 227114 234723
rect 227062 234659 227114 234665
rect 227458 232133 227486 239686
rect 227856 239672 228062 239700
rect 228192 239672 228446 239700
rect 228576 239672 228830 239700
rect 227830 235309 227882 235315
rect 227830 235251 227882 235257
rect 227446 232127 227498 232133
rect 227446 232069 227498 232075
rect 227842 221482 227870 235251
rect 228034 227545 228062 239672
rect 228418 235315 228446 239672
rect 228406 235309 228458 235315
rect 228406 235251 228458 235257
rect 228502 235161 228554 235167
rect 228502 235103 228554 235109
rect 228022 227539 228074 227545
rect 228022 227481 228074 227487
rect 228514 221792 228542 235103
rect 228802 234575 228830 239672
rect 228790 234569 228842 234575
rect 228790 234511 228842 234517
rect 228898 228803 228926 239686
rect 229296 239672 229598 239700
rect 229270 235975 229322 235981
rect 229270 235917 229322 235923
rect 228886 228797 228938 228803
rect 228886 228739 228938 228745
rect 228514 221764 228590 221792
rect 228562 221482 228590 221764
rect 229282 221482 229310 235917
rect 229570 227323 229598 239672
rect 229558 227317 229610 227323
rect 229558 227259 229610 227265
rect 229762 227249 229790 239686
rect 230112 239672 230366 239700
rect 230496 239672 230750 239700
rect 230880 239672 231134 239700
rect 230038 235901 230090 235907
rect 230038 235843 230090 235849
rect 229750 227243 229802 227249
rect 229750 227185 229802 227191
rect 230050 221482 230078 235843
rect 230338 228581 230366 239672
rect 230722 236174 230750 239672
rect 230722 236146 230846 236174
rect 230710 235679 230762 235685
rect 230710 235621 230762 235627
rect 230326 228575 230378 228581
rect 230326 228517 230378 228523
rect 230722 221792 230750 235621
rect 230818 228729 230846 236146
rect 230806 228723 230858 228729
rect 230806 228665 230858 228671
rect 231106 227175 231134 239672
rect 231202 236129 231230 239686
rect 231586 236174 231614 239686
rect 231586 236146 231710 236174
rect 231190 236123 231242 236129
rect 231190 236065 231242 236071
rect 231574 235531 231626 235537
rect 231574 235473 231626 235479
rect 231094 227169 231146 227175
rect 231094 227111 231146 227117
rect 230722 221764 230798 221792
rect 230770 221482 230798 221764
rect 231586 221482 231614 235473
rect 231682 228655 231710 236146
rect 231970 229247 231998 239686
rect 232320 239672 232574 239700
rect 232704 239672 232958 239700
rect 233088 239672 233246 239700
rect 232342 235827 232394 235833
rect 232342 235769 232394 235775
rect 231958 229241 232010 229247
rect 231958 229183 232010 229189
rect 231670 228649 231722 228655
rect 231670 228591 231722 228597
rect 232354 221482 232382 235769
rect 232546 227027 232574 239672
rect 232930 235167 232958 239672
rect 233014 235753 233066 235759
rect 233014 235695 233066 235701
rect 232918 235161 232970 235167
rect 232918 235103 232970 235109
rect 232918 227391 232970 227397
rect 232918 227333 232970 227339
rect 232534 227021 232586 227027
rect 232534 226963 232586 226969
rect 232930 226065 232958 227333
rect 232918 226059 232970 226065
rect 232918 226001 232970 226007
rect 233026 221792 233054 235695
rect 233218 232059 233246 239672
rect 233506 235833 233534 239686
rect 233494 235827 233546 235833
rect 233494 235769 233546 235775
rect 233206 232053 233258 232059
rect 233206 231995 233258 232001
rect 233890 227101 233918 239686
rect 234274 235537 234302 239686
rect 234624 239672 234878 239700
rect 235008 239672 235262 239700
rect 235392 239672 235646 239700
rect 234262 235531 234314 235537
rect 234262 235473 234314 235479
rect 234850 231985 234878 239672
rect 234838 231979 234890 231985
rect 234838 231921 234890 231927
rect 235234 229173 235262 239672
rect 235318 235605 235370 235611
rect 235318 235547 235370 235553
rect 235222 229167 235274 229173
rect 235222 229109 235274 229115
rect 233878 227095 233930 227101
rect 233878 227037 233930 227043
rect 233782 226873 233834 226879
rect 233782 226815 233834 226821
rect 233026 221764 233102 221792
rect 233074 221482 233102 221764
rect 233794 221482 233822 226815
rect 234550 226577 234602 226583
rect 234550 226519 234602 226525
rect 234562 221779 234590 226519
rect 235330 221833 235358 235547
rect 235618 226953 235646 239672
rect 235714 235241 235742 239686
rect 235894 235457 235946 235463
rect 235894 235399 235946 235405
rect 235990 235457 236042 235463
rect 235990 235399 236042 235405
rect 235702 235235 235754 235241
rect 235702 235177 235754 235183
rect 235906 235093 235934 235399
rect 235798 235087 235850 235093
rect 235798 235029 235850 235035
rect 235894 235087 235946 235093
rect 235894 235029 235946 235035
rect 235810 227534 235838 235029
rect 236002 234649 236030 235399
rect 235990 234643 236042 234649
rect 235990 234585 236042 234591
rect 236098 231837 236126 239686
rect 236086 231831 236138 231837
rect 236086 231773 236138 231779
rect 235810 227506 236126 227534
rect 235606 226947 235658 226953
rect 235606 226889 235658 226895
rect 235330 221799 235378 221833
rect 234542 221743 234590 221779
rect 234542 221482 234570 221743
rect 235350 221496 235378 221799
rect 235350 221468 235392 221496
rect 236098 221482 236126 227506
rect 236482 225621 236510 239686
rect 236832 239672 237086 239700
rect 237312 239672 237470 239700
rect 236854 226725 236906 226731
rect 236854 226667 236906 226673
rect 236470 225615 236522 225621
rect 236470 225557 236522 225563
rect 236866 221496 236894 226667
rect 237058 226583 237086 239672
rect 237442 226879 237470 239672
rect 237634 231911 237662 239686
rect 238018 235833 238046 239686
rect 238006 235827 238058 235833
rect 238006 235769 238058 235775
rect 237622 231905 237674 231911
rect 237622 231847 237674 231853
rect 237430 226873 237482 226879
rect 237430 226815 237482 226821
rect 238402 226805 238430 239686
rect 237526 226799 237578 226805
rect 237526 226741 237578 226747
rect 238390 226799 238442 226805
rect 238390 226741 238442 226747
rect 237046 226577 237098 226583
rect 237046 226519 237098 226525
rect 236832 221468 236894 221496
rect 237538 221496 237566 226741
rect 238390 226355 238442 226361
rect 238390 226297 238442 226303
rect 237538 221468 237600 221496
rect 238402 221482 238430 226297
rect 238786 225769 238814 239686
rect 239136 239672 239390 239700
rect 239520 239672 239774 239700
rect 239856 239672 240158 239700
rect 239362 231319 239390 239672
rect 239350 231313 239402 231319
rect 239350 231255 239402 231261
rect 239746 229099 239774 239672
rect 239734 229093 239786 229099
rect 239734 229035 239786 229041
rect 239062 229019 239114 229025
rect 239062 228961 239114 228967
rect 238774 225763 238826 225769
rect 238774 225705 238826 225711
rect 239074 221792 239102 228961
rect 240130 226657 240158 239672
rect 239830 226651 239882 226657
rect 239830 226593 239882 226599
rect 240118 226651 240170 226657
rect 240118 226593 240170 226599
rect 239074 221764 239150 221792
rect 239122 221482 239150 221764
rect 239842 221482 239870 226593
rect 240226 226435 240254 239686
rect 240610 231541 240638 239686
rect 240694 235457 240746 235463
rect 240694 235399 240746 235405
rect 240598 231535 240650 231541
rect 240598 231477 240650 231483
rect 240214 226429 240266 226435
rect 240214 226371 240266 226377
rect 240598 226133 240650 226139
rect 240598 226075 240650 226081
rect 240610 221482 240638 226075
rect 240706 224733 240734 235399
rect 241090 228951 241118 239686
rect 241440 239672 241694 239700
rect 241666 235981 241694 239672
rect 241810 239404 241838 239686
rect 241810 239376 241886 239404
rect 241654 235975 241706 235981
rect 241654 235917 241706 235923
rect 241078 228945 241130 228951
rect 241078 228887 241130 228893
rect 241270 226355 241322 226361
rect 241270 226297 241322 226303
rect 240694 224727 240746 224733
rect 240694 224669 240746 224675
rect 241282 221792 241310 226297
rect 241858 226139 241886 239376
rect 242146 231393 242174 239686
rect 242544 239672 242846 239700
rect 242928 239672 243230 239700
rect 242134 231387 242186 231393
rect 242134 231329 242186 231335
rect 242818 229395 242846 239672
rect 242134 229389 242186 229395
rect 242134 229331 242186 229337
rect 242806 229389 242858 229395
rect 242806 229331 242858 229337
rect 241846 226133 241898 226139
rect 241846 226075 241898 226081
rect 242146 221828 242174 229331
rect 243202 228877 243230 239672
rect 243190 228871 243242 228877
rect 243190 228813 243242 228819
rect 243298 226361 243326 239686
rect 243648 239672 243902 239700
rect 244032 239672 244190 239700
rect 243874 231615 243902 239672
rect 243862 231609 243914 231615
rect 243862 231551 243914 231557
rect 244162 229025 244190 239672
rect 244354 235907 244382 239686
rect 244848 239672 245054 239700
rect 245026 236174 245054 239672
rect 244930 236146 245054 236174
rect 244342 235901 244394 235907
rect 244342 235843 244394 235849
rect 244534 235383 244586 235389
rect 244534 235325 244586 235331
rect 244150 229019 244202 229025
rect 244150 228961 244202 228967
rect 243286 226355 243338 226361
rect 243286 226297 243338 226303
rect 243574 226281 243626 226287
rect 243574 226223 243626 226229
rect 242902 224727 242954 224733
rect 242902 224669 242954 224675
rect 241282 221764 241358 221792
rect 242146 221791 242184 221828
rect 241330 221482 241358 221764
rect 242156 221482 242184 221791
rect 242914 221482 242942 224669
rect 243586 221792 243614 226223
rect 244342 225911 244394 225917
rect 244342 225853 244394 225859
rect 243586 221764 243662 221792
rect 243634 221482 243662 221764
rect 244354 221482 244382 225853
rect 244546 224733 244574 235325
rect 244930 226287 244958 236146
rect 245218 235463 245246 239686
rect 245568 239672 245726 239700
rect 245952 239672 246206 239700
rect 246336 239672 246590 239700
rect 245206 235457 245258 235463
rect 245206 235399 245258 235405
rect 245014 235087 245066 235093
rect 245014 235029 245066 235035
rect 244918 226281 244970 226287
rect 244918 226223 244970 226229
rect 245026 224807 245054 235029
rect 245110 232497 245162 232503
rect 245110 232439 245162 232445
rect 245014 224801 245066 224807
rect 245014 224743 245066 224749
rect 244534 224727 244586 224733
rect 244534 224669 244586 224675
rect 245122 221482 245150 232439
rect 245698 229765 245726 239672
rect 246178 230431 246206 239672
rect 246562 234649 246590 239672
rect 246658 235093 246686 239686
rect 246646 235087 246698 235093
rect 246646 235029 246698 235035
rect 246550 234643 246602 234649
rect 246550 234585 246602 234591
rect 246166 230425 246218 230431
rect 246166 230367 246218 230373
rect 247042 229987 247070 239686
rect 247426 234353 247454 239686
rect 247776 239672 248030 239700
rect 248160 239672 248414 239700
rect 248640 239672 248798 239700
rect 247414 234347 247466 234353
rect 247414 234289 247466 234295
rect 247030 229981 247082 229987
rect 247030 229923 247082 229929
rect 245686 229759 245738 229765
rect 245686 229701 245738 229707
rect 247714 226657 247934 226676
rect 247702 226651 247946 226657
rect 247754 226648 247894 226651
rect 247702 226593 247754 226599
rect 247894 226593 247946 226599
rect 248002 226583 248030 239672
rect 248086 232571 248138 232577
rect 248086 232513 248138 232519
rect 247990 226577 248042 226583
rect 247990 226519 248042 226525
rect 246646 226207 246698 226213
rect 246646 226149 246698 226155
rect 245878 224727 245930 224733
rect 245878 224669 245930 224675
rect 245890 221792 245918 224669
rect 245890 221764 245966 221792
rect 245938 221482 245966 221764
rect 246658 221482 246686 226149
rect 247414 225837 247466 225843
rect 247414 225779 247466 225785
rect 247426 221482 247454 225779
rect 248098 221792 248126 232513
rect 248386 231467 248414 239672
rect 248374 231461 248426 231467
rect 248374 231403 248426 231409
rect 248770 228211 248798 239672
rect 248962 230357 248990 239686
rect 249346 234501 249374 239686
rect 249730 235611 249758 239686
rect 250080 239672 250334 239700
rect 249718 235605 249770 235611
rect 249718 235547 249770 235553
rect 249334 234495 249386 234501
rect 249334 234437 249386 234443
rect 248950 230351 249002 230357
rect 248950 230293 249002 230299
rect 250306 230061 250334 239672
rect 250450 239404 250478 239686
rect 250848 239672 251102 239700
rect 250450 239376 250526 239404
rect 250498 236055 250526 239376
rect 250486 236049 250538 236055
rect 250486 235991 250538 235997
rect 250582 235013 250634 235019
rect 250582 234955 250634 234961
rect 250486 234865 250538 234871
rect 250486 234807 250538 234813
rect 250294 230055 250346 230061
rect 250294 229997 250346 230003
rect 249718 229611 249770 229617
rect 249718 229553 249770 229559
rect 248758 228205 248810 228211
rect 248758 228147 248810 228153
rect 248854 224801 248906 224807
rect 248854 224743 248906 224749
rect 248098 221764 248174 221792
rect 248146 221482 248174 221764
rect 248866 221482 248894 224743
rect 249730 221482 249758 229553
rect 250390 226503 250442 226509
rect 250390 226445 250442 226451
rect 250402 221792 250430 226445
rect 250498 224881 250526 234807
rect 250594 225769 250622 234955
rect 250774 234791 250826 234797
rect 250774 234733 250826 234739
rect 250786 226065 250814 234733
rect 250870 226355 250922 226361
rect 250870 226297 250922 226303
rect 250774 226059 250826 226065
rect 250774 226001 250826 226007
rect 250882 225843 250910 226297
rect 251074 225843 251102 239672
rect 251170 235389 251198 239686
rect 251158 235383 251210 235389
rect 251158 235325 251210 235331
rect 251158 232423 251210 232429
rect 251158 232365 251210 232371
rect 250870 225837 250922 225843
rect 250870 225779 250922 225785
rect 251062 225837 251114 225843
rect 251062 225779 251114 225785
rect 250582 225763 250634 225769
rect 250582 225705 250634 225711
rect 250486 224875 250538 224881
rect 250486 224817 250538 224823
rect 250402 221764 250478 221792
rect 250450 221482 250478 221764
rect 251170 221482 251198 232365
rect 251554 229691 251582 239686
rect 251938 230283 251966 239686
rect 252384 239672 252638 239700
rect 252768 239672 253022 239700
rect 252610 234427 252638 239672
rect 252598 234421 252650 234427
rect 252598 234363 252650 234369
rect 252994 231171 253022 239672
rect 252982 231165 253034 231171
rect 252982 231107 253034 231113
rect 251926 230277 251978 230283
rect 251926 230219 251978 230225
rect 251542 229685 251594 229691
rect 251542 229627 251594 229633
rect 252598 229463 252650 229469
rect 252598 229405 252650 229411
rect 252214 226799 252266 226805
rect 252214 226741 252266 226747
rect 252226 226583 252254 226741
rect 252406 226725 252458 226731
rect 252406 226667 252458 226673
rect 252214 226577 252266 226583
rect 252214 226519 252266 226525
rect 252418 225621 252446 226667
rect 252406 225615 252458 225621
rect 252406 225557 252458 225563
rect 251926 224875 251978 224881
rect 251926 224817 251978 224823
rect 251938 221482 251966 224817
rect 252610 221792 252638 229405
rect 253090 227989 253118 239686
rect 253474 234279 253502 239686
rect 253558 236123 253610 236129
rect 253558 236065 253610 236071
rect 253462 234273 253514 234279
rect 253462 234215 253514 234221
rect 253078 227983 253130 227989
rect 253078 227925 253130 227931
rect 253570 225695 253598 236065
rect 253858 225917 253886 239686
rect 254242 235019 254270 239686
rect 254592 239672 254846 239700
rect 254976 239672 255230 239700
rect 254230 235013 254282 235019
rect 254230 234955 254282 234961
rect 254230 232349 254282 232355
rect 254230 232291 254282 232297
rect 253846 225911 253898 225917
rect 253846 225853 253898 225859
rect 253462 225689 253514 225695
rect 253462 225631 253514 225637
rect 253558 225689 253610 225695
rect 253558 225631 253610 225637
rect 252610 221764 252686 221792
rect 252658 221482 252686 221764
rect 253474 221482 253502 225631
rect 254242 221482 254270 232291
rect 254818 229839 254846 239672
rect 255202 229913 255230 239672
rect 255298 236129 255326 239686
rect 255286 236123 255338 236129
rect 255286 236065 255338 236071
rect 255778 234797 255806 239686
rect 255766 234791 255818 234797
rect 255766 234733 255818 234739
rect 255190 229907 255242 229913
rect 255190 229849 255242 229855
rect 254806 229833 254858 229839
rect 254806 229775 254858 229781
rect 255670 229537 255722 229543
rect 255670 229479 255722 229485
rect 254902 226059 254954 226065
rect 254902 226001 254954 226007
rect 254914 221792 254942 226001
rect 254914 221764 254990 221792
rect 254962 221482 254990 221764
rect 255682 221482 255710 229479
rect 256162 229469 256190 239686
rect 256546 233539 256574 239686
rect 256896 239672 257150 239700
rect 257280 239672 257534 239700
rect 256534 233533 256586 233539
rect 256534 233475 256586 233481
rect 256150 229463 256202 229469
rect 256150 229405 256202 229411
rect 257122 225991 257150 239672
rect 257206 232275 257258 232281
rect 257206 232217 257258 232223
rect 256438 225985 256490 225991
rect 256438 225927 256490 225933
rect 257110 225985 257162 225991
rect 257110 225927 257162 225933
rect 256450 221757 256478 225927
rect 257218 221792 257246 232217
rect 257506 231689 257534 239672
rect 257494 231683 257546 231689
rect 257494 231625 257546 231631
rect 257602 229617 257630 239686
rect 257986 235759 258014 239686
rect 257974 235753 258026 235759
rect 257974 235695 258026 235701
rect 258370 233983 258398 239686
rect 258754 234871 258782 239686
rect 259104 239672 259166 239700
rect 259584 239672 259838 239700
rect 259030 235161 259082 235167
rect 259030 235103 259082 235109
rect 258742 234865 258794 234871
rect 258742 234807 258794 234813
rect 258358 233977 258410 233983
rect 258358 233919 258410 233925
rect 258742 232201 258794 232207
rect 258742 232143 258794 232149
rect 257590 229611 257642 229617
rect 257590 229553 257642 229559
rect 257974 225763 258026 225769
rect 257974 225705 258026 225711
rect 257218 221764 257294 221792
rect 256440 221726 256478 221757
rect 256440 221482 256468 221726
rect 257266 221482 257294 221764
rect 257986 221482 258014 225705
rect 258754 221482 258782 232143
rect 259042 225621 259070 235103
rect 259138 233243 259166 239672
rect 259126 233237 259178 233243
rect 259126 233179 259178 233185
rect 259810 229543 259838 239672
rect 259798 229537 259850 229543
rect 259798 229479 259850 229485
rect 259414 227465 259466 227471
rect 259414 227407 259466 227413
rect 259030 225615 259082 225621
rect 259030 225557 259082 225563
rect 259426 221792 259454 227407
rect 259906 225103 259934 239686
rect 260182 234939 260234 234945
rect 260182 234881 260234 234887
rect 259894 225097 259946 225103
rect 259894 225039 259946 225045
rect 259426 221764 259502 221792
rect 259474 221482 259502 221764
rect 260194 221482 260222 234881
rect 260290 231763 260318 239686
rect 260278 231757 260330 231763
rect 260278 231699 260330 231705
rect 260674 230579 260702 239686
rect 261024 239672 261278 239700
rect 261408 239672 261662 239700
rect 261792 239672 261950 239700
rect 261250 234057 261278 239672
rect 261238 234051 261290 234057
rect 261238 233993 261290 233999
rect 261634 233835 261662 239672
rect 261922 234945 261950 239672
rect 262006 235679 262058 235685
rect 262006 235621 262058 235627
rect 261910 234939 261962 234945
rect 261910 234881 261962 234887
rect 261622 233829 261674 233835
rect 261622 233771 261674 233777
rect 260662 230573 260714 230579
rect 260662 230515 260714 230521
rect 261718 229315 261770 229321
rect 261718 229257 261770 229263
rect 261046 227391 261098 227397
rect 261046 227333 261098 227339
rect 261058 221482 261086 227333
rect 261730 221792 261758 229257
rect 262018 228359 262046 235621
rect 262114 233095 262142 239686
rect 262512 239672 262814 239700
rect 262102 233089 262154 233095
rect 262102 233031 262154 233037
rect 262786 229321 262814 239672
rect 262882 233391 262910 239686
rect 263328 239672 263582 239700
rect 263712 239672 263966 239700
rect 264096 239672 264350 239700
rect 263254 234717 263306 234723
rect 263254 234659 263306 234665
rect 262870 233385 262922 233391
rect 262870 233327 262922 233333
rect 262774 229315 262826 229321
rect 262774 229257 262826 229263
rect 262006 228353 262058 228359
rect 262006 228295 262058 228301
rect 262486 227539 262538 227545
rect 262486 227481 262538 227487
rect 261730 221764 261806 221792
rect 261778 221482 261806 221764
rect 262498 221482 262526 227481
rect 263266 221782 263294 234659
rect 263554 233169 263582 239672
rect 263542 233163 263594 233169
rect 263542 233105 263594 233111
rect 263938 230653 263966 239672
rect 264022 235309 264074 235315
rect 264022 235251 264074 235257
rect 263926 230647 263978 230653
rect 263926 230589 263978 230595
rect 263246 221734 263294 221782
rect 264034 221778 264062 235251
rect 264322 234131 264350 239672
rect 264418 234723 264446 239686
rect 264610 239672 264816 239700
rect 264406 234717 264458 234723
rect 264406 234659 264458 234665
rect 264310 234125 264362 234131
rect 264310 234067 264362 234073
rect 264610 223623 264638 239672
rect 264694 235827 264746 235833
rect 264694 235769 264746 235775
rect 264706 228285 264734 235769
rect 264886 235531 264938 235537
rect 264886 235473 264938 235479
rect 264790 232127 264842 232133
rect 264790 232069 264842 232075
rect 264694 228279 264746 228285
rect 264694 228221 264746 228227
rect 264598 223617 264650 223623
rect 264598 223559 264650 223565
rect 264034 221745 264082 221778
rect 263246 221482 263274 221734
rect 264054 221496 264082 221745
rect 264054 221468 264096 221496
rect 264802 221482 264830 232069
rect 264898 226065 264926 235473
rect 265186 232947 265214 239686
rect 265536 239672 265790 239700
rect 265920 239672 266174 239700
rect 266304 239672 266558 239700
rect 265762 235833 265790 239672
rect 265750 235827 265802 235833
rect 265750 235769 265802 235775
rect 266146 233317 266174 239672
rect 266326 235975 266378 235981
rect 266326 235917 266378 235923
rect 266230 234569 266282 234575
rect 266230 234511 266282 234517
rect 266134 233311 266186 233317
rect 266134 233253 266186 233259
rect 265174 232941 265226 232947
rect 265174 232883 265226 232889
rect 265558 227317 265610 227323
rect 265558 227259 265610 227265
rect 264886 226059 264938 226065
rect 264886 226001 264938 226007
rect 265570 221496 265598 227259
rect 265536 221468 265598 221496
rect 266242 221496 266270 234511
rect 266338 228433 266366 235917
rect 266326 228427 266378 228433
rect 266326 228369 266378 228375
rect 266530 223697 266558 239672
rect 266626 232725 266654 239686
rect 267106 234575 267134 239686
rect 267490 235315 267518 239686
rect 267840 239672 268094 239700
rect 268224 239672 268478 239700
rect 267478 235309 267530 235315
rect 267478 235251 267530 235257
rect 267958 234643 268010 234649
rect 267958 234585 268010 234591
rect 267094 234569 267146 234575
rect 267094 234511 267146 234517
rect 266614 232719 266666 232725
rect 266614 232661 266666 232667
rect 267862 228797 267914 228803
rect 267862 228739 267914 228745
rect 266998 227243 267050 227249
rect 266998 227185 267050 227191
rect 266518 223691 266570 223697
rect 266518 223633 266570 223639
rect 266242 221468 266304 221496
rect 267010 221482 267038 227185
rect 267874 221792 267902 228739
rect 267970 227323 267998 234585
rect 267958 227317 268010 227323
rect 267958 227259 268010 227265
rect 268066 223549 268094 239672
rect 268150 235901 268202 235907
rect 268150 235843 268202 235849
rect 268162 228507 268190 235843
rect 268450 232799 268478 239672
rect 268546 234205 268574 239686
rect 268534 234199 268586 234205
rect 268534 234141 268586 234147
rect 268930 233465 268958 239686
rect 269328 239672 269630 239700
rect 269398 234347 269450 234353
rect 269398 234289 269450 234295
rect 268918 233459 268970 233465
rect 268918 233401 268970 233407
rect 268438 232793 268490 232799
rect 268438 232735 268490 232741
rect 269410 228581 269438 234289
rect 269302 228575 269354 228581
rect 269302 228517 269354 228523
rect 269398 228575 269450 228581
rect 269398 228517 269450 228523
rect 268150 228501 268202 228507
rect 268150 228443 268202 228449
rect 268534 227169 268586 227175
rect 268534 227111 268586 227117
rect 268054 223543 268106 223549
rect 268054 223485 268106 223491
rect 267826 221764 267902 221792
rect 267826 221482 267854 221764
rect 268546 221482 268574 227111
rect 269314 221482 269342 228517
rect 269602 223475 269630 239672
rect 269698 232429 269726 239686
rect 270048 239672 270302 239700
rect 270432 239672 270686 239700
rect 270274 234353 270302 239672
rect 270262 234347 270314 234353
rect 270262 234289 270314 234295
rect 269686 232423 269738 232429
rect 269686 232365 269738 232371
rect 270658 227175 270686 239672
rect 270850 236174 270878 239686
rect 270850 236146 270974 236174
rect 270838 234273 270890 234279
rect 270838 234215 270890 234221
rect 270850 228729 270878 234215
rect 270742 228723 270794 228729
rect 270742 228665 270794 228671
rect 270838 228723 270890 228729
rect 270838 228665 270890 228671
rect 270646 227169 270698 227175
rect 270646 227111 270698 227117
rect 269974 225689 270026 225695
rect 269974 225631 270026 225637
rect 269590 223469 269642 223475
rect 269590 223411 269642 223417
rect 269986 221792 270014 225631
rect 269986 221764 270062 221792
rect 270034 221482 270062 221764
rect 270754 221482 270782 228665
rect 270946 223401 270974 236146
rect 271126 235235 271178 235241
rect 271126 235177 271178 235183
rect 271030 234495 271082 234501
rect 271030 234437 271082 234443
rect 271042 225325 271070 234437
rect 271138 225843 271166 235177
rect 271234 232503 271262 239686
rect 271618 232651 271646 239686
rect 272002 235907 272030 239686
rect 272352 239672 272606 239700
rect 272736 239672 272990 239700
rect 272374 236049 272426 236055
rect 272374 235991 272426 235997
rect 271990 235901 272042 235907
rect 271990 235843 272042 235849
rect 271606 232645 271658 232651
rect 271606 232587 271658 232593
rect 271222 232497 271274 232503
rect 271222 232439 271274 232445
rect 272386 228655 272414 235991
rect 272278 228649 272330 228655
rect 272278 228591 272330 228597
rect 272374 228649 272426 228655
rect 272374 228591 272426 228597
rect 271606 227021 271658 227027
rect 271606 226963 271658 226969
rect 271126 225837 271178 225843
rect 271126 225779 271178 225785
rect 271030 225319 271082 225325
rect 271030 225261 271082 225267
rect 270934 223395 270986 223401
rect 270934 223337 270986 223343
rect 271618 221482 271646 226963
rect 272290 221792 272318 228591
rect 272578 223327 272606 239672
rect 272962 232355 272990 239672
rect 273058 234279 273086 239686
rect 273442 235537 273470 239686
rect 273840 239672 274142 239700
rect 273718 236123 273770 236129
rect 273718 236065 273770 236071
rect 273430 235531 273482 235537
rect 273430 235473 273482 235479
rect 273622 234421 273674 234427
rect 273622 234363 273674 234369
rect 273046 234273 273098 234279
rect 273046 234215 273098 234221
rect 273430 233459 273482 233465
rect 273430 233401 273482 233407
rect 272950 232349 273002 232355
rect 272950 232291 273002 232297
rect 273442 227249 273470 233401
rect 273430 227243 273482 227249
rect 273430 227185 273482 227191
rect 273046 225615 273098 225621
rect 273046 225557 273098 225563
rect 272566 223321 272618 223327
rect 272566 223263 272618 223269
rect 272290 221764 272366 221792
rect 272338 221482 272366 221764
rect 273058 221482 273086 225557
rect 273634 225473 273662 234363
rect 273730 225547 273758 236065
rect 273814 229241 273866 229247
rect 273814 229183 273866 229189
rect 273718 225541 273770 225547
rect 273718 225483 273770 225489
rect 273622 225467 273674 225473
rect 273622 225409 273674 225415
rect 273826 221482 273854 229183
rect 274114 223253 274142 239672
rect 274210 232281 274238 239686
rect 274656 239672 274910 239700
rect 275040 239672 275294 239700
rect 275376 239672 275678 239700
rect 274678 233533 274730 233539
rect 274678 233475 274730 233481
rect 274198 232275 274250 232281
rect 274198 232217 274250 232223
rect 274690 228803 274718 233475
rect 274882 232577 274910 239672
rect 275266 235241 275294 239672
rect 275254 235235 275306 235241
rect 275254 235177 275306 235183
rect 274870 232571 274922 232577
rect 274870 232513 274922 232519
rect 275350 232053 275402 232059
rect 275350 231995 275402 232001
rect 274678 228797 274730 228803
rect 274678 228739 274730 228745
rect 274486 227095 274538 227101
rect 274486 227037 274538 227043
rect 274102 223247 274154 223253
rect 274102 223189 274154 223195
rect 274498 221792 274526 227037
rect 275362 221797 275390 231995
rect 275650 224289 275678 239672
rect 275746 232133 275774 239686
rect 276130 234427 276158 239686
rect 276480 239672 276734 239700
rect 276864 239672 277118 239700
rect 277248 239672 277502 239700
rect 276118 234421 276170 234427
rect 276118 234363 276170 234369
rect 275734 232127 275786 232133
rect 275734 232069 275786 232075
rect 276706 227101 276734 239672
rect 276790 228353 276842 228359
rect 276790 228295 276842 228301
rect 276694 227095 276746 227101
rect 276694 227037 276746 227043
rect 276118 226059 276170 226065
rect 276118 226001 276170 226007
rect 275638 224283 275690 224289
rect 275638 224225 275690 224231
rect 274498 221764 274574 221792
rect 274546 221482 274574 221764
rect 275362 221762 275410 221797
rect 275382 221482 275410 221762
rect 276130 221482 276158 226001
rect 276802 221792 276830 228295
rect 277090 222661 277118 239672
rect 277474 232873 277502 239672
rect 277570 234649 277598 239686
rect 277558 234643 277610 234649
rect 277558 234585 277610 234591
rect 277954 233465 277982 239686
rect 278434 236721 278462 239686
rect 278784 239672 279038 239700
rect 279168 239672 279326 239700
rect 279552 239672 279806 239700
rect 278422 236715 278474 236721
rect 278422 236657 278474 236663
rect 278230 235457 278282 235463
rect 278230 235399 278282 235405
rect 278134 233977 278186 233983
rect 278134 233919 278186 233925
rect 277942 233459 277994 233465
rect 277942 233401 277994 233407
rect 277462 232867 277514 232873
rect 277462 232809 277514 232815
rect 277558 226947 277610 226953
rect 277558 226889 277610 226895
rect 277078 222655 277130 222661
rect 277078 222597 277130 222603
rect 276802 221764 276878 221792
rect 276850 221482 276878 221764
rect 277570 221482 277598 226889
rect 278146 225399 278174 233919
rect 278242 231097 278270 235399
rect 279010 232207 279038 239672
rect 279190 235753 279242 235759
rect 279190 235695 279242 235701
rect 278998 232201 279050 232207
rect 278998 232143 279050 232149
rect 278326 231979 278378 231985
rect 278326 231921 278378 231927
rect 278230 231091 278282 231097
rect 278230 231033 278282 231039
rect 278134 225393 278186 225399
rect 278134 225335 278186 225341
rect 278338 221482 278366 231921
rect 279202 228359 279230 235695
rect 279298 235685 279326 239672
rect 279286 235679 279338 235685
rect 279286 235621 279338 235627
rect 279670 234051 279722 234057
rect 279670 233993 279722 233999
rect 279286 233829 279338 233835
rect 279286 233771 279338 233777
rect 279190 228353 279242 228359
rect 279190 228295 279242 228301
rect 279094 225837 279146 225843
rect 279094 225779 279146 225785
rect 279106 221792 279134 225779
rect 279298 225621 279326 233771
rect 279682 227619 279710 233993
rect 279670 227613 279722 227619
rect 279670 227555 279722 227561
rect 279778 227027 279806 239672
rect 279874 236647 279902 239686
rect 279862 236641 279914 236647
rect 279862 236583 279914 236589
rect 280258 232059 280286 239686
rect 280642 234501 280670 239686
rect 280992 239672 281246 239700
rect 281376 239672 281630 239700
rect 281760 239672 282014 239700
rect 280630 234495 280682 234501
rect 280630 234437 280682 234443
rect 281218 234057 281246 239672
rect 281602 236795 281630 239672
rect 281590 236789 281642 236795
rect 281590 236731 281642 236737
rect 281206 234051 281258 234057
rect 281206 233993 281258 233999
rect 281206 233385 281258 233391
rect 281206 233327 281258 233333
rect 280918 233311 280970 233317
rect 280918 233253 280970 233259
rect 280246 232053 280298 232059
rect 280246 231995 280298 232001
rect 279862 229167 279914 229173
rect 279862 229109 279914 229115
rect 279766 227021 279818 227027
rect 279766 226963 279818 226969
rect 279286 225615 279338 225621
rect 279286 225557 279338 225563
rect 279106 221764 279182 221792
rect 279154 221482 279182 221764
rect 279874 221482 279902 229109
rect 280630 226799 280682 226805
rect 280630 226741 280682 226747
rect 280642 221482 280670 226741
rect 280930 225843 280958 233253
rect 280918 225837 280970 225843
rect 280918 225779 280970 225785
rect 281218 225695 281246 233327
rect 281986 231837 282014 239672
rect 282178 236055 282206 239686
rect 282166 236049 282218 236055
rect 282166 235991 282218 235997
rect 282358 235901 282410 235907
rect 282358 235843 282410 235849
rect 281302 231831 281354 231837
rect 281302 231773 281354 231779
rect 281974 231831 282026 231837
rect 281974 231773 282026 231779
rect 281206 225689 281258 225695
rect 281206 225631 281258 225637
rect 281314 221792 281342 231773
rect 282370 227471 282398 235843
rect 282358 227465 282410 227471
rect 282358 227407 282410 227413
rect 282562 226953 282590 239686
rect 282960 239672 283166 239700
rect 283296 239672 283550 239700
rect 283680 239672 283934 239700
rect 282550 226947 282602 226953
rect 282550 226889 282602 226895
rect 282070 226873 282122 226879
rect 282070 226815 282122 226821
rect 281314 221764 281390 221792
rect 281362 221482 281390 221764
rect 282082 221482 282110 226815
rect 282934 226725 282986 226731
rect 282934 226667 282986 226673
rect 282946 221482 282974 226667
rect 283138 222143 283166 239672
rect 283522 231985 283550 239672
rect 283906 235759 283934 239672
rect 283894 235753 283946 235759
rect 283894 235695 283946 235701
rect 283510 231979 283562 231985
rect 283510 231921 283562 231927
rect 284002 226731 284030 239686
rect 284400 239672 284702 239700
rect 284374 231905 284426 231911
rect 284374 231847 284426 231853
rect 283990 226725 284042 226731
rect 283990 226667 284042 226673
rect 283606 226577 283658 226583
rect 283606 226519 283658 226525
rect 283126 222137 283178 222143
rect 283126 222079 283178 222085
rect 283618 221792 283646 226519
rect 283618 221764 283694 221792
rect 283666 221482 283694 221764
rect 284386 221482 284414 231847
rect 284674 222291 284702 239672
rect 284770 235463 284798 239686
rect 285154 236129 285182 239686
rect 285504 239672 285758 239700
rect 285984 239672 286238 239700
rect 285142 236123 285194 236129
rect 285142 236065 285194 236071
rect 284758 235457 284810 235463
rect 284758 235399 284810 235405
rect 285730 233391 285758 239672
rect 286210 236869 286238 239672
rect 286198 236863 286250 236869
rect 286198 236805 286250 236811
rect 285718 233385 285770 233391
rect 285718 233327 285770 233333
rect 286306 229173 286334 239686
rect 286690 235981 286718 239686
rect 286678 235975 286730 235981
rect 286678 235917 286730 235923
rect 287074 233983 287102 239686
rect 287458 235907 287486 239686
rect 287808 239672 287966 239700
rect 288192 239672 288446 239700
rect 287446 235901 287498 235907
rect 287446 235843 287498 235849
rect 287062 233977 287114 233983
rect 287062 233919 287114 233925
rect 287446 231313 287498 231319
rect 287446 231255 287498 231261
rect 286294 229167 286346 229173
rect 286294 229109 286346 229115
rect 285910 228279 285962 228285
rect 285910 228221 285962 228227
rect 285142 226355 285194 226361
rect 285142 226297 285194 226303
rect 284662 222285 284714 222291
rect 284662 222227 284714 222233
rect 285154 221774 285182 226297
rect 285144 221729 285182 221774
rect 285922 221792 285950 228221
rect 286678 226651 286730 226657
rect 286678 226593 286730 226599
rect 285922 221764 285998 221792
rect 285144 221482 285172 221729
rect 285970 221482 285998 221764
rect 286690 221482 286718 226593
rect 287458 221482 287486 231255
rect 287938 229247 287966 239672
rect 287926 229241 287978 229247
rect 287926 229183 287978 229189
rect 288418 228063 288446 239672
rect 288514 233317 288542 239686
rect 288912 239672 289118 239700
rect 288502 233311 288554 233317
rect 288502 233253 288554 233259
rect 288886 229093 288938 229099
rect 288886 229035 288938 229041
rect 288406 228057 288458 228063
rect 288406 227999 288458 228005
rect 288118 226429 288170 226435
rect 288118 226371 288170 226377
rect 288130 221792 288158 226371
rect 288130 221764 288206 221792
rect 288178 221482 288206 221764
rect 288898 221482 288926 229035
rect 289090 224659 289118 239672
rect 289378 229173 289406 239686
rect 289728 239672 289982 239700
rect 290112 239672 290366 239700
rect 290496 239672 290750 239700
rect 289846 234125 289898 234131
rect 289846 234067 289898 234073
rect 289750 231609 289802 231615
rect 289750 231551 289802 231557
rect 289762 231023 289790 231551
rect 289750 231017 289802 231023
rect 289750 230959 289802 230965
rect 289366 229167 289418 229173
rect 289366 229109 289418 229115
rect 289858 228433 289886 234067
rect 289954 231541 289982 239672
rect 290338 233613 290366 239672
rect 290722 235167 290750 239672
rect 290710 235161 290762 235167
rect 290710 235103 290762 235109
rect 290326 233607 290378 233613
rect 290326 233549 290378 233555
rect 290710 233385 290762 233391
rect 290710 233327 290762 233333
rect 290422 231609 290474 231615
rect 290422 231551 290474 231557
rect 289942 231535 289994 231541
rect 289942 231477 289994 231483
rect 289750 228427 289802 228433
rect 289750 228369 289802 228375
rect 289846 228427 289898 228433
rect 289846 228369 289898 228375
rect 289078 224653 289130 224659
rect 289078 224595 289130 224601
rect 289762 221482 289790 228369
rect 290434 221792 290462 231551
rect 290722 226805 290750 233327
rect 290818 231319 290846 239686
rect 291216 239672 291518 239700
rect 290998 235827 291050 235833
rect 290998 235769 291050 235775
rect 290902 235087 290954 235093
rect 290902 235029 290954 235035
rect 290914 231393 290942 235029
rect 290902 231387 290954 231393
rect 290902 231329 290954 231335
rect 290806 231313 290858 231319
rect 290806 231255 290858 231261
rect 291010 230135 291038 235769
rect 291094 235235 291146 235241
rect 291094 235177 291146 235183
rect 290998 230129 291050 230135
rect 290998 230071 291050 230077
rect 291106 227545 291134 235177
rect 291490 228285 291518 239672
rect 291586 233391 291614 239686
rect 291936 239672 292190 239700
rect 292320 239672 292574 239700
rect 292704 239672 292958 239700
rect 291574 233385 291626 233391
rect 291574 233327 291626 233333
rect 291958 228945 292010 228951
rect 291958 228887 292010 228893
rect 291478 228279 291530 228285
rect 291478 228221 291530 228227
rect 291094 227539 291146 227545
rect 291094 227481 291146 227487
rect 290710 226799 290762 226805
rect 290710 226741 290762 226747
rect 291190 226133 291242 226139
rect 291190 226075 291242 226081
rect 290434 221764 290510 221792
rect 290482 221482 290510 221764
rect 291202 221482 291230 226075
rect 291970 221482 291998 228887
rect 292162 227767 292190 239672
rect 292546 227915 292574 239672
rect 292930 233835 292958 239672
rect 292918 233829 292970 233835
rect 292918 233771 292970 233777
rect 292822 233311 292874 233317
rect 292822 233253 292874 233259
rect 292630 228871 292682 228877
rect 292630 228813 292682 228819
rect 292534 227909 292586 227915
rect 292534 227851 292586 227857
rect 292150 227761 292202 227767
rect 292150 227703 292202 227709
rect 292642 221792 292670 228813
rect 292834 226657 292862 233253
rect 292822 226651 292874 226657
rect 292822 226593 292874 226599
rect 293122 226583 293150 239686
rect 293506 235241 293534 239686
rect 293782 235605 293834 235611
rect 293782 235547 293834 235553
rect 293494 235235 293546 235241
rect 293494 235177 293546 235183
rect 293494 231239 293546 231245
rect 293494 231181 293546 231187
rect 293110 226577 293162 226583
rect 293110 226519 293162 226525
rect 292642 221764 292718 221792
rect 292690 221482 292718 221764
rect 293506 221482 293534 231181
rect 293794 230949 293822 235547
rect 293890 231245 293918 239686
rect 294240 239672 294494 239700
rect 294624 239672 294878 239700
rect 295008 239672 295262 239700
rect 294466 235833 294494 239672
rect 294454 235827 294506 235833
rect 294454 235769 294506 235775
rect 293974 234199 294026 234205
rect 293974 234141 294026 234147
rect 293878 231239 293930 231245
rect 293878 231181 293930 231187
rect 293782 230943 293834 230949
rect 293782 230885 293834 230891
rect 293986 227693 294014 234141
rect 294454 233459 294506 233465
rect 294454 233401 294506 233407
rect 293974 227687 294026 227693
rect 293974 227629 294026 227635
rect 294466 227397 294494 233401
rect 294454 227391 294506 227397
rect 294454 227333 294506 227339
rect 294850 226435 294878 239672
rect 294934 229389 294986 229395
rect 294934 229331 294986 229337
rect 294838 226429 294890 226435
rect 294838 226371 294890 226377
rect 294262 226281 294314 226287
rect 294262 226223 294314 226229
rect 294274 221496 294302 226223
rect 294240 221468 294302 221496
rect 294946 221496 294974 229331
rect 295234 226287 295262 239672
rect 295330 228877 295358 239686
rect 295714 234205 295742 239686
rect 296098 235093 296126 239686
rect 296448 239672 296606 239700
rect 296928 239672 297182 239700
rect 296086 235087 296138 235093
rect 296086 235029 296138 235035
rect 295702 234199 295754 234205
rect 295702 234141 295754 234147
rect 295606 232867 295658 232873
rect 295606 232809 295658 232815
rect 295618 232207 295646 232809
rect 295510 232201 295562 232207
rect 295510 232143 295562 232149
rect 295606 232201 295658 232207
rect 295606 232143 295658 232149
rect 295522 231985 295550 232143
rect 295510 231979 295562 231985
rect 295510 231921 295562 231927
rect 296470 231017 296522 231023
rect 296470 230959 296522 230965
rect 295318 228871 295370 228877
rect 295318 228813 295370 228819
rect 295702 228501 295754 228507
rect 295702 228443 295754 228449
rect 295222 226281 295274 226287
rect 295222 226223 295274 226229
rect 294946 221468 295008 221496
rect 295714 221482 295742 228443
rect 296482 221785 296510 230959
rect 296578 229395 296606 239672
rect 297154 231615 297182 239672
rect 297250 233391 297278 239686
rect 297238 233385 297290 233391
rect 297238 233327 297290 233333
rect 297142 231609 297194 231615
rect 297142 231551 297194 231557
rect 296566 229389 296618 229395
rect 296566 229331 296618 229337
rect 297634 226361 297662 239686
rect 298018 235611 298046 239686
rect 298006 235605 298058 235611
rect 298006 235547 298058 235553
rect 298198 234569 298250 234575
rect 298198 234511 298250 234517
rect 298210 230209 298238 234511
rect 298198 230203 298250 230209
rect 298198 230145 298250 230151
rect 298006 229019 298058 229025
rect 298006 228961 298058 228967
rect 297622 226355 297674 226361
rect 297622 226297 297674 226303
rect 297238 226207 297290 226213
rect 297238 226149 297290 226155
rect 296462 221751 296510 221785
rect 297250 221804 297278 226149
rect 297250 221752 297298 221804
rect 296462 221496 296490 221751
rect 296448 221468 296490 221496
rect 297270 221482 297298 221752
rect 298018 221482 298046 228961
rect 298402 228951 298430 239686
rect 298752 239672 299006 239700
rect 299136 239672 299390 239700
rect 298978 234131 299006 239672
rect 299254 235383 299306 235389
rect 299254 235325 299306 235331
rect 298966 234125 299018 234131
rect 298966 234067 299018 234073
rect 299266 230727 299294 235325
rect 299362 233909 299390 239672
rect 299350 233903 299402 233909
rect 299350 233845 299402 233851
rect 299458 231264 299486 239686
rect 299842 233761 299870 239686
rect 299830 233755 299882 233761
rect 299830 233697 299882 233703
rect 299458 231236 299582 231264
rect 299554 231097 299582 231236
rect 299446 231091 299498 231097
rect 299446 231033 299498 231039
rect 299542 231091 299594 231097
rect 299542 231033 299594 231039
rect 299254 230721 299306 230727
rect 299254 230663 299306 230669
rect 298678 230425 298730 230431
rect 298678 230367 298730 230373
rect 298390 228945 298442 228951
rect 298390 228887 298442 228893
rect 298690 221792 298718 230367
rect 298690 221764 298766 221792
rect 298738 221482 298766 221764
rect 299458 221482 299486 231033
rect 300226 230431 300254 239686
rect 300720 239672 300926 239700
rect 301056 239672 301214 239700
rect 301440 239672 301694 239700
rect 300790 234051 300842 234057
rect 300790 233993 300842 233999
rect 300214 230425 300266 230431
rect 300214 230367 300266 230373
rect 300802 227323 300830 233993
rect 300214 227317 300266 227323
rect 300214 227259 300266 227265
rect 300790 227317 300842 227323
rect 300790 227259 300842 227265
rect 300226 221482 300254 227259
rect 300898 226139 300926 239672
rect 300982 229759 301034 229765
rect 300982 229701 301034 229707
rect 300886 226133 300938 226139
rect 300886 226075 300938 226081
rect 300994 221792 301022 229701
rect 301186 227841 301214 239672
rect 301666 233317 301694 239672
rect 301762 236943 301790 239686
rect 301750 236937 301802 236943
rect 301750 236879 301802 236885
rect 301558 233311 301610 233317
rect 301558 233253 301610 233259
rect 301654 233311 301706 233317
rect 301654 233253 301706 233259
rect 301174 227835 301226 227841
rect 301174 227777 301226 227783
rect 301570 226879 301598 233253
rect 301750 228575 301802 228581
rect 301750 228517 301802 228523
rect 301558 226873 301610 226879
rect 301558 226815 301610 226821
rect 300994 221764 301070 221792
rect 301042 221482 301070 221764
rect 301762 221482 301790 228517
rect 302146 226213 302174 239686
rect 302544 239672 302846 239700
rect 302518 231387 302570 231393
rect 302518 231329 302570 231335
rect 302134 226207 302186 226213
rect 302134 226149 302186 226155
rect 302530 221482 302558 231329
rect 302818 222439 302846 239672
rect 302914 228475 302942 239686
rect 303264 239672 303518 239700
rect 303648 239672 303902 239700
rect 303984 239672 304286 239700
rect 303490 234575 303518 239672
rect 303478 234569 303530 234575
rect 303478 234511 303530 234517
rect 303574 234199 303626 234205
rect 303574 234141 303626 234147
rect 302900 228466 302956 228475
rect 302900 228401 302956 228410
rect 303586 228137 303614 234141
rect 303574 228131 303626 228137
rect 303574 228073 303626 228079
rect 303190 226503 303242 226509
rect 303190 226445 303242 226451
rect 302806 222433 302858 222439
rect 302806 222375 302858 222381
rect 303202 221792 303230 226445
rect 303874 225177 303902 239672
rect 303958 229981 304010 229987
rect 303958 229923 304010 229929
rect 303862 225171 303914 225177
rect 303862 225113 303914 225119
rect 303202 221764 303278 221792
rect 303250 221482 303278 221764
rect 303970 221482 303998 229923
rect 304258 226509 304286 239672
rect 304342 234347 304394 234353
rect 304342 234289 304394 234295
rect 304354 229987 304382 234289
rect 304450 233539 304478 239686
rect 304834 237017 304862 239686
rect 305184 239672 305246 239700
rect 305568 239672 305822 239700
rect 305952 239672 306206 239700
rect 306288 239672 306590 239700
rect 304822 237011 304874 237017
rect 304822 236953 304874 236959
rect 305110 235013 305162 235019
rect 305110 234955 305162 234961
rect 304438 233533 304490 233539
rect 304438 233475 304490 233481
rect 305122 230505 305150 234955
rect 305218 233687 305246 239672
rect 305794 236174 305822 239672
rect 305794 236146 305918 236174
rect 305782 234791 305834 234797
rect 305782 234733 305834 234739
rect 305206 233681 305258 233687
rect 305206 233623 305258 233629
rect 305494 231461 305546 231467
rect 305494 231403 305546 231409
rect 305110 230499 305162 230505
rect 305110 230441 305162 230447
rect 304822 230351 304874 230357
rect 304822 230293 304874 230299
rect 304342 229981 304394 229987
rect 304342 229923 304394 229929
rect 304246 226503 304298 226509
rect 304246 226445 304298 226451
rect 304834 221482 304862 230293
rect 305506 221792 305534 231403
rect 305794 230875 305822 234733
rect 305782 230869 305834 230875
rect 305782 230811 305834 230817
rect 305890 222365 305918 236146
rect 306178 228507 306206 239672
rect 306166 228501 306218 228507
rect 306166 228443 306218 228449
rect 306262 225319 306314 225325
rect 306262 225261 306314 225267
rect 305878 222359 305930 222365
rect 305878 222301 305930 222307
rect 305506 221764 305582 221792
rect 305554 221482 305582 221764
rect 306274 221482 306302 225261
rect 306562 222513 306590 239672
rect 306658 236174 306686 239686
rect 307042 237091 307070 239686
rect 307392 239672 307646 239700
rect 307776 239672 307934 239700
rect 308256 239672 308510 239700
rect 308592 239672 308894 239700
rect 307030 237085 307082 237091
rect 307030 237027 307082 237033
rect 306658 236146 306782 236174
rect 306646 234273 306698 234279
rect 306646 234215 306698 234221
rect 306658 229765 306686 234215
rect 306646 229759 306698 229765
rect 306646 229701 306698 229707
rect 306646 229241 306698 229247
rect 306646 229183 306698 229189
rect 306658 229025 306686 229183
rect 306646 229019 306698 229025
rect 306646 228961 306698 228967
rect 306754 225251 306782 236146
rect 307618 231393 307646 239672
rect 307606 231387 307658 231393
rect 307606 231329 307658 231335
rect 307702 228649 307754 228655
rect 307702 228591 307754 228597
rect 307030 228205 307082 228211
rect 307030 228147 307082 228153
rect 306742 225245 306794 225251
rect 306742 225187 306794 225193
rect 306550 222507 306602 222513
rect 306550 222449 306602 222455
rect 307042 221482 307070 228147
rect 307714 221792 307742 228591
rect 307906 222587 307934 239672
rect 308182 234865 308234 234871
rect 308182 234807 308234 234813
rect 308194 230949 308222 234807
rect 308482 234205 308510 239672
rect 308470 234199 308522 234205
rect 308470 234141 308522 234147
rect 308182 230943 308234 230949
rect 308182 230885 308234 230891
rect 308566 230795 308618 230801
rect 308566 230737 308618 230743
rect 307894 222581 307946 222587
rect 307894 222523 307946 222529
rect 307714 221764 307790 221792
rect 307762 221482 307790 221764
rect 308578 221773 308606 230737
rect 308866 222809 308894 239672
rect 308962 228581 308990 239686
rect 309346 234797 309374 239686
rect 309696 239672 309950 239700
rect 310080 239672 310334 239700
rect 310464 239672 310718 239700
rect 309334 234791 309386 234797
rect 309334 234733 309386 234739
rect 308950 228575 309002 228581
rect 308950 228517 309002 228523
rect 309334 225763 309386 225769
rect 309334 225705 309386 225711
rect 308854 222803 308906 222809
rect 308854 222745 308906 222751
rect 308578 221741 308616 221773
rect 308588 221482 308616 221741
rect 309346 221482 309374 225705
rect 309922 225325 309950 239672
rect 310198 233311 310250 233317
rect 310198 233253 310250 233259
rect 310006 230055 310058 230061
rect 310006 229997 310058 230003
rect 309910 225319 309962 225325
rect 309910 225261 309962 225267
rect 310018 221792 310046 229997
rect 310210 228211 310238 233253
rect 310198 228205 310250 228211
rect 310198 228147 310250 228153
rect 310306 222883 310334 239672
rect 310690 228623 310718 239672
rect 310786 237165 310814 239686
rect 310774 237159 310826 237165
rect 310774 237101 310826 237107
rect 311062 234939 311114 234945
rect 311062 234881 311114 234887
rect 311074 231023 311102 234881
rect 311170 234057 311198 239686
rect 311554 235389 311582 239686
rect 312000 239672 312254 239700
rect 312384 239672 312638 239700
rect 312720 239672 313022 239700
rect 311542 235383 311594 235389
rect 311542 235325 311594 235331
rect 311158 234051 311210 234057
rect 311158 233993 311210 233999
rect 312226 231467 312254 239672
rect 312214 231461 312266 231467
rect 312214 231403 312266 231409
rect 311062 231017 311114 231023
rect 311062 230959 311114 230965
rect 311638 230721 311690 230727
rect 311638 230663 311690 230669
rect 310774 230277 310826 230283
rect 310774 230219 310826 230225
rect 310676 228614 310732 228623
rect 310676 228549 310732 228558
rect 310294 222877 310346 222883
rect 310294 222819 310346 222825
rect 310018 221764 310094 221792
rect 310066 221482 310094 221764
rect 310786 221482 310814 230219
rect 311650 221482 311678 230663
rect 312310 225467 312362 225473
rect 312310 225409 312362 225415
rect 312322 221792 312350 225409
rect 312610 222735 312638 239672
rect 312694 233385 312746 233391
rect 312694 233327 312746 233333
rect 312706 229025 312734 233327
rect 312694 229019 312746 229025
rect 312694 228961 312746 228967
rect 312994 225473 313022 239672
rect 313090 234945 313118 239686
rect 313078 234939 313130 234945
rect 313078 234881 313130 234887
rect 313270 230425 313322 230431
rect 313270 230367 313322 230373
rect 313282 229765 313310 230367
rect 313270 229759 313322 229765
rect 313270 229701 313322 229707
rect 313078 229685 313130 229691
rect 313078 229627 313130 229633
rect 312982 225467 313034 225473
rect 312982 225409 313034 225415
rect 312598 222729 312650 222735
rect 312598 222671 312650 222677
rect 312322 221764 312398 221792
rect 312370 221482 312398 221764
rect 313090 221482 313118 229627
rect 313474 228655 313502 239686
rect 313858 237239 313886 239686
rect 314208 239672 314462 239700
rect 314592 239672 314846 239700
rect 313846 237233 313898 237239
rect 313846 237175 313898 237181
rect 313942 234421 313994 234427
rect 313942 234363 313994 234369
rect 313954 230061 313982 234363
rect 314434 234353 314462 239672
rect 314818 237313 314846 239672
rect 314806 237307 314858 237313
rect 314806 237249 314858 237255
rect 314422 234347 314474 234353
rect 314422 234289 314474 234295
rect 314518 231165 314570 231171
rect 314518 231107 314570 231113
rect 313942 230055 313994 230061
rect 313942 229997 313994 230003
rect 313846 228723 313898 228729
rect 313846 228665 313898 228671
rect 313462 228649 313514 228655
rect 313462 228591 313514 228597
rect 313858 221482 313886 228665
rect 314530 221792 314558 231107
rect 314914 228771 314942 239686
rect 314900 228762 314956 228771
rect 314900 228697 314956 228706
rect 315298 222957 315326 239686
rect 315778 233465 315806 239686
rect 316176 239672 316382 239700
rect 316512 239672 316766 239700
rect 316896 239672 317150 239700
rect 315766 233459 315818 233465
rect 315766 233401 315818 233407
rect 316246 229019 316298 229025
rect 316246 228961 316298 228967
rect 316258 227989 316286 228961
rect 316150 227983 316202 227989
rect 316150 227925 316202 227931
rect 316246 227983 316298 227989
rect 316246 227925 316298 227931
rect 315382 225911 315434 225917
rect 315382 225853 315434 225859
rect 315286 222951 315338 222957
rect 315286 222893 315338 222899
rect 314530 221764 314606 221792
rect 314578 221482 314606 221764
rect 315394 221482 315422 225853
rect 316162 221482 316190 227925
rect 316354 223031 316382 239672
rect 316738 231287 316766 239672
rect 317122 234871 317150 239672
rect 317110 234865 317162 234871
rect 317110 234807 317162 234813
rect 317218 234279 317246 239686
rect 317602 237387 317630 239686
rect 317590 237381 317642 237387
rect 317590 237323 317642 237329
rect 317206 234273 317258 234279
rect 317206 234215 317258 234221
rect 316724 231278 316780 231287
rect 316724 231213 316780 231222
rect 317590 230499 317642 230505
rect 317590 230441 317642 230447
rect 316822 229907 316874 229913
rect 316822 229849 316874 229855
rect 316342 223025 316394 223031
rect 316342 222967 316394 222973
rect 316834 221792 316862 229849
rect 316834 221764 316910 221792
rect 316882 221482 316910 221764
rect 317602 221482 317630 230441
rect 317986 229913 318014 239686
rect 318370 235019 318398 239686
rect 318720 239672 318974 239700
rect 319200 239672 319454 239700
rect 318358 235013 318410 235019
rect 318358 234955 318410 234961
rect 318166 234643 318218 234649
rect 318166 234585 318218 234591
rect 318178 230727 318206 234585
rect 318166 230721 318218 230727
rect 318166 230663 318218 230669
rect 317974 229907 318026 229913
rect 317974 229849 318026 229855
rect 318946 225547 318974 239672
rect 319126 229833 319178 229839
rect 319126 229775 319178 229781
rect 318358 225541 318410 225547
rect 318358 225483 318410 225489
rect 318934 225541 318986 225547
rect 318934 225483 318986 225489
rect 318370 221832 318398 225483
rect 318350 221800 318398 221832
rect 318350 221482 318378 221800
rect 319138 221792 319166 229775
rect 319426 223105 319454 239672
rect 319522 231435 319550 239686
rect 319906 234723 319934 239686
rect 319606 234717 319658 234723
rect 319606 234659 319658 234665
rect 319894 234717 319946 234723
rect 319894 234659 319946 234665
rect 319508 231426 319564 231435
rect 319508 231361 319564 231370
rect 319618 225769 319646 234659
rect 320290 234427 320318 239686
rect 320640 239672 320894 239700
rect 321024 239672 321278 239700
rect 321408 239672 321662 239700
rect 320866 237461 320894 239672
rect 320854 237455 320906 237461
rect 320854 237397 320906 237403
rect 320278 234421 320330 234427
rect 320278 234363 320330 234369
rect 321142 233977 321194 233983
rect 321142 233919 321194 233925
rect 320662 230869 320714 230875
rect 320662 230811 320714 230817
rect 319894 228797 319946 228803
rect 319894 228739 319946 228745
rect 319606 225763 319658 225769
rect 319606 225705 319658 225711
rect 319414 223099 319466 223105
rect 319414 223041 319466 223047
rect 319138 221764 319214 221792
rect 319186 221482 319214 221764
rect 319906 221482 319934 228739
rect 320674 221482 320702 230811
rect 321154 225991 321182 233919
rect 321250 228729 321278 239672
rect 321634 230117 321662 239672
rect 321730 233391 321758 239686
rect 322128 239672 322334 239700
rect 322198 234495 322250 234501
rect 322198 234437 322250 234443
rect 321718 233385 321770 233391
rect 321718 233327 321770 233333
rect 322210 230505 322238 234437
rect 322198 230499 322250 230505
rect 322198 230441 322250 230447
rect 321634 230089 321758 230117
rect 321622 230055 321674 230061
rect 321622 229997 321674 230003
rect 321430 229537 321482 229543
rect 321430 229479 321482 229485
rect 321442 229321 321470 229479
rect 321634 229469 321662 229997
rect 321622 229463 321674 229469
rect 321622 229405 321674 229411
rect 321334 229315 321386 229321
rect 321334 229257 321386 229263
rect 321430 229315 321482 229321
rect 321430 229257 321482 229263
rect 321346 228951 321374 229257
rect 321334 228945 321386 228951
rect 321334 228887 321386 228893
rect 321238 228723 321290 228729
rect 321238 228665 321290 228671
rect 321334 226059 321386 226065
rect 321334 226001 321386 226007
rect 321142 225985 321194 225991
rect 321142 225927 321194 225933
rect 321346 221792 321374 226001
rect 321730 223179 321758 230089
rect 322102 229537 322154 229543
rect 322102 229479 322154 229485
rect 321718 223173 321770 223179
rect 321718 223115 321770 223121
rect 321346 221764 321422 221792
rect 321394 221482 321422 221764
rect 322114 221482 322142 229479
rect 322306 224585 322334 239672
rect 322498 236174 322526 239686
rect 322944 239672 323198 239700
rect 323328 239672 323582 239700
rect 323712 239672 323966 239700
rect 323170 237535 323198 239672
rect 323158 237529 323210 237535
rect 323158 237471 323210 237477
rect 322402 236146 322526 236174
rect 322402 228803 322430 236146
rect 322486 235679 322538 235685
rect 322486 235621 322538 235627
rect 322498 232873 322526 235621
rect 323446 234939 323498 234945
rect 323446 234881 323498 234887
rect 322486 232867 322538 232873
rect 322486 232809 322538 232815
rect 323458 229839 323486 234881
rect 323554 234501 323582 239672
rect 323938 239015 323966 239672
rect 323926 239009 323978 239015
rect 323926 238951 323978 238957
rect 323542 234495 323594 234501
rect 323542 234437 323594 234443
rect 323638 231683 323690 231689
rect 323638 231625 323690 231631
rect 323446 229833 323498 229839
rect 323446 229775 323498 229781
rect 322390 228797 322442 228803
rect 322390 228739 322442 228745
rect 322966 228353 323018 228359
rect 322966 228295 323018 228301
rect 322294 224579 322346 224585
rect 322294 224521 322346 224527
rect 322978 221496 323006 228295
rect 322944 221468 323006 221496
rect 323650 221496 323678 231625
rect 324034 231583 324062 239686
rect 324418 234945 324446 239686
rect 324406 234939 324458 234945
rect 324406 234881 324458 234887
rect 324020 231574 324076 231583
rect 324020 231509 324076 231518
rect 324802 225515 324830 239686
rect 325152 239672 325310 239700
rect 325536 239672 325790 239700
rect 325920 239672 326174 239700
rect 325282 236174 325310 239672
rect 325090 236146 325310 236174
rect 324788 225506 324844 225515
rect 324788 225441 324844 225450
rect 324406 225393 324458 225399
rect 324406 225335 324458 225341
rect 323650 221468 323712 221496
rect 324418 221482 324446 225335
rect 325090 224511 325118 236146
rect 325366 236049 325418 236055
rect 325366 235991 325418 235997
rect 325270 235383 325322 235389
rect 325270 235325 325322 235331
rect 325174 233607 325226 233613
rect 325174 233549 325226 233555
rect 325186 233317 325214 233549
rect 325174 233311 325226 233317
rect 325174 233253 325226 233259
rect 325282 229617 325310 235325
rect 325378 233021 325406 235991
rect 325462 233829 325514 233835
rect 325462 233771 325514 233777
rect 325474 233613 325502 233771
rect 325462 233607 325514 233613
rect 325462 233549 325514 233555
rect 325366 233015 325418 233021
rect 325366 232957 325418 232963
rect 325762 230431 325790 239672
rect 325846 235753 325898 235759
rect 325846 235695 325898 235701
rect 325858 230801 325886 235695
rect 326146 233983 326174 239672
rect 326242 234649 326270 239686
rect 326722 238867 326750 239686
rect 326710 238861 326762 238867
rect 326710 238803 326762 238809
rect 326806 236123 326858 236129
rect 326806 236065 326858 236071
rect 326230 234643 326282 234649
rect 326230 234585 326282 234591
rect 326134 233977 326186 233983
rect 326134 233919 326186 233925
rect 326818 230949 326846 236065
rect 326902 233311 326954 233317
rect 326902 233253 326954 233259
rect 326710 230943 326762 230949
rect 326710 230885 326762 230891
rect 326806 230943 326858 230949
rect 326806 230885 326858 230891
rect 325846 230795 325898 230801
rect 325846 230737 325898 230743
rect 325750 230425 325802 230431
rect 325750 230367 325802 230373
rect 325174 229611 325226 229617
rect 325174 229553 325226 229559
rect 325270 229611 325322 229617
rect 325270 229553 325322 229559
rect 325078 224505 325130 224511
rect 325078 224447 325130 224453
rect 325186 221496 325214 229553
rect 325846 229315 325898 229321
rect 325846 229257 325898 229263
rect 325152 221468 325214 221496
rect 325858 221496 325886 229257
rect 325858 221468 325920 221496
rect 326722 221482 326750 230885
rect 326914 226065 326942 233253
rect 327106 231731 327134 239686
rect 327456 239672 327710 239700
rect 327840 239672 328094 239700
rect 327682 238941 327710 239672
rect 327670 238935 327722 238941
rect 327670 238877 327722 238883
rect 327092 231722 327148 231731
rect 327092 231657 327148 231666
rect 326902 226059 326954 226065
rect 326902 226001 326954 226007
rect 328066 225663 328094 239672
rect 328162 236174 328190 239686
rect 328162 236146 328286 236174
rect 328150 233237 328202 233243
rect 328150 233179 328202 233185
rect 328052 225654 328108 225663
rect 328052 225589 328108 225598
rect 327382 225097 327434 225103
rect 327382 225039 327434 225045
rect 327394 221792 327422 225039
rect 327394 221764 327470 221792
rect 327442 221482 327470 221764
rect 328162 221482 328190 233179
rect 328258 224363 328286 236146
rect 328342 235309 328394 235315
rect 328342 235251 328394 235257
rect 328354 225103 328382 235251
rect 328546 229543 328574 239686
rect 328930 235759 328958 239686
rect 328918 235753 328970 235759
rect 328918 235695 328970 235701
rect 329314 233317 329342 239686
rect 329664 239672 329918 239700
rect 330048 239672 330302 239700
rect 329890 238793 329918 239672
rect 329878 238787 329930 238793
rect 329878 238729 329930 238735
rect 329302 233311 329354 233317
rect 329302 233253 329354 233259
rect 329590 231757 329642 231763
rect 329590 231699 329642 231705
rect 328534 229537 328586 229543
rect 328534 229479 328586 229485
rect 328918 227613 328970 227619
rect 328918 227555 328970 227561
rect 328342 225097 328394 225103
rect 328342 225039 328394 225045
rect 328246 224357 328298 224363
rect 328246 224299 328298 224305
rect 328930 221482 328958 227555
rect 329602 221792 329630 231699
rect 330274 230357 330302 239672
rect 330466 235315 330494 239686
rect 330454 235309 330506 235315
rect 330454 235251 330506 235257
rect 330262 230351 330314 230357
rect 330262 230293 330314 230299
rect 330850 225811 330878 239686
rect 331248 239672 331550 239700
rect 331126 235975 331178 235981
rect 331126 235917 331178 235923
rect 331138 230672 331166 235917
rect 331138 230644 331358 230672
rect 331330 230579 331358 230644
rect 331222 230573 331274 230579
rect 331222 230515 331274 230521
rect 331318 230573 331370 230579
rect 331318 230515 331370 230521
rect 330836 225802 330892 225811
rect 330836 225737 330892 225746
rect 330454 225615 330506 225621
rect 330454 225557 330506 225563
rect 330466 221824 330494 225557
rect 329602 221764 329678 221792
rect 330466 221790 330514 221824
rect 329650 221482 329678 221764
rect 330486 221482 330514 221790
rect 331234 221482 331262 230515
rect 331522 224437 331550 239672
rect 331618 233243 331646 239686
rect 331968 239672 332222 239700
rect 332352 239672 332606 239700
rect 332194 235389 332222 239672
rect 332182 235383 332234 235389
rect 332182 235325 332234 235331
rect 332086 233385 332138 233391
rect 332086 233327 332138 233333
rect 331606 233237 331658 233243
rect 331606 233179 331658 233185
rect 331894 228945 331946 228951
rect 331894 228887 331946 228893
rect 331510 224431 331562 224437
rect 331510 224373 331562 224379
rect 331906 221792 331934 228887
rect 332098 225399 332126 233327
rect 332468 228910 332524 228919
rect 332468 228845 332470 228854
rect 332522 228845 332524 228854
rect 332470 228813 332522 228819
rect 332578 225959 332606 239672
rect 332674 238719 332702 239686
rect 332662 238713 332714 238719
rect 332662 238655 332714 238661
rect 332662 231017 332714 231023
rect 332662 230959 332714 230965
rect 332564 225950 332620 225959
rect 332564 225885 332620 225894
rect 332086 225393 332138 225399
rect 332086 225335 332138 225341
rect 331906 221764 331982 221792
rect 331954 221482 331982 221764
rect 332674 221482 332702 230959
rect 333058 229321 333086 239686
rect 333442 233391 333470 239686
rect 333826 236055 333854 239686
rect 334272 239672 334526 239700
rect 334656 239672 334910 239700
rect 333814 236049 333866 236055
rect 333814 235991 333866 235997
rect 334006 233533 334058 233539
rect 334006 233475 334058 233481
rect 333430 233385 333482 233391
rect 333430 233327 333482 233333
rect 334018 231171 334046 233475
rect 334198 233089 334250 233095
rect 334198 233031 334250 233037
rect 334294 233089 334346 233095
rect 334294 233031 334346 233037
rect 334006 231165 334058 231171
rect 334006 231107 334058 231113
rect 333046 229315 333098 229321
rect 333046 229257 333098 229263
rect 333526 225689 333578 225695
rect 333526 225631 333578 225637
rect 333538 221482 333566 225631
rect 334210 221792 334238 233031
rect 334306 232799 334334 233031
rect 334294 232793 334346 232799
rect 334294 232735 334346 232741
rect 334498 224141 334526 239672
rect 334882 231689 334910 239672
rect 334978 233761 335006 239686
rect 334966 233755 335018 233761
rect 334966 233697 335018 233703
rect 334870 231683 334922 231689
rect 334870 231625 334922 231631
rect 334966 228427 335018 228433
rect 334966 228369 335018 228375
rect 334486 224135 334538 224141
rect 334486 224077 334538 224083
rect 334210 221764 334286 221792
rect 334258 221482 334286 221764
rect 334978 221482 335006 228369
rect 335362 227439 335390 239686
rect 335746 238645 335774 239686
rect 336096 239672 336254 239700
rect 336480 239672 336734 239700
rect 335734 238639 335786 238645
rect 335734 238581 335786 238587
rect 335734 233163 335786 233169
rect 335734 233105 335786 233111
rect 335446 232941 335498 232947
rect 335446 232883 335498 232889
rect 335348 227430 335404 227439
rect 335348 227365 335404 227374
rect 335458 225917 335486 232883
rect 335446 225911 335498 225917
rect 335446 225853 335498 225859
rect 335746 221482 335774 233105
rect 336226 230283 336254 239672
rect 336502 235531 336554 235537
rect 336502 235473 336554 235479
rect 336310 233607 336362 233613
rect 336310 233549 336362 233555
rect 336322 230875 336350 233549
rect 336310 230869 336362 230875
rect 336310 230811 336362 230817
rect 336214 230277 336266 230283
rect 336214 230219 336266 230225
rect 336514 225769 336542 235473
rect 336706 233539 336734 239672
rect 336802 239672 336864 239700
rect 336802 236171 336830 239672
rect 336788 236162 336844 236171
rect 336788 236097 336844 236106
rect 336694 233533 336746 233539
rect 336694 233475 336746 233481
rect 336406 225763 336458 225769
rect 336406 225705 336458 225711
rect 336502 225763 336554 225769
rect 336502 225705 336554 225711
rect 336418 221792 336446 225705
rect 337186 224215 337214 239686
rect 337270 230647 337322 230653
rect 337270 230589 337322 230595
rect 337174 224209 337226 224215
rect 337174 224151 337226 224157
rect 337282 221799 337310 230589
rect 337570 230061 337598 239686
rect 338064 239672 338174 239700
rect 338400 239672 338654 239700
rect 338784 239672 339038 239700
rect 339168 239672 339422 239700
rect 337942 233163 337994 233169
rect 337942 233105 337994 233111
rect 337954 232355 337982 233105
rect 338038 232941 338090 232947
rect 338038 232883 338090 232889
rect 338050 232503 338078 232883
rect 338038 232497 338090 232503
rect 338038 232439 338090 232445
rect 337942 232349 337994 232355
rect 337942 232291 337994 232297
rect 338038 230129 338090 230135
rect 338038 230071 338090 230077
rect 337558 230055 337610 230061
rect 337558 229997 337610 230003
rect 336418 221764 336494 221792
rect 337282 221764 337320 221799
rect 336466 221482 336494 221764
rect 337292 221482 337320 221764
rect 338050 221482 338078 230071
rect 338146 224067 338174 239672
rect 338518 235827 338570 235833
rect 338518 235769 338570 235775
rect 338326 235605 338378 235611
rect 338326 235547 338378 235553
rect 338338 233687 338366 235547
rect 338326 233681 338378 233687
rect 338326 233623 338378 233629
rect 338230 232719 338282 232725
rect 338230 232661 338282 232667
rect 338326 232719 338378 232725
rect 338326 232661 338378 232667
rect 338242 231763 338270 232661
rect 338338 232577 338366 232661
rect 338326 232571 338378 232577
rect 338326 232513 338378 232519
rect 338422 232571 338474 232577
rect 338422 232513 338474 232519
rect 338434 232337 338462 232513
rect 338338 232309 338462 232337
rect 338338 232281 338366 232309
rect 338326 232275 338378 232281
rect 338326 232217 338378 232223
rect 338422 232275 338474 232281
rect 338422 232217 338474 232223
rect 338230 231757 338282 231763
rect 338230 231699 338282 231705
rect 338326 230943 338378 230949
rect 338326 230885 338378 230891
rect 338338 230579 338366 230885
rect 338434 230727 338462 232217
rect 338530 230949 338558 235769
rect 338518 230943 338570 230949
rect 338518 230885 338570 230891
rect 338422 230721 338474 230727
rect 338422 230663 338474 230669
rect 338326 230573 338378 230579
rect 338326 230515 338378 230521
rect 338518 229907 338570 229913
rect 338518 229849 338570 229855
rect 338422 229833 338474 229839
rect 338422 229775 338474 229781
rect 338326 229611 338378 229617
rect 338326 229553 338378 229559
rect 338338 228359 338366 229553
rect 338326 228353 338378 228359
rect 338326 228295 338378 228301
rect 338434 227619 338462 229775
rect 338530 228729 338558 229849
rect 338518 228723 338570 228729
rect 338518 228665 338570 228671
rect 338422 227613 338474 227619
rect 338422 227555 338474 227561
rect 338626 227291 338654 239672
rect 339010 238571 339038 239672
rect 338998 238565 339050 238571
rect 338998 238507 339050 238513
rect 339394 233211 339422 239672
rect 339490 235833 339518 239686
rect 339874 235981 339902 239686
rect 340272 239672 340478 239700
rect 340608 239672 340862 239700
rect 340992 239672 341246 239700
rect 341376 239672 341630 239700
rect 339862 235975 339914 235981
rect 339862 235917 339914 235923
rect 339478 235827 339530 235833
rect 339478 235769 339530 235775
rect 339862 233829 339914 233835
rect 339862 233771 339914 233777
rect 339380 233202 339436 233211
rect 339380 233137 339436 233146
rect 338710 232497 338762 232503
rect 338710 232439 338762 232445
rect 338722 232133 338750 232439
rect 338710 232127 338762 232133
rect 338710 232069 338762 232075
rect 339874 231023 339902 233771
rect 339862 231017 339914 231023
rect 339862 230959 339914 230965
rect 338708 228910 338764 228919
rect 338708 228845 338710 228854
rect 338762 228845 338764 228854
rect 338710 228813 338762 228819
rect 338612 227282 338668 227291
rect 338612 227217 338668 227226
rect 340246 225911 340298 225917
rect 340246 225853 340298 225859
rect 339478 225837 339530 225843
rect 339478 225779 339530 225785
rect 338134 224061 338186 224067
rect 338134 224003 338186 224009
rect 338710 223617 338762 223623
rect 338710 223559 338762 223565
rect 338722 221792 338750 223559
rect 338722 221764 338798 221792
rect 338770 221482 338798 221764
rect 339490 221482 339518 225779
rect 340258 221786 340286 225853
rect 340450 223993 340478 239672
rect 340834 228433 340862 239672
rect 341218 235537 341246 239672
rect 341206 235531 341258 235537
rect 341206 235473 341258 235479
rect 341014 230203 341066 230209
rect 341014 230145 341066 230151
rect 340822 228427 340874 228433
rect 340822 228369 340874 228375
rect 340438 223987 340490 223993
rect 340438 223929 340490 223935
rect 340248 221758 340286 221786
rect 341026 221792 341054 230145
rect 341602 226995 341630 239672
rect 341794 238497 341822 239686
rect 341782 238491 341834 238497
rect 341782 238433 341834 238439
rect 341974 235901 342026 235907
rect 341974 235843 342026 235849
rect 341588 226986 341644 226995
rect 341588 226921 341644 226930
rect 341986 225917 342014 235843
rect 342178 233063 342206 239686
rect 342562 234691 342590 239686
rect 342912 239672 343166 239700
rect 343296 239672 343550 239700
rect 343138 235907 343166 239672
rect 343126 235901 343178 235907
rect 343126 235843 343178 235849
rect 342548 234682 342604 234691
rect 342548 234617 342604 234626
rect 343522 233613 343550 239672
rect 342934 233607 342986 233613
rect 342934 233549 342986 233555
rect 343510 233607 343562 233613
rect 343510 233549 343562 233555
rect 342164 233054 342220 233063
rect 342164 232989 342220 232998
rect 341974 225911 342026 225917
rect 341974 225853 342026 225859
rect 342946 225103 342974 233549
rect 343414 233237 343466 233243
rect 343414 233179 343466 233185
rect 343222 231757 343274 231763
rect 343222 231699 343274 231705
rect 342550 225097 342602 225103
rect 342550 225039 342602 225045
rect 342934 225097 342986 225103
rect 342934 225039 342986 225045
rect 341782 223691 341834 223697
rect 341782 223633 341834 223639
rect 341026 221764 341102 221792
rect 340248 221482 340276 221758
rect 341074 221482 341102 221764
rect 341794 221482 341822 223633
rect 342562 221482 342590 225039
rect 343234 221792 343262 231699
rect 343426 231689 343454 233179
rect 343414 231683 343466 231689
rect 343414 231625 343466 231631
rect 343618 222217 343646 239686
rect 343702 230351 343754 230357
rect 343702 230293 343754 230299
rect 343714 229543 343742 230293
rect 344002 229913 344030 239686
rect 344386 236023 344414 239686
rect 344372 236014 344428 236023
rect 344372 235949 344428 235958
rect 344662 233903 344714 233909
rect 344662 233845 344714 233851
rect 343990 229907 344042 229913
rect 343990 229849 344042 229855
rect 343702 229537 343754 229543
rect 343702 229479 343754 229485
rect 344566 228427 344618 228433
rect 344566 228369 344618 228375
rect 344578 227693 344606 228369
rect 343990 227687 344042 227693
rect 343990 227629 344042 227635
rect 344566 227687 344618 227693
rect 344566 227629 344618 227635
rect 343606 222211 343658 222217
rect 343606 222153 343658 222159
rect 343234 221764 343310 221792
rect 343282 221482 343310 221764
rect 344002 221482 344030 227629
rect 344674 225029 344702 233845
rect 344770 233359 344798 239686
rect 345120 239672 345374 239700
rect 345346 238349 345374 239672
rect 345538 239672 345600 239700
rect 345334 238343 345386 238349
rect 345334 238285 345386 238291
rect 344756 233350 344812 233359
rect 344756 233285 344812 233294
rect 345538 232799 345566 239672
rect 345922 238423 345950 239686
rect 345910 238417 345962 238423
rect 345910 238359 345962 238365
rect 346306 236203 346334 239686
rect 346294 236197 346346 236203
rect 346294 236139 346346 236145
rect 345622 235457 345674 235463
rect 345622 235399 345674 235405
rect 345526 232793 345578 232799
rect 345526 232735 345578 232741
rect 345634 232429 345662 235399
rect 346294 233089 346346 233095
rect 346294 233031 346346 233037
rect 345622 232423 345674 232429
rect 345622 232365 345674 232371
rect 344758 229315 344810 229321
rect 344758 229257 344810 229263
rect 344770 228433 344798 229257
rect 344758 228427 344810 228433
rect 344758 228369 344810 228375
rect 345526 227243 345578 227249
rect 345526 227185 345578 227191
rect 344662 225023 344714 225029
rect 344662 224965 344714 224971
rect 344854 223543 344906 223549
rect 344854 223485 344906 223491
rect 344866 221482 344894 223485
rect 345538 221792 345566 227185
rect 345538 221764 345614 221792
rect 345586 221482 345614 221764
rect 346306 221482 346334 233031
rect 346690 223919 346718 239686
rect 347074 229839 347102 239686
rect 347424 239672 347678 239700
rect 347808 239672 347966 239700
rect 347650 235463 347678 239672
rect 347638 235457 347690 235463
rect 347638 235399 347690 235405
rect 347158 229981 347210 229987
rect 347158 229923 347210 229929
rect 347062 229833 347114 229839
rect 347062 229775 347114 229781
rect 347170 225492 347198 229923
rect 347074 225464 347198 225492
rect 346678 223913 346730 223919
rect 346678 223855 346730 223861
rect 347074 221482 347102 225464
rect 347938 223771 347966 239672
rect 348130 238275 348158 239686
rect 348528 239672 348830 239700
rect 348118 238269 348170 238275
rect 348118 238211 348170 238217
rect 348502 234125 348554 234131
rect 348502 234067 348554 234073
rect 348514 230727 348542 234067
rect 348694 233607 348746 233613
rect 348694 233549 348746 233555
rect 348502 230721 348554 230727
rect 348502 230663 348554 230669
rect 348598 227169 348650 227175
rect 348706 227143 348734 233549
rect 348802 230399 348830 239672
rect 348898 235685 348926 239686
rect 349344 239672 349598 239700
rect 349728 239672 349982 239700
rect 350112 239672 350366 239700
rect 348886 235679 348938 235685
rect 348886 235621 348938 235627
rect 349366 232349 349418 232355
rect 349366 232291 349418 232297
rect 348788 230390 348844 230399
rect 348788 230325 348844 230334
rect 348598 227111 348650 227117
rect 348692 227134 348748 227143
rect 347926 223765 347978 223771
rect 347926 223707 347978 223713
rect 347734 223469 347786 223475
rect 347734 223411 347786 223417
rect 347746 221792 347774 223411
rect 347746 221764 347822 221792
rect 347794 221482 347822 221764
rect 348610 221482 348638 227111
rect 348692 227069 348748 227078
rect 349378 221482 349406 232291
rect 349570 222069 349598 239672
rect 349954 223697 349982 239672
rect 350338 233243 350366 239672
rect 350434 236129 350462 239686
rect 350422 236123 350474 236129
rect 350422 236065 350474 236071
rect 350326 233237 350378 233243
rect 350326 233179 350378 233185
rect 350038 232645 350090 232651
rect 350038 232587 350090 232593
rect 349942 223691 349994 223697
rect 349942 223633 349994 223639
rect 349558 222063 349610 222069
rect 349558 222005 349610 222011
rect 350050 221792 350078 232587
rect 350818 223549 350846 239686
rect 351202 238201 351230 239686
rect 351552 239672 351806 239700
rect 351936 239672 352190 239700
rect 352320 239672 352574 239700
rect 352752 239672 353054 239700
rect 351190 238195 351242 238201
rect 351190 238137 351242 238143
rect 351778 229691 351806 239672
rect 352162 234131 352190 239672
rect 352150 234125 352202 234131
rect 352150 234067 352202 234073
rect 352342 232941 352394 232947
rect 352342 232883 352394 232889
rect 351766 229685 351818 229691
rect 351766 229627 351818 229633
rect 351574 227465 351626 227471
rect 351574 227407 351626 227413
rect 350806 223543 350858 223549
rect 350806 223485 350858 223491
rect 350806 223395 350858 223401
rect 350806 223337 350858 223343
rect 350050 221764 350126 221792
rect 350098 221482 350126 221764
rect 350818 221482 350846 223337
rect 351586 221808 351614 227407
rect 351566 221756 351614 221808
rect 352354 221829 352382 232883
rect 352546 223401 352574 239672
rect 352822 239601 352874 239607
rect 352822 239543 352874 239549
rect 352834 233465 352862 239543
rect 352822 233459 352874 233465
rect 352822 233401 352874 233407
rect 352726 230203 352778 230209
rect 352726 230145 352778 230151
rect 352738 230061 352766 230145
rect 352726 230055 352778 230061
rect 352726 229997 352778 230003
rect 353026 223475 353054 239672
rect 353122 233095 353150 239686
rect 353506 234987 353534 239686
rect 353856 239672 354110 239700
rect 353492 234978 353548 234987
rect 353492 234913 353548 234922
rect 353110 233089 353162 233095
rect 353110 233031 353162 233037
rect 353110 229611 353162 229617
rect 353110 229553 353162 229559
rect 353014 223469 353066 223475
rect 353014 223411 353066 223417
rect 352534 223395 352586 223401
rect 352534 223337 352586 223343
rect 352354 221794 352402 221829
rect 351566 221482 351594 221756
rect 352374 221496 352402 221794
rect 352374 221468 352416 221496
rect 353122 221482 353150 229553
rect 353878 223321 353930 223327
rect 353878 223263 353930 223269
rect 353890 221496 353918 223263
rect 354082 222851 354110 239672
rect 354226 239404 354254 239686
rect 354624 239672 354878 239700
rect 354178 239376 354254 239404
rect 354178 238127 354206 239376
rect 354166 238121 354218 238127
rect 354166 238063 354218 238069
rect 354358 235161 354410 235167
rect 354358 235103 354410 235109
rect 354262 234569 354314 234575
rect 354262 234511 354314 234517
rect 354274 232133 354302 234511
rect 354262 232127 354314 232133
rect 354262 232069 354314 232075
rect 354262 227761 354314 227767
rect 354262 227703 354314 227709
rect 354274 227471 354302 227703
rect 354262 227465 354314 227471
rect 354262 227407 354314 227413
rect 354370 227249 354398 235103
rect 354850 229617 354878 239672
rect 354946 233909 354974 239686
rect 355344 239672 355646 239700
rect 354934 233903 354986 233909
rect 354934 233845 354986 233851
rect 355318 233163 355370 233169
rect 355318 233105 355370 233111
rect 354838 229611 354890 229617
rect 354838 229553 354890 229559
rect 354358 227243 354410 227249
rect 354358 227185 354410 227191
rect 354550 225763 354602 225769
rect 354550 225705 354602 225711
rect 354068 222842 354124 222851
rect 354068 222777 354124 222786
rect 353856 221468 353918 221496
rect 354562 221496 354590 225705
rect 354562 221468 354624 221496
rect 355330 221482 355358 233105
rect 355618 223327 355646 239672
rect 355606 223321 355658 223327
rect 355606 223263 355658 223269
rect 355714 222999 355742 239686
rect 356064 239672 356318 239700
rect 356544 239672 356798 239700
rect 356086 232719 356138 232725
rect 356086 232661 356138 232667
rect 355700 222990 355756 222999
rect 355700 222925 355756 222934
rect 356098 221792 356126 232661
rect 356290 230251 356318 239672
rect 356770 233835 356798 239672
rect 356758 233829 356810 233835
rect 356758 233771 356810 233777
rect 356276 230242 356332 230251
rect 356276 230177 356332 230186
rect 356866 226847 356894 239686
rect 357250 229987 357278 239686
rect 357634 232355 357662 239686
rect 358018 235611 358046 239686
rect 358368 239672 358622 239700
rect 358752 239672 359006 239700
rect 358006 235605 358058 235611
rect 358006 235547 358058 235553
rect 358594 233687 358622 239672
rect 358486 233681 358538 233687
rect 358486 233623 358538 233629
rect 358582 233681 358634 233687
rect 358582 233623 358634 233629
rect 358294 232571 358346 232577
rect 358294 232513 358346 232519
rect 357622 232349 357674 232355
rect 357622 232291 357674 232297
rect 357238 229981 357290 229987
rect 357238 229923 357290 229929
rect 357622 227539 357674 227545
rect 357622 227481 357674 227487
rect 356852 226838 356908 226847
rect 356852 226773 356908 226782
rect 356854 223247 356906 223253
rect 356854 223189 356906 223195
rect 356098 221764 356174 221792
rect 356146 221482 356174 221764
rect 356866 221482 356894 223189
rect 357634 221482 357662 227481
rect 358306 221792 358334 232513
rect 358498 227534 358526 233623
rect 358498 227506 358622 227534
rect 358486 226725 358538 226731
rect 358486 226667 358538 226673
rect 358498 225769 358526 226667
rect 358486 225763 358538 225769
rect 358486 225705 358538 225711
rect 358594 224881 358622 227506
rect 358582 224875 358634 224881
rect 358582 224817 358634 224823
rect 358978 224627 359006 239672
rect 359074 230103 359102 239686
rect 359458 235431 359486 239686
rect 359444 235422 359500 235431
rect 359444 235357 359500 235366
rect 359060 230094 359116 230103
rect 359060 230029 359116 230038
rect 359158 229463 359210 229469
rect 359158 229405 359210 229411
rect 358964 224618 359020 224627
rect 358964 224553 359020 224562
rect 358774 223913 358826 223919
rect 358774 223855 358826 223861
rect 358786 222217 358814 223855
rect 358774 222211 358826 222217
rect 358774 222153 358826 222159
rect 359170 221798 359198 229405
rect 359842 224479 359870 239686
rect 360322 237905 360350 239686
rect 360672 239672 360926 239700
rect 361056 239672 361310 239700
rect 360310 237899 360362 237905
rect 360310 237841 360362 237847
rect 359926 235235 359978 235241
rect 359926 235177 359978 235183
rect 359938 227175 359966 235177
rect 360898 233021 360926 239672
rect 361282 233465 361310 239672
rect 361378 238053 361406 239686
rect 361366 238047 361418 238053
rect 361366 237989 361418 237995
rect 361654 236197 361706 236203
rect 361654 236139 361706 236145
rect 361270 233459 361322 233465
rect 361270 233401 361322 233407
rect 360790 233015 360842 233021
rect 360790 232957 360842 232963
rect 360886 233015 360938 233021
rect 360886 232957 360938 232963
rect 360802 232651 360830 232957
rect 360790 232645 360842 232651
rect 360790 232587 360842 232593
rect 361270 232497 361322 232503
rect 361270 232439 361322 232445
rect 359926 227169 359978 227175
rect 359926 227111 359978 227117
rect 360598 227095 360650 227101
rect 360598 227037 360650 227043
rect 359828 224470 359884 224479
rect 359828 224405 359884 224414
rect 359926 224283 359978 224289
rect 359926 224225 359978 224231
rect 358306 221764 358382 221792
rect 358354 221482 358382 221764
rect 359170 221762 359218 221798
rect 359190 221482 359218 221762
rect 359938 221482 359966 224225
rect 360610 221792 360638 227037
rect 361282 223420 361310 232439
rect 361366 229389 361418 229395
rect 361366 229331 361418 229337
rect 361378 224807 361406 229331
rect 361366 224801 361418 224807
rect 361366 224743 361418 224749
rect 361666 223771 361694 236139
rect 361762 229955 361790 239686
rect 362038 232275 362090 232281
rect 362038 232217 362090 232223
rect 361748 229946 361804 229955
rect 361748 229881 361804 229890
rect 362050 227534 362078 232217
rect 362146 229543 362174 239686
rect 362530 234543 362558 239686
rect 362880 239672 363134 239700
rect 363106 237979 363134 239672
rect 363250 239533 363278 239686
rect 363238 239527 363290 239533
rect 363238 239469 363290 239475
rect 363094 237973 363146 237979
rect 363094 237915 363146 237921
rect 363586 236351 363614 239686
rect 363574 236345 363626 236351
rect 363574 236287 363626 236293
rect 362710 235087 362762 235093
rect 362710 235029 362762 235035
rect 362516 234534 362572 234543
rect 362516 234469 362572 234478
rect 362134 229537 362186 229543
rect 362134 229479 362186 229485
rect 362050 227506 362174 227534
rect 361654 223765 361706 223771
rect 361654 223707 361706 223713
rect 361282 223392 361406 223420
rect 360610 221764 360686 221792
rect 360658 221482 360686 221764
rect 361378 221482 361406 223392
rect 362146 221482 362174 227506
rect 362722 224733 362750 235029
rect 364066 233539 364094 239686
rect 364450 237831 364478 239686
rect 364800 239672 364958 239700
rect 365184 239672 365438 239700
rect 365568 239672 365726 239700
rect 364438 237825 364490 237831
rect 364438 237767 364490 237773
rect 363958 233533 364010 233539
rect 363958 233475 364010 233481
rect 364054 233533 364106 233539
rect 364054 233475 364106 233481
rect 362804 233350 362860 233359
rect 362804 233285 362860 233294
rect 362710 224727 362762 224733
rect 362710 224669 362762 224675
rect 362818 224289 362846 233285
rect 363382 232867 363434 232873
rect 363382 232809 363434 232815
rect 363190 232275 363242 232281
rect 363190 232217 363242 232223
rect 363202 231911 363230 232217
rect 363190 231905 363242 231911
rect 363190 231847 363242 231853
rect 363394 231837 363422 232809
rect 363382 231831 363434 231837
rect 363382 231773 363434 231779
rect 363286 227835 363338 227841
rect 363286 227777 363338 227783
rect 363298 224955 363326 227777
rect 363670 227391 363722 227397
rect 363670 227333 363722 227339
rect 363286 224949 363338 224955
rect 363286 224891 363338 224897
rect 362806 224283 362858 224289
rect 362806 224225 362858 224231
rect 362902 222655 362954 222661
rect 362902 222597 362954 222603
rect 362914 221792 362942 222597
rect 362914 221764 362990 221792
rect 362962 221482 362990 221764
rect 363682 221482 363710 227333
rect 363970 222661 363998 233475
rect 364930 232577 364958 239672
rect 365014 239379 365066 239385
rect 365014 239321 365066 239327
rect 365026 235685 365054 239321
rect 365014 235679 365066 235685
rect 365014 235621 365066 235627
rect 364918 232571 364970 232577
rect 364918 232513 364970 232519
rect 364438 232201 364490 232207
rect 364438 232143 364490 232149
rect 363958 222655 364010 222661
rect 363958 222597 364010 222603
rect 364450 221482 364478 232143
rect 365110 231831 365162 231837
rect 365110 231773 365162 231779
rect 364534 223543 364586 223549
rect 364534 223485 364586 223491
rect 364630 223543 364682 223549
rect 364630 223485 364682 223491
rect 364546 223401 364574 223485
rect 364534 223395 364586 223401
rect 364534 223337 364586 223343
rect 364642 222069 364670 223485
rect 364630 222063 364682 222069
rect 364630 222005 364682 222011
rect 365122 221792 365150 231773
rect 365410 229469 365438 239672
rect 365698 233613 365726 239672
rect 365890 237757 365918 239686
rect 365878 237751 365930 237757
rect 365878 237693 365930 237699
rect 365686 233607 365738 233613
rect 365686 233549 365738 233555
rect 366274 232503 366302 239686
rect 366658 232725 366686 239686
rect 367008 239672 367262 239700
rect 367392 239672 367646 239700
rect 367872 239672 368126 239700
rect 367234 239163 367262 239672
rect 367222 239157 367274 239163
rect 367222 239099 367274 239105
rect 367618 237683 367646 239672
rect 367606 237677 367658 237683
rect 367606 237619 367658 237625
rect 366742 236715 366794 236721
rect 366742 236657 366794 236663
rect 366646 232719 366698 232725
rect 366646 232661 366698 232667
rect 366262 232497 366314 232503
rect 366262 232439 366314 232445
rect 365398 229463 365450 229469
rect 365398 229405 365450 229411
rect 366754 228600 366782 236657
rect 367222 233237 367274 233243
rect 367222 233179 367274 233185
rect 367234 232799 367262 233179
rect 367222 232793 367274 232799
rect 367222 232735 367274 232741
rect 368098 232281 368126 239672
rect 368086 232275 368138 232281
rect 368086 232217 368138 232223
rect 367126 232127 367178 232133
rect 367126 232069 367178 232075
rect 366934 231905 366986 231911
rect 366934 231847 366986 231853
rect 366946 230579 366974 231847
rect 366934 230573 366986 230579
rect 366934 230515 366986 230521
rect 367138 230505 367166 232069
rect 367414 231979 367466 231985
rect 367414 231921 367466 231927
rect 367126 230499 367178 230505
rect 367126 230441 367178 230447
rect 367030 229241 367082 229247
rect 367030 229183 367082 229189
rect 365890 228572 366782 228600
rect 365122 221764 365198 221792
rect 365170 221482 365198 221764
rect 365890 221482 365918 228572
rect 366742 227021 366794 227027
rect 366742 226963 366794 226969
rect 366754 221482 366782 226963
rect 367042 225621 367070 229183
rect 367030 225615 367082 225621
rect 367030 225557 367082 225563
rect 367426 221792 367454 231921
rect 368086 230573 368138 230579
rect 368086 230515 368138 230521
rect 368098 227534 368126 230515
rect 368194 229395 368222 239686
rect 368578 234099 368606 239686
rect 368976 239672 369182 239700
rect 368950 236641 369002 236647
rect 368950 236583 369002 236589
rect 368564 234090 368620 234099
rect 368564 234025 368620 234034
rect 368662 231091 368714 231097
rect 368662 231033 368714 231039
rect 368182 229389 368234 229395
rect 368182 229331 368234 229337
rect 368098 227506 368222 227534
rect 367426 221764 367502 221792
rect 367474 221482 367502 221764
rect 368194 221482 368222 227506
rect 368674 227027 368702 231033
rect 368662 227021 368714 227027
rect 368662 226963 368714 226969
rect 368962 221482 368990 236583
rect 369154 224331 369182 239672
rect 369298 239459 369326 239686
rect 369696 239672 369950 239700
rect 370080 239672 370334 239700
rect 369286 239453 369338 239459
rect 369286 239395 369338 239401
rect 369922 232207 369950 239672
rect 369910 232201 369962 232207
rect 369910 232143 369962 232149
rect 369622 227317 369674 227323
rect 369622 227259 369674 227265
rect 369140 224322 369196 224331
rect 369140 224257 369196 224266
rect 369634 221792 369662 227259
rect 370306 224183 370334 239672
rect 370402 237609 370430 239686
rect 370390 237603 370442 237609
rect 370390 237545 370442 237551
rect 370390 232053 370442 232059
rect 370390 231995 370442 232001
rect 370402 226528 370430 231995
rect 370786 231097 370814 239686
rect 370774 231091 370826 231097
rect 370774 231033 370826 231039
rect 371170 229807 371198 239686
rect 371616 239672 371870 239700
rect 372000 239672 372254 239700
rect 371842 232651 371870 239672
rect 372118 239305 372170 239311
rect 372118 239247 372170 239253
rect 372130 235611 372158 239247
rect 372226 236319 372254 239672
rect 372212 236310 372268 236319
rect 372212 236245 372268 236254
rect 372118 235605 372170 235611
rect 372118 235547 372170 235553
rect 371254 232645 371306 232651
rect 371254 232587 371306 232593
rect 371830 232645 371882 232651
rect 371830 232587 371882 232593
rect 371156 229798 371212 229807
rect 371156 229733 371212 229742
rect 370402 226500 370526 226528
rect 370292 224174 370348 224183
rect 370292 224109 370348 224118
rect 369634 221764 369710 221792
rect 369682 221482 369710 221764
rect 370498 221482 370526 226500
rect 371266 221482 371294 232587
rect 372322 232059 372350 239686
rect 372406 236789 372458 236795
rect 372406 236731 372458 236737
rect 372310 232053 372362 232059
rect 372310 231995 372362 232001
rect 371542 229315 371594 229321
rect 371542 229257 371594 229263
rect 371554 227323 371582 229257
rect 371542 227317 371594 227323
rect 371542 227259 371594 227265
rect 372418 221792 372446 236731
rect 372706 229247 372734 239686
rect 373090 235389 373118 239686
rect 373474 236911 373502 239686
rect 373824 239672 374078 239700
rect 374208 239672 374366 239700
rect 373460 236902 373516 236911
rect 373460 236837 373516 236846
rect 372886 235383 372938 235389
rect 372886 235325 372938 235331
rect 373078 235383 373130 235389
rect 373078 235325 373130 235331
rect 372898 235093 372926 235325
rect 372886 235087 372938 235093
rect 372886 235029 372938 235035
rect 374050 232619 374078 239672
rect 374338 232767 374366 239672
rect 374530 235685 374558 239686
rect 374518 235679 374570 235685
rect 374518 235621 374570 235627
rect 374614 233977 374666 233983
rect 374614 233919 374666 233925
rect 374324 232758 374380 232767
rect 374324 232693 374380 232702
rect 374036 232610 374092 232619
rect 374036 232545 374092 232554
rect 373462 231831 373514 231837
rect 373462 231773 373514 231779
rect 372694 229241 372746 229247
rect 372694 229183 372746 229189
rect 372694 226947 372746 226953
rect 372694 226889 372746 226895
rect 371986 221764 372446 221792
rect 371986 221482 372014 221764
rect 372706 221482 372734 226889
rect 373474 221825 373502 231773
rect 374518 231313 374570 231319
rect 374518 231255 374570 231261
rect 374230 230795 374282 230801
rect 374230 230737 374282 230743
rect 373454 221792 373502 221825
rect 374242 221792 374270 230737
rect 374422 229167 374474 229173
rect 374422 229109 374474 229115
rect 374434 225843 374462 229109
rect 374530 226953 374558 231255
rect 374518 226947 374570 226953
rect 374518 226889 374570 226895
rect 374422 225837 374474 225843
rect 374422 225779 374474 225785
rect 374626 222217 374654 233919
rect 374914 224035 374942 239686
rect 375394 232873 375422 239686
rect 375382 232867 375434 232873
rect 375382 232809 375434 232815
rect 375778 229173 375806 239686
rect 376128 239672 376382 239700
rect 376512 239672 376766 239700
rect 376150 239453 376202 239459
rect 376150 239395 376202 239401
rect 376162 230801 376190 239395
rect 376354 235875 376382 239672
rect 376738 236467 376766 239672
rect 376724 236458 376780 236467
rect 376724 236393 376780 236402
rect 376340 235866 376396 235875
rect 376340 235801 376396 235810
rect 376438 232127 376490 232133
rect 376438 232069 376490 232075
rect 376150 230795 376202 230801
rect 376150 230737 376202 230743
rect 375766 229167 375818 229173
rect 375766 229109 375818 229115
rect 375766 225763 375818 225769
rect 375766 225705 375818 225711
rect 374900 224026 374956 224035
rect 374900 223961 374956 223970
rect 374614 222211 374666 222217
rect 374614 222153 374666 222159
rect 374998 222137 375050 222143
rect 374998 222079 375050 222085
rect 373454 221482 373482 221792
rect 374242 221764 374318 221792
rect 374290 221482 374318 221764
rect 375010 221482 375038 222079
rect 375778 221482 375806 225705
rect 376450 221792 376478 232069
rect 376834 231837 376862 239686
rect 377218 231985 377246 239686
rect 377602 239089 377630 239686
rect 377590 239083 377642 239089
rect 377590 239025 377642 239031
rect 377986 237059 378014 239686
rect 378336 239672 378590 239700
rect 377972 237050 378028 237059
rect 377972 236985 378028 236994
rect 378454 232867 378506 232873
rect 378454 232809 378506 232815
rect 378466 232059 378494 232809
rect 378454 232053 378506 232059
rect 378454 231995 378506 232001
rect 377206 231979 377258 231985
rect 377206 231921 377258 231927
rect 378562 231911 378590 239672
rect 378706 239404 378734 239686
rect 378838 239527 378890 239533
rect 378838 239469 378890 239475
rect 378706 239376 378782 239404
rect 378646 235753 378698 235759
rect 378646 235695 378698 235701
rect 378658 235463 378686 235695
rect 378646 235457 378698 235463
rect 378646 235399 378698 235405
rect 377110 231905 377162 231911
rect 377110 231847 377162 231853
rect 378550 231905 378602 231911
rect 378550 231847 378602 231853
rect 376822 231831 376874 231837
rect 376822 231773 376874 231779
rect 377122 225788 377150 231847
rect 378754 229099 378782 239376
rect 378850 232799 378878 239469
rect 379138 234395 379166 239686
rect 379536 239672 379838 239700
rect 379124 234386 379180 234395
rect 379124 234321 379180 234330
rect 378934 233015 378986 233021
rect 378934 232957 378986 232963
rect 378838 232793 378890 232799
rect 378838 232735 378890 232741
rect 378946 232355 378974 232957
rect 379510 232423 379562 232429
rect 379510 232365 379562 232371
rect 378934 232349 378986 232355
rect 378934 232291 378986 232297
rect 378934 229981 378986 229987
rect 378934 229923 378986 229929
rect 378946 229543 378974 229923
rect 378934 229537 378986 229543
rect 378934 229479 378986 229485
rect 378742 229093 378794 229099
rect 378742 229035 378794 229041
rect 378742 226725 378794 226731
rect 378742 226667 378794 226673
rect 377122 225760 377246 225788
rect 376450 221764 376526 221792
rect 376498 221482 376526 221764
rect 377218 221482 377246 225760
rect 378070 222285 378122 222291
rect 378070 222227 378122 222233
rect 378082 221482 378110 222227
rect 378754 221792 378782 226667
rect 378754 221764 378830 221792
rect 378802 221482 378830 221764
rect 379522 221482 379550 232365
rect 379810 223887 379838 239672
rect 379906 232027 379934 239686
rect 380256 239672 380510 239700
rect 380640 239672 380894 239700
rect 381024 239672 381278 239700
rect 380182 232645 380234 232651
rect 380182 232587 380234 232593
rect 380278 232645 380330 232651
rect 380278 232587 380330 232593
rect 380194 232355 380222 232587
rect 380182 232349 380234 232355
rect 380182 232291 380234 232297
rect 380290 232207 380318 232587
rect 380482 232471 380510 239672
rect 380866 236615 380894 239672
rect 381046 236863 381098 236869
rect 381046 236805 381098 236811
rect 380852 236606 380908 236615
rect 380852 236541 380908 236550
rect 380468 232462 380524 232471
rect 380468 232397 380524 232406
rect 380278 232201 380330 232207
rect 380278 232143 380330 232149
rect 380662 232127 380714 232133
rect 380662 232069 380714 232075
rect 379892 232018 379948 232027
rect 379892 231953 379948 231962
rect 379990 231239 380042 231245
rect 379990 231181 380042 231187
rect 380002 226731 380030 231181
rect 380674 231097 380702 232069
rect 380662 231091 380714 231097
rect 380662 231033 380714 231039
rect 380278 230647 380330 230653
rect 380278 230589 380330 230595
rect 380086 227909 380138 227915
rect 380086 227851 380138 227857
rect 379990 226725 380042 226731
rect 379990 226667 380042 226673
rect 380098 225695 380126 227851
rect 380086 225689 380138 225695
rect 380086 225631 380138 225637
rect 379796 223878 379852 223887
rect 379796 223813 379852 223822
rect 380290 221760 380318 230589
rect 381058 221827 381086 236805
rect 381250 236763 381278 239672
rect 381236 236754 381292 236763
rect 381236 236689 381292 236698
rect 381346 232175 381374 239686
rect 381430 236345 381482 236351
rect 381430 236287 381482 236293
rect 381442 232873 381470 236287
rect 381430 232867 381482 232873
rect 381430 232809 381482 232815
rect 381332 232166 381388 232175
rect 381332 232101 381388 232110
rect 381730 229511 381758 239686
rect 382114 234247 382142 239686
rect 382560 239672 382814 239700
rect 382100 234238 382156 234247
rect 382100 234173 382156 234182
rect 381716 229502 381772 229511
rect 381716 229437 381772 229446
rect 381814 225985 381866 225991
rect 381814 225927 381866 225933
rect 381058 221794 381106 221827
rect 380270 221727 380318 221760
rect 380270 221482 380298 221727
rect 381078 221496 381106 221794
rect 381078 221468 381120 221496
rect 381826 221482 381854 225927
rect 382582 225615 382634 225621
rect 382582 225557 382634 225563
rect 382594 221496 382622 225557
rect 382786 223591 382814 239672
rect 382930 239404 382958 239686
rect 383062 239675 383114 239681
rect 383328 239672 383582 239700
rect 383062 239617 383114 239623
rect 382882 239376 382958 239404
rect 382882 223739 382910 239376
rect 383074 235611 383102 239617
rect 383158 239527 383210 239533
rect 383158 239469 383210 239475
rect 383062 235605 383114 235611
rect 383062 235547 383114 235553
rect 383062 235457 383114 235463
rect 383062 235399 383114 235405
rect 383074 231319 383102 235399
rect 383170 233391 383198 239469
rect 383158 233385 383210 233391
rect 383158 233327 383210 233333
rect 383554 232323 383582 239672
rect 383540 232314 383596 232323
rect 383540 232249 383596 232258
rect 383062 231313 383114 231319
rect 383062 231255 383114 231261
rect 383650 229363 383678 239686
rect 384034 236911 384062 239686
rect 383828 236902 383884 236911
rect 383828 236837 383884 236846
rect 384020 236902 384076 236911
rect 384020 236837 384076 236846
rect 383842 236203 383870 236837
rect 383830 236197 383882 236203
rect 383830 236139 383882 236145
rect 384418 235389 384446 239686
rect 384768 239672 385022 239700
rect 385152 239672 385406 239700
rect 385536 239672 385790 239700
rect 384406 235383 384458 235389
rect 384406 235325 384458 235331
rect 383636 229354 383692 229363
rect 383636 229289 383692 229298
rect 384994 229215 385022 239672
rect 385378 233835 385406 239672
rect 385762 235727 385790 239672
rect 385748 235718 385804 235727
rect 385748 235653 385804 235662
rect 385366 233829 385418 233835
rect 385366 233771 385418 233777
rect 384980 229206 385036 229215
rect 384980 229141 385036 229150
rect 383254 228057 383306 228063
rect 383254 227999 383306 228005
rect 382868 223730 382924 223739
rect 382868 223665 382924 223674
rect 382772 223582 382828 223591
rect 382772 223517 382828 223526
rect 382560 221468 382622 221496
rect 383266 221496 383294 227999
rect 385858 227767 385886 239686
rect 386352 239672 386654 239700
rect 386326 231535 386378 231541
rect 386326 231477 386378 231483
rect 385846 227761 385898 227767
rect 385846 227703 385898 227709
rect 385558 227317 385610 227323
rect 385558 227259 385610 227265
rect 384790 226651 384842 226657
rect 384790 226593 384842 226599
rect 384022 225911 384074 225917
rect 384022 225853 384074 225859
rect 383266 221468 383328 221496
rect 384034 221482 384062 225853
rect 384802 221792 384830 226593
rect 384802 221764 384878 221792
rect 384850 221482 384878 221764
rect 385570 221482 385598 227259
rect 386338 221482 386366 231477
rect 386626 225621 386654 239672
rect 386614 225615 386666 225621
rect 386614 225557 386666 225563
rect 386722 223443 386750 239686
rect 387072 239672 387326 239700
rect 387456 239672 387710 239700
rect 387190 233977 387242 233983
rect 387190 233919 387242 233925
rect 387202 227534 387230 233919
rect 387298 233632 387326 239672
rect 387298 233604 387422 233632
rect 387202 227506 387326 227534
rect 387298 224659 387326 227506
rect 387394 225917 387422 233604
rect 387682 225991 387710 239672
rect 387778 231245 387806 239686
rect 387766 231239 387818 231245
rect 387766 231181 387818 231187
rect 388162 226805 388190 239686
rect 388354 239672 388560 239700
rect 388354 227534 388382 239672
rect 388534 239231 388586 239237
rect 388534 239173 388586 239179
rect 388546 236319 388574 239173
rect 388628 237050 388684 237059
rect 388628 236985 388684 236994
rect 388642 236647 388670 236985
rect 388822 236715 388874 236721
rect 388822 236657 388874 236663
rect 388630 236641 388682 236647
rect 388834 236615 388862 236657
rect 388630 236583 388682 236589
rect 388820 236606 388876 236615
rect 388820 236541 388876 236550
rect 388532 236310 388588 236319
rect 388532 236245 388588 236254
rect 388724 236310 388780 236319
rect 388724 236245 388780 236254
rect 388738 236203 388766 236245
rect 388726 236197 388778 236203
rect 388726 236139 388778 236145
rect 388354 227506 388574 227534
rect 388150 226799 388202 226805
rect 388150 226741 388202 226747
rect 388546 226657 388574 227506
rect 388534 226651 388586 226657
rect 388534 226593 388586 226599
rect 387766 226059 387818 226065
rect 387766 226001 387818 226007
rect 387670 225985 387722 225991
rect 387670 225927 387722 225933
rect 387382 225911 387434 225917
rect 387382 225853 387434 225859
rect 386998 224653 387050 224659
rect 386998 224595 387050 224601
rect 387286 224653 387338 224659
rect 387286 224595 387338 224601
rect 386708 223434 386764 223443
rect 386708 223369 386764 223378
rect 387010 221792 387038 224595
rect 387010 221764 387086 221792
rect 387058 221482 387086 221764
rect 387778 221482 387806 226001
rect 388930 225917 388958 239686
rect 389280 239672 389534 239700
rect 389664 239672 389822 239700
rect 389014 236641 389066 236647
rect 389012 236606 389014 236615
rect 389066 236606 389068 236615
rect 389012 236541 389068 236550
rect 389302 228279 389354 228285
rect 389302 228221 389354 228227
rect 388918 225911 388970 225917
rect 388918 225853 388970 225859
rect 388630 225837 388682 225843
rect 388630 225779 388682 225785
rect 388642 221482 388670 225779
rect 389314 221792 389342 228221
rect 389506 225991 389534 239672
rect 389794 235167 389822 239672
rect 389782 235161 389834 235167
rect 389782 235103 389834 235109
rect 390082 227397 390110 239686
rect 390356 236754 390412 236763
rect 390356 236689 390358 236698
rect 390410 236689 390412 236698
rect 390358 236657 390410 236663
rect 390358 236567 390410 236573
rect 390358 236509 390410 236515
rect 390370 233761 390398 236509
rect 390358 233755 390410 233761
rect 390358 233697 390410 233703
rect 390466 227397 390494 239686
rect 390850 235241 390878 239686
rect 390838 235235 390890 235241
rect 390838 235177 390890 235183
rect 391234 234575 391262 239686
rect 391584 239672 391646 239700
rect 391968 239672 392222 239700
rect 391414 234939 391466 234945
rect 391414 234881 391466 234887
rect 391222 234569 391274 234575
rect 391222 234511 391274 234517
rect 391426 227915 391454 234881
rect 391510 234865 391562 234871
rect 391510 234807 391562 234813
rect 391414 227909 391466 227915
rect 391414 227851 391466 227857
rect 391522 227841 391550 234807
rect 391510 227835 391562 227841
rect 391510 227777 391562 227783
rect 390070 227391 390122 227397
rect 390070 227333 390122 227339
rect 390454 227391 390506 227397
rect 390454 227333 390506 227339
rect 390070 227243 390122 227249
rect 390070 227185 390122 227191
rect 389494 225985 389546 225991
rect 389494 225927 389546 225933
rect 389314 221764 389390 221792
rect 389362 221482 389390 221764
rect 390082 221482 390110 227185
rect 390742 226947 390794 226953
rect 390742 226889 390794 226895
rect 390754 225769 390782 226889
rect 390838 226873 390890 226879
rect 390838 226815 390890 226821
rect 390742 225763 390794 225769
rect 390742 225705 390794 225711
rect 390850 221482 390878 226815
rect 391618 226551 391646 239672
rect 392086 235087 392138 235093
rect 392086 235029 392138 235035
rect 392098 233909 392126 235029
rect 392086 233903 392138 233909
rect 392086 233845 392138 233851
rect 392194 227545 392222 239672
rect 392290 235093 392318 239686
rect 392278 235087 392330 235093
rect 392278 235029 392330 235035
rect 392674 234871 392702 239686
rect 392854 235309 392906 235315
rect 392854 235251 392906 235257
rect 392662 234865 392714 234871
rect 392662 234807 392714 234813
rect 392866 231245 392894 235251
rect 393058 234945 393086 239686
rect 393046 234939 393098 234945
rect 393046 234881 393098 234887
rect 392566 231239 392618 231245
rect 392566 231181 392618 231187
rect 392854 231239 392906 231245
rect 392854 231181 392906 231187
rect 392374 230869 392426 230875
rect 392374 230811 392426 230817
rect 392182 227539 392234 227545
rect 392182 227481 392234 227487
rect 391604 226542 391660 226551
rect 391604 226477 391660 226486
rect 391510 225763 391562 225769
rect 391510 225705 391562 225711
rect 391522 221792 391550 225705
rect 392386 221845 392414 230811
rect 392578 225769 392606 231181
rect 393142 227465 393194 227471
rect 393142 227407 393194 227413
rect 392566 225763 392618 225769
rect 392566 225705 392618 225711
rect 392386 221797 392424 221845
rect 391522 221764 391598 221792
rect 391570 221482 391598 221764
rect 392396 221482 392424 221797
rect 393154 221482 393182 227407
rect 393442 226699 393470 239686
rect 393888 239672 394142 239700
rect 394272 239672 394430 239700
rect 394608 239672 394910 239700
rect 394114 235283 394142 239672
rect 394100 235274 394156 235283
rect 394100 235209 394156 235218
rect 393910 235013 393962 235019
rect 393910 234955 393962 234961
rect 393922 230875 393950 234955
rect 394402 234797 394430 239672
rect 394486 239453 394538 239459
rect 394486 239395 394538 239401
rect 394498 236023 394526 239395
rect 394484 236014 394540 236023
rect 394484 235949 394540 235958
rect 394198 234791 394250 234797
rect 394198 234733 394250 234739
rect 394390 234791 394442 234797
rect 394390 234733 394442 234739
rect 393910 230869 393962 230875
rect 393910 230811 393962 230817
rect 394210 230579 394238 234733
rect 394198 230573 394250 230579
rect 394198 230515 394250 230521
rect 394582 228871 394634 228877
rect 394582 228813 394634 228819
rect 393428 226690 393484 226699
rect 393428 226625 393484 226634
rect 393814 226577 393866 226583
rect 393814 226519 393866 226525
rect 393826 221792 393854 226519
rect 394390 225689 394442 225695
rect 394390 225631 394442 225637
rect 394402 225344 394430 225631
rect 394594 225621 394622 228813
rect 394882 227101 394910 239672
rect 394978 227249 395006 239686
rect 395362 235579 395390 239686
rect 395712 239672 395966 239700
rect 396096 239672 396350 239700
rect 396480 239672 396734 239700
rect 395348 235570 395404 235579
rect 395348 235505 395404 235514
rect 395350 230943 395402 230949
rect 395350 230885 395402 230891
rect 395062 227539 395114 227545
rect 395062 227481 395114 227487
rect 394966 227243 395018 227249
rect 394966 227185 395018 227191
rect 394870 227095 394922 227101
rect 394870 227037 394922 227043
rect 395074 226805 395102 227481
rect 395062 226799 395114 226805
rect 395062 226741 395114 226747
rect 394870 225763 394922 225769
rect 394870 225705 394922 225711
rect 394486 225615 394538 225621
rect 394486 225557 394538 225563
rect 394582 225615 394634 225621
rect 394582 225557 394634 225563
rect 394498 225492 394526 225557
rect 394882 225492 394910 225705
rect 394498 225464 394910 225492
rect 394402 225316 394622 225344
rect 393826 221764 393902 221792
rect 393874 221482 393902 221764
rect 394594 221482 394622 225316
rect 395362 221482 395390 230885
rect 395938 229067 395966 239672
rect 396322 235315 396350 239672
rect 396310 235309 396362 235315
rect 396310 235251 396362 235257
rect 396706 235019 396734 239672
rect 396694 235013 396746 235019
rect 396694 234955 396746 234961
rect 395924 229058 395980 229067
rect 395924 228993 395980 229002
rect 396118 227169 396170 227175
rect 396118 227111 396170 227117
rect 396130 221792 396158 227111
rect 396802 226403 396830 239686
rect 396982 233903 397034 233909
rect 396982 233845 397034 233851
rect 396994 228063 397022 233845
rect 396982 228057 397034 228063
rect 396982 227999 397034 228005
rect 396886 226429 396938 226435
rect 396788 226394 396844 226403
rect 396886 226371 396938 226377
rect 396788 226329 396844 226338
rect 396130 221764 396206 221792
rect 396178 221482 396206 221764
rect 396898 221482 396926 226371
rect 397186 223295 397214 239686
rect 397366 236493 397418 236499
rect 397366 236435 397418 236441
rect 397378 235833 397406 236435
rect 397366 235827 397418 235833
rect 397366 235769 397418 235775
rect 397666 235537 397694 239686
rect 398016 239672 398270 239700
rect 398400 239672 398654 239700
rect 398784 239672 398942 239700
rect 398242 235833 398270 239672
rect 398230 235827 398282 235833
rect 398230 235769 398282 235775
rect 398626 235759 398654 239672
rect 398518 235753 398570 235759
rect 398518 235695 398570 235701
rect 398614 235753 398666 235759
rect 398614 235695 398666 235701
rect 397654 235531 397706 235537
rect 397654 235473 397706 235479
rect 397364 234386 397420 234395
rect 397364 234321 397420 234330
rect 397378 232915 397406 234321
rect 397364 232906 397420 232915
rect 397364 232841 397420 232850
rect 398326 228131 398378 228137
rect 398326 228073 398378 228079
rect 397654 226725 397706 226731
rect 397654 226667 397706 226673
rect 397558 226429 397610 226435
rect 397558 226371 397610 226377
rect 397570 226213 397598 226371
rect 397558 226207 397610 226213
rect 397558 226149 397610 226155
rect 397172 223286 397228 223295
rect 397172 223221 397228 223230
rect 397666 221482 397694 226667
rect 397750 226133 397802 226139
rect 397750 226075 397802 226081
rect 397762 225177 397790 226075
rect 397846 225615 397898 225621
rect 397846 225557 397898 225563
rect 397858 225177 397886 225557
rect 397750 225171 397802 225177
rect 397750 225113 397802 225119
rect 397846 225171 397898 225177
rect 397846 225113 397898 225119
rect 398338 221792 398366 228073
rect 398530 222291 398558 235695
rect 398806 235383 398858 235389
rect 398806 235325 398858 235331
rect 398710 231017 398762 231023
rect 398710 230959 398762 230965
rect 398722 230727 398750 230959
rect 398710 230721 398762 230727
rect 398710 230663 398762 230669
rect 398818 229659 398846 235325
rect 398914 231879 398942 239672
rect 399106 236023 399134 239686
rect 399092 236014 399148 236023
rect 399092 235949 399148 235958
rect 399490 233761 399518 239686
rect 399478 233755 399530 233761
rect 399478 233697 399530 233703
rect 398900 231870 398956 231879
rect 398900 231805 398956 231814
rect 398804 229650 398860 229659
rect 398804 229585 398860 229594
rect 399094 226281 399146 226287
rect 399094 226223 399146 226229
rect 398518 222285 398570 222291
rect 398518 222227 398570 222233
rect 398338 221764 398414 221792
rect 398386 221482 398414 221764
rect 399106 221482 399134 226223
rect 399874 224863 399902 239686
rect 399970 239672 400224 239700
rect 400608 239672 400862 239700
rect 400992 239672 401246 239700
rect 401424 239672 401726 239700
rect 399970 227249 399998 239672
rect 400246 236123 400298 236129
rect 400246 236065 400298 236071
rect 400258 235833 400286 236065
rect 400246 235827 400298 235833
rect 400246 235769 400298 235775
rect 400342 235827 400394 235833
rect 400342 235769 400394 235775
rect 400354 235704 400382 235769
rect 400258 235676 400382 235704
rect 400258 235537 400286 235676
rect 400246 235531 400298 235537
rect 400246 235473 400298 235479
rect 400628 234682 400684 234691
rect 400628 234617 400684 234626
rect 400438 234125 400490 234131
rect 400438 234067 400490 234073
rect 400342 233459 400394 233465
rect 400342 233401 400394 233407
rect 400246 231609 400298 231615
rect 400246 231551 400298 231557
rect 399958 227243 400010 227249
rect 399958 227185 400010 227191
rect 400258 226287 400286 231551
rect 400354 231541 400382 233401
rect 400342 231535 400394 231541
rect 400342 231477 400394 231483
rect 400450 228285 400478 234067
rect 400438 228279 400490 228285
rect 400438 228221 400490 228227
rect 400642 228137 400670 234617
rect 400630 228131 400682 228137
rect 400630 228073 400682 228079
rect 400834 226805 400862 239672
rect 401218 233909 401246 239672
rect 401206 233903 401258 233909
rect 401206 233845 401258 233851
rect 401398 227983 401450 227989
rect 401398 227925 401450 227931
rect 400822 226799 400874 226805
rect 400822 226741 400874 226747
rect 400246 226281 400298 226287
rect 400246 226223 400298 226229
rect 400630 225171 400682 225177
rect 400630 225113 400682 225119
rect 399874 224835 400094 224863
rect 400066 224733 400094 224835
rect 399958 224727 400010 224733
rect 399958 224669 400010 224675
rect 400054 224727 400106 224733
rect 400054 224669 400106 224675
rect 399970 221482 399998 224669
rect 400642 221792 400670 225113
rect 400642 221764 400718 221792
rect 400690 221482 400718 221764
rect 401410 221482 401438 227925
rect 401698 226879 401726 239672
rect 401794 235537 401822 239686
rect 401782 235531 401834 235537
rect 401782 235473 401834 235479
rect 402178 235135 402206 239686
rect 402528 239672 402782 239700
rect 402164 235126 402220 235135
rect 402164 235061 402220 235070
rect 402754 234395 402782 239672
rect 402850 239672 402912 239700
rect 403248 239672 403550 239700
rect 402740 234386 402796 234395
rect 402740 234321 402796 234330
rect 401974 227761 402026 227767
rect 401974 227703 402026 227709
rect 401986 226953 402014 227703
rect 401974 226947 402026 226953
rect 401974 226889 402026 226895
rect 401686 226873 401738 226879
rect 401686 226815 401738 226821
rect 402850 226731 402878 239672
rect 403318 236345 403370 236351
rect 403318 236287 403370 236293
rect 403222 236271 403274 236277
rect 403222 236213 403274 236219
rect 403234 235431 403262 236213
rect 403220 235422 403276 235431
rect 403220 235357 403276 235366
rect 403220 234978 403276 234987
rect 403220 234913 403276 234922
rect 403234 231319 403262 234913
rect 403330 233983 403358 236287
rect 403414 234717 403466 234723
rect 403414 234659 403466 234665
rect 403318 233977 403370 233983
rect 403318 233919 403370 233925
rect 403222 231313 403274 231319
rect 403222 231255 403274 231261
rect 403426 230949 403454 234659
rect 403522 234131 403550 239672
rect 403618 235389 403646 239686
rect 403606 235383 403658 235389
rect 403606 235325 403658 235331
rect 403510 234125 403562 234131
rect 403510 234067 403562 234073
rect 403414 230943 403466 230949
rect 403414 230885 403466 230891
rect 404002 228919 404030 239686
rect 404386 234839 404414 239686
rect 404736 239672 404990 239700
rect 405216 239672 405470 239700
rect 404372 234830 404428 234839
rect 404372 234765 404428 234774
rect 404962 234543 404990 239672
rect 405442 234987 405470 239672
rect 405428 234978 405484 234987
rect 405428 234913 405484 234922
rect 404756 234534 404812 234543
rect 404756 234469 404812 234478
rect 404948 234534 405004 234543
rect 404948 234469 405004 234478
rect 404470 230647 404522 230653
rect 404470 230589 404522 230595
rect 403988 228910 404044 228919
rect 403988 228845 404044 228854
rect 402838 226725 402890 226731
rect 402838 226667 402890 226673
rect 402838 226355 402890 226361
rect 402838 226297 402890 226303
rect 402166 224801 402218 224807
rect 402166 224743 402218 224749
rect 402178 221482 402206 224743
rect 402850 221792 402878 226297
rect 403702 226281 403754 226287
rect 403702 226223 403754 226229
rect 402850 221764 402926 221792
rect 402898 221482 402926 221764
rect 403714 221482 403742 226223
rect 404482 221482 404510 230589
rect 404770 222703 404798 234469
rect 405538 224881 405566 239686
rect 405922 234691 405950 239686
rect 405908 234682 405964 234691
rect 405908 234617 405964 234626
rect 406198 233903 406250 233909
rect 406198 233845 406250 233851
rect 406210 233761 406238 233845
rect 406198 233755 406250 233761
rect 406198 233697 406250 233703
rect 406102 233533 406154 233539
rect 406102 233475 406154 233481
rect 406006 229019 406058 229025
rect 406006 228961 406058 228967
rect 406018 225029 406046 228961
rect 406114 228877 406142 233475
rect 406306 233391 406334 239686
rect 406294 233385 406346 233391
rect 406294 233327 406346 233333
rect 406102 228871 406154 228877
rect 406102 228813 406154 228819
rect 406486 226947 406538 226953
rect 406486 226889 406538 226895
rect 406498 225769 406526 226889
rect 406690 226583 406718 239686
rect 407040 239672 407294 239700
rect 407424 239672 407678 239700
rect 407158 227761 407210 227767
rect 407158 227703 407210 227709
rect 407170 227323 407198 227703
rect 407158 227317 407210 227323
rect 407158 227259 407210 227265
rect 406678 226577 406730 226583
rect 406678 226519 406730 226525
rect 407266 226361 407294 239672
rect 407446 229759 407498 229765
rect 407446 229701 407498 229707
rect 407350 227243 407402 227249
rect 407350 227185 407402 227191
rect 407362 226953 407390 227185
rect 407350 226947 407402 226953
rect 407350 226889 407402 226895
rect 407254 226355 407306 226361
rect 407254 226297 407306 226303
rect 406486 225763 406538 225769
rect 406486 225705 406538 225711
rect 405910 225023 405962 225029
rect 405910 224965 405962 224971
rect 406006 225023 406058 225029
rect 406006 224965 406058 224971
rect 406774 225023 406826 225029
rect 406774 224965 406826 224971
rect 405142 224875 405194 224881
rect 405142 224817 405194 224823
rect 405526 224875 405578 224881
rect 405526 224817 405578 224823
rect 404756 222694 404812 222703
rect 404756 222629 404812 222638
rect 405154 221792 405182 224817
rect 405154 221764 405230 221792
rect 405202 221482 405230 221764
rect 405922 221482 405950 224965
rect 406786 221482 406814 224965
rect 407458 221792 407486 229701
rect 407650 227534 407678 239672
rect 407746 234723 407774 239686
rect 407734 234717 407786 234723
rect 407734 234659 407786 234665
rect 407650 227506 407774 227534
rect 407638 227391 407690 227397
rect 407638 227333 407690 227339
rect 407650 227249 407678 227333
rect 407638 227243 407690 227249
rect 407638 227185 407690 227191
rect 407746 226657 407774 227506
rect 407830 227391 407882 227397
rect 407830 227333 407882 227339
rect 407638 226651 407690 226657
rect 407638 226593 407690 226599
rect 407734 226651 407786 226657
rect 407734 226593 407786 226599
rect 407650 226565 407678 226593
rect 407842 226565 407870 227333
rect 407650 226537 407870 226565
rect 408130 226255 408158 239686
rect 408310 235013 408362 235019
rect 408310 234955 408362 234961
rect 408322 229025 408350 234955
rect 408310 229019 408362 229025
rect 408310 228961 408362 228967
rect 408214 227021 408266 227027
rect 408214 226963 408266 226969
rect 408116 226246 408172 226255
rect 408116 226181 408172 226190
rect 407458 221764 407534 221792
rect 407506 221482 407534 221764
rect 408226 221482 408254 226963
rect 408514 226107 408542 239686
rect 408960 239672 409214 239700
rect 409344 239672 409598 239700
rect 409728 239672 409982 239700
rect 409186 235463 409214 239672
rect 409174 235457 409226 235463
rect 409174 235399 409226 235405
rect 409570 233835 409598 239672
rect 409654 236937 409706 236943
rect 409654 236879 409706 236885
rect 409666 236174 409694 236879
rect 409666 236146 409886 236174
rect 409558 233829 409610 233835
rect 409558 233771 409610 233777
rect 408982 233607 409034 233613
rect 408982 233549 409034 233555
rect 408994 231615 409022 233549
rect 409174 233385 409226 233391
rect 409174 233327 409226 233333
rect 408982 231609 409034 231615
rect 408982 231551 409034 231557
rect 408982 226207 409034 226213
rect 408982 226149 409034 226155
rect 408500 226098 408556 226107
rect 408500 226033 408556 226042
rect 408994 221482 409022 226149
rect 409186 223147 409214 233327
rect 409654 230721 409706 230727
rect 409654 230663 409706 230669
rect 409558 226503 409610 226509
rect 409558 226445 409610 226451
rect 409570 225029 409598 226445
rect 409558 225023 409610 225029
rect 409558 224965 409610 224971
rect 409172 223138 409228 223147
rect 409172 223073 409228 223082
rect 409666 221792 409694 230663
rect 409858 228600 409886 236146
rect 409954 233391 409982 239672
rect 410050 233465 410078 239686
rect 410434 235019 410462 239686
rect 410710 236937 410762 236943
rect 410710 236879 410762 236885
rect 410722 235685 410750 236879
rect 410818 235685 410846 239686
rect 411168 239672 411422 239700
rect 411552 239672 411806 239700
rect 411936 239672 412190 239700
rect 410710 235679 410762 235685
rect 410710 235621 410762 235627
rect 410806 235679 410858 235685
rect 410806 235621 410858 235627
rect 410614 235531 410666 235537
rect 410614 235473 410666 235479
rect 410422 235013 410474 235019
rect 410422 234955 410474 234961
rect 410038 233459 410090 233465
rect 410038 233401 410090 233407
rect 409942 233385 409994 233391
rect 409942 233327 409994 233333
rect 409858 228572 410558 228600
rect 409750 226429 409802 226435
rect 409750 226371 409802 226377
rect 409762 224881 409790 226371
rect 409750 224875 409802 224881
rect 409750 224817 409802 224823
rect 409666 221764 409742 221792
rect 409714 221482 409742 221764
rect 410530 221482 410558 228572
rect 410626 227027 410654 235473
rect 411394 235431 411422 239672
rect 411574 237011 411626 237017
rect 411574 236953 411626 236959
rect 411586 235611 411614 236953
rect 411670 236197 411722 236203
rect 411670 236139 411722 236145
rect 411574 235605 411626 235611
rect 411574 235547 411626 235553
rect 411380 235422 411436 235431
rect 411380 235357 411436 235366
rect 411682 234099 411710 236139
rect 411778 235537 411806 239672
rect 411766 235531 411818 235537
rect 411766 235473 411818 235479
rect 411668 234090 411724 234099
rect 411668 234025 411724 234034
rect 411670 233459 411722 233465
rect 411670 233401 411722 233407
rect 411682 228327 411710 233401
rect 411766 233385 411818 233391
rect 411766 233327 411818 233333
rect 411668 228318 411724 228327
rect 411668 228253 411724 228262
rect 410614 227021 410666 227027
rect 410614 226963 410666 226969
rect 411778 226139 411806 233327
rect 411958 226503 412010 226509
rect 411958 226445 412010 226451
rect 411766 226133 411818 226139
rect 411766 226075 411818 226081
rect 411286 224949 411338 224955
rect 411286 224891 411338 224897
rect 411298 221496 411326 224891
rect 411264 221468 411326 221496
rect 411970 221496 411998 226445
rect 412162 226213 412190 239672
rect 420418 239237 420446 241129
rect 464758 239675 464810 239681
rect 464758 239617 464810 239623
rect 439126 239601 439178 239607
rect 439126 239543 439178 239549
rect 413398 239231 413450 239237
rect 413398 239173 413450 239179
rect 420406 239231 420458 239237
rect 420406 239173 420458 239179
rect 413410 238983 413438 239173
rect 413396 238974 413452 238983
rect 413396 238909 413452 238918
rect 413684 238678 413740 238687
rect 413684 238613 413740 238622
rect 413698 236943 413726 238613
rect 413972 238382 414028 238391
rect 413972 238317 414028 238326
rect 413986 237017 414014 238317
rect 438358 237307 438410 237313
rect 438358 237249 438410 237255
rect 434614 237233 434666 237239
rect 434614 237175 434666 237181
rect 428662 237159 428714 237165
rect 428662 237101 428714 237107
rect 423286 237085 423338 237091
rect 423286 237027 423338 237033
rect 413974 237011 414026 237017
rect 413974 236953 414026 236959
rect 413686 236937 413738 236943
rect 413686 236879 413738 236885
rect 416470 236863 416522 236869
rect 416470 236805 416522 236811
rect 413494 230499 413546 230505
rect 413494 230441 413546 230447
rect 412726 228205 412778 228211
rect 412726 228147 412778 228153
rect 412150 226207 412202 226213
rect 412150 226149 412202 226155
rect 411970 221468 412032 221496
rect 412738 221482 412766 228147
rect 413206 227761 413258 227767
rect 413206 227703 413258 227709
rect 413218 227323 413246 227703
rect 413206 227317 413258 227323
rect 413206 227259 413258 227265
rect 413206 226799 413258 226805
rect 413206 226741 413258 226747
rect 413218 226509 413246 226741
rect 413206 226503 413258 226509
rect 413206 226445 413258 226451
rect 413506 221778 413534 230441
rect 415700 228466 415756 228475
rect 415700 228401 415756 228410
rect 415412 228318 415468 228327
rect 415412 228253 415468 228262
rect 415030 226281 415082 226287
rect 415030 226223 415082 226229
rect 414262 222433 414314 222439
rect 414262 222375 414314 222381
rect 413486 221743 413534 221778
rect 414274 221787 414302 222375
rect 414274 221755 414322 221787
rect 413486 221496 413514 221743
rect 413472 221468 413514 221496
rect 414294 221482 414322 221755
rect 415042 221482 415070 226223
rect 415426 225177 415454 228253
rect 415414 225171 415466 225177
rect 415414 225113 415466 225119
rect 415714 221792 415742 228401
rect 415714 221764 415790 221792
rect 415762 221482 415790 221764
rect 416482 221482 416510 236805
rect 416948 234238 417004 234247
rect 416948 234173 417004 234182
rect 416962 229765 416990 234173
rect 420406 234051 420458 234057
rect 420406 233993 420458 233999
rect 418774 231017 418826 231023
rect 418774 230959 418826 230965
rect 416950 229759 417002 229765
rect 416950 229701 417002 229707
rect 418006 225097 418058 225103
rect 418006 225039 418058 225045
rect 417238 225023 417290 225029
rect 417238 224965 417290 224971
rect 417250 221482 417278 224965
rect 418018 221792 418046 225039
rect 418018 221764 418094 221792
rect 418066 221482 418094 221764
rect 418786 221482 418814 230959
rect 420418 230505 420446 233993
rect 420406 230499 420458 230505
rect 420406 230441 420458 230447
rect 421846 228501 421898 228507
rect 421846 228443 421898 228449
rect 418978 226981 419198 227009
rect 418978 226953 419006 226981
rect 418966 226947 419018 226953
rect 418966 226889 419018 226895
rect 419170 226805 419198 226981
rect 419254 226947 419306 226953
rect 419254 226889 419306 226895
rect 419158 226799 419210 226805
rect 419158 226741 419210 226747
rect 419062 226725 419114 226731
rect 419062 226667 419114 226673
rect 418870 226651 418922 226657
rect 418870 226593 418922 226599
rect 418882 226287 418910 226593
rect 418870 226281 418922 226287
rect 418870 226223 418922 226229
rect 419074 224733 419102 226667
rect 419266 226509 419294 226889
rect 419254 226503 419306 226509
rect 419254 226445 419306 226451
rect 420982 225245 421034 225251
rect 420982 225187 421034 225193
rect 419062 224727 419114 224733
rect 419062 224669 419114 224675
rect 419542 222507 419594 222513
rect 419542 222449 419594 222455
rect 419554 221482 419582 222449
rect 420214 222359 420266 222365
rect 420214 222301 420266 222307
rect 420226 221792 420254 222301
rect 420226 221764 420302 221792
rect 420274 221482 420302 221764
rect 420994 221482 421022 225187
rect 421858 221482 421886 228443
rect 422518 222581 422570 222587
rect 422518 222523 422570 222529
rect 422530 221792 422558 222523
rect 422530 221764 422606 221792
rect 422578 221482 422606 221764
rect 423298 221482 423326 237027
rect 424054 234199 424106 234205
rect 424054 234141 424106 234147
rect 424066 221482 424094 234141
rect 424726 231387 424778 231393
rect 424726 231329 424778 231335
rect 424738 221792 424766 231329
rect 425590 230647 425642 230653
rect 425590 230589 425642 230595
rect 424738 221764 424814 221792
rect 424786 221482 424814 221764
rect 425602 221788 425630 230589
rect 427798 228575 427850 228581
rect 427798 228517 427850 228523
rect 427030 225319 427082 225325
rect 427030 225261 427082 225267
rect 426358 222803 426410 222809
rect 426358 222745 426410 222751
rect 425602 221759 425640 221788
rect 425612 221482 425640 221759
rect 426370 221482 426398 222745
rect 427042 221792 427070 225261
rect 427042 221764 427118 221792
rect 427090 221482 427118 221764
rect 427810 221482 427838 228517
rect 428674 221482 428702 237101
rect 429142 233681 429194 233687
rect 429142 233623 429194 233629
rect 429154 228581 429182 233623
rect 433846 231461 433898 231467
rect 433846 231403 433898 231409
rect 430102 230499 430154 230505
rect 430102 230441 430154 230447
rect 429142 228575 429194 228581
rect 429142 228517 429194 228523
rect 429334 222877 429386 222883
rect 429334 222819 429386 222825
rect 429346 221792 429374 222819
rect 429346 221764 429422 221792
rect 429394 221482 429422 221764
rect 430114 221482 430142 230441
rect 430868 228614 430924 228623
rect 430868 228549 430924 228558
rect 430882 221482 430910 228549
rect 432406 228353 432458 228359
rect 432406 228295 432458 228301
rect 431542 222729 431594 222735
rect 431542 222671 431594 222677
rect 431554 221792 431582 222671
rect 431554 221764 431630 221792
rect 431602 221482 431630 221764
rect 432418 221482 432446 228295
rect 433174 225467 433226 225473
rect 433174 225409 433226 225415
rect 433186 221482 433214 225409
rect 433858 221792 433886 231403
rect 433858 221764 433934 221792
rect 433906 221482 433934 221764
rect 434626 221482 434654 237175
rect 436150 234347 436202 234353
rect 436150 234289 436202 234295
rect 434902 234273 434954 234279
rect 434902 234215 434954 234221
rect 434914 227989 434942 234215
rect 434902 227983 434954 227989
rect 434902 227925 434954 227931
rect 435382 227613 435434 227619
rect 435382 227555 435434 227561
rect 435394 221809 435422 227555
rect 435384 221776 435422 221809
rect 436162 221792 436190 234289
rect 436918 228649 436970 228655
rect 436918 228591 436970 228597
rect 435384 221482 435412 221776
rect 436162 221764 436238 221792
rect 436210 221482 436238 221764
rect 436930 221482 436958 228591
rect 437686 222951 437738 222957
rect 437686 222893 437738 222899
rect 437698 221482 437726 222893
rect 438370 221792 438398 237249
rect 438370 221764 438446 221792
rect 438418 221482 438446 221764
rect 439138 221482 439166 239543
rect 455062 239009 455114 239015
rect 455062 238951 455114 238957
rect 452758 237529 452810 237535
rect 452758 237471 452810 237477
rect 450454 237455 450506 237461
rect 450454 237397 450506 237403
rect 444502 237381 444554 237387
rect 444502 237323 444554 237329
rect 443446 234421 443498 234427
rect 443446 234363 443498 234369
rect 442868 231278 442924 231287
rect 442868 231213 442924 231222
rect 439988 228762 440044 228771
rect 439988 228697 440044 228706
rect 440002 221496 440030 228697
rect 442198 227983 442250 227989
rect 442198 227925 442250 227931
rect 440662 227835 440714 227841
rect 440662 227777 440714 227783
rect 439968 221468 440030 221496
rect 440674 221496 440702 227777
rect 441430 223025 441482 223031
rect 441430 222967 441482 222973
rect 440674 221468 440736 221496
rect 441442 221482 441470 222967
rect 442210 221496 442238 227925
rect 442176 221468 442238 221496
rect 442882 221496 442910 231213
rect 443458 227619 443486 234363
rect 443734 230869 443786 230875
rect 443734 230811 443786 230817
rect 443446 227613 443498 227619
rect 443446 227555 443498 227561
rect 442882 221468 442944 221496
rect 443746 221482 443774 230811
rect 444514 221792 444542 237323
rect 449302 234643 449354 234649
rect 449302 234585 449354 234591
rect 446326 234495 446378 234501
rect 446326 234437 446378 234443
rect 445942 228723 445994 228729
rect 445942 228665 445994 228671
rect 445174 225541 445226 225547
rect 445174 225483 445226 225489
rect 444466 221764 444542 221792
rect 444466 221482 444494 221764
rect 445186 221482 445214 225483
rect 445954 221482 445982 228665
rect 446338 227767 446366 234437
rect 448916 231426 448972 231435
rect 448916 231361 448972 231370
rect 446614 230943 446666 230949
rect 446614 230885 446666 230891
rect 446326 227761 446378 227767
rect 446326 227703 446378 227709
rect 446626 221792 446654 230885
rect 448246 227613 448298 227619
rect 448246 227555 448298 227561
rect 447478 223099 447530 223105
rect 447478 223041 447530 223047
rect 446626 221764 446702 221792
rect 446674 221482 446702 221764
rect 447490 221767 447518 223041
rect 447490 221725 447538 221767
rect 447510 221482 447538 221725
rect 448258 221482 448286 227555
rect 448930 221792 448958 231361
rect 449314 228359 449342 234585
rect 449302 228353 449354 228359
rect 449302 228295 449354 228301
rect 449686 223173 449738 223179
rect 449686 223115 449738 223121
rect 448930 221764 449006 221792
rect 448978 221482 449006 221764
rect 449698 221482 449726 223115
rect 450466 221482 450494 237397
rect 451990 228797 452042 228803
rect 451990 228739 452042 228745
rect 451222 225393 451274 225399
rect 451222 225335 451274 225341
rect 451234 221792 451262 225335
rect 451234 221764 451310 221792
rect 451282 221482 451310 221764
rect 452002 221482 452030 228739
rect 452770 221482 452798 237471
rect 455074 228507 455102 238951
rect 461878 238935 461930 238941
rect 461878 238877 461930 238883
rect 455254 233755 455306 233761
rect 455254 233697 455306 233703
rect 455266 228951 455294 233697
rect 460726 233311 460778 233317
rect 460726 233253 460778 233259
rect 458036 231574 458092 231583
rect 458036 231509 458092 231518
rect 455158 228945 455210 228951
rect 455158 228887 455210 228893
rect 455254 228945 455306 228951
rect 455254 228887 455306 228893
rect 455062 228501 455114 228507
rect 455062 228443 455114 228449
rect 454294 227761 454346 227767
rect 454294 227703 454346 227709
rect 453430 224579 453482 224585
rect 453430 224521 453482 224527
rect 453442 221792 453470 224521
rect 453442 221764 453518 221792
rect 453490 221482 453518 221764
rect 454306 221743 454334 227703
rect 455170 224900 455198 228887
rect 456502 228501 456554 228507
rect 456502 228443 456554 228449
rect 455734 227909 455786 227915
rect 455734 227851 455786 227857
rect 455074 224872 455198 224900
rect 454306 221707 454344 221743
rect 454316 221482 454344 221707
rect 455074 221482 455102 224872
rect 455746 221792 455774 227851
rect 455746 221764 455822 221792
rect 455794 221482 455822 221764
rect 456514 221482 456542 228443
rect 457268 225506 457324 225515
rect 457268 225441 457324 225450
rect 457282 221773 457310 225441
rect 457272 221731 457310 221773
rect 458050 221792 458078 231509
rect 460246 228353 460298 228359
rect 460246 228295 460298 228301
rect 459574 224505 459626 224511
rect 459574 224447 459626 224453
rect 458806 222211 458858 222217
rect 458806 222153 458858 222159
rect 458050 221764 458126 221792
rect 457272 221482 457300 221731
rect 458098 221482 458126 221764
rect 458818 221482 458846 222153
rect 459586 221482 459614 224447
rect 460258 221792 460286 228295
rect 460738 227619 460766 233253
rect 461014 230425 461066 230431
rect 461014 230367 461066 230373
rect 460726 227613 460778 227619
rect 460726 227555 460778 227561
rect 460258 221764 460334 221792
rect 460306 221482 460334 221764
rect 461026 221482 461054 230367
rect 461890 221482 461918 238877
rect 462550 238861 462602 238867
rect 462550 238803 462602 238809
rect 462562 221792 462590 238803
rect 464084 231722 464140 231731
rect 464084 231657 464140 231666
rect 463316 225654 463372 225663
rect 463316 225589 463372 225598
rect 462562 221764 462638 221792
rect 462610 221482 462638 221764
rect 463330 221482 463358 225589
rect 464098 221482 464126 231657
rect 464770 221792 464798 239617
rect 473878 239527 473930 239533
rect 473878 239469 473930 239475
rect 468598 238787 468650 238793
rect 468598 238729 468650 238735
rect 466486 236049 466538 236055
rect 466486 235991 466538 235997
rect 466498 228507 466526 235991
rect 467830 231091 467882 231097
rect 467830 231033 467882 231039
rect 467062 230351 467114 230357
rect 467062 230293 467114 230299
rect 466486 228501 466538 228507
rect 466486 228443 466538 228449
rect 466390 227613 466442 227619
rect 466390 227555 466442 227561
rect 465622 224357 465674 224363
rect 465622 224299 465674 224305
rect 464770 221764 464846 221792
rect 464818 221482 464846 221764
rect 465634 221482 465662 224299
rect 466402 221482 466430 227555
rect 467074 221792 467102 230293
rect 467074 221764 467150 221792
rect 467122 221482 467150 221764
rect 467842 221482 467870 231033
rect 468610 221728 468638 238729
rect 471284 236162 471340 236171
rect 471284 236097 471340 236106
rect 471298 230431 471326 236097
rect 473110 231683 473162 231689
rect 473110 231625 473162 231631
rect 471286 230425 471338 230431
rect 471286 230367 471338 230373
rect 470134 230277 470186 230283
rect 470134 230219 470186 230225
rect 469364 225802 469420 225811
rect 469364 225737 469420 225746
rect 469378 221778 469406 225737
rect 469378 221736 469426 221778
rect 468585 221682 468638 221728
rect 468585 221546 468618 221682
rect 468590 221482 468618 221546
rect 469398 221496 469426 221736
rect 469398 221468 469440 221496
rect 470146 221482 470174 230219
rect 470902 228057 470954 228063
rect 470902 227999 470954 228005
rect 470914 221496 470942 227999
rect 472340 225950 472396 225959
rect 472340 225885 472396 225894
rect 471574 224431 471626 224437
rect 471574 224373 471626 224379
rect 470880 221468 470942 221496
rect 471586 221496 471614 224373
rect 471586 221468 471648 221496
rect 472354 221482 472382 225885
rect 473122 221792 473150 231625
rect 473122 221764 473198 221792
rect 473170 221482 473198 221764
rect 473890 221482 473918 239469
rect 496534 239453 496586 239459
rect 496534 239395 496586 239401
rect 474646 238713 474698 238719
rect 474646 238655 474698 238661
rect 474658 221482 474686 238655
rect 480694 238639 480746 238645
rect 480694 238581 480746 238587
rect 476950 236567 477002 236573
rect 476950 236509 477002 236515
rect 475222 235975 475274 235981
rect 475222 235917 475274 235923
rect 475234 230357 475262 235917
rect 475222 230351 475274 230357
rect 475222 230293 475274 230299
rect 475318 228501 475370 228507
rect 475318 228443 475370 228449
rect 475330 221792 475358 228443
rect 476182 228427 476234 228433
rect 476182 228369 476234 228375
rect 475330 221764 475406 221792
rect 475378 221482 475406 221764
rect 476194 221780 476222 228369
rect 476194 221744 476242 221780
rect 476214 221482 476242 221744
rect 476962 221482 476990 236509
rect 479158 231757 479210 231763
rect 479158 231699 479210 231705
rect 478388 227430 478444 227439
rect 478388 227365 478444 227374
rect 477622 224135 477674 224141
rect 477622 224077 477674 224083
rect 477634 221792 477662 224077
rect 477634 221764 477710 221792
rect 477682 221482 477710 221764
rect 478402 221482 478430 227365
rect 479170 221482 479198 231699
rect 479926 222655 479978 222661
rect 479926 222597 479978 222603
rect 479938 221792 479966 222597
rect 479938 221764 480014 221792
rect 479986 221482 480014 221764
rect 480706 221482 480734 238581
rect 486742 238565 486794 238571
rect 486742 238507 486794 238513
rect 483862 236493 483914 236499
rect 483862 236435 483914 236441
rect 483766 235901 483818 235907
rect 483766 235843 483818 235849
rect 481462 230425 481514 230431
rect 481462 230367 481514 230373
rect 481474 221482 481502 230367
rect 482134 230055 482186 230061
rect 482134 229997 482186 230003
rect 482146 221792 482174 229997
rect 483778 228433 483806 235843
rect 483874 228507 483902 236435
rect 485590 236123 485642 236129
rect 485590 236065 485642 236071
rect 485206 230129 485258 230135
rect 485206 230071 485258 230077
rect 483862 228501 483914 228507
rect 483862 228443 483914 228449
rect 483766 228427 483818 228433
rect 483766 228369 483818 228375
rect 484436 227282 484492 227291
rect 484436 227217 484492 227226
rect 483766 224209 483818 224215
rect 483766 224151 483818 224157
rect 482902 224061 482954 224067
rect 482902 224003 482954 224009
rect 482146 221764 482222 221792
rect 482194 221482 482222 221764
rect 482914 221482 482942 224003
rect 483778 221482 483806 224151
rect 484450 221792 484478 227217
rect 484450 221764 484526 221792
rect 484498 221482 484526 221764
rect 485218 221482 485246 230071
rect 485602 230061 485630 236065
rect 485590 230055 485642 230061
rect 485590 229997 485642 230003
rect 485974 228501 486026 228507
rect 485974 228443 486026 228449
rect 485986 221482 486014 228443
rect 486754 221792 486782 238507
rect 492790 238491 492842 238497
rect 492790 238433 492842 238439
rect 492502 233977 492554 233983
rect 492502 233919 492554 233925
rect 489622 233903 489674 233909
rect 489622 233845 489674 233851
rect 488276 233202 488332 233211
rect 488276 233137 488332 233146
rect 487510 230351 487562 230357
rect 487510 230293 487562 230299
rect 486706 221764 486782 221792
rect 486706 221482 486734 221764
rect 487522 221482 487550 230293
rect 488290 221482 488318 233137
rect 488950 231239 489002 231245
rect 488950 231181 489002 231187
rect 488962 221792 488990 231181
rect 489634 229987 489662 233845
rect 492514 230209 492542 233919
rect 492502 230203 492554 230209
rect 492502 230145 492554 230151
rect 489622 229981 489674 229987
rect 489622 229923 489674 229929
rect 492022 228131 492074 228137
rect 492022 228073 492074 228079
rect 491254 227687 491306 227693
rect 491254 227629 491306 227635
rect 490484 226986 490540 226995
rect 490484 226921 490540 226930
rect 489718 223987 489770 223993
rect 489718 223929 489770 223935
rect 488962 221764 489038 221792
rect 489010 221482 489038 221764
rect 489730 221482 489758 223929
rect 490498 221740 490526 226921
rect 491266 221792 491294 227629
rect 491266 221764 491342 221792
rect 490488 221704 490526 221740
rect 490488 221482 490516 221704
rect 491314 221482 491342 221764
rect 492034 221482 492062 228073
rect 492802 221482 492830 238433
rect 494228 233054 494284 233063
rect 494228 232989 494284 232998
rect 493462 228427 493514 228433
rect 493462 228369 493514 228375
rect 493474 221792 493502 228369
rect 493474 221764 493550 221792
rect 493522 221482 493550 221764
rect 494242 221482 494270 232989
rect 495094 229907 495146 229913
rect 495094 229849 495146 229855
rect 495106 221482 495134 229849
rect 495764 227134 495820 227143
rect 495764 227069 495820 227078
rect 495778 221792 495806 227069
rect 495778 221764 495854 221792
rect 495826 221482 495854 221764
rect 496546 221482 496574 239395
rect 505654 239379 505706 239385
rect 505654 239321 505706 239327
rect 498262 238417 498314 238423
rect 498262 238359 498314 238365
rect 497974 233237 498026 233243
rect 497974 233179 498026 233185
rect 497302 223913 497354 223919
rect 497302 223855 497354 223861
rect 497314 221482 497342 223855
rect 497986 221792 498014 233179
rect 497986 221764 498062 221792
rect 498274 221773 498302 238359
rect 500278 238343 500330 238349
rect 500278 238285 500330 238291
rect 498838 224283 498890 224289
rect 498838 224225 498890 224231
rect 498034 221482 498062 221764
rect 498262 221767 498314 221773
rect 498262 221709 498314 221715
rect 498850 221482 498878 224225
rect 499558 221767 499610 221773
rect 499558 221709 499610 221715
rect 499570 221482 499598 221709
rect 500290 221496 500318 238285
rect 504118 238269 504170 238275
rect 504118 238211 504170 238217
rect 501044 234386 501100 234395
rect 501044 234321 501100 234330
rect 501058 230135 501086 234321
rect 504020 230390 504076 230399
rect 504020 230325 504076 230334
rect 501046 230129 501098 230135
rect 501046 230071 501098 230077
rect 501046 229833 501098 229839
rect 501046 229775 501098 229781
rect 500290 221468 500352 221496
rect 501058 221482 501086 229775
rect 503350 223839 503402 223845
rect 503350 223781 503402 223787
rect 501814 223765 501866 223771
rect 501814 223707 501866 223713
rect 501826 221792 501854 223707
rect 502582 222285 502634 222291
rect 502582 222227 502634 222233
rect 501826 221764 501902 221792
rect 501874 221482 501902 221764
rect 502594 221482 502622 222227
rect 503362 221482 503390 223781
rect 504034 221792 504062 230325
rect 504130 227534 504158 238211
rect 504130 227506 504254 227534
rect 504034 221764 504110 221792
rect 504226 221773 504254 227506
rect 504790 223617 504842 223623
rect 504790 223559 504842 223565
rect 504082 221482 504110 221764
rect 504214 221767 504266 221773
rect 504214 221709 504266 221715
rect 504802 221482 504830 223559
rect 505666 221482 505694 239321
rect 523798 239305 523850 239311
rect 523798 239247 523850 239253
rect 512374 238195 512426 238201
rect 512374 238137 512426 238143
rect 508630 236419 508682 236425
rect 508630 236361 508682 236367
rect 507094 233163 507146 233169
rect 507094 233105 507146 233111
rect 506134 229833 506186 229839
rect 506134 229775 506186 229781
rect 506146 229617 506174 229775
rect 506134 229611 506186 229617
rect 506134 229553 506186 229559
rect 506374 221767 506426 221773
rect 506374 221709 506426 221715
rect 506386 221482 506414 221709
rect 507106 221482 507134 233105
rect 507862 223543 507914 223549
rect 507862 223485 507914 223491
rect 507874 221482 507902 223485
rect 508642 221792 508670 236361
rect 509782 234125 509834 234131
rect 509782 234067 509834 234073
rect 509794 229691 509822 234067
rect 509782 229685 509834 229691
rect 509782 229627 509834 229633
rect 510166 229611 510218 229617
rect 510166 229553 510218 229559
rect 509398 223691 509450 223697
rect 509398 223633 509450 223639
rect 508594 221764 508670 221792
rect 509410 221814 509438 223633
rect 509410 221771 509448 221814
rect 508594 221482 508622 221764
rect 509420 221482 509448 221771
rect 510178 221482 510206 229553
rect 511606 228279 511658 228285
rect 511606 228221 511658 228227
rect 510838 223395 510890 223401
rect 510838 223337 510890 223343
rect 510850 221792 510878 223337
rect 510850 221764 510926 221792
rect 510898 221482 510926 221764
rect 511618 221482 511646 228221
rect 512386 221482 512414 238137
rect 518518 238121 518570 238127
rect 518518 238063 518570 238069
rect 518530 236174 518558 238063
rect 520726 236345 520778 236351
rect 520726 236287 520778 236293
rect 518434 236146 518558 236174
rect 512662 234569 512714 234575
rect 512662 234511 512714 234517
rect 516212 234534 516268 234543
rect 512674 233095 512702 234511
rect 516212 234469 516268 234478
rect 513142 233163 513194 233169
rect 513142 233105 513194 233111
rect 512662 233089 512714 233095
rect 512662 233031 512714 233037
rect 513154 221792 513182 233105
rect 514678 231313 514730 231319
rect 514678 231255 514730 231261
rect 513910 223321 513962 223327
rect 513910 223263 513962 223269
rect 513154 221764 513230 221792
rect 513202 221482 513230 221764
rect 513922 221482 513950 223263
rect 514690 221482 514718 231255
rect 516118 229833 516170 229839
rect 516118 229775 516170 229781
rect 515350 223469 515402 223475
rect 515350 223411 515402 223417
rect 515362 221792 515390 223411
rect 515362 221764 515438 221792
rect 515410 221482 515438 221764
rect 516130 221482 516158 229775
rect 516226 229617 516254 234469
rect 516214 229611 516266 229617
rect 516214 229553 516266 229559
rect 517654 224653 517706 224659
rect 517654 224595 517706 224601
rect 516980 222842 517036 222851
rect 516980 222777 517036 222786
rect 516994 221482 517022 222777
rect 517666 221792 517694 224595
rect 517666 221764 517742 221792
rect 517714 221482 517742 221764
rect 518434 221482 518462 236146
rect 519188 230242 519244 230251
rect 519188 230177 519244 230186
rect 519202 221482 519230 230177
rect 519862 223247 519914 223253
rect 519862 223189 519914 223195
rect 519874 221681 519902 223189
rect 519874 221653 519950 221681
rect 519922 221482 519950 221653
rect 520738 221482 520766 236287
rect 522166 233015 522218 233021
rect 522166 232957 522218 232963
rect 521492 222990 521548 222999
rect 521492 222925 521548 222934
rect 521506 221482 521534 222925
rect 522178 221681 522206 232957
rect 522932 226838 522988 226847
rect 522932 226773 522988 226782
rect 522178 221653 522254 221681
rect 522226 221482 522254 221653
rect 522946 221482 522974 226773
rect 523810 221482 523838 239247
rect 596182 239231 596234 239237
rect 596182 239173 596234 239179
rect 542614 239157 542666 239163
rect 542614 239099 542666 239105
rect 532054 238047 532106 238053
rect 532054 237989 532106 237995
rect 530518 237899 530570 237905
rect 530518 237841 530570 237847
rect 526678 236271 526730 236277
rect 526678 236213 526730 236219
rect 525236 230094 525292 230103
rect 525236 230029 525292 230038
rect 524470 229537 524522 229543
rect 524470 229479 524522 229485
rect 524482 221681 524510 229479
rect 524482 221653 524558 221681
rect 524530 221482 524558 221653
rect 525250 221482 525278 230029
rect 526006 228575 526058 228581
rect 526006 228517 526058 228523
rect 526018 221482 526046 228517
rect 526690 221792 526718 236213
rect 528310 232941 528362 232947
rect 528310 232883 528362 232889
rect 527540 224618 527596 224627
rect 527540 224553 527596 224562
rect 526690 221764 526766 221792
rect 526738 221482 526766 221764
rect 527554 221482 527582 224553
rect 528322 221496 528350 232883
rect 529750 231535 529802 231541
rect 529750 231477 529802 231483
rect 528980 224470 529036 224479
rect 528980 224405 529036 224414
rect 528288 221468 528350 221496
rect 528994 221496 529022 224405
rect 528994 221468 529056 221496
rect 529762 221482 529790 231477
rect 530530 221825 530558 237841
rect 531286 229463 531338 229469
rect 531286 229405 531338 229411
rect 530510 221782 530558 221825
rect 531298 221799 531326 229405
rect 530510 221496 530538 221782
rect 531298 221761 531346 221799
rect 530496 221468 530538 221496
rect 531318 221482 531346 221761
rect 532066 221482 532094 237989
rect 535126 237973 535178 237979
rect 535126 237915 535178 237921
rect 534262 232867 534314 232873
rect 534262 232809 534314 232815
rect 533492 229946 533548 229955
rect 533492 229881 533548 229890
rect 532820 222694 532876 222703
rect 532820 222629 532876 222638
rect 532834 221755 532862 222629
rect 532738 221727 532862 221755
rect 532738 221681 532766 221727
rect 532738 221653 532814 221681
rect 532786 221482 532814 221653
rect 533506 221482 533534 229881
rect 534274 221482 534302 232809
rect 535138 221792 535166 237915
rect 538006 237825 538058 237831
rect 538006 237767 538058 237773
rect 536566 232793 536618 232799
rect 536566 232735 536618 232741
rect 535798 228871 535850 228877
rect 535798 228813 535850 228819
rect 535090 221764 535166 221792
rect 535090 221482 535118 221764
rect 535810 221482 535838 228813
rect 536578 221482 536606 232735
rect 537238 229389 537290 229395
rect 537238 229331 537290 229337
rect 537250 221681 537278 229331
rect 537250 221653 537326 221681
rect 537298 221482 537326 221653
rect 538018 221482 538046 237767
rect 538582 237751 538634 237757
rect 538582 237693 538634 237699
rect 538594 228581 538622 237693
rect 541558 237677 541610 237683
rect 541558 237619 541610 237625
rect 540310 232719 540362 232725
rect 540310 232661 540362 232667
rect 539542 232571 539594 232577
rect 539542 232513 539594 232519
rect 538870 231609 538922 231615
rect 538870 231551 538922 231557
rect 538582 228575 538634 228581
rect 538582 228517 538634 228523
rect 538882 221482 538910 231551
rect 539554 221792 539582 232513
rect 539554 221764 539630 221792
rect 539602 221482 539630 221764
rect 540322 221482 540350 232661
rect 541078 228575 541130 228581
rect 541078 228517 541130 228523
rect 541090 221482 541118 228517
rect 541570 221773 541598 237619
rect 542626 236174 542654 239099
rect 561718 239083 561770 239089
rect 561718 239025 561770 239031
rect 555380 238974 555436 238983
rect 555380 238909 555436 238918
rect 553940 238382 553996 238391
rect 553940 238317 553996 238326
rect 550870 237603 550922 237609
rect 550870 237545 550922 237551
rect 541858 236146 542654 236174
rect 544342 236197 544394 236203
rect 541858 221792 541886 236146
rect 550882 236174 550910 237545
rect 544394 236146 544862 236174
rect 544342 236139 544394 236145
rect 542614 232497 542666 232503
rect 542614 232439 542666 232445
rect 541558 221767 541610 221773
rect 541558 221709 541610 221715
rect 541810 221764 541886 221792
rect 541810 221482 541838 221764
rect 542626 221704 542654 232439
rect 543382 229315 543434 229321
rect 543382 229257 543434 229263
rect 542626 221672 542664 221704
rect 542636 221482 542664 221672
rect 543394 221482 543422 229257
rect 544102 221767 544154 221773
rect 544102 221709 544154 221715
rect 544114 221482 544142 221709
rect 544834 221482 544862 236146
rect 550210 236146 550910 236174
rect 546358 232645 546410 232651
rect 546358 232587 546410 232593
rect 545590 232275 545642 232281
rect 545590 232217 545642 232223
rect 545602 221740 545630 232217
rect 546370 221792 546398 232587
rect 548566 230795 548618 230801
rect 548566 230737 548618 230743
rect 547124 224322 547180 224331
rect 547124 224257 547180 224266
rect 546370 221764 546446 221792
rect 545592 221705 545630 221740
rect 545592 221482 545620 221705
rect 546418 221482 546446 221764
rect 547138 221482 547166 224257
rect 547892 224174 547948 224183
rect 547892 224109 547948 224118
rect 547906 221482 547934 224109
rect 548578 221792 548606 230737
rect 549428 229798 549484 229807
rect 549428 229733 549484 229742
rect 548578 221764 548654 221792
rect 548626 221482 548654 221764
rect 549442 221482 549470 229733
rect 550210 221482 550238 236146
rect 550870 232349 550922 232355
rect 550870 232291 550922 232297
rect 550882 221792 550910 232291
rect 551638 232127 551690 232133
rect 551638 232069 551690 232075
rect 550882 221764 550958 221792
rect 550930 221482 550958 221764
rect 551650 221482 551678 232069
rect 552406 229241 552458 229247
rect 552406 229183 552458 229189
rect 552418 221785 552446 229183
rect 552398 221749 552446 221785
rect 553222 221767 553274 221773
rect 552398 221482 552426 221749
rect 553222 221709 553274 221715
rect 553234 221482 553262 221709
rect 553954 221482 553982 238317
rect 555394 236174 555422 238909
rect 557012 238678 557068 238687
rect 557012 238613 557068 238622
rect 556148 236310 556204 236319
rect 556148 236245 556204 236254
rect 555298 236146 555422 236174
rect 554710 232201 554762 232207
rect 554710 232143 554762 232149
rect 554722 221482 554750 232143
rect 555298 221773 555326 236146
rect 555476 232758 555532 232767
rect 555476 232693 555532 232702
rect 555490 221792 555518 232693
rect 555286 221767 555338 221773
rect 555286 221709 555338 221715
rect 555442 221764 555518 221792
rect 555442 221482 555470 221764
rect 556162 221482 556190 236245
rect 557026 221496 557054 238613
rect 559892 235866 559948 235875
rect 559222 235827 559274 235833
rect 559892 235801 559948 235810
rect 559222 235769 559274 235775
rect 557684 232610 557740 232619
rect 557684 232545 557740 232554
rect 556992 221468 557054 221496
rect 557698 221496 557726 232545
rect 559234 229247 559262 235769
rect 559222 229241 559274 229247
rect 559222 229183 559274 229189
rect 558454 229167 558506 229173
rect 558454 229109 558506 229115
rect 557698 221468 557760 221496
rect 558466 221482 558494 229109
rect 559220 224026 559276 224035
rect 559220 223961 559276 223970
rect 559234 221496 559262 223961
rect 559200 221468 559262 221496
rect 559906 221496 559934 235801
rect 560758 232053 560810 232059
rect 560758 231995 560810 232001
rect 559906 221468 559968 221496
rect 560770 221482 560798 231995
rect 561430 231979 561482 231985
rect 561430 231921 561482 231927
rect 561442 221792 561470 231921
rect 561730 228581 561758 239025
rect 576020 237050 576076 237059
rect 576020 236985 576076 236994
rect 570260 236902 570316 236911
rect 570260 236837 570316 236846
rect 567380 236754 567436 236763
rect 567380 236689 567436 236698
rect 565268 236606 565324 236615
rect 565268 236541 565324 236550
rect 562196 236458 562252 236467
rect 562196 236393 562252 236402
rect 561718 228575 561770 228581
rect 561718 228517 561770 228523
rect 561442 221764 561518 221792
rect 561490 221482 561518 221764
rect 562210 221482 562238 236393
rect 564404 236014 564460 236023
rect 564404 235949 564460 235958
rect 564310 235753 564362 235759
rect 564310 235695 564362 235701
rect 563638 231831 563690 231837
rect 563638 231773 563690 231779
rect 562966 228575 563018 228581
rect 562966 228517 563018 228523
rect 562978 221482 563006 228517
rect 563650 221792 563678 231773
rect 564322 229173 564350 235695
rect 564418 229321 564446 235949
rect 564406 229315 564458 229321
rect 564406 229257 564458 229263
rect 564310 229167 564362 229173
rect 564310 229109 564362 229115
rect 564502 229093 564554 229099
rect 564502 229035 564554 229041
rect 564514 221817 564542 229035
rect 563650 221764 563726 221792
rect 564514 221777 564562 221817
rect 563698 221482 563726 221764
rect 564534 221482 564562 221777
rect 565282 221482 565310 236541
rect 565940 232906 565996 232915
rect 565940 232841 565996 232850
rect 565954 221792 565982 232841
rect 566710 231905 566762 231911
rect 566710 231847 566762 231853
rect 565954 221764 566030 221792
rect 566002 221482 566030 221764
rect 566722 221482 566750 231847
rect 567394 228581 567422 236689
rect 570274 236174 570302 236837
rect 570274 236146 571358 236174
rect 567476 232462 567532 232471
rect 567476 232397 567532 232406
rect 567382 228575 567434 228581
rect 567382 228517 567434 228523
rect 567490 221482 567518 232397
rect 569780 232018 569836 232027
rect 569780 231953 569836 231962
rect 569014 228575 569066 228581
rect 569014 228517 569066 228523
rect 568244 223878 568300 223887
rect 568244 223813 568300 223822
rect 568258 221792 568286 223813
rect 568258 221764 568334 221792
rect 568306 221482 568334 221764
rect 569026 221482 569054 228517
rect 569794 221482 569822 231953
rect 570452 229502 570508 229511
rect 570452 229437 570508 229446
rect 570466 221792 570494 229437
rect 571330 221819 571358 236146
rect 573524 232314 573580 232323
rect 573524 232249 573580 232258
rect 572756 232166 572812 232175
rect 572756 232101 572812 232110
rect 572086 229759 572138 229765
rect 572086 229701 572138 229707
rect 570466 221764 570542 221792
rect 571330 221782 571368 221819
rect 570514 221482 570542 221764
rect 571340 221482 571368 221782
rect 572098 221482 572126 229701
rect 572770 221792 572798 232101
rect 572770 221764 572846 221792
rect 572818 221482 572846 221764
rect 573538 221482 573566 232249
rect 575060 229354 575116 229363
rect 575060 229289 575116 229298
rect 574292 223582 574348 223591
rect 574292 223517 574348 223526
rect 574306 221801 574334 223517
rect 574296 221766 574334 221801
rect 575074 221792 575102 229289
rect 575828 223730 575884 223739
rect 575828 223665 575884 223674
rect 574296 221482 574324 221766
rect 575074 221764 575150 221792
rect 575122 221482 575150 221764
rect 575842 221482 575870 223665
rect 576034 221773 576062 236985
rect 579572 235718 579628 235727
rect 579572 235653 579628 235662
rect 585238 235679 585290 235685
rect 578900 229650 578956 229659
rect 578900 229585 578956 229594
rect 576596 229206 576652 229215
rect 576596 229141 576652 229150
rect 576022 221767 576074 221773
rect 576022 221709 576074 221715
rect 576610 221482 576638 229141
rect 578038 228945 578090 228951
rect 578038 228887 578090 228893
rect 577318 221767 577370 221773
rect 577318 221709 577370 221715
rect 577330 221482 577358 221709
rect 578050 221482 578078 228887
rect 578914 221482 578942 229585
rect 579586 221792 579614 235653
rect 585238 235621 585290 235627
rect 585142 235383 585194 235389
rect 585142 235325 585194 235331
rect 582550 233829 582602 233835
rect 582550 233771 582602 233777
rect 580342 225763 580394 225769
rect 580342 225705 580394 225711
rect 579586 221764 579662 221792
rect 579634 221482 579662 221764
rect 580354 221482 580382 225705
rect 581110 225689 581162 225695
rect 581110 225631 581162 225637
rect 581122 221482 581150 225631
rect 582562 225547 582590 233771
rect 584854 227539 584906 227545
rect 584854 227481 584906 227487
rect 583414 226059 583466 226065
rect 583414 226001 583466 226007
rect 582646 225837 582698 225843
rect 582646 225779 582698 225785
rect 582550 225541 582602 225547
rect 582550 225483 582602 225489
rect 581780 223434 581836 223443
rect 581780 223369 581836 223378
rect 581794 221792 581822 223369
rect 581794 221764 581870 221792
rect 581842 221482 581870 221764
rect 582658 221482 582686 225779
rect 583426 221482 583454 226001
rect 584086 225615 584138 225621
rect 584086 225557 584138 225563
rect 584098 221792 584126 225557
rect 584098 221764 584174 221792
rect 584146 221482 584174 221764
rect 584866 221482 584894 227481
rect 585154 225695 585182 235325
rect 585250 227545 585278 235621
rect 588980 235570 589036 235579
rect 587446 235531 587498 235537
rect 588980 235505 589036 235514
rect 587446 235473 587498 235479
rect 587350 235309 587402 235315
rect 587350 235251 587402 235257
rect 585238 227539 585290 227545
rect 585238 227481 585290 227487
rect 585622 227391 585674 227397
rect 585622 227333 585674 227339
rect 585142 225689 585194 225695
rect 585142 225631 585194 225637
rect 585634 221788 585662 227333
rect 587158 225985 587210 225991
rect 587158 225927 587210 225933
rect 586390 225911 586442 225917
rect 586390 225853 586442 225859
rect 585614 221751 585662 221788
rect 586402 221774 586430 225853
rect 585614 221482 585642 221751
rect 586402 221742 586450 221774
rect 586422 221496 586450 221742
rect 586422 221468 586464 221496
rect 587170 221482 587198 225927
rect 587362 225621 587390 235251
rect 587458 226065 587486 235473
rect 588886 235457 588938 235463
rect 588886 235399 588938 235405
rect 587926 235161 587978 235167
rect 587926 235103 587978 235109
rect 587446 226059 587498 226065
rect 587446 226001 587498 226007
rect 587350 225615 587402 225621
rect 587350 225557 587402 225563
rect 587938 221496 587966 235103
rect 588598 227317 588650 227323
rect 588598 227259 588650 227265
rect 587904 221468 587966 221496
rect 588610 221496 588638 227259
rect 588898 226509 588926 235399
rect 588994 227397 589022 235505
rect 590134 235235 590186 235241
rect 590134 235177 590186 235183
rect 588982 227391 589034 227397
rect 588982 227333 589034 227339
rect 589366 227243 589418 227249
rect 589366 227185 589418 227191
rect 588886 226503 588938 226509
rect 588886 226445 588938 226451
rect 588610 221468 588672 221496
rect 589378 221482 589406 227185
rect 590146 221792 590174 235177
rect 593110 235087 593162 235093
rect 593110 235029 593162 235035
rect 590902 233089 590954 233095
rect 590902 233031 590954 233037
rect 590146 221764 590222 221792
rect 590194 221482 590222 221764
rect 590914 221482 590942 233031
rect 592342 227465 592394 227471
rect 592342 227407 592394 227413
rect 591668 226542 591724 226551
rect 591668 226477 591724 226486
rect 591682 221482 591710 226477
rect 592354 221792 592382 227407
rect 592354 221764 592430 221792
rect 592402 221482 592430 221764
rect 593122 221482 593150 235029
rect 594646 234939 594698 234945
rect 594646 234881 594698 234887
rect 593974 234865 594026 234871
rect 593974 234807 594026 234813
rect 593986 221482 594014 234807
rect 594658 221792 594686 234881
rect 596194 227249 596222 239173
rect 596276 235274 596332 235283
rect 596276 235209 596332 235218
rect 596182 227243 596234 227249
rect 596182 227185 596234 227191
rect 596290 227120 596318 235209
rect 596950 234791 597002 234797
rect 596950 234733 597002 234739
rect 596194 227092 596318 227120
rect 595412 226690 595468 226699
rect 595412 226625 595468 226634
rect 594658 221764 594734 221792
rect 594706 221482 594734 221764
rect 595426 221482 595454 226625
rect 596194 221482 596222 227092
rect 596962 221792 596990 234733
rect 599924 229058 599980 229067
rect 599924 228993 599980 229002
rect 599158 227391 599210 227397
rect 599158 227333 599210 227339
rect 598486 227169 598538 227175
rect 598486 227111 598538 227117
rect 597718 227095 597770 227101
rect 597718 227037 597770 227043
rect 596962 221764 597038 221792
rect 597010 221482 597038 221764
rect 597730 221482 597758 227037
rect 598498 221482 598526 227111
rect 599170 221792 599198 227333
rect 599170 221764 599246 221792
rect 599218 221482 599246 221764
rect 599938 221482 599966 228993
rect 600418 225991 600446 247757
rect 600502 241969 600554 241975
rect 600502 241911 600554 241917
rect 600514 227323 600542 241911
rect 601462 229019 601514 229025
rect 601462 228961 601514 228967
rect 600502 227317 600554 227323
rect 600502 227259 600554 227265
rect 600406 225985 600458 225991
rect 600406 225927 600458 225933
rect 600790 225615 600842 225621
rect 600790 225557 600842 225563
rect 600802 221482 600830 225557
rect 601474 221792 601502 228961
rect 602228 226394 602284 226403
rect 602228 226329 602284 226338
rect 601474 221764 601550 221792
rect 601522 221482 601550 221764
rect 602242 221482 602270 226329
rect 603298 225917 603326 259227
rect 603382 256399 603434 256405
rect 603382 256341 603434 256347
rect 603394 227175 603422 256341
rect 603478 253513 603530 253519
rect 603478 253455 603530 253461
rect 603382 227169 603434 227175
rect 603382 227111 603434 227117
rect 603286 225911 603338 225917
rect 603286 225853 603338 225859
rect 603490 225769 603518 253455
rect 603574 250627 603626 250633
rect 603574 250569 603626 250575
rect 603586 225843 603614 250569
rect 605972 231870 606028 231879
rect 605972 231805 606028 231814
rect 604534 230055 604586 230061
rect 604534 229997 604586 230003
rect 603670 229241 603722 229247
rect 603670 229183 603722 229189
rect 603574 225837 603626 225843
rect 603574 225779 603626 225785
rect 603478 225763 603530 225769
rect 603478 225705 603530 225711
rect 602996 223286 603052 223295
rect 602996 223221 603052 223230
rect 603010 221482 603038 223221
rect 603682 221792 603710 229183
rect 603682 221764 603758 221792
rect 603730 221482 603758 221764
rect 604546 221482 604574 229997
rect 605302 229167 605354 229173
rect 605302 229109 605354 229115
rect 605314 221482 605342 229109
rect 605986 221792 606014 231805
rect 606178 227471 606206 262113
rect 646486 256399 646538 256405
rect 646486 256341 646538 256347
rect 626326 247741 626378 247747
rect 626326 247683 626378 247689
rect 609140 235422 609196 235431
rect 609140 235357 609196 235366
rect 609046 235013 609098 235019
rect 609046 234955 609098 234961
rect 607510 229981 607562 229987
rect 607510 229923 607562 229929
rect 606742 229315 606794 229321
rect 606742 229257 606794 229263
rect 606166 227465 606218 227471
rect 606166 227407 606218 227413
rect 605986 221764 606062 221792
rect 606034 221482 606062 221764
rect 606754 221482 606782 229257
rect 607522 221781 607550 229923
rect 609058 226805 609086 234955
rect 608950 226799 609002 226805
rect 608950 226741 609002 226747
rect 609046 226799 609098 226805
rect 609046 226741 609098 226747
rect 608278 226725 608330 226731
rect 608278 226667 608330 226673
rect 607512 221744 607550 221781
rect 608290 221792 608318 226667
rect 608962 223864 608990 226741
rect 609154 226731 609182 235357
rect 612788 235126 612844 235135
rect 612788 235061 612844 235070
rect 610486 230203 610538 230209
rect 610486 230145 610538 230151
rect 609814 226947 609866 226953
rect 609814 226889 609866 226895
rect 609142 226725 609194 226731
rect 609142 226667 609194 226673
rect 608962 223836 609086 223864
rect 608290 221764 608366 221792
rect 607512 221482 607540 221744
rect 608338 221482 608366 221764
rect 609058 221482 609086 223836
rect 609826 221482 609854 226889
rect 610498 221792 610526 230145
rect 612118 227021 612170 227027
rect 612118 226963 612170 226969
rect 611254 226873 611306 226879
rect 611254 226815 611306 226821
rect 610498 221764 610574 221792
rect 610546 221482 610574 221764
rect 611266 221482 611294 226815
rect 612130 221482 612158 226963
rect 612802 221792 612830 235061
rect 618836 234978 618892 234987
rect 618836 234913 618892 234922
rect 617300 234830 617356 234839
rect 617300 234765 617356 234774
rect 613558 230129 613610 230135
rect 613558 230071 613610 230077
rect 612802 221764 612878 221792
rect 612850 221482 612878 221764
rect 613570 221482 613598 230071
rect 614998 229685 615050 229691
rect 614998 229627 615050 229633
rect 614326 226651 614378 226657
rect 614326 226593 614378 226599
rect 614338 221482 614366 226593
rect 615010 221792 615038 229627
rect 616628 228910 616684 228919
rect 616628 228845 616684 228854
rect 615862 225689 615914 225695
rect 615862 225631 615914 225637
rect 615010 221764 615086 221792
rect 615058 221482 615086 221764
rect 615874 221482 615902 225631
rect 616642 221496 616670 228845
rect 616608 221468 616670 221496
rect 617314 221496 617342 234765
rect 618070 229611 618122 229617
rect 618070 229553 618122 229559
rect 617314 221468 617376 221496
rect 618082 221482 618110 229553
rect 618850 221792 618878 234913
rect 624118 234717 624170 234723
rect 620372 234682 620428 234691
rect 624118 234659 624170 234665
rect 620372 234617 620428 234626
rect 619606 226429 619658 226435
rect 619606 226371 619658 226377
rect 618850 221764 618926 221792
rect 618898 221482 618926 221764
rect 619618 221482 619646 226371
rect 620386 221482 620414 234617
rect 621814 226577 621866 226583
rect 621814 226519 621866 226525
rect 621044 223138 621100 223147
rect 621044 223073 621100 223082
rect 621058 221792 621086 223073
rect 621058 221764 621134 221792
rect 621106 221482 621134 221764
rect 621826 221482 621854 226519
rect 622678 226355 622730 226361
rect 622678 226297 622730 226303
rect 622690 221482 622718 226297
rect 623350 226281 623402 226287
rect 623350 226223 623402 226229
rect 623362 221792 623390 226223
rect 623362 221764 623438 221792
rect 623410 221482 623438 221764
rect 624130 221482 624158 234659
rect 624884 226246 624940 226255
rect 624884 226181 624940 226190
rect 624898 221482 624926 226181
rect 625556 226098 625612 226107
rect 625556 226033 625612 226042
rect 625570 221792 625598 226033
rect 626338 225769 626366 247683
rect 629206 244855 629258 244861
rect 629206 244797 629258 244803
rect 629218 226509 629246 244797
rect 630166 227539 630218 227545
rect 630166 227481 630218 227487
rect 629398 226799 629450 226805
rect 629398 226741 629450 226747
rect 626422 226503 626474 226509
rect 626422 226445 626474 226451
rect 629206 226503 629258 226509
rect 629206 226445 629258 226451
rect 626326 225763 626378 225769
rect 626326 225705 626378 225711
rect 626434 221857 626462 226445
rect 627862 226133 627914 226139
rect 627862 226075 627914 226081
rect 627190 225541 627242 225547
rect 627190 225483 627242 225489
rect 626434 221818 626472 221857
rect 625570 221764 625646 221792
rect 625618 221482 625646 221764
rect 626444 221482 626472 221818
rect 627202 221482 627230 225483
rect 627874 221792 627902 226075
rect 628630 225171 628682 225177
rect 628630 225113 628682 225119
rect 627874 221764 627950 221792
rect 627922 221482 627950 221764
rect 628642 221482 628670 225113
rect 629410 221482 629438 226741
rect 630178 221792 630206 227481
rect 639958 227391 640010 227397
rect 639958 227333 640010 227339
rect 634678 227317 634730 227323
rect 634678 227259 634730 227265
rect 633142 227243 633194 227249
rect 633142 227185 633194 227191
rect 630934 226725 630986 226731
rect 630934 226667 630986 226673
rect 630178 221764 630254 221792
rect 630226 221482 630254 221764
rect 630946 221482 630974 226667
rect 632374 226207 632426 226213
rect 632374 226149 632426 226155
rect 631702 226059 631754 226065
rect 631702 226001 631754 226007
rect 631714 221482 631742 226001
rect 632386 221792 632414 226149
rect 632386 221764 632462 221792
rect 632434 221482 632462 221764
rect 633154 221482 633182 227185
rect 634006 226503 634058 226509
rect 634006 226445 634058 226451
rect 634018 221482 634046 226445
rect 634690 221792 634718 227259
rect 638518 227169 638570 227175
rect 638518 227111 638570 227117
rect 636214 225985 636266 225991
rect 636214 225927 636266 225933
rect 635446 225763 635498 225769
rect 635446 225705 635498 225711
rect 634690 221764 634766 221792
rect 634738 221482 634766 221764
rect 635458 221482 635486 225705
rect 636226 221482 636254 225927
rect 636886 225837 636938 225843
rect 636886 225779 636938 225785
rect 636898 221792 636926 225779
rect 637750 225689 637802 225695
rect 637750 225631 637802 225637
rect 636898 221764 636974 221792
rect 636946 221482 636974 221764
rect 637762 221482 637790 225631
rect 638530 221482 638558 227111
rect 639190 225911 639242 225917
rect 639190 225853 639242 225859
rect 639202 221792 639230 225853
rect 639202 221764 639278 221792
rect 639250 221482 639278 221764
rect 639970 221482 639998 227333
rect 645142 221323 645194 221329
rect 645142 221265 645194 221271
rect 645154 221223 645182 221265
rect 645140 221214 645196 221223
rect 645140 221149 645196 221158
rect 645142 216883 645194 216889
rect 645142 216825 645194 216831
rect 645154 216014 645182 216825
rect 645058 215986 645182 216014
rect 645058 215895 645086 215986
rect 645044 215886 645100 215895
rect 645044 215821 645100 215830
rect 645142 212961 645194 212967
rect 645140 212926 645142 212935
rect 645194 212926 645196 212935
rect 645140 212861 645196 212870
rect 645142 209853 645194 209859
rect 645142 209795 645194 209801
rect 645154 209679 645182 209795
rect 645140 209670 645196 209679
rect 645140 209605 645196 209614
rect 645142 206079 645194 206085
rect 645142 206021 645194 206027
rect 645154 205979 645182 206021
rect 645140 205970 645196 205979
rect 645140 205905 645196 205914
rect 645142 201565 645194 201571
rect 645140 201530 645142 201539
rect 645194 201530 645196 201539
rect 645140 201465 645196 201474
rect 187220 199162 187276 199171
rect 187220 199097 187276 199106
rect 645142 198531 645194 198537
rect 645142 198473 645194 198479
rect 645154 198283 645182 198473
rect 645140 198274 645196 198283
rect 645140 198209 645196 198218
rect 185986 195826 186206 195854
rect 186178 174751 186206 195826
rect 645142 194017 645194 194023
rect 645140 193982 645142 193991
rect 645194 193982 645196 193991
rect 645140 193917 645196 193926
rect 645142 190465 645194 190471
rect 645142 190407 645194 190413
rect 645154 190143 645182 190407
rect 645140 190134 645196 190143
rect 645140 190069 645196 190078
rect 646198 184619 646250 184625
rect 646198 184561 646250 184567
rect 646210 184371 646238 184561
rect 646196 184362 646252 184371
rect 646196 184297 646252 184306
rect 645910 183139 645962 183145
rect 645910 183081 645962 183087
rect 645922 183039 645950 183081
rect 645908 183030 645964 183039
rect 645908 182965 645964 182974
rect 646006 179439 646058 179445
rect 646006 179381 646058 179387
rect 646018 179339 646046 179381
rect 646004 179330 646060 179339
rect 646004 179265 646060 179274
rect 645142 174925 645194 174931
rect 645140 174890 645142 174899
rect 645194 174890 645196 174899
rect 645140 174825 645196 174834
rect 186164 174742 186220 174751
rect 186164 174677 186220 174686
rect 185780 173262 185836 173271
rect 185780 173197 185836 173206
rect 645142 171447 645194 171453
rect 645142 171389 645194 171395
rect 645154 171051 645182 171389
rect 645140 171042 645196 171051
rect 645140 170977 645196 170986
rect 645142 168043 645194 168049
rect 645142 167985 645194 167991
rect 645154 167795 645182 167985
rect 645140 167786 645196 167795
rect 645140 167721 645196 167730
rect 645526 161827 645578 161833
rect 645526 161769 645578 161775
rect 645538 161431 645566 161769
rect 645524 161422 645580 161431
rect 645524 161357 645580 161366
rect 645526 158497 645578 158503
rect 645526 158439 645578 158445
rect 645538 157583 645566 158439
rect 645524 157574 645580 157583
rect 645524 157509 645580 157518
rect 645142 155907 645194 155913
rect 645142 155849 645194 155855
rect 645154 155511 645182 155849
rect 645140 155502 645196 155511
rect 645140 155437 645196 155446
rect 646006 152577 646058 152583
rect 646004 152542 646006 152551
rect 646058 152542 646060 152551
rect 646004 152477 646060 152486
rect 645142 149395 645194 149401
rect 645142 149337 645194 149343
rect 645154 148111 645182 149337
rect 645140 148102 645196 148111
rect 645140 148037 645196 148046
rect 185782 146879 185834 146885
rect 185782 146821 185834 146827
rect 185794 146631 185822 146821
rect 185780 146622 185836 146631
rect 185780 146557 185836 146566
rect 646498 144263 646526 256341
rect 646582 210297 646634 210303
rect 646582 210239 646634 210245
rect 646484 144254 646540 144263
rect 646484 144189 646540 144198
rect 646594 141007 646622 210239
rect 649378 194023 649406 987017
rect 649474 198537 649502 987387
rect 649570 201571 649598 989459
rect 649654 989443 649706 989449
rect 649654 989385 649706 989391
rect 649666 206085 649694 989385
rect 658006 989369 658058 989375
rect 658006 989311 658058 989317
rect 649750 989295 649802 989301
rect 649750 989237 649802 989243
rect 649762 209859 649790 989237
rect 650902 987815 650954 987821
rect 650902 987757 650954 987763
rect 649846 986853 649898 986859
rect 649846 986795 649898 986801
rect 649858 212967 649886 986795
rect 649942 986557 649994 986563
rect 649942 986499 649994 986505
rect 649954 216889 649982 986499
rect 650038 983523 650090 983529
rect 650038 983465 650090 983471
rect 650050 221329 650078 983465
rect 650038 221323 650090 221329
rect 650038 221265 650090 221271
rect 649942 216883 649994 216889
rect 649942 216825 649994 216831
rect 649846 212961 649898 212967
rect 649846 212903 649898 212909
rect 649750 209853 649802 209859
rect 649750 209795 649802 209801
rect 649654 206079 649706 206085
rect 649654 206021 649706 206027
rect 649558 201565 649610 201571
rect 649558 201507 649610 201513
rect 649462 198531 649514 198537
rect 649462 198473 649514 198479
rect 649366 194017 649418 194023
rect 649366 193959 649418 193965
rect 646678 167303 646730 167309
rect 646678 167245 646730 167251
rect 646580 140998 646636 141007
rect 185686 140959 185738 140965
rect 646580 140933 646636 140942
rect 185686 140901 185738 140907
rect 184628 138334 184684 138343
rect 184628 138269 184684 138278
rect 184534 138221 184586 138227
rect 184534 138163 184586 138169
rect 184342 138147 184394 138153
rect 184342 138089 184394 138095
rect 184354 137455 184382 138089
rect 184438 138073 184490 138079
rect 184438 138015 184490 138021
rect 184340 137446 184396 137455
rect 184340 137381 184396 137390
rect 184450 135975 184478 138015
rect 184546 136863 184574 138163
rect 184532 136854 184588 136863
rect 184532 136789 184588 136798
rect 184436 135966 184492 135975
rect 184436 135901 184492 135910
rect 184438 135335 184490 135341
rect 184438 135277 184490 135283
rect 184342 135261 184394 135267
rect 184340 135226 184342 135235
rect 184394 135226 184396 135235
rect 184340 135161 184396 135170
rect 184342 135113 184394 135119
rect 184342 135055 184394 135061
rect 184354 133755 184382 135055
rect 184450 134495 184478 135277
rect 184534 135187 184586 135193
rect 184534 135129 184586 135135
rect 184436 134486 184492 134495
rect 184436 134421 184492 134430
rect 184340 133746 184396 133755
rect 184340 133681 184396 133690
rect 184546 133015 184574 135129
rect 184532 133006 184588 133015
rect 184532 132941 184588 132950
rect 646582 132523 646634 132529
rect 646582 132465 646634 132471
rect 184630 132449 184682 132455
rect 184630 132391 184682 132397
rect 184534 132375 184586 132381
rect 184534 132317 184586 132323
rect 184438 132301 184490 132307
rect 184340 132266 184396 132275
rect 184438 132243 184490 132249
rect 184340 132201 184342 132210
rect 184394 132201 184396 132210
rect 184342 132169 184394 132175
rect 184450 131535 184478 132243
rect 184436 131526 184492 131535
rect 184436 131461 184492 131470
rect 184546 130647 184574 132317
rect 184532 130638 184588 130647
rect 184532 130573 184588 130582
rect 184642 129907 184670 132391
rect 184628 129898 184684 129907
rect 184628 129833 184684 129842
rect 184342 129563 184394 129569
rect 184342 129505 184394 129511
rect 184354 129167 184382 129505
rect 184438 129489 184490 129495
rect 184438 129431 184490 129437
rect 184340 129158 184396 129167
rect 184340 129093 184396 129102
rect 184450 128427 184478 129431
rect 184534 129415 184586 129421
rect 184534 129357 184586 129363
rect 184436 128418 184492 128427
rect 184436 128353 184492 128362
rect 184546 127687 184574 129357
rect 184726 129341 184778 129347
rect 184726 129283 184778 129289
rect 184532 127678 184588 127687
rect 184532 127613 184588 127622
rect 184738 126947 184766 129283
rect 646594 129019 646622 132465
rect 646580 129010 646636 129019
rect 646580 128945 646636 128954
rect 184724 126938 184780 126947
rect 184724 126873 184780 126882
rect 184342 126677 184394 126683
rect 184342 126619 184394 126625
rect 182998 126529 183050 126535
rect 182998 126471 183050 126477
rect 184354 126059 184382 126619
rect 184438 126603 184490 126609
rect 184438 126545 184490 126551
rect 184340 126050 184396 126059
rect 184340 125985 184396 125994
rect 184450 124579 184478 126545
rect 186838 126529 186890 126535
rect 186838 126471 186890 126477
rect 186850 125467 186878 126471
rect 646690 125763 646718 167245
rect 646870 167229 646922 167235
rect 646870 167171 646922 167177
rect 646774 167155 646826 167161
rect 646774 167097 646826 167103
rect 646786 127687 646814 167097
rect 646882 134791 646910 167171
rect 646868 134782 646924 134791
rect 646868 134717 646924 134726
rect 647828 130934 647884 130943
rect 647828 130869 647884 130878
rect 647734 129711 647786 129717
rect 647734 129653 647786 129659
rect 646772 127678 646828 127687
rect 646772 127613 646828 127622
rect 646676 125754 646732 125763
rect 646676 125689 646732 125698
rect 186836 125458 186892 125467
rect 186836 125393 186892 125402
rect 184436 124570 184492 124579
rect 184436 124505 184492 124514
rect 184630 123865 184682 123871
rect 184340 123830 184396 123839
rect 184630 123807 184682 123813
rect 184340 123765 184396 123774
rect 184438 123791 184490 123797
rect 184354 123649 184382 123765
rect 184438 123733 184490 123739
rect 184342 123643 184394 123649
rect 184342 123585 184394 123591
rect 184450 122211 184478 123733
rect 184534 123717 184586 123723
rect 184534 123659 184586 123665
rect 184436 122202 184492 122211
rect 184436 122137 184492 122146
rect 184546 121619 184574 123659
rect 184642 123099 184670 123807
rect 184628 123090 184684 123099
rect 184628 123025 184684 123034
rect 647746 122063 647774 129653
rect 647732 122054 647788 122063
rect 647732 121989 647788 121998
rect 184532 121610 184588 121619
rect 184532 121545 184588 121554
rect 646678 121275 646730 121281
rect 646678 121217 646730 121223
rect 184534 120979 184586 120985
rect 184534 120921 184586 120927
rect 184342 120831 184394 120837
rect 184342 120773 184394 120779
rect 184354 120731 184382 120773
rect 184438 120757 184490 120763
rect 184340 120722 184396 120731
rect 184438 120699 184490 120705
rect 184340 120657 184396 120666
rect 184450 118659 184478 120699
rect 184546 120139 184574 120921
rect 184630 120905 184682 120911
rect 184630 120847 184682 120853
rect 184532 120130 184588 120139
rect 184532 120065 184588 120074
rect 184642 119251 184670 120847
rect 184628 119242 184684 119251
rect 184628 119177 184684 119186
rect 184436 118650 184492 118659
rect 184436 118585 184492 118594
rect 184630 118093 184682 118099
rect 184630 118035 184682 118041
rect 184342 118019 184394 118025
rect 184342 117961 184394 117967
rect 151894 117871 151946 117877
rect 151894 117813 151946 117819
rect 184354 117771 184382 117961
rect 184438 117945 184490 117951
rect 184438 117887 184490 117893
rect 184340 117762 184396 117771
rect 184340 117697 184396 117706
rect 184450 117031 184478 117887
rect 184534 117871 184586 117877
rect 184534 117813 184586 117819
rect 184436 117022 184492 117031
rect 184436 116957 184492 116966
rect 184546 115403 184574 117813
rect 184642 116291 184670 118035
rect 646690 117623 646718 121217
rect 647842 121133 647870 130869
rect 650914 129643 650942 987757
rect 650998 987741 651050 987747
rect 650998 987683 651050 987689
rect 651010 129865 651038 987683
rect 652246 987371 652298 987377
rect 652246 987313 652298 987319
rect 652258 175935 652286 987313
rect 652438 987297 652490 987303
rect 652438 987239 652490 987245
rect 652342 982857 652394 982863
rect 652342 982799 652394 982805
rect 652354 616415 652382 982799
rect 652342 616409 652394 616415
rect 652342 616351 652394 616357
rect 652342 613523 652394 613529
rect 652342 613465 652394 613471
rect 652244 175926 652300 175935
rect 652244 175861 652300 175870
rect 652354 171453 652382 613465
rect 652450 175787 652478 987239
rect 653782 986705 653834 986711
rect 653782 986647 653834 986653
rect 652630 983449 652682 983455
rect 652630 983391 652682 983397
rect 652534 983301 652586 983307
rect 652534 983243 652586 983249
rect 652546 751761 652574 983243
rect 652534 751755 652586 751761
rect 652534 751697 652586 751703
rect 652534 715717 652586 715723
rect 652534 715659 652586 715665
rect 652546 278457 652574 715659
rect 652642 550259 652670 983391
rect 652918 983375 652970 983381
rect 652918 983317 652970 983323
rect 652822 983227 652874 983233
rect 652822 983169 652874 983175
rect 652726 982931 652778 982937
rect 652726 982873 652778 982879
rect 652738 559879 652766 982873
rect 652834 582005 652862 983169
rect 652930 789131 652958 983317
rect 653014 983153 653066 983159
rect 653014 983095 653066 983101
rect 653026 797863 653054 983095
rect 653014 797857 653066 797863
rect 653014 797799 653066 797805
rect 652918 789125 652970 789131
rect 652918 789067 652970 789073
rect 652918 607751 652970 607757
rect 652918 607693 652970 607699
rect 652822 581999 652874 582005
rect 652822 581941 652874 581947
rect 652822 567421 652874 567427
rect 652822 567363 652874 567369
rect 652726 559873 652778 559879
rect 652726 559815 652778 559821
rect 652630 550253 652682 550259
rect 652630 550195 652682 550201
rect 652630 370137 652682 370143
rect 652630 370079 652682 370085
rect 652534 278451 652586 278457
rect 652534 278393 652586 278399
rect 652642 278055 652670 370079
rect 652726 362885 652778 362891
rect 652726 362827 652778 362833
rect 652738 278605 652766 362827
rect 652726 278599 652778 278605
rect 652726 278541 652778 278547
rect 652628 278046 652684 278055
rect 652628 277981 652684 277990
rect 652436 175778 652492 175787
rect 652436 175713 652492 175722
rect 652342 171447 652394 171453
rect 652342 171389 652394 171395
rect 652834 168049 652862 567363
rect 652930 278679 652958 607693
rect 653014 602053 653066 602059
rect 653014 601995 653066 602001
rect 652918 278673 652970 278679
rect 652918 278615 652970 278621
rect 653026 278531 653054 601995
rect 653014 278525 653066 278531
rect 653014 278467 653066 278473
rect 653794 190471 653822 986647
rect 655126 986631 655178 986637
rect 655126 986573 655178 986579
rect 654452 909562 654508 909571
rect 654452 909497 654508 909506
rect 654466 908789 654494 909497
rect 654454 908783 654506 908789
rect 654454 908725 654506 908731
rect 654452 896242 654508 896251
rect 654452 896177 654508 896186
rect 654466 895765 654494 896177
rect 654454 895759 654506 895765
rect 654454 895701 654506 895707
rect 654452 869750 654508 869759
rect 654452 869685 654508 869694
rect 654466 869347 654494 869685
rect 654454 869341 654506 869347
rect 654454 869283 654506 869289
rect 654452 856430 654508 856439
rect 654452 856365 654508 856374
rect 654466 855435 654494 856365
rect 654454 855429 654506 855435
rect 654454 855371 654506 855377
rect 654452 842962 654508 842971
rect 654452 842897 654508 842906
rect 654466 841005 654494 842897
rect 654454 840999 654506 841005
rect 654454 840941 654506 840947
rect 654740 829790 654796 829799
rect 654740 829725 654796 829734
rect 654754 829535 654782 829725
rect 654742 829529 654794 829535
rect 654742 829471 654794 829477
rect 654452 803150 654508 803159
rect 654452 803085 654508 803094
rect 654466 800675 654494 803085
rect 654454 800669 654506 800675
rect 654454 800611 654506 800617
rect 654452 763338 654508 763347
rect 654452 763273 654454 763282
rect 654506 763273 654508 763282
rect 654454 763241 654506 763247
rect 654452 750166 654508 750175
rect 654452 750101 654508 750110
rect 654466 748949 654494 750101
rect 654454 748943 654506 748949
rect 654454 748885 654506 748891
rect 654452 736846 654508 736855
rect 654452 736781 654508 736790
rect 654466 735925 654494 736781
rect 654454 735919 654506 735925
rect 654454 735861 654506 735867
rect 654452 710354 654508 710363
rect 654452 710289 654454 710298
rect 654506 710289 654508 710298
rect 654454 710257 654506 710263
rect 654452 697034 654508 697043
rect 654452 696969 654454 696978
rect 654506 696969 654508 696978
rect 654454 696937 654506 696943
rect 654452 683566 654508 683575
rect 654452 683501 654508 683510
rect 654466 682645 654494 683501
rect 654454 682639 654506 682645
rect 654454 682581 654506 682587
rect 654452 657074 654508 657083
rect 654452 657009 654508 657018
rect 654466 656745 654494 657009
rect 654454 656739 654506 656745
rect 654454 656681 654506 656687
rect 654452 643754 654508 643763
rect 654452 643689 654508 643698
rect 654466 642315 654494 643689
rect 654454 642309 654506 642315
rect 654454 642251 654506 642257
rect 654452 630582 654508 630591
rect 654452 630517 654508 630526
rect 654466 627885 654494 630517
rect 654454 627879 654506 627885
rect 654454 627821 654506 627827
rect 654548 617262 654604 617271
rect 654548 617197 654604 617206
rect 653878 614559 653930 614565
rect 653878 614501 653930 614507
rect 653890 607757 653918 614501
rect 653878 607751 653930 607757
rect 653878 607693 653930 607699
rect 654452 603942 654508 603951
rect 654452 603877 654508 603886
rect 654466 601985 654494 603877
rect 654562 603391 654590 617197
rect 654550 603385 654602 603391
rect 654550 603327 654602 603333
rect 654454 601979 654506 601985
rect 654454 601921 654506 601927
rect 654452 590770 654508 590779
rect 654452 590705 654508 590714
rect 654466 590441 654494 590705
rect 654454 590435 654506 590441
rect 654454 590377 654506 590383
rect 654452 577450 654508 577459
rect 654452 577385 654508 577394
rect 654466 577343 654494 577385
rect 654454 577337 654506 577343
rect 654454 577279 654506 577285
rect 654836 550958 654892 550967
rect 654836 550893 654892 550902
rect 654850 550185 654878 550893
rect 654838 550179 654890 550185
rect 654838 550121 654890 550127
rect 654452 537638 654508 537647
rect 654452 537573 654508 537582
rect 654466 537531 654494 537573
rect 654454 537525 654506 537531
rect 654454 537467 654506 537473
rect 654452 524318 654508 524327
rect 654452 524253 654454 524262
rect 654506 524253 654508 524262
rect 654454 524221 654506 524227
rect 654452 510998 654508 511007
rect 654452 510933 654508 510942
rect 654466 509855 654494 510933
rect 654454 509849 654506 509855
rect 654454 509791 654506 509797
rect 654452 497678 654508 497687
rect 654452 497613 654508 497622
rect 654466 495425 654494 497613
rect 654454 495419 654506 495425
rect 654454 495361 654506 495367
rect 654452 484358 654508 484367
rect 654452 484293 654508 484302
rect 654466 484103 654494 484293
rect 654454 484097 654506 484103
rect 654454 484039 654506 484045
rect 654452 471186 654508 471195
rect 654452 471121 654508 471130
rect 654466 469525 654494 471121
rect 654454 469519 654506 469525
rect 654454 469461 654506 469467
rect 654452 457866 654508 457875
rect 654452 457801 654508 457810
rect 654466 455095 654494 457801
rect 654454 455089 654506 455095
rect 654454 455031 654506 455037
rect 654452 444546 654508 444555
rect 654452 444481 654508 444490
rect 654466 443625 654494 444481
rect 654454 443619 654506 443625
rect 654454 443561 654506 443567
rect 654452 431374 654508 431383
rect 654452 431309 654508 431318
rect 654466 429195 654494 431309
rect 654454 429189 654506 429195
rect 654454 429131 654506 429137
rect 654452 418054 654508 418063
rect 654452 417989 654508 417998
rect 654466 417651 654494 417989
rect 654454 417645 654506 417651
rect 654454 417587 654506 417593
rect 654452 404734 654508 404743
rect 654452 404669 654508 404678
rect 654466 403295 654494 404669
rect 654454 403289 654506 403295
rect 654454 403231 654506 403237
rect 654836 391562 654892 391571
rect 654836 391497 654892 391506
rect 654850 390789 654878 391497
rect 654838 390783 654890 390789
rect 654838 390725 654890 390731
rect 654452 378242 654508 378251
rect 654452 378177 654508 378186
rect 654466 377321 654494 378177
rect 654454 377315 654506 377321
rect 654454 377257 654506 377263
rect 654452 364922 654508 364931
rect 654452 364857 654454 364866
rect 654506 364857 654508 364866
rect 654454 364825 654506 364831
rect 654452 351602 654508 351611
rect 654452 351537 654508 351546
rect 654466 351421 654494 351537
rect 654454 351415 654506 351421
rect 654454 351357 654506 351363
rect 654836 324962 654892 324971
rect 654836 324897 654892 324906
rect 654850 323301 654878 324897
rect 654838 323295 654890 323301
rect 654838 323237 654890 323243
rect 654452 311790 654508 311799
rect 654452 311725 654508 311734
rect 654466 311091 654494 311725
rect 655138 311207 655166 986573
rect 655414 983079 655466 983085
rect 655414 983021 655466 983027
rect 655318 983005 655370 983011
rect 655318 982947 655370 982953
rect 655220 975866 655276 975875
rect 655220 975801 655276 975810
rect 655234 939129 655262 975801
rect 655222 939123 655274 939129
rect 655222 939065 655274 939071
rect 655220 776658 655276 776667
rect 655220 776593 655276 776602
rect 655234 738737 655262 776593
rect 655222 738731 655274 738737
rect 655222 738673 655274 738679
rect 655220 723526 655276 723535
rect 655220 723461 655276 723470
rect 655234 692635 655262 723461
rect 655222 692629 655274 692635
rect 655222 692571 655274 692577
rect 655222 659551 655274 659557
rect 655222 659493 655274 659499
rect 655124 311198 655180 311207
rect 655124 311133 655180 311142
rect 654454 311085 654506 311091
rect 654454 311027 654506 311033
rect 655124 298470 655180 298479
rect 655124 298405 655180 298414
rect 653782 190465 653834 190471
rect 653782 190407 653834 190413
rect 652822 168043 652874 168049
rect 652822 167985 652874 167991
rect 655138 132677 655166 298405
rect 655234 174931 655262 659493
rect 655330 627811 655358 982947
rect 655426 662369 655454 983021
rect 655508 962546 655564 962555
rect 655508 962481 655564 962490
rect 655522 939277 655550 962481
rect 655606 959177 655658 959183
rect 655606 959119 655658 959125
rect 655510 939271 655562 939277
rect 655510 939213 655562 939219
rect 655618 936211 655646 959119
rect 655700 949374 655756 949383
rect 655700 949309 655756 949318
rect 655714 939425 655742 949309
rect 655702 939419 655754 939425
rect 655702 939361 655754 939367
rect 655604 936202 655660 936211
rect 655604 936137 655660 936146
rect 656372 922734 656428 922743
rect 656372 922669 656428 922678
rect 656386 921665 656414 922669
rect 656374 921659 656426 921665
rect 656374 921601 656426 921607
rect 656564 882922 656620 882931
rect 656564 882857 656620 882866
rect 656578 871197 656606 882857
rect 656566 871191 656618 871197
rect 656566 871133 656618 871139
rect 655508 816470 655564 816479
rect 655508 816405 655564 816414
rect 655522 815105 655550 816405
rect 655510 815099 655562 815105
rect 655510 815041 655562 815047
rect 657910 797783 657962 797789
rect 657910 797725 657962 797731
rect 655604 789978 655660 789987
rect 655604 789913 655660 789922
rect 655618 789205 655646 789913
rect 655606 789199 655658 789205
rect 655606 789141 655658 789147
rect 657922 789131 657950 797725
rect 655510 789125 655562 789131
rect 655510 789067 655562 789073
rect 657910 789125 657962 789131
rect 657910 789067 657962 789073
rect 655522 761825 655550 789067
rect 655510 761819 655562 761825
rect 655510 761761 655562 761767
rect 655510 751755 655562 751761
rect 655510 751697 655562 751703
rect 655522 731929 655550 751697
rect 655510 731923 655562 731929
rect 655510 731865 655562 731871
rect 655508 670394 655564 670403
rect 655508 670329 655564 670338
rect 655414 662363 655466 662369
rect 655414 662305 655466 662311
rect 655522 646607 655550 670329
rect 655510 646601 655562 646607
rect 655510 646543 655562 646549
rect 655318 627805 655370 627811
rect 655318 627747 655370 627753
rect 655318 616409 655370 616415
rect 655318 616351 655370 616357
rect 655330 588665 655358 616351
rect 655318 588659 655370 588665
rect 655318 588601 655370 588607
rect 656564 564130 656620 564139
rect 656564 564065 656620 564074
rect 656578 557289 656606 564065
rect 656566 557283 656618 557289
rect 656566 557225 656618 557231
rect 656566 550253 656618 550259
rect 656566 550195 656618 550201
rect 656578 544432 656606 550195
rect 656578 544404 656702 544432
rect 656674 541601 656702 544404
rect 656662 541595 656714 541601
rect 656662 541537 656714 541543
rect 655318 378721 655370 378727
rect 655318 378663 655370 378669
rect 655330 362891 655358 378663
rect 655318 362885 655370 362891
rect 655318 362827 655370 362833
rect 655316 338282 655372 338291
rect 655316 338217 655372 338226
rect 655330 178705 655358 338217
rect 655412 285298 655468 285307
rect 655412 285233 655468 285242
rect 655318 178699 655370 178705
rect 655318 178641 655370 178647
rect 655222 174925 655274 174931
rect 655222 174867 655274 174873
rect 655426 132825 655454 285233
rect 658018 219003 658046 989311
rect 658102 987223 658154 987229
rect 658102 987165 658154 987171
rect 658114 221815 658142 987165
rect 658198 987001 658250 987007
rect 658198 986943 658250 986949
rect 658210 265031 658238 986943
rect 658390 986927 658442 986933
rect 658390 986869 658442 986875
rect 658294 748869 658346 748875
rect 658294 748811 658346 748817
rect 658196 265022 658252 265031
rect 658196 264957 658252 264966
rect 658100 221806 658156 221815
rect 658100 221741 658156 221750
rect 658004 218994 658060 219003
rect 658004 218929 658060 218938
rect 658306 183145 658334 748811
rect 658402 265179 658430 986869
rect 660898 939795 660926 989533
rect 669622 986483 669674 986489
rect 669622 986425 669674 986431
rect 660982 983745 661034 983751
rect 660982 983687 661034 983693
rect 660886 939789 660938 939795
rect 660886 939731 660938 939737
rect 660886 927431 660938 927437
rect 660886 927373 660938 927379
rect 658870 731923 658922 731929
rect 658870 731865 658922 731871
rect 658882 728599 658910 731865
rect 658870 728593 658922 728599
rect 658870 728535 658922 728541
rect 658486 702767 658538 702773
rect 658486 702709 658538 702715
rect 658388 265170 658444 265179
rect 658388 265105 658444 265114
rect 658294 183139 658346 183145
rect 658294 183081 658346 183087
rect 658498 179445 658526 702709
rect 659062 662363 659114 662369
rect 659062 662305 659114 662311
rect 659074 653859 659102 662305
rect 659062 653853 659114 653859
rect 659062 653795 659114 653801
rect 660598 607973 660650 607979
rect 660598 607915 660650 607921
rect 660610 602059 660638 607915
rect 660598 602053 660650 602059
rect 660598 601995 660650 602001
rect 658870 588659 658922 588665
rect 658870 588601 658922 588607
rect 658882 586075 658910 588601
rect 658870 586069 658922 586075
rect 658870 586011 658922 586017
rect 658582 345643 658634 345649
rect 658582 345585 658634 345591
rect 658486 179439 658538 179445
rect 658486 179381 658538 179387
rect 658594 152583 658622 345585
rect 658678 302575 658730 302581
rect 658678 302517 658730 302523
rect 658582 152577 658634 152583
rect 658582 152519 658634 152525
rect 658690 149401 658718 302517
rect 660898 184625 660926 927373
rect 660994 311059 661022 983687
rect 666646 921659 666698 921665
rect 666646 921601 666698 921607
rect 661078 908783 661130 908789
rect 661078 908725 661130 908731
rect 661090 762935 661118 908725
rect 663766 869341 663818 869347
rect 663766 869283 663818 869289
rect 661270 829529 661322 829535
rect 661270 829471 661322 829477
rect 661174 815099 661226 815105
rect 661174 815041 661226 815047
rect 661078 762929 661130 762935
rect 661078 762871 661130 762877
rect 661186 672359 661214 815041
rect 661282 783359 661310 829471
rect 662326 789125 662378 789131
rect 662326 789067 662378 789073
rect 662338 783729 662366 789067
rect 662326 783723 662378 783729
rect 662326 783665 662378 783671
rect 661270 783353 661322 783359
rect 661270 783295 661322 783301
rect 661270 735919 661322 735925
rect 661270 735861 661322 735867
rect 661174 672353 661226 672359
rect 661174 672295 661226 672301
rect 661078 656739 661130 656745
rect 661078 656681 661130 656687
rect 661090 536939 661118 656681
rect 661282 626627 661310 735861
rect 662134 728593 662186 728599
rect 662134 728535 662186 728541
rect 662146 720977 662174 728535
rect 662134 720971 662186 720977
rect 662134 720913 662186 720919
rect 663382 720971 663434 720977
rect 663382 720913 663434 720919
rect 663394 717203 663422 720913
rect 663778 717351 663806 869283
rect 663862 789199 663914 789205
rect 663862 789141 663914 789147
rect 663766 717345 663818 717351
rect 663766 717287 663818 717293
rect 663382 717197 663434 717203
rect 663382 717139 663434 717145
rect 663766 710315 663818 710321
rect 663766 710257 663818 710263
rect 661270 626621 661322 626627
rect 661270 626563 661322 626569
rect 661172 625106 661228 625115
rect 661172 625041 661228 625050
rect 661186 614565 661214 625041
rect 661174 614559 661226 614565
rect 661174 614501 661226 614507
rect 663778 582005 663806 710257
rect 663874 671619 663902 789141
rect 666658 762343 666686 921601
rect 669526 866973 669578 866979
rect 669526 866915 669578 866921
rect 666742 840999 666794 841005
rect 666742 840941 666794 840947
rect 666646 762337 666698 762343
rect 666646 762279 666698 762285
rect 666358 761819 666410 761825
rect 666358 761761 666410 761767
rect 666370 758865 666398 761761
rect 666358 758859 666410 758865
rect 666358 758801 666410 758807
rect 666646 748943 666698 748949
rect 666646 748885 666698 748891
rect 663862 671613 663914 671619
rect 663862 671555 663914 671561
rect 665014 653779 665066 653785
rect 665014 653721 665066 653727
rect 665026 640465 665054 653721
rect 665014 640459 665066 640465
rect 665014 640401 665066 640407
rect 663958 627879 664010 627885
rect 663958 627821 664010 627827
rect 663766 581999 663818 582005
rect 663766 581941 663818 581947
rect 661174 577337 661226 577343
rect 661174 577279 661226 577285
rect 661078 536933 661130 536939
rect 661078 536875 661130 536881
rect 661078 524205 661130 524211
rect 661078 524147 661130 524153
rect 660980 311050 661036 311059
rect 660980 310985 661036 310994
rect 660886 184619 660938 184625
rect 660886 184561 660938 184567
rect 661090 161833 661118 524147
rect 661186 492391 661214 577279
rect 663766 559873 663818 559879
rect 663766 559815 663818 559821
rect 663778 541379 663806 559815
rect 663766 541373 663818 541379
rect 663766 541315 663818 541321
rect 663862 537525 663914 537531
rect 663862 537467 663914 537473
rect 661174 492385 661226 492391
rect 661174 492327 661226 492333
rect 661462 484097 661514 484103
rect 661462 484039 661514 484045
rect 661174 479509 661226 479515
rect 661174 479451 661226 479457
rect 661078 161827 661130 161833
rect 661078 161769 661130 161775
rect 661186 158503 661214 479451
rect 661270 391745 661322 391751
rect 661270 391687 661322 391693
rect 661174 158497 661226 158503
rect 661174 158439 661226 158445
rect 661282 155913 661310 391687
rect 661366 390783 661418 390789
rect 661366 390725 661418 390731
rect 661378 224363 661406 390725
rect 661474 359043 661502 484039
rect 661558 455089 661610 455095
rect 661558 455031 661610 455037
rect 661462 359037 661514 359043
rect 661462 358979 661514 358985
rect 661462 323295 661514 323301
rect 661462 323237 661514 323243
rect 661366 224357 661418 224363
rect 661366 224299 661418 224305
rect 661474 178853 661502 323237
rect 661570 315087 661598 455031
rect 663766 429189 663818 429195
rect 663766 429131 663818 429137
rect 661558 315081 661610 315087
rect 661558 315023 661610 315029
rect 663778 269799 663806 429131
rect 663874 405515 663902 537467
rect 663970 536643 663998 627821
rect 665206 627805 665258 627811
rect 665206 627747 665258 627753
rect 665218 623593 665246 627747
rect 666658 627737 666686 748885
rect 666754 717055 666782 840941
rect 666838 783723 666890 783729
rect 666838 783665 666890 783671
rect 666850 731263 666878 783665
rect 666838 731257 666890 731263
rect 666838 731199 666890 731205
rect 666742 717049 666794 717055
rect 666742 716991 666794 716997
rect 666742 682639 666794 682645
rect 666742 682581 666794 682587
rect 666646 627731 666698 627737
rect 666646 627673 666698 627679
rect 665206 623587 665258 623593
rect 665206 623529 665258 623535
rect 665878 581777 665930 581783
rect 665878 581719 665930 581725
rect 665890 578453 665918 581719
rect 666754 581635 666782 682581
rect 667990 669615 668042 669621
rect 667990 669557 668042 669563
rect 668002 625115 668030 669557
rect 668086 640459 668138 640465
rect 668086 640401 668138 640407
rect 668098 627811 668126 640401
rect 668086 627805 668138 627811
rect 668086 627747 668138 627753
rect 667988 625106 668044 625115
rect 667988 625041 668044 625050
rect 666836 624218 666892 624227
rect 666836 624153 666892 624162
rect 666850 607979 666878 624153
rect 666838 607973 666890 607979
rect 666838 607915 666890 607921
rect 666838 590435 666890 590441
rect 666838 590377 666890 590383
rect 666742 581629 666794 581635
rect 666742 581571 666794 581577
rect 665878 578447 665930 578453
rect 665878 578389 665930 578395
rect 666646 550179 666698 550185
rect 666646 550121 666698 550127
rect 663958 536637 664010 536643
rect 663958 536579 664010 536585
rect 663958 524279 664010 524285
rect 663958 524221 664010 524227
rect 663862 405509 663914 405515
rect 663862 405451 663914 405457
rect 663970 404257 663998 524221
rect 666658 404775 666686 550121
rect 666850 493723 666878 590377
rect 668086 586069 668138 586075
rect 668086 586011 668138 586017
rect 668098 581857 668126 586011
rect 668086 581851 668138 581857
rect 668086 581793 668138 581799
rect 666838 493717 666890 493723
rect 666838 493659 666890 493665
rect 666742 469519 666794 469525
rect 666742 469461 666794 469467
rect 666646 404769 666698 404775
rect 666646 404711 666698 404717
rect 663958 404251 664010 404257
rect 663958 404193 664010 404199
rect 666646 401291 666698 401297
rect 666646 401233 666698 401239
rect 666658 378727 666686 401233
rect 666646 378721 666698 378727
rect 666646 378663 666698 378669
rect 663862 364883 663914 364889
rect 663862 364825 663914 364831
rect 663766 269793 663818 269799
rect 663766 269735 663818 269741
rect 663874 223845 663902 364825
rect 666646 351415 666698 351421
rect 666646 351357 666698 351363
rect 663862 223839 663914 223845
rect 663862 223781 663914 223787
rect 666658 179371 666686 351357
rect 666754 314791 666782 469461
rect 666838 403289 666890 403295
rect 666838 403231 666890 403237
rect 666742 314785 666794 314791
rect 666742 314727 666794 314733
rect 666850 269207 666878 403231
rect 666838 269201 666890 269207
rect 666838 269143 666890 269149
rect 666646 179365 666698 179371
rect 666646 179307 666698 179313
rect 661462 178847 661514 178853
rect 661462 178789 661514 178795
rect 661270 155907 661322 155913
rect 661270 155849 661322 155855
rect 658678 149395 658730 149401
rect 658678 149337 658730 149343
rect 655414 132819 655466 132825
rect 655414 132761 655466 132767
rect 655126 132671 655178 132677
rect 655126 132613 655178 132619
rect 650998 129859 651050 129865
rect 650998 129801 651050 129807
rect 651010 129717 651038 129801
rect 650998 129711 651050 129717
rect 650998 129653 651050 129659
rect 647926 129637 647978 129643
rect 647926 129579 647978 129585
rect 650902 129637 650954 129643
rect 650902 129579 650954 129585
rect 647938 123839 647966 129579
rect 647924 123830 647980 123839
rect 647924 123765 647980 123774
rect 647926 121201 647978 121207
rect 647926 121143 647978 121149
rect 647830 121127 647882 121133
rect 647830 121069 647882 121075
rect 647938 119547 647966 121143
rect 647924 119538 647980 119547
rect 647924 119473 647980 119482
rect 646676 117614 646732 117623
rect 646676 117549 646732 117558
rect 184628 116282 184684 116291
rect 184628 116217 184684 116226
rect 647924 115690 647980 115699
rect 647924 115625 647980 115634
rect 184532 115394 184588 115403
rect 184532 115329 184588 115338
rect 647938 115287 647966 115625
rect 647926 115281 647978 115287
rect 647926 115223 647978 115229
rect 665206 115281 665258 115287
rect 665206 115223 665258 115229
rect 184534 115207 184586 115213
rect 184534 115149 184586 115155
rect 665218 115158 665246 115223
rect 184438 115059 184490 115065
rect 184438 115001 184490 115007
rect 151510 114985 151562 114991
rect 151510 114927 151562 114933
rect 184342 114985 184394 114991
rect 184342 114927 184394 114933
rect 184354 114811 184382 114927
rect 184340 114802 184396 114811
rect 184340 114737 184396 114746
rect 184450 113923 184478 115001
rect 184436 113914 184492 113923
rect 184436 113849 184492 113858
rect 184546 113183 184574 115149
rect 184630 115133 184682 115139
rect 665218 115130 665342 115158
rect 184630 115075 184682 115081
rect 184532 113174 184588 113183
rect 184532 113109 184588 113118
rect 184642 112443 184670 115075
rect 646580 113174 646636 113183
rect 646580 113109 646636 113118
rect 184628 112434 184684 112443
rect 184628 112369 184684 112378
rect 184438 112321 184490 112327
rect 184438 112263 184490 112269
rect 184342 112173 184394 112179
rect 184342 112115 184394 112121
rect 184354 110963 184382 112115
rect 184450 111703 184478 112263
rect 184534 112247 184586 112253
rect 184534 112189 184586 112195
rect 184436 111694 184492 111703
rect 184436 111629 184492 111638
rect 184340 110954 184396 110963
rect 184340 110889 184396 110898
rect 184546 110223 184574 112189
rect 184532 110214 184588 110223
rect 184532 110149 184588 110158
rect 184534 109435 184586 109441
rect 184534 109377 184586 109383
rect 184438 109361 184490 109367
rect 184438 109303 184490 109309
rect 184342 109287 184394 109293
rect 184342 109229 184394 109235
rect 184354 107855 184382 109229
rect 184450 108743 184478 109303
rect 184436 108734 184492 108743
rect 184436 108669 184492 108678
rect 184340 107846 184396 107855
rect 184340 107781 184396 107790
rect 184546 107115 184574 109377
rect 184532 107106 184588 107115
rect 184532 107041 184588 107050
rect 184630 106549 184682 106555
rect 184630 106491 184682 106497
rect 184438 106475 184490 106481
rect 184438 106417 184490 106423
rect 184450 106375 184478 106417
rect 184534 106401 184586 106407
rect 184436 106366 184492 106375
rect 184342 106327 184394 106333
rect 184534 106343 184586 106349
rect 184436 106301 184492 106310
rect 184342 106269 184394 106275
rect 184354 105635 184382 106269
rect 184340 105626 184396 105635
rect 184340 105561 184396 105570
rect 184546 104895 184574 106343
rect 184532 104886 184588 104895
rect 184532 104821 184588 104830
rect 184642 104007 184670 106491
rect 645908 106070 645964 106079
rect 645908 106005 645964 106014
rect 184628 103998 184684 104007
rect 184628 103933 184684 103942
rect 645922 103743 645950 106005
rect 645910 103737 645962 103743
rect 645910 103679 645962 103685
rect 184534 103663 184586 103669
rect 184534 103605 184586 103611
rect 184438 103515 184490 103521
rect 184438 103457 184490 103463
rect 184342 103441 184394 103447
rect 184340 103406 184342 103415
rect 184394 103406 184396 103415
rect 184340 103341 184396 103350
rect 184450 101935 184478 103457
rect 184546 102527 184574 103605
rect 184630 103589 184682 103595
rect 184630 103531 184682 103537
rect 184532 102518 184588 102527
rect 184532 102453 184588 102462
rect 184436 101926 184492 101935
rect 184436 101861 184492 101870
rect 184642 101047 184670 103531
rect 645140 102222 645196 102231
rect 645140 102157 645196 102166
rect 645154 102115 645182 102157
rect 645142 102109 645194 102115
rect 645142 102051 645194 102057
rect 184628 101038 184684 101047
rect 149698 100996 149822 101024
rect 149684 100890 149740 100899
rect 149684 100825 149740 100834
rect 149590 94783 149642 94789
rect 149590 94725 149642 94731
rect 149698 83393 149726 100825
rect 149794 100561 149822 100996
rect 184628 100973 184684 100982
rect 184438 100777 184490 100783
rect 184438 100719 184490 100725
rect 149782 100555 149834 100561
rect 149782 100497 149834 100503
rect 184342 100555 184394 100561
rect 184342 100497 184394 100503
rect 184354 100307 184382 100497
rect 184340 100298 184396 100307
rect 184340 100233 184396 100242
rect 184450 99567 184478 100719
rect 184534 100703 184586 100709
rect 184534 100645 184586 100651
rect 184436 99558 184492 99567
rect 184436 99493 184492 99502
rect 184546 98679 184574 100645
rect 184630 100629 184682 100635
rect 184630 100571 184682 100577
rect 184532 98670 184588 98679
rect 184532 98605 184588 98614
rect 184642 98087 184670 100571
rect 184628 98078 184684 98087
rect 184628 98013 184684 98022
rect 184534 97891 184586 97897
rect 184534 97833 184586 97839
rect 184342 97817 184394 97823
rect 184342 97759 184394 97765
rect 184354 97199 184382 97759
rect 184438 97743 184490 97749
rect 184438 97685 184490 97691
rect 184340 97190 184396 97199
rect 184340 97125 184396 97134
rect 184450 96459 184478 97685
rect 184436 96450 184492 96459
rect 184436 96385 184492 96394
rect 184546 95719 184574 97833
rect 645428 96006 645484 96015
rect 645428 95941 645430 95950
rect 645482 95941 645484 95950
rect 645430 95909 645482 95915
rect 184532 95710 184588 95719
rect 184532 95645 184588 95654
rect 184534 95005 184586 95011
rect 184340 94970 184396 94979
rect 184534 94947 184586 94953
rect 184340 94905 184342 94914
rect 184394 94905 184396 94914
rect 184342 94873 184394 94879
rect 184438 94857 184490 94863
rect 184438 94799 184490 94805
rect 184342 94783 184394 94789
rect 184342 94725 184394 94731
rect 184354 92759 184382 94725
rect 184450 93499 184478 94799
rect 184546 94239 184574 94947
rect 184532 94230 184588 94239
rect 184532 94165 184588 94174
rect 184436 93490 184492 93499
rect 184436 93425 184492 93434
rect 184340 92750 184396 92759
rect 184340 92685 184396 92694
rect 646486 92415 646538 92421
rect 646486 92357 646538 92363
rect 645526 92341 645578 92347
rect 645526 92283 645578 92289
rect 184534 92119 184586 92125
rect 184534 92061 184586 92067
rect 184438 91971 184490 91977
rect 184438 91913 184490 91919
rect 184342 91897 184394 91903
rect 184340 91862 184342 91871
rect 184394 91862 184396 91871
rect 184340 91797 184396 91806
rect 184450 91131 184478 91913
rect 184436 91122 184492 91131
rect 184436 91057 184492 91066
rect 184546 90391 184574 92061
rect 184630 92045 184682 92051
rect 184630 91987 184682 91993
rect 184532 90382 184588 90391
rect 184532 90317 184588 90326
rect 184642 89651 184670 91987
rect 184628 89642 184684 89651
rect 184628 89577 184684 89586
rect 184630 89233 184682 89239
rect 184630 89175 184682 89181
rect 184534 89159 184586 89165
rect 184534 89101 184586 89107
rect 184342 89085 184394 89091
rect 184342 89027 184394 89033
rect 184354 88911 184382 89027
rect 184438 89011 184490 89017
rect 184438 88953 184490 88959
rect 184340 88902 184396 88911
rect 184340 88837 184396 88846
rect 184450 87283 184478 88953
rect 184546 88171 184574 89101
rect 184532 88162 184588 88171
rect 184532 88097 184588 88106
rect 184436 87274 184492 87283
rect 184436 87209 184492 87218
rect 184642 86691 184670 89175
rect 184628 86682 184684 86691
rect 184628 86617 184684 86626
rect 184342 86421 184394 86427
rect 184342 86363 184394 86369
rect 184354 85803 184382 86363
rect 184438 86347 184490 86353
rect 184438 86289 184490 86295
rect 184340 85794 184396 85803
rect 184340 85729 184396 85738
rect 184450 85211 184478 86289
rect 184534 86273 184586 86279
rect 184534 86215 184586 86221
rect 184436 85202 184492 85211
rect 184436 85137 184492 85146
rect 184546 84323 184574 86215
rect 184532 84314 184588 84323
rect 184532 84249 184588 84258
rect 640726 83683 640778 83689
rect 640726 83625 640778 83631
rect 184534 83535 184586 83541
rect 184534 83477 184586 83483
rect 184340 83426 184396 83435
rect 149686 83387 149738 83393
rect 184340 83361 184342 83370
rect 149686 83329 149738 83335
rect 184394 83361 184396 83370
rect 184342 83329 184394 83335
rect 184438 83313 184490 83319
rect 184438 83255 184490 83261
rect 149588 82390 149644 82399
rect 149588 82325 149644 82334
rect 149494 80575 149546 80581
rect 149494 80517 149546 80523
rect 149398 77615 149450 77621
rect 149398 77557 149450 77563
rect 149302 77541 149354 77547
rect 149302 77483 149354 77489
rect 149108 76766 149164 76775
rect 149108 76701 149164 76710
rect 148822 74877 148874 74883
rect 148822 74819 148874 74825
rect 149012 73066 149068 73075
rect 149012 73001 149068 73010
rect 148726 71917 148778 71923
rect 148726 71859 148778 71865
rect 148630 69105 148682 69111
rect 148630 69047 148682 69053
rect 149026 66077 149054 73001
rect 149122 68963 149150 76701
rect 149396 75582 149452 75591
rect 149396 75517 149452 75526
rect 149410 74894 149438 75517
rect 149410 74866 149534 74894
rect 149204 72030 149260 72039
rect 149204 71965 149260 71974
rect 149110 68957 149162 68963
rect 149110 68899 149162 68905
rect 149218 66151 149246 71965
rect 149396 70846 149452 70855
rect 149396 70781 149452 70790
rect 149300 69514 149356 69523
rect 149300 69449 149356 69458
rect 149206 66145 149258 66151
rect 149206 66087 149258 66093
rect 149014 66071 149066 66077
rect 149014 66013 149066 66019
rect 149314 66003 149342 69449
rect 149410 66225 149438 70781
rect 149506 69037 149534 74866
rect 149602 74661 149630 82325
rect 184450 81955 184478 83255
rect 184546 82843 184574 83477
rect 184630 83461 184682 83467
rect 184630 83403 184682 83409
rect 184532 82834 184588 82843
rect 184532 82769 184588 82778
rect 184436 81946 184492 81955
rect 184436 81881 184492 81890
rect 184642 81363 184670 83403
rect 184628 81354 184684 81363
rect 184628 81289 184684 81298
rect 184630 80649 184682 80655
rect 184630 80591 184682 80597
rect 184342 80575 184394 80581
rect 184342 80517 184394 80523
rect 184354 80475 184382 80517
rect 184438 80501 184490 80507
rect 184340 80466 184396 80475
rect 184438 80443 184490 80449
rect 184340 80401 184396 80410
rect 184450 79883 184478 80443
rect 184534 80427 184586 80433
rect 184534 80369 184586 80375
rect 184436 79874 184492 79883
rect 184436 79809 184492 79818
rect 149684 79282 149740 79291
rect 149684 79217 149740 79226
rect 149590 74655 149642 74661
rect 149590 74597 149642 74603
rect 149588 73806 149644 73815
rect 149588 73741 149644 73750
rect 149494 69031 149546 69037
rect 149494 68973 149546 68979
rect 149602 68889 149630 73741
rect 149698 71849 149726 79217
rect 184546 78255 184574 80369
rect 184642 78995 184670 80591
rect 184628 78986 184684 78995
rect 184628 78921 184684 78930
rect 184532 78246 184588 78255
rect 184532 78181 184588 78190
rect 184438 77763 184490 77769
rect 184438 77705 184490 77711
rect 184342 77541 184394 77547
rect 184450 77515 184478 77705
rect 184534 77689 184586 77695
rect 184534 77631 184586 77637
rect 184342 77483 184394 77489
rect 184436 77506 184492 77515
rect 184354 76035 184382 77483
rect 184436 77441 184492 77450
rect 184546 76775 184574 77631
rect 184630 77615 184682 77621
rect 184630 77557 184682 77563
rect 184532 76766 184588 76775
rect 184532 76701 184588 76710
rect 184340 76026 184396 76035
rect 184340 75961 184396 75970
rect 184642 75147 184670 77557
rect 184628 75138 184684 75147
rect 184628 75073 184684 75082
rect 184342 74877 184394 74883
rect 184342 74819 184394 74825
rect 184354 74407 184382 74819
rect 184438 74803 184490 74809
rect 184438 74745 184490 74751
rect 184340 74398 184396 74407
rect 184340 74333 184396 74342
rect 184450 73667 184478 74745
rect 184534 74729 184586 74735
rect 184534 74671 184586 74677
rect 184436 73658 184492 73667
rect 184436 73593 184492 73602
rect 184546 72927 184574 74671
rect 184630 74655 184682 74661
rect 184630 74597 184682 74603
rect 184532 72918 184588 72927
rect 184532 72853 184588 72862
rect 184642 72187 184670 74597
rect 184628 72178 184684 72187
rect 184628 72113 184684 72122
rect 184342 71991 184394 71997
rect 184342 71933 184394 71939
rect 149686 71843 149738 71849
rect 149686 71785 149738 71791
rect 184354 71447 184382 71933
rect 184438 71917 184490 71923
rect 184438 71859 184490 71865
rect 184340 71438 184396 71447
rect 184340 71373 184396 71382
rect 184450 70559 184478 71859
rect 184534 71843 184586 71849
rect 184534 71785 184586 71791
rect 184436 70550 184492 70559
rect 184436 70485 184492 70494
rect 184546 69967 184574 71785
rect 184532 69958 184588 69967
rect 184532 69893 184588 69902
rect 184342 69105 184394 69111
rect 184340 69070 184342 69079
rect 184394 69070 184396 69079
rect 184340 69005 184396 69014
rect 184534 69031 184586 69037
rect 184534 68973 184586 68979
rect 184342 68957 184394 68963
rect 184342 68899 184394 68905
rect 149590 68883 149642 68889
rect 149590 68825 149642 68831
rect 184354 68487 184382 68899
rect 184438 68883 184490 68889
rect 184438 68825 184490 68831
rect 184340 68478 184396 68487
rect 184340 68413 184396 68422
rect 149588 68330 149644 68339
rect 149588 68265 149644 68274
rect 149492 67146 149548 67155
rect 149492 67081 149548 67090
rect 149398 66219 149450 66225
rect 149398 66161 149450 66167
rect 149302 65997 149354 66003
rect 149302 65939 149354 65945
rect 149396 64630 149452 64639
rect 149396 64565 149452 64574
rect 149300 63446 149356 63455
rect 149300 63381 149356 63390
rect 149314 60305 149342 63381
rect 149410 63117 149438 64565
rect 149506 63265 149534 67081
rect 149494 63259 149546 63265
rect 149494 63201 149546 63207
rect 149602 63191 149630 68265
rect 184450 66859 184478 68825
rect 184546 67599 184574 68973
rect 184532 67590 184588 67599
rect 184532 67525 184588 67534
rect 184436 66850 184492 66859
rect 184436 66785 184492 66794
rect 184630 66219 184682 66225
rect 184630 66161 184682 66167
rect 184534 66145 184586 66151
rect 184340 66110 184396 66119
rect 184534 66087 184586 66093
rect 184340 66045 184342 66054
rect 184394 66045 184396 66054
rect 184342 66013 184394 66019
rect 184438 65997 184490 66003
rect 184438 65939 184490 65945
rect 149684 65370 149740 65379
rect 149684 65305 149740 65314
rect 149698 63339 149726 65305
rect 184450 63751 184478 65939
rect 184546 65231 184574 66087
rect 184532 65222 184588 65231
rect 184532 65157 184588 65166
rect 184642 64639 184670 66161
rect 184628 64630 184684 64639
rect 184628 64565 184684 64574
rect 184436 63742 184492 63751
rect 184436 63677 184492 63686
rect 149686 63333 149738 63339
rect 149686 63275 149738 63281
rect 184630 63333 184682 63339
rect 184630 63275 184682 63281
rect 184438 63259 184490 63265
rect 184438 63201 184490 63207
rect 149590 63185 149642 63191
rect 184342 63185 184394 63191
rect 149590 63127 149642 63133
rect 184340 63150 184342 63159
rect 184394 63150 184396 63159
rect 149398 63111 149450 63117
rect 184340 63085 184396 63094
rect 149398 63053 149450 63059
rect 184450 62271 184478 63201
rect 184534 63111 184586 63117
rect 184534 63053 184586 63059
rect 149396 62262 149452 62271
rect 149396 62197 149452 62206
rect 184436 62262 184492 62271
rect 184436 62197 184492 62206
rect 149410 60453 149438 62197
rect 184546 60791 184574 63053
rect 184642 61531 184670 63275
rect 184628 61522 184684 61531
rect 184628 61457 184684 61466
rect 184532 60782 184588 60791
rect 184532 60717 184588 60726
rect 149492 60634 149548 60643
rect 149492 60569 149548 60578
rect 149398 60447 149450 60453
rect 149398 60389 149450 60395
rect 149506 60379 149534 60569
rect 184438 60447 184490 60453
rect 184438 60389 184490 60395
rect 149494 60373 149546 60379
rect 149494 60315 149546 60321
rect 149302 60299 149354 60305
rect 149302 60241 149354 60247
rect 184342 60299 184394 60305
rect 184342 60241 184394 60247
rect 184354 60051 184382 60241
rect 184340 60042 184396 60051
rect 184340 59977 184396 59986
rect 149396 59746 149452 59755
rect 149396 59681 149452 59690
rect 149410 59047 149438 59681
rect 184450 59311 184478 60389
rect 184534 60373 184586 60379
rect 184534 60315 184586 60321
rect 184436 59302 184492 59311
rect 184436 59237 184492 59246
rect 149398 59041 149450 59047
rect 149398 58983 149450 58989
rect 184342 59041 184394 59047
rect 184342 58983 184394 58989
rect 149396 58562 149452 58571
rect 149396 58497 149452 58506
rect 149410 57567 149438 58497
rect 184354 57683 184382 58983
rect 184546 58423 184574 60315
rect 184532 58414 184588 58423
rect 184532 58349 184588 58358
rect 184340 57674 184396 57683
rect 184340 57609 184396 57618
rect 149398 57561 149450 57567
rect 149398 57503 149450 57509
rect 184342 57561 184394 57567
rect 184342 57503 184394 57509
rect 149492 57378 149548 57387
rect 149492 57313 149548 57322
rect 149398 56229 149450 56235
rect 149396 56194 149398 56203
rect 149450 56194 149452 56203
rect 149506 56161 149534 57313
rect 184354 56943 184382 57503
rect 184340 56934 184396 56943
rect 184340 56869 184396 56878
rect 184438 56229 184490 56235
rect 184340 56194 184396 56203
rect 149396 56129 149452 56138
rect 149494 56155 149546 56161
rect 184438 56171 184490 56177
rect 184340 56129 184342 56138
rect 149494 56097 149546 56103
rect 184394 56129 184396 56138
rect 184342 56097 184394 56103
rect 184450 55463 184478 56171
rect 184436 55454 184492 55463
rect 184436 55389 184492 55398
rect 149684 54862 149740 54871
rect 149684 54797 149740 54806
rect 149698 54681 149726 54797
rect 184340 54714 184396 54723
rect 149686 54675 149738 54681
rect 184340 54649 184342 54658
rect 149686 54617 149738 54623
rect 184394 54649 184396 54658
rect 184342 54617 184394 54623
rect 184340 53974 184396 53983
rect 184340 53909 184396 53918
rect 149396 53826 149452 53835
rect 149396 53761 149452 53770
rect 149410 53275 149438 53761
rect 184354 53275 184382 53909
rect 149398 53269 149450 53275
rect 149398 53211 149450 53217
rect 184342 53269 184394 53275
rect 184342 53211 184394 53217
rect 145104 49788 145406 49816
rect 145378 47133 145406 49788
rect 199138 47133 199166 53650
rect 145366 47127 145418 47133
rect 145366 47069 145418 47075
rect 199126 47127 199178 47133
rect 199126 47069 199178 47075
rect 142306 46680 142416 46708
rect 142306 40219 142334 46680
rect 187604 41838 187660 41847
rect 187344 41796 187604 41824
rect 194324 41838 194380 41847
rect 194064 41796 194324 41824
rect 187604 41773 187660 41782
rect 194324 41773 194380 41782
rect 216418 40413 216446 53650
rect 233698 47651 233726 53650
rect 233686 47645 233738 47651
rect 233686 47587 233738 47593
rect 250978 47577 251006 53650
rect 268320 53636 268574 53664
rect 285600 53636 285854 53664
rect 268546 47725 268574 53636
rect 285826 47873 285854 53636
rect 285814 47867 285866 47873
rect 285814 47809 285866 47815
rect 302914 47799 302942 53650
rect 311062 48015 311114 48021
rect 311062 47957 311114 47963
rect 302902 47793 302954 47799
rect 302902 47735 302954 47741
rect 268534 47719 268586 47725
rect 268534 47661 268586 47667
rect 250966 47571 251018 47577
rect 250966 47513 251018 47519
rect 311074 42268 311102 47957
rect 320194 47947 320222 53650
rect 331222 48089 331274 48095
rect 331222 48031 331274 48037
rect 320182 47941 320234 47947
rect 320182 47883 320234 47889
rect 310498 42240 311102 42268
rect 310498 42120 310526 42240
rect 310128 42092 310526 42120
rect 302900 41838 302956 41847
rect 302688 41796 302900 41824
rect 307220 41838 307276 41847
rect 307008 41796 307220 41824
rect 302900 41773 302956 41782
rect 307220 41773 307276 41782
rect 331234 40811 331262 48031
rect 337474 40963 337502 53650
rect 354850 48095 354878 53650
rect 371938 53636 372192 53664
rect 389218 53636 389472 53664
rect 354838 48089 354890 48095
rect 354838 48031 354890 48037
rect 362038 48089 362090 48095
rect 362038 48031 362090 48037
rect 357716 42134 357772 42143
rect 357456 42092 357716 42120
rect 362050 42120 362078 48031
rect 371938 48021 371966 53636
rect 389218 48095 389246 53636
rect 389206 48089 389258 48095
rect 389206 48031 389258 48037
rect 371926 48015 371978 48021
rect 371926 47957 371978 47963
rect 405526 48015 405578 48021
rect 405526 47957 405578 47963
rect 398902 42391 398954 42397
rect 398902 42333 398954 42339
rect 365314 42240 365726 42268
rect 365314 42120 365342 42240
rect 361776 42092 362078 42120
rect 364944 42092 365342 42120
rect 357716 42069 357772 42078
rect 365698 41824 365726 42240
rect 365698 41796 365918 41824
rect 337460 40954 337516 40963
rect 337460 40889 337516 40898
rect 331220 40802 331276 40811
rect 331220 40737 331276 40746
rect 216404 40404 216460 40413
rect 216404 40339 216460 40348
rect 142292 40210 142348 40219
rect 142292 40145 142348 40154
rect 365890 38356 365918 41796
rect 365890 38328 365948 38356
rect 365920 37439 365948 38328
rect 398914 37439 398942 42333
rect 405538 42106 405566 47957
rect 406786 47471 406814 53650
rect 424066 48095 424094 53650
rect 411862 48089 411914 48095
rect 411862 48031 411914 48037
rect 424054 48089 424106 48095
rect 424054 48031 424106 48037
rect 434902 48089 434954 48095
rect 434902 48031 434954 48037
rect 406772 47462 406828 47471
rect 406772 47397 406828 47406
rect 411874 42397 411902 48031
rect 419732 47610 419788 47619
rect 419732 47545 419788 47554
rect 419746 44608 419774 47545
rect 411862 42391 411914 42397
rect 411862 42333 411914 42339
rect 434914 41995 434942 48031
rect 441346 48021 441374 53650
rect 441334 48015 441386 48021
rect 441334 47957 441386 47963
rect 458626 46985 458654 53650
rect 475714 53636 475968 53664
rect 492994 53636 493248 53664
rect 510370 53636 510624 53664
rect 475714 48095 475742 53636
rect 475702 48089 475754 48095
rect 475702 48031 475754 48037
rect 460342 48015 460394 48021
rect 460342 47957 460394 47963
rect 455062 46979 455114 46985
rect 455062 46921 455114 46927
rect 458614 46979 458666 46985
rect 458614 46921 458666 46927
rect 415508 41986 415564 41995
rect 415440 41944 415508 41972
rect 415508 41921 415564 41930
rect 434900 41986 434956 41995
rect 434900 41921 434956 41930
rect 416852 41838 416908 41847
rect 416592 41796 416852 41824
rect 416852 41773 416908 41782
rect 420692 40654 420748 40663
rect 420692 40589 420748 40598
rect 420706 37439 420734 40589
rect 455074 37439 455102 46921
rect 460354 42106 460382 47957
rect 475606 47645 475658 47651
rect 492994 47619 493022 53636
rect 510370 48021 510398 53636
rect 510358 48015 510410 48021
rect 510358 47957 510410 47963
rect 515542 47941 515594 47947
rect 515542 47883 515594 47889
rect 493942 47867 493994 47873
rect 493942 47809 493994 47815
rect 475606 47587 475658 47593
rect 492980 47610 493036 47619
rect 474452 47462 474508 47471
rect 474452 47397 474508 47406
rect 474466 44312 474494 47397
rect 470324 41838 470380 41847
rect 470160 41796 470324 41824
rect 471408 41805 471710 41824
rect 471408 41799 471722 41805
rect 471408 41796 471670 41799
rect 470324 41773 470380 41782
rect 471670 41741 471722 41747
rect 475510 41799 475562 41805
rect 475510 41741 475562 41747
rect 475522 37439 475550 41741
rect 365908 37433 365960 37439
rect 365908 37375 365960 37381
rect 398902 37433 398954 37439
rect 398902 37375 398954 37381
rect 420694 37433 420746 37439
rect 420694 37375 420746 37381
rect 455062 37433 455114 37439
rect 455062 37375 455114 37381
rect 475510 37433 475562 37439
rect 475510 37375 475562 37381
rect 475618 37365 475646 47587
rect 492980 47545 493036 47554
rect 493954 40811 493982 47809
rect 503926 47719 503978 47725
rect 503926 47661 503978 47667
rect 493940 40802 493996 40811
rect 493940 40737 493996 40746
rect 503938 40325 503966 47661
rect 515554 45135 515582 47883
rect 525910 47793 525962 47799
rect 525910 47735 525962 47741
rect 521206 47571 521258 47577
rect 521206 47513 521258 47519
rect 515542 45129 515594 45135
rect 515542 45071 515594 45077
rect 509782 43205 509834 43211
rect 509782 43147 509834 43153
rect 521218 43156 521246 47513
rect 521494 46387 521546 46393
rect 521494 46329 521546 46335
rect 521506 43285 521534 46329
rect 521494 43279 521546 43285
rect 521494 43221 521546 43227
rect 503926 40319 503978 40325
rect 503926 40261 503978 40267
rect 506806 40319 506858 40325
rect 506806 40261 506858 40267
rect 506818 40219 506846 40261
rect 506804 40210 506860 40219
rect 506804 40145 506860 40154
rect 509794 37439 509822 43147
rect 521218 43128 521534 43156
rect 521506 42120 521534 43128
rect 525922 42120 525950 47735
rect 527938 46393 527966 53650
rect 527926 46387 527978 46393
rect 527926 46329 527978 46335
rect 529270 45129 529322 45135
rect 529270 45071 529322 45077
rect 521506 42092 521856 42120
rect 525922 42092 526176 42120
rect 529282 42106 529310 45071
rect 518708 41838 518764 41847
rect 514882 41805 515136 41824
rect 514006 41799 514058 41805
rect 514006 41741 514058 41747
rect 514870 41799 515136 41805
rect 514922 41796 515136 41799
rect 520340 41838 520396 41847
rect 518764 41796 518832 41824
rect 518708 41773 518764 41782
rect 520396 41796 520656 41824
rect 520340 41773 520396 41782
rect 514870 41741 514922 41747
rect 509782 37433 509834 37439
rect 509782 37375 509834 37381
rect 514018 37365 514046 41741
rect 545218 40663 545246 53650
rect 562498 47471 562526 53650
rect 579796 53602 579852 54402
rect 597092 53602 597148 54402
rect 614388 53602 614444 54402
rect 631684 53602 631740 54402
rect 562484 47462 562540 47471
rect 562484 47397 562540 47406
rect 640738 43285 640766 83625
rect 645538 79439 645566 92283
rect 645908 88902 645964 88911
rect 645908 88837 645964 88846
rect 645922 87537 645950 88837
rect 645910 87531 645962 87537
rect 645910 87473 645962 87479
rect 645908 84462 645964 84471
rect 645908 84397 645964 84406
rect 645922 84207 645950 84397
rect 645910 84201 645962 84207
rect 645910 84143 645962 84149
rect 645524 79430 645580 79439
rect 645524 79365 645580 79374
rect 646006 76135 646058 76141
rect 646006 76077 646058 76083
rect 646018 75591 646046 76077
rect 646004 75582 646060 75591
rect 646004 75517 646060 75526
rect 646004 66258 646060 66267
rect 646004 66193 646006 66202
rect 646058 66193 646060 66202
rect 646006 66161 646058 66167
rect 646006 59115 646058 59121
rect 646006 59057 646058 59063
rect 646018 59015 646046 59057
rect 646004 59006 646060 59015
rect 646004 58941 646060 58950
rect 646498 54723 646526 92357
rect 646594 77695 646622 113109
rect 647060 111398 647116 111407
rect 647060 111333 647116 111342
rect 646676 109474 646732 109483
rect 646676 109409 646732 109418
rect 646582 77689 646634 77695
rect 646582 77631 646634 77637
rect 646690 77621 646718 109409
rect 646772 107994 646828 108003
rect 646772 107929 646828 107938
rect 646786 92717 646814 107929
rect 646964 98078 647020 98087
rect 646964 98013 647020 98022
rect 646774 92711 646826 92717
rect 646774 92653 646826 92659
rect 646870 92267 646922 92273
rect 646870 92209 646922 92215
rect 646774 83609 646826 83615
rect 646774 83551 646826 83557
rect 646678 77615 646730 77621
rect 646678 77557 646730 77563
rect 646786 57091 646814 83551
rect 646882 68635 646910 92209
rect 646978 77769 647006 98013
rect 647074 87093 647102 111333
rect 665314 105191 665342 115130
rect 669538 106375 669566 866915
rect 669634 356199 669662 986425
rect 669814 986409 669866 986415
rect 669814 986351 669866 986357
rect 669718 985077 669770 985083
rect 669718 985019 669770 985025
rect 669730 937797 669758 985019
rect 669718 937791 669770 937797
rect 669718 937733 669770 937739
rect 669718 757601 669770 757607
rect 669718 757543 669770 757549
rect 669620 356190 669676 356199
rect 669620 356125 669676 356134
rect 669730 278203 669758 757543
rect 669826 357087 669854 986351
rect 669910 985003 669962 985009
rect 669910 984945 669962 984951
rect 669922 938907 669950 984945
rect 675394 966255 675422 966736
rect 675380 966246 675436 966255
rect 675380 966181 675436 966190
rect 675490 965811 675518 966070
rect 675476 965802 675532 965811
rect 675476 965737 675532 965746
rect 675490 965071 675518 965435
rect 675476 965062 675532 965071
rect 675476 964997 675532 965006
rect 675394 963443 675422 963595
rect 675380 963434 675436 963443
rect 675380 963369 675436 963378
rect 675490 962703 675518 963036
rect 675476 962694 675532 962703
rect 675476 962629 675532 962638
rect 675778 962259 675806 962399
rect 675764 962250 675820 962259
rect 675764 962185 675820 962194
rect 675394 961329 675422 961778
rect 674710 961323 674762 961329
rect 674710 961265 674762 961271
rect 675382 961323 675434 961329
rect 675382 961265 675434 961271
rect 674722 953379 674750 961265
rect 674806 959177 674858 959183
rect 675490 959151 675518 959262
rect 674806 959119 674858 959125
rect 675476 959142 675532 959151
rect 674818 955483 674846 959119
rect 675476 959077 675532 959086
rect 675778 958411 675806 958744
rect 675764 958402 675820 958411
rect 675764 958337 675820 958346
rect 675394 957671 675422 958078
rect 675380 957662 675436 957671
rect 675380 957597 675436 957606
rect 675778 957079 675806 957412
rect 675764 957070 675820 957079
rect 675764 957005 675820 957014
rect 675586 956043 675614 956228
rect 675572 956034 675628 956043
rect 675572 955969 675628 955978
rect 674806 955477 674858 955483
rect 674806 955419 674858 955425
rect 675382 955477 675434 955483
rect 675382 955419 675434 955425
rect 675394 955132 675422 955419
rect 675394 955104 675432 955132
rect 675404 955030 675432 955104
rect 675490 953971 675518 954378
rect 675476 953962 675532 953971
rect 675476 953897 675532 953906
rect 674708 953370 674764 953379
rect 674708 953305 674764 953314
rect 675778 952047 675806 952528
rect 675764 952038 675820 952047
rect 675764 951973 675820 951982
rect 676148 941086 676204 941095
rect 676148 941021 676204 941030
rect 676054 939789 676106 939795
rect 676052 939754 676054 939763
rect 676106 939754 676108 939763
rect 676052 939689 676108 939698
rect 676052 939310 676108 939319
rect 676162 939277 676190 941021
rect 676340 940494 676396 940503
rect 676340 940429 676396 940438
rect 676244 940050 676300 940059
rect 676244 939985 676300 939994
rect 676258 939425 676286 939985
rect 676246 939419 676298 939425
rect 676246 939361 676298 939367
rect 676052 939245 676108 939254
rect 676150 939271 676202 939277
rect 676066 939203 676094 939245
rect 676150 939213 676202 939219
rect 670774 939197 670826 939203
rect 670774 939139 670826 939145
rect 676054 939197 676106 939203
rect 676054 939139 676106 939145
rect 669910 938901 669962 938907
rect 669910 938843 669962 938849
rect 670006 800669 670058 800675
rect 670006 800611 670058 800617
rect 669910 757527 669962 757533
rect 669910 757469 669962 757475
rect 669812 357078 669868 357087
rect 669812 357013 669868 357022
rect 669922 278499 669950 757469
rect 670018 672729 670046 800611
rect 670786 761603 670814 939139
rect 676354 939129 676382 940429
rect 676342 939123 676394 939129
rect 676342 939065 676394 939071
rect 676246 938901 676298 938907
rect 676244 938866 676246 938875
rect 676298 938866 676300 938875
rect 676244 938801 676300 938810
rect 676244 938126 676300 938135
rect 670870 938087 670922 938093
rect 676244 938061 676246 938070
rect 670870 938029 670922 938035
rect 676298 938061 676300 938070
rect 676246 938029 676298 938035
rect 670774 761597 670826 761603
rect 670774 761539 670826 761545
rect 670882 760345 670910 938029
rect 676054 937791 676106 937797
rect 676052 937756 676054 937765
rect 676106 937756 676108 937765
rect 676052 937691 676108 937700
rect 676052 937238 676108 937247
rect 670966 937199 671018 937205
rect 676052 937173 676054 937182
rect 670966 937141 671018 937147
rect 676106 937173 676108 937182
rect 676054 937141 676106 937147
rect 670870 760339 670922 760345
rect 670870 760281 670922 760287
rect 670678 759895 670730 759901
rect 670678 759837 670730 759843
rect 670102 731257 670154 731263
rect 670102 731199 670154 731205
rect 670114 714909 670142 731199
rect 670390 717197 670442 717203
rect 670390 717139 670442 717145
rect 670102 714903 670154 714909
rect 670102 714845 670154 714851
rect 670402 713799 670430 717139
rect 670690 715723 670718 759837
rect 670774 758859 670826 758865
rect 670774 758801 670826 758807
rect 670678 715717 670730 715723
rect 670678 715659 670730 715665
rect 670690 715353 670718 715659
rect 670678 715347 670730 715353
rect 670678 715289 670730 715295
rect 670786 714391 670814 758801
rect 670882 757607 670910 760281
rect 670978 759383 671006 937141
rect 679796 929542 679852 929551
rect 679796 929477 679852 929486
rect 679810 928959 679838 929477
rect 679796 928950 679852 928959
rect 679796 928885 679852 928894
rect 685460 928950 685516 928959
rect 685460 928885 685516 928894
rect 679810 927437 679838 928885
rect 685474 928515 685502 928885
rect 685460 928506 685516 928515
rect 685460 928441 685516 928450
rect 679798 927431 679850 927437
rect 679798 927373 679850 927379
rect 672598 895759 672650 895765
rect 672598 895701 672650 895707
rect 672502 855429 672554 855435
rect 672502 855371 672554 855377
rect 672406 763299 672458 763305
rect 672406 763241 672458 763247
rect 670966 759377 671018 759383
rect 670966 759319 671018 759325
rect 670870 757601 670922 757607
rect 670870 757543 670922 757549
rect 670978 757533 671006 759319
rect 670966 757527 671018 757533
rect 670966 757469 671018 757475
rect 670966 714903 671018 714909
rect 670966 714845 671018 714851
rect 670774 714385 670826 714391
rect 670774 714327 670826 714333
rect 670390 713793 670442 713799
rect 670390 713735 670442 713741
rect 670870 713793 670922 713799
rect 670870 713735 670922 713741
rect 670102 696995 670154 697001
rect 670102 696937 670154 696943
rect 670006 672723 670058 672729
rect 670006 672665 670058 672671
rect 670114 582523 670142 696937
rect 670882 669399 670910 713735
rect 670978 670139 671006 714845
rect 672310 670651 672362 670657
rect 672310 670593 672362 670599
rect 670966 670133 671018 670139
rect 670966 670075 671018 670081
rect 670870 669393 670922 669399
rect 670870 669335 670922 669341
rect 672322 635655 672350 670593
rect 672310 635649 672362 635655
rect 672310 635591 672362 635597
rect 670870 627805 670922 627811
rect 670870 627747 670922 627753
rect 670882 624703 670910 627747
rect 672418 627367 672446 763241
rect 672514 718091 672542 855371
rect 672610 762047 672638 895701
rect 675298 877509 675408 877537
rect 673750 876593 673802 876599
rect 673750 876535 673802 876541
rect 673558 873485 673610 873491
rect 673558 873427 673610 873433
rect 672790 872153 672842 872159
rect 672790 872095 672842 872101
rect 672598 762041 672650 762047
rect 672598 761983 672650 761989
rect 672598 760635 672650 760641
rect 672598 760577 672650 760583
rect 672610 722975 672638 760577
rect 672802 752871 672830 872095
rect 673462 869193 673514 869199
rect 673462 869135 673514 869141
rect 673366 867861 673418 867867
rect 673366 867803 673418 867809
rect 673270 787349 673322 787355
rect 673270 787291 673322 787297
rect 673174 784315 673226 784321
rect 673174 784257 673226 784263
rect 673078 783501 673130 783507
rect 673078 783443 673130 783449
rect 672982 782983 673034 782989
rect 672982 782925 673034 782931
rect 672886 778617 672938 778623
rect 672886 778559 672938 778565
rect 672790 752865 672842 752871
rect 672790 752807 672842 752813
rect 672790 733625 672842 733631
rect 672790 733567 672842 733573
rect 672694 732367 672746 732373
rect 672694 732309 672746 732315
rect 672598 722969 672650 722975
rect 672598 722911 672650 722917
rect 672502 718085 672554 718091
rect 672502 718027 672554 718033
rect 672706 663923 672734 732309
rect 672694 663917 672746 663923
rect 672694 663859 672746 663865
rect 672802 661703 672830 733567
rect 672898 706917 672926 778559
rect 672994 708027 673022 782925
rect 673090 709359 673118 783443
rect 673186 710099 673214 784257
rect 673282 710469 673310 787291
rect 673378 751909 673406 867803
rect 673474 752427 673502 869135
rect 673570 755091 673598 873427
rect 673654 779949 673706 779955
rect 673654 779891 673706 779897
rect 673558 755085 673610 755091
rect 673558 755027 673610 755033
rect 673462 752421 673514 752427
rect 673462 752363 673514 752369
rect 673366 751903 673418 751909
rect 673366 751845 673418 751851
rect 673462 738509 673514 738515
rect 673462 738451 673514 738457
rect 673366 737917 673418 737923
rect 673366 737859 673418 737865
rect 673270 710463 673322 710469
rect 673270 710405 673322 710411
rect 673174 710093 673226 710099
rect 673174 710035 673226 710041
rect 673078 709353 673130 709359
rect 673078 709295 673130 709301
rect 672982 708021 673034 708027
rect 672982 707963 673034 707969
rect 672886 706911 672938 706917
rect 672886 706853 672938 706859
rect 673174 699881 673226 699887
rect 673174 699823 673226 699829
rect 672886 689817 672938 689823
rect 672886 689759 672938 689765
rect 672790 661697 672842 661703
rect 672790 661639 672842 661645
rect 672502 656739 672554 656745
rect 672502 656681 672554 656687
rect 672406 627361 672458 627367
rect 672406 627303 672458 627309
rect 672022 625659 672074 625665
rect 672022 625601 672074 625607
rect 670870 624697 670922 624703
rect 670870 624639 670922 624645
rect 670102 582517 670154 582523
rect 670102 582459 670154 582465
rect 670774 581851 670826 581857
rect 670774 581793 670826 581799
rect 670582 580223 670634 580229
rect 670582 580165 670634 580171
rect 670594 558788 670622 580165
rect 670786 579489 670814 581793
rect 670882 580007 670910 624639
rect 670966 623587 671018 623593
rect 670966 623529 671018 623535
rect 670870 580001 670922 580007
rect 670870 579943 670922 579949
rect 670774 579483 670826 579489
rect 670774 579425 670826 579431
rect 670786 578894 670814 579425
rect 670978 578971 671006 623529
rect 672034 581043 672062 625601
rect 672514 624227 672542 656681
rect 672790 644825 672842 644831
rect 672790 644767 672842 644773
rect 672694 643419 672746 643425
rect 672694 643361 672746 643367
rect 672598 642309 672650 642315
rect 672598 642251 672650 642257
rect 672500 624218 672556 624227
rect 672500 624153 672556 624162
rect 672214 607085 672266 607091
rect 672214 607027 672266 607033
rect 672118 599833 672170 599839
rect 672118 599775 672170 599781
rect 672022 581037 672074 581043
rect 672022 580979 672074 580985
rect 670966 578965 671018 578971
rect 670966 578907 671018 578913
rect 670786 578866 670910 578894
rect 670678 578447 670730 578453
rect 670678 578389 670730 578395
rect 670690 568556 670718 578389
rect 670882 568852 670910 578866
rect 670882 568824 671006 568852
rect 670690 568528 670910 568556
rect 670594 558760 670814 558788
rect 670786 547225 670814 558760
rect 670774 547219 670826 547225
rect 670774 547161 670826 547167
rect 670774 541447 670826 541453
rect 670774 541389 670826 541395
rect 670786 537383 670814 541389
rect 670774 537377 670826 537383
rect 670774 537319 670826 537325
rect 670882 533979 670910 568528
rect 670978 534941 671006 568824
rect 670966 534935 671018 534941
rect 670966 534877 671018 534883
rect 670870 533973 670922 533979
rect 670870 533915 670922 533921
rect 672130 527023 672158 599775
rect 672226 530057 672254 607027
rect 672310 602719 672362 602725
rect 672310 602661 672362 602667
rect 672214 530051 672266 530057
rect 672214 529993 672266 529999
rect 672322 527467 672350 602661
rect 672502 601979 672554 601985
rect 672502 601921 672554 601927
rect 672406 597169 672458 597175
rect 672406 597111 672458 597117
rect 672418 528503 672446 597111
rect 672406 528497 672458 528503
rect 672406 528439 672458 528445
rect 672310 527461 672362 527467
rect 672310 527403 672362 527409
rect 672118 527017 672170 527023
rect 672118 526959 672170 526965
rect 672406 509849 672458 509855
rect 672406 509791 672458 509797
rect 670102 495419 670154 495425
rect 670102 495361 670154 495367
rect 670006 377315 670058 377321
rect 670006 377257 670058 377263
rect 669908 278490 669964 278499
rect 669908 278425 669964 278434
rect 669716 278194 669772 278203
rect 669716 278129 669772 278138
rect 670018 225103 670046 377257
rect 670114 360079 670142 495361
rect 670870 402253 670922 402259
rect 670870 402195 670922 402201
rect 670198 385899 670250 385905
rect 670198 385841 670250 385847
rect 670210 370143 670238 385841
rect 670198 370137 670250 370143
rect 670198 370079 670250 370085
rect 670102 360073 670154 360079
rect 670102 360015 670154 360021
rect 670882 357785 670910 402195
rect 670966 400995 671018 401001
rect 670966 400937 671018 400943
rect 670102 357779 670154 357785
rect 670102 357721 670154 357727
rect 670870 357779 670922 357785
rect 670870 357721 670922 357727
rect 670114 278351 670142 357721
rect 670978 356601 671006 400937
rect 672418 359783 672446 509791
rect 672514 492983 672542 601921
rect 672610 537531 672638 642251
rect 672706 571719 672734 643361
rect 672802 572015 672830 644767
rect 672898 617451 672926 689759
rect 672982 688633 673034 688639
rect 672982 688575 673034 688581
rect 672886 617445 672938 617451
rect 672886 617387 672938 617393
rect 672994 616711 673022 688575
rect 673186 671249 673214 699823
rect 673270 689151 673322 689157
rect 673270 689093 673322 689099
rect 673174 671243 673226 671249
rect 673174 671185 673226 671191
rect 673078 649117 673130 649123
rect 673078 649059 673130 649065
rect 672982 616705 673034 616711
rect 672982 616647 673034 616653
rect 672886 599315 672938 599321
rect 672886 599257 672938 599263
rect 672790 572009 672842 572015
rect 672790 571951 672842 571957
rect 672694 571713 672746 571719
rect 672694 571655 672746 571661
rect 672598 537525 672650 537531
rect 672598 537467 672650 537473
rect 672898 528207 672926 599257
rect 672982 598427 673034 598433
rect 672982 598369 673034 598375
rect 672886 528201 672938 528207
rect 672886 528143 672938 528149
rect 672994 526727 673022 598369
rect 673090 574679 673118 649059
rect 673174 648303 673226 648309
rect 673174 648245 673226 648251
rect 673078 574673 673130 574679
rect 673078 574615 673130 574621
rect 673186 573939 673214 648245
rect 673282 618191 673310 689093
rect 673378 662665 673406 737859
rect 673474 664367 673502 738451
rect 673666 707435 673694 779891
rect 673762 755461 673790 876535
rect 675298 876419 675326 877509
rect 675394 876599 675422 876900
rect 675382 876593 675434 876599
rect 675382 876535 675434 876541
rect 675284 876410 675340 876419
rect 675284 876345 675340 876354
rect 675284 876262 675340 876271
rect 675340 876220 675408 876248
rect 675284 876197 675340 876206
rect 675490 874051 675518 874384
rect 675476 874042 675532 874051
rect 675476 873977 675532 873986
rect 675394 873491 675422 873866
rect 675382 873485 675434 873491
rect 675382 873427 675434 873433
rect 675394 872677 675422 873200
rect 673846 872671 673898 872677
rect 673846 872613 673898 872619
rect 675382 872671 675434 872677
rect 675382 872613 675434 872619
rect 673750 755455 673802 755461
rect 673750 755397 673802 755403
rect 673858 754351 673886 872613
rect 675490 872159 675518 872534
rect 675478 872153 675530 872159
rect 675478 872095 675530 872101
rect 674710 871191 674762 871197
rect 674710 871133 674762 871139
rect 674614 868379 674666 868385
rect 674614 868321 674666 868327
rect 674230 866529 674282 866535
rect 674230 866471 674282 866477
rect 674242 774891 674270 866471
rect 674626 777555 674654 868321
rect 674722 866313 674750 871133
rect 675394 869907 675422 870092
rect 675380 869898 675436 869907
rect 675380 869833 675436 869842
rect 675490 869199 675518 869500
rect 675478 869193 675530 869199
rect 675478 869135 675530 869141
rect 675394 868385 675422 868875
rect 675382 868379 675434 868385
rect 675382 868321 675434 868327
rect 675394 867867 675422 868242
rect 675382 867861 675434 867867
rect 675382 867803 675434 867809
rect 675208 866973 675260 866979
rect 675208 866915 675260 866921
rect 675220 866910 675248 866915
rect 675394 866535 675422 867058
rect 675382 866529 675434 866535
rect 675382 866471 675434 866477
rect 674710 866307 674762 866313
rect 674710 866249 674762 866255
rect 675382 866307 675434 866313
rect 675382 866249 675434 866255
rect 675394 865839 675422 866249
rect 675778 864727 675806 865208
rect 675764 864718 675820 864727
rect 675764 864653 675820 864662
rect 675394 862951 675422 863358
rect 675380 862942 675436 862951
rect 675380 862877 675436 862886
rect 675394 787915 675422 788322
rect 675380 787906 675436 787915
rect 675380 787841 675436 787850
rect 675490 787355 675518 787656
rect 675478 787349 675530 787355
rect 675478 787291 675530 787297
rect 675394 786731 675422 787035
rect 675380 786722 675436 786731
rect 675380 786657 675436 786666
rect 675490 784807 675518 785214
rect 675476 784798 675532 784807
rect 675476 784733 675532 784742
rect 675490 784321 675518 784622
rect 675478 784315 675530 784321
rect 675478 784257 675530 784263
rect 675394 783507 675422 783999
rect 675382 783501 675434 783507
rect 675382 783443 675434 783449
rect 674710 783353 674762 783359
rect 674710 783295 674762 783301
rect 674612 777546 674668 777555
rect 674612 777481 674668 777490
rect 674722 777069 674750 783295
rect 675490 782989 675518 783364
rect 675478 782983 675530 782989
rect 675478 782925 675530 782931
rect 675778 780663 675806 780848
rect 675764 780654 675820 780663
rect 675764 780589 675820 780598
rect 675394 779955 675422 780330
rect 675382 779949 675434 779955
rect 675382 779891 675434 779897
rect 675778 779183 675806 779664
rect 675764 779174 675820 779183
rect 675764 779109 675820 779118
rect 675394 778623 675422 779031
rect 675382 778617 675434 778623
rect 675382 778559 675434 778565
rect 675778 777407 675806 777814
rect 675764 777398 675820 777407
rect 675764 777333 675820 777342
rect 674710 777063 674762 777069
rect 674710 777005 674762 777011
rect 675382 777063 675434 777069
rect 675382 777005 675434 777011
rect 675394 776630 675422 777005
rect 675778 775483 675806 775995
rect 675764 775474 675820 775483
rect 675764 775409 675820 775418
rect 674228 774882 674284 774891
rect 674228 774817 674284 774826
rect 675490 773707 675518 774155
rect 675476 773698 675532 773707
rect 675476 773633 675532 773642
rect 676054 762929 676106 762935
rect 676052 762894 676054 762903
rect 676106 762894 676108 762903
rect 676052 762829 676108 762838
rect 676054 762337 676106 762343
rect 676052 762302 676054 762311
rect 676106 762302 676108 762311
rect 676052 762237 676108 762246
rect 676246 762041 676298 762047
rect 676244 762006 676246 762015
rect 676298 762006 676300 762015
rect 676244 761941 676300 761950
rect 676246 761597 676298 761603
rect 676244 761562 676246 761571
rect 676298 761562 676300 761571
rect 676244 761497 676300 761506
rect 676244 760674 676300 760683
rect 676244 760609 676246 760618
rect 676298 760609 676300 760618
rect 676246 760577 676298 760583
rect 676054 760339 676106 760345
rect 676052 760304 676054 760313
rect 676106 760304 676108 760313
rect 676052 760239 676108 760248
rect 676052 759934 676108 759943
rect 676052 759869 676054 759878
rect 676106 759869 676108 759878
rect 676054 759837 676106 759843
rect 676054 759377 676106 759383
rect 676052 759342 676054 759351
rect 676106 759342 676108 759351
rect 676052 759277 676108 759286
rect 676054 758859 676106 758865
rect 676052 758824 676054 758833
rect 676106 758824 676108 758833
rect 676052 758759 676108 758768
rect 676054 755455 676106 755461
rect 676052 755420 676054 755429
rect 676106 755420 676108 755429
rect 676052 755355 676108 755364
rect 676246 755085 676298 755091
rect 676244 755050 676246 755059
rect 676298 755050 676300 755059
rect 676244 754985 676300 754994
rect 673846 754345 673898 754351
rect 676054 754345 676106 754351
rect 673846 754287 673898 754293
rect 676052 754310 676054 754319
rect 676106 754310 676108 754319
rect 676052 754245 676108 754254
rect 676054 752865 676106 752871
rect 676052 752830 676054 752839
rect 676106 752830 676108 752839
rect 676052 752765 676108 752774
rect 676054 752421 676106 752427
rect 676052 752386 676054 752395
rect 676106 752386 676108 752395
rect 676052 752321 676108 752330
rect 676054 751903 676106 751909
rect 676052 751868 676054 751877
rect 676106 751868 676108 751877
rect 676052 751803 676108 751812
rect 679796 751498 679852 751507
rect 679796 751433 679852 751442
rect 679810 750619 679838 751433
rect 679796 750610 679852 750619
rect 679796 750545 679852 750554
rect 685460 750610 685516 750619
rect 685460 750545 685516 750554
rect 679810 748875 679838 750545
rect 685474 750175 685502 750545
rect 685460 750166 685516 750175
rect 685460 750101 685516 750110
rect 679798 748869 679850 748875
rect 679798 748811 679850 748817
rect 675394 743219 675422 743330
rect 675380 743210 675436 743219
rect 675380 743145 675436 743154
rect 675778 742183 675806 742664
rect 675764 742174 675820 742183
rect 675764 742109 675820 742118
rect 675394 741739 675422 742035
rect 675380 741730 675436 741739
rect 675380 741665 675436 741674
rect 675476 740398 675532 740407
rect 675476 740333 675532 740342
rect 675490 740222 675518 740333
rect 675490 739181 675518 739630
rect 673846 739175 673898 739181
rect 673846 739117 673898 739123
rect 675478 739175 675530 739181
rect 675478 739117 675530 739123
rect 673750 734957 673802 734963
rect 673750 734899 673802 734905
rect 673654 707429 673706 707435
rect 673654 707371 673706 707377
rect 673654 693517 673706 693523
rect 673654 693459 673706 693465
rect 673558 692925 673610 692931
rect 673558 692867 673610 692873
rect 673462 664361 673514 664367
rect 673462 664303 673514 664309
rect 673366 662659 673418 662665
rect 673366 662601 673418 662607
rect 673462 644011 673514 644017
rect 673462 643953 673514 643959
rect 673366 642309 673418 642315
rect 673366 642251 673418 642257
rect 673270 618185 673322 618191
rect 673270 618127 673322 618133
rect 673270 603311 673322 603317
rect 673270 603253 673322 603259
rect 673174 573933 673226 573939
rect 673174 573875 673226 573881
rect 673078 553953 673130 553959
rect 673078 553895 673130 553901
rect 672982 526721 673034 526727
rect 672982 526663 673034 526669
rect 672502 492977 672554 492983
rect 672502 492919 672554 492925
rect 673090 484029 673118 553895
rect 673174 553213 673226 553219
rect 673174 553155 673226 553161
rect 673078 484023 673130 484029
rect 673078 483965 673130 483971
rect 673186 482475 673214 553155
rect 673282 528947 673310 603253
rect 673378 573569 673406 642251
rect 673366 573563 673418 573569
rect 673366 573505 673418 573511
rect 673474 573051 673502 643953
rect 673570 617673 673598 692867
rect 673666 619227 673694 693459
rect 673762 662295 673790 734899
rect 673858 664663 673886 739117
rect 674710 738731 674762 738737
rect 674710 738673 674762 738679
rect 674722 732077 674750 738673
rect 675394 738515 675422 738999
rect 675382 738509 675434 738515
rect 675382 738451 675434 738457
rect 675394 737923 675422 738372
rect 675382 737917 675434 737923
rect 675382 737859 675434 737865
rect 675682 735523 675710 735856
rect 675668 735514 675724 735523
rect 675668 735449 675724 735458
rect 675394 734963 675422 735338
rect 675382 734957 675434 734963
rect 675382 734899 675434 734905
rect 675778 734487 675806 734672
rect 675764 734478 675820 734487
rect 675764 734413 675820 734422
rect 675490 733631 675518 734006
rect 675478 733625 675530 733631
rect 675478 733567 675530 733573
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 674710 732071 674762 732077
rect 674710 732013 674762 732019
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 674326 730517 674378 730523
rect 674326 730459 674378 730465
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 674230 685525 674282 685531
rect 674230 685467 674282 685473
rect 673846 664657 673898 664663
rect 673846 664599 673898 664605
rect 673750 662289 673802 662295
rect 673750 662231 673802 662237
rect 673750 652151 673802 652157
rect 673750 652093 673802 652099
rect 673654 619221 673706 619227
rect 673654 619163 673706 619169
rect 673558 617667 673610 617673
rect 673558 617609 673610 617615
rect 673558 603977 673610 603983
rect 673558 603919 673610 603925
rect 673462 573045 673514 573051
rect 673462 572987 673514 572993
rect 673570 529687 673598 603919
rect 673762 575049 673790 652093
rect 673846 647933 673898 647939
rect 673846 647875 673898 647881
rect 673750 575043 673802 575049
rect 673750 574985 673802 574991
rect 673858 572459 673886 647875
rect 674242 624925 674270 685467
rect 674338 668141 674366 730459
rect 675490 728673 675518 729155
rect 674518 728667 674570 728673
rect 674518 728609 674570 728615
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 674422 683675 674474 683681
rect 674422 683617 674474 683623
rect 674326 668135 674378 668141
rect 674326 668077 674378 668083
rect 674230 624919 674282 624925
rect 674230 624861 674282 624867
rect 674434 622039 674462 683617
rect 674530 668067 674558 728609
rect 679702 722969 679754 722975
rect 679702 722911 679754 722917
rect 676246 718085 676298 718091
rect 676244 718050 676246 718059
rect 676298 718050 676300 718059
rect 676244 717985 676300 717994
rect 676054 717345 676106 717351
rect 676052 717310 676054 717319
rect 676106 717310 676108 717319
rect 676052 717245 676108 717254
rect 676246 717049 676298 717055
rect 676244 717014 676246 717023
rect 676298 717014 676300 717023
rect 676244 716949 676300 716958
rect 679714 716579 679742 722911
rect 679700 716570 679756 716579
rect 679700 716505 679756 716514
rect 679700 715534 679756 715543
rect 679700 715469 679756 715478
rect 676054 715347 676106 715353
rect 676052 715312 676054 715321
rect 676106 715312 676108 715321
rect 676052 715247 676108 715256
rect 676052 714942 676108 714951
rect 676052 714877 676054 714886
rect 676106 714877 676108 714886
rect 676054 714845 676106 714851
rect 676054 714385 676106 714391
rect 676052 714350 676054 714359
rect 676106 714350 676108 714359
rect 676052 714285 676108 714294
rect 676054 713793 676106 713799
rect 676052 713758 676054 713767
rect 676106 713758 676108 713767
rect 676052 713693 676108 713702
rect 676054 710463 676106 710469
rect 676052 710428 676054 710437
rect 676106 710428 676108 710437
rect 676052 710363 676108 710372
rect 676246 710093 676298 710099
rect 676244 710058 676246 710067
rect 676298 710058 676300 710067
rect 676244 709993 676300 710002
rect 676054 709353 676106 709359
rect 676052 709318 676054 709327
rect 676106 709318 676108 709327
rect 676052 709253 676108 709262
rect 676246 708021 676298 708027
rect 676244 707986 676246 707995
rect 676298 707986 676300 707995
rect 676244 707921 676300 707930
rect 676054 707429 676106 707435
rect 676052 707394 676054 707403
rect 676106 707394 676108 707403
rect 676052 707329 676108 707338
rect 676054 706911 676106 706917
rect 676052 706876 676054 706885
rect 676106 706876 676108 706885
rect 676052 706811 676108 706820
rect 679714 699887 679742 715469
rect 679988 706506 680044 706515
rect 679988 706441 680044 706450
rect 680002 705627 680030 706441
rect 679796 705618 679852 705627
rect 679796 705553 679852 705562
rect 679988 705618 680044 705627
rect 679988 705553 680044 705562
rect 679810 705183 679838 705553
rect 679796 705174 679852 705183
rect 679796 705109 679852 705118
rect 680002 702773 680030 705553
rect 679990 702767 680042 702773
rect 679990 702709 680042 702715
rect 679702 699881 679754 699887
rect 679702 699823 679754 699829
rect 675394 697931 675422 698338
rect 675380 697922 675436 697931
rect 675380 697857 675436 697866
rect 675778 697339 675806 697672
rect 675764 697330 675820 697339
rect 675764 697265 675820 697274
rect 675586 696895 675614 697035
rect 675572 696886 675628 696895
rect 675572 696821 675628 696830
rect 675394 694823 675422 695195
rect 675380 694814 675436 694823
rect 675380 694749 675436 694758
rect 675778 694231 675806 694638
rect 675764 694222 675820 694231
rect 675764 694157 675820 694166
rect 675490 693523 675518 693972
rect 675478 693517 675530 693523
rect 675478 693459 675530 693465
rect 675490 692931 675518 693380
rect 675478 692925 675530 692931
rect 675478 692867 675530 692873
rect 674710 692629 674762 692635
rect 674710 692571 674762 692577
rect 674722 687085 674750 692571
rect 675490 690531 675518 690864
rect 675476 690522 675532 690531
rect 675476 690457 675532 690466
rect 675394 689823 675422 690346
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675394 689157 675422 689680
rect 675382 689151 675434 689157
rect 675382 689093 675434 689099
rect 675490 688639 675518 689014
rect 675478 688633 675530 688639
rect 675478 688575 675530 688581
rect 675778 687423 675806 687830
rect 675764 687414 675820 687423
rect 675764 687349 675820 687358
rect 674710 687079 674762 687085
rect 674710 687021 674762 687027
rect 675478 687079 675530 687085
rect 675478 687021 675530 687027
rect 675490 686646 675518 687021
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 676054 672723 676106 672729
rect 676052 672688 676054 672697
rect 676106 672688 676108 672697
rect 676052 672623 676108 672632
rect 676246 672353 676298 672359
rect 676244 672318 676246 672327
rect 676298 672318 676300 672327
rect 676244 672253 676300 672262
rect 676054 671613 676106 671619
rect 676052 671578 676054 671587
rect 676106 671578 676108 671587
rect 676052 671513 676108 671522
rect 676054 671243 676106 671249
rect 676052 671208 676054 671217
rect 676106 671208 676108 671217
rect 676052 671143 676108 671152
rect 676052 670690 676108 670699
rect 676052 670625 676054 670634
rect 676106 670625 676108 670634
rect 676054 670593 676106 670599
rect 676054 670133 676106 670139
rect 676052 670098 676054 670107
rect 676106 670098 676108 670107
rect 676052 670033 676108 670042
rect 676052 669654 676108 669663
rect 676052 669589 676054 669598
rect 676106 669589 676108 669598
rect 676054 669557 676106 669563
rect 676246 669393 676298 669399
rect 676244 669358 676246 669367
rect 676298 669358 676300 669367
rect 676244 669293 676300 669302
rect 679892 668914 679948 668923
rect 679892 668849 679948 668858
rect 676054 668135 676106 668141
rect 676054 668077 676106 668083
rect 674518 668061 674570 668067
rect 674518 668003 674570 668009
rect 676066 667665 676094 668077
rect 676246 668061 676298 668067
rect 676246 668003 676298 668009
rect 676052 667656 676108 667665
rect 676052 667591 676108 667600
rect 676258 665815 676286 668003
rect 676244 665806 676300 665815
rect 676244 665741 676300 665750
rect 676054 664657 676106 664663
rect 676052 664622 676054 664631
rect 676106 664622 676108 664631
rect 676052 664557 676108 664566
rect 676246 664361 676298 664367
rect 676244 664326 676246 664335
rect 676298 664326 676300 664335
rect 676244 664261 676300 664270
rect 676246 663917 676298 663923
rect 676244 663882 676246 663891
rect 676298 663882 676300 663891
rect 676244 663817 676300 663826
rect 676054 662659 676106 662665
rect 676052 662624 676054 662633
rect 676106 662624 676108 662633
rect 676052 662559 676108 662568
rect 676054 662289 676106 662295
rect 676052 662254 676054 662263
rect 676106 662254 676108 662263
rect 676052 662189 676108 662198
rect 676054 661697 676106 661703
rect 676052 661662 676054 661671
rect 676106 661662 676108 661671
rect 676052 661597 676108 661606
rect 679796 660922 679852 660931
rect 679796 660857 679852 660866
rect 679810 660487 679838 660857
rect 679796 660478 679852 660487
rect 679796 660413 679852 660422
rect 679810 659557 679838 660413
rect 679798 659551 679850 659557
rect 679798 659493 679850 659499
rect 679906 656745 679934 668849
rect 685556 660478 685612 660487
rect 685556 660413 685612 660422
rect 685570 659895 685598 660413
rect 685556 659886 685612 659895
rect 685556 659821 685612 659830
rect 679894 656739 679946 656745
rect 679894 656681 679946 656687
rect 675394 652643 675422 653124
rect 675380 652634 675436 652643
rect 675380 652569 675436 652578
rect 675490 652157 675518 652458
rect 675478 652151 675530 652157
rect 675478 652093 675530 652099
rect 675394 651607 675422 651835
rect 675380 651598 675436 651607
rect 675380 651533 675436 651542
rect 675682 649683 675710 650016
rect 675668 649674 675724 649683
rect 675668 649609 675724 649618
rect 675490 649123 675518 649424
rect 675478 649117 675530 649123
rect 675478 649059 675530 649065
rect 675394 648309 675422 648799
rect 675382 648303 675434 648309
rect 675382 648245 675434 648251
rect 675490 647939 675518 648166
rect 675478 647933 675530 647939
rect 675478 647875 675530 647881
rect 674710 646601 674762 646607
rect 674710 646543 674762 646549
rect 674722 641871 674750 646543
rect 675490 645391 675518 645650
rect 675476 645382 675532 645391
rect 675476 645317 675532 645326
rect 675394 644831 675422 645132
rect 675382 644825 675434 644831
rect 675382 644767 675434 644773
rect 675490 644017 675518 644466
rect 675478 644011 675530 644017
rect 675478 643953 675530 643959
rect 675394 643425 675422 643831
rect 675382 643419 675434 643425
rect 675382 643361 675434 643367
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 674710 641865 674762 641871
rect 674710 641807 674762 641813
rect 675382 641865 675434 641871
rect 675382 641807 675434 641813
rect 675394 641432 675422 641807
rect 675778 640359 675806 640795
rect 675764 640350 675820 640359
rect 675764 640285 675820 640294
rect 675490 638583 675518 638955
rect 675476 638574 675532 638583
rect 675476 638509 675532 638518
rect 679702 635649 679754 635655
rect 679702 635591 679754 635597
rect 676054 627731 676106 627737
rect 676052 627696 676054 627705
rect 676106 627696 676108 627705
rect 676052 627631 676108 627640
rect 676246 627361 676298 627367
rect 676244 627326 676246 627335
rect 676298 627326 676300 627335
rect 676244 627261 676300 627270
rect 676054 626621 676106 626627
rect 676052 626586 676054 626595
rect 676106 626586 676108 626595
rect 676052 626521 676108 626530
rect 679714 626447 679742 635591
rect 679700 626438 679756 626447
rect 679700 626373 679756 626382
rect 676052 625698 676108 625707
rect 676052 625633 676054 625642
rect 676106 625633 676108 625642
rect 676054 625601 676106 625607
rect 676054 624919 676106 624925
rect 676054 624861 676106 624867
rect 675958 624697 676010 624703
rect 675956 624662 675958 624671
rect 676010 624662 676012 624671
rect 675956 624597 676012 624606
rect 675956 623626 676012 623635
rect 675956 623561 675958 623570
rect 676010 623561 676012 623570
rect 675958 623529 676010 623535
rect 676066 622673 676094 624861
rect 676052 622664 676108 622673
rect 676052 622599 676108 622608
rect 674422 622033 674474 622039
rect 674422 621975 674474 621981
rect 676246 622033 676298 622039
rect 676246 621975 676298 621981
rect 676258 620823 676286 621975
rect 676244 620814 676300 620823
rect 676244 620749 676300 620758
rect 676054 619221 676106 619227
rect 676052 619186 676054 619195
rect 676106 619186 676108 619195
rect 676052 619121 676108 619130
rect 676054 618185 676106 618191
rect 676052 618150 676054 618159
rect 676106 618150 676108 618159
rect 676052 618085 676108 618094
rect 676054 617667 676106 617673
rect 676052 617632 676054 617641
rect 676106 617632 676108 617641
rect 676052 617567 676108 617576
rect 676246 617445 676298 617451
rect 676244 617410 676246 617419
rect 676298 617410 676300 617419
rect 676244 617345 676300 617354
rect 676054 616705 676106 616711
rect 676052 616670 676054 616679
rect 676106 616670 676108 616679
rect 676052 616605 676108 616614
rect 679796 615930 679852 615939
rect 679796 615865 679852 615874
rect 679810 615347 679838 615865
rect 679796 615338 679852 615347
rect 679796 615273 679852 615282
rect 685460 615338 685516 615347
rect 685460 615273 685516 615282
rect 679810 613529 679838 615273
rect 685474 614903 685502 615273
rect 685460 614894 685516 614903
rect 685460 614829 685516 614838
rect 679798 613523 679850 613529
rect 679798 613465 679850 613471
rect 675394 607799 675422 608132
rect 675380 607790 675436 607799
rect 675380 607725 675436 607734
rect 675490 607091 675518 607466
rect 675478 607085 675530 607091
rect 675478 607027 675530 607033
rect 675394 606467 675422 606835
rect 675380 606458 675436 606467
rect 675380 606393 675436 606402
rect 675394 604839 675422 604995
rect 675380 604830 675436 604839
rect 675380 604765 675436 604774
rect 675490 603983 675518 604432
rect 675478 603977 675530 603983
rect 675478 603919 675530 603925
rect 674614 603385 674666 603391
rect 674614 603327 674666 603333
rect 674626 596879 674654 603327
rect 675394 603317 675422 603799
rect 675382 603311 675434 603317
rect 675382 603253 675434 603259
rect 675394 602725 675422 603174
rect 675382 602719 675434 602725
rect 675382 602661 675434 602667
rect 675490 600251 675518 600658
rect 675476 600242 675532 600251
rect 675476 600177 675532 600186
rect 675394 599839 675422 600140
rect 675382 599833 675434 599839
rect 675382 599775 675434 599781
rect 675394 599321 675422 599474
rect 675382 599315 675434 599321
rect 675382 599257 675434 599263
rect 675490 598433 675518 598808
rect 675478 598427 675530 598433
rect 675478 598369 675530 598375
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 674614 596873 674666 596879
rect 674614 596815 674666 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675778 595367 675806 595774
rect 675764 595358 675820 595367
rect 675764 595293 675820 595302
rect 675490 593443 675518 593955
rect 675476 593434 675532 593443
rect 675476 593369 675532 593378
rect 676054 582517 676106 582523
rect 676052 582482 676054 582491
rect 676106 582482 676108 582491
rect 676052 582417 676108 582426
rect 676054 581999 676106 582005
rect 676052 581964 676054 581973
rect 676106 581964 676108 581973
rect 676052 581899 676108 581908
rect 676246 581629 676298 581635
rect 676244 581594 676246 581603
rect 676298 581594 676300 581603
rect 676244 581529 676300 581538
rect 676054 581037 676106 581043
rect 676052 581002 676054 581011
rect 676106 581002 676108 581011
rect 676052 580937 676108 580946
rect 676244 580262 676300 580271
rect 676244 580197 676246 580206
rect 676298 580197 676300 580206
rect 676246 580165 676298 580171
rect 676054 580001 676106 580007
rect 676052 579966 676054 579975
rect 676106 579966 676108 579975
rect 676052 579901 676108 579910
rect 676052 579522 676108 579531
rect 676052 579457 676054 579466
rect 676106 579457 676108 579466
rect 676054 579425 676106 579431
rect 676054 578965 676106 578971
rect 676052 578930 676054 578939
rect 676106 578930 676108 578939
rect 676052 578865 676108 578874
rect 676054 578447 676106 578453
rect 676052 578412 676054 578421
rect 676106 578412 676108 578421
rect 676052 578347 676108 578356
rect 676054 575043 676106 575049
rect 676052 575008 676054 575017
rect 676106 575008 676108 575017
rect 676052 574943 676108 574952
rect 676246 574673 676298 574679
rect 676244 574638 676246 574647
rect 676298 574638 676300 574647
rect 676244 574573 676300 574582
rect 676054 573933 676106 573939
rect 676052 573898 676054 573907
rect 676106 573898 676108 573907
rect 676052 573833 676108 573842
rect 676054 573563 676106 573569
rect 676052 573528 676054 573537
rect 676106 573528 676108 573537
rect 676052 573463 676108 573472
rect 676054 573045 676106 573051
rect 676052 573010 676054 573019
rect 676106 573010 676108 573019
rect 676052 572945 676108 572954
rect 673846 572453 673898 572459
rect 676054 572453 676106 572459
rect 673846 572395 673898 572401
rect 676052 572418 676054 572427
rect 676106 572418 676108 572427
rect 676052 572353 676108 572362
rect 676054 572009 676106 572015
rect 676052 571974 676054 571983
rect 676106 571974 676108 571983
rect 676052 571909 676108 571918
rect 676246 571713 676298 571719
rect 676244 571678 676246 571687
rect 676298 571678 676300 571687
rect 676244 571613 676300 571622
rect 679988 571234 680044 571243
rect 679988 571169 680044 571178
rect 680002 570207 680030 571169
rect 679796 570198 679852 570207
rect 679796 570133 679852 570142
rect 679988 570198 680044 570207
rect 679988 570133 680044 570142
rect 679810 569763 679838 570133
rect 679796 569754 679852 569763
rect 679796 569689 679852 569698
rect 680002 567427 680030 570133
rect 679990 567421 680042 567427
rect 679990 567363 680042 567369
rect 675490 562659 675518 562918
rect 675476 562650 675532 562659
rect 675476 562585 675532 562594
rect 675490 561771 675518 562252
rect 675476 561762 675532 561771
rect 675476 561697 675532 561706
rect 675490 561475 675518 561660
rect 675476 561466 675532 561475
rect 675476 561401 675532 561410
rect 675394 559435 675422 559810
rect 674614 559429 674666 559435
rect 674614 559371 674666 559377
rect 675382 559429 675434 559435
rect 675382 559371 675434 559377
rect 674518 558985 674570 558991
rect 674518 558927 674570 558933
rect 673846 558097 673898 558103
rect 673846 558039 673898 558045
rect 673750 554397 673802 554403
rect 673750 554339 673802 554345
rect 673654 551955 673706 551961
rect 673654 551897 673706 551903
rect 673558 529681 673610 529687
rect 673558 529623 673610 529629
rect 673270 528941 673322 528947
rect 673270 528883 673322 528889
rect 673666 484547 673694 551897
rect 673654 484541 673706 484547
rect 673654 484483 673706 484489
rect 673762 483067 673790 554339
rect 673858 485139 673886 558039
rect 674422 548921 674474 548927
rect 674422 548863 674474 548869
rect 674326 548255 674378 548261
rect 674326 548197 674378 548203
rect 674338 486619 674366 548197
rect 674434 489431 674462 548863
rect 674422 489425 674474 489431
rect 674422 489367 674474 489373
rect 674530 486693 674558 558927
rect 674626 489505 674654 559371
rect 675490 558991 675518 559218
rect 675478 558985 675530 558991
rect 675478 558927 675530 558933
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675778 557627 675806 557960
rect 675764 557618 675820 557627
rect 675764 557553 675820 557562
rect 675286 557283 675338 557289
rect 675286 557225 675338 557231
rect 674710 555285 674762 555291
rect 674710 555227 674762 555233
rect 674722 528577 674750 555227
rect 675298 551240 675326 557225
rect 675490 555291 675518 555444
rect 675478 555285 675530 555291
rect 675478 555227 675530 555233
rect 675394 554403 675422 554926
rect 675382 554397 675434 554403
rect 675382 554339 675434 554345
rect 675490 553959 675518 554260
rect 675478 553953 675530 553959
rect 675478 553895 675530 553901
rect 675394 553219 675422 553631
rect 675382 553213 675434 553219
rect 675382 553155 675434 553161
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 675298 551212 675408 551240
rect 675298 550581 675408 550609
rect 675298 548927 675326 550581
rect 675286 548921 675338 548927
rect 675286 548863 675338 548869
rect 675298 548741 675408 548769
rect 675298 548261 675326 548741
rect 675286 548255 675338 548261
rect 675286 548197 675338 548203
rect 679702 547219 679754 547225
rect 679702 547161 679754 547167
rect 676726 541373 676778 541379
rect 676726 541315 676778 541321
rect 676054 537525 676106 537531
rect 676052 537490 676054 537499
rect 676106 537490 676108 537499
rect 676052 537425 676108 537434
rect 676630 537377 676682 537383
rect 676630 537319 676682 537325
rect 676054 536933 676106 536939
rect 676052 536898 676054 536907
rect 676106 536898 676108 536907
rect 676052 536833 676108 536842
rect 676246 536637 676298 536643
rect 676244 536602 676246 536611
rect 676298 536602 676300 536611
rect 676244 536537 676300 536546
rect 676532 535270 676588 535279
rect 676532 535205 676588 535214
rect 676054 534935 676106 534941
rect 676052 534900 676054 534909
rect 676106 534900 676108 534909
rect 676052 534835 676108 534844
rect 676054 533973 676106 533979
rect 676052 533938 676054 533947
rect 676106 533938 676108 533947
rect 676052 533873 676108 533882
rect 676054 530051 676106 530057
rect 676052 530016 676054 530025
rect 676106 530016 676108 530025
rect 676052 529951 676108 529960
rect 676246 529681 676298 529687
rect 676244 529646 676246 529655
rect 676298 529646 676300 529655
rect 676244 529581 676300 529590
rect 676054 528941 676106 528947
rect 676052 528906 676054 528915
rect 676106 528906 676108 528915
rect 676052 528841 676108 528850
rect 674710 528571 674762 528577
rect 674710 528513 674762 528519
rect 674998 528571 675050 528577
rect 674998 528513 675050 528519
rect 675010 489579 675038 528513
rect 676054 528497 676106 528503
rect 676052 528462 676054 528471
rect 676106 528462 676108 528471
rect 676052 528397 676108 528406
rect 676246 528201 676298 528207
rect 676244 528166 676246 528175
rect 676298 528166 676300 528175
rect 676244 528101 676300 528110
rect 676054 527461 676106 527467
rect 676052 527426 676054 527435
rect 676106 527426 676108 527435
rect 676052 527361 676108 527370
rect 676054 527017 676106 527023
rect 676052 526982 676054 526991
rect 676106 526982 676108 526991
rect 676052 526917 676108 526926
rect 676246 526721 676298 526727
rect 676244 526686 676246 526695
rect 676298 526686 676300 526695
rect 676244 526621 676300 526630
rect 676546 498311 676574 535205
rect 676642 534243 676670 537319
rect 676628 534234 676684 534243
rect 676628 534169 676684 534178
rect 676534 498305 676586 498311
rect 676534 498247 676586 498253
rect 676246 493717 676298 493723
rect 676244 493682 676246 493691
rect 676298 493682 676300 493691
rect 676244 493617 676300 493626
rect 676054 492977 676106 492983
rect 676052 492942 676054 492951
rect 676106 492942 676108 492951
rect 676052 492877 676108 492886
rect 676054 492385 676106 492391
rect 676052 492350 676054 492359
rect 676106 492350 676108 492359
rect 676052 492285 676108 492294
rect 676532 491610 676588 491619
rect 676532 491545 676588 491554
rect 674998 489573 675050 489579
rect 674998 489515 675050 489521
rect 676246 489573 676298 489579
rect 676246 489515 676298 489521
rect 674614 489499 674666 489505
rect 674614 489441 674666 489447
rect 676054 489499 676106 489505
rect 676054 489441 676106 489447
rect 676066 487475 676094 489441
rect 676150 489425 676202 489431
rect 676150 489367 676202 489373
rect 676162 488659 676190 489367
rect 676148 488650 676204 488659
rect 676148 488585 676204 488594
rect 676052 487466 676108 487475
rect 676052 487401 676108 487410
rect 676258 487179 676286 489515
rect 676244 487170 676300 487179
rect 676244 487105 676300 487114
rect 674518 486687 674570 486693
rect 674518 486629 674570 486635
rect 676054 486687 676106 486693
rect 676054 486629 676106 486635
rect 674326 486613 674378 486619
rect 674326 486555 674378 486561
rect 676066 485477 676094 486629
rect 676246 486613 676298 486619
rect 676244 486578 676246 486587
rect 676298 486578 676300 486587
rect 676244 486513 676300 486522
rect 676052 485468 676108 485477
rect 676052 485403 676108 485412
rect 673846 485133 673898 485139
rect 676246 485133 676298 485139
rect 673846 485075 673898 485081
rect 676244 485098 676246 485107
rect 676298 485098 676300 485107
rect 676244 485033 676300 485042
rect 676054 484541 676106 484547
rect 676052 484506 676054 484515
rect 676106 484506 676108 484515
rect 676052 484441 676108 484450
rect 676054 484023 676106 484029
rect 676052 483988 676054 483997
rect 676106 483988 676108 483997
rect 676052 483923 676108 483932
rect 673750 483061 673802 483067
rect 676054 483061 676106 483067
rect 673750 483003 673802 483009
rect 676052 483026 676054 483035
rect 676106 483026 676108 483035
rect 676052 482961 676108 482970
rect 673174 482469 673226 482475
rect 676054 482469 676106 482475
rect 673174 482411 673226 482417
rect 676052 482434 676054 482443
rect 676106 482434 676108 482443
rect 676052 482369 676108 482378
rect 672598 443619 672650 443625
rect 672598 443561 672650 443567
rect 672502 417645 672554 417651
rect 672502 417587 672554 417593
rect 672406 359777 672458 359783
rect 672406 359719 672458 359725
rect 670966 356595 671018 356601
rect 670966 356537 671018 356543
rect 670978 354307 671006 356537
rect 670294 354301 670346 354307
rect 670294 354243 670346 354249
rect 670966 354301 671018 354307
rect 670966 354243 671018 354249
rect 670306 278647 670334 354243
rect 672406 311085 672458 311091
rect 672406 311027 672458 311033
rect 670292 278638 670348 278647
rect 670292 278573 670348 278582
rect 670100 278342 670156 278351
rect 670100 278277 670156 278286
rect 670006 225097 670058 225103
rect 670006 225039 670058 225045
rect 672418 134379 672446 311027
rect 672514 270095 672542 417587
rect 672610 314051 672638 443561
rect 676246 405509 676298 405515
rect 676244 405474 676246 405483
rect 676298 405474 676300 405483
rect 676244 405409 676300 405418
rect 676054 404769 676106 404775
rect 676052 404734 676054 404743
rect 676106 404734 676108 404743
rect 676052 404669 676108 404678
rect 676054 404251 676106 404257
rect 676052 404216 676054 404225
rect 676106 404216 676108 404225
rect 676052 404151 676108 404160
rect 676546 404003 676574 491545
rect 676642 491175 676670 534169
rect 676738 533207 676766 541315
rect 679714 536167 679742 547161
rect 679700 536158 679756 536167
rect 679700 536093 679756 536102
rect 676724 533198 676780 533207
rect 676724 533133 676780 533142
rect 676628 491166 676684 491175
rect 676628 491101 676684 491110
rect 676628 490278 676684 490287
rect 676628 490213 676684 490222
rect 676642 489376 676670 490213
rect 676738 490139 676766 533133
rect 679796 526094 679852 526103
rect 679796 526029 679852 526038
rect 679810 525215 679838 526029
rect 679796 525206 679852 525215
rect 679796 525141 679852 525150
rect 685460 525206 685516 525215
rect 685460 525141 685516 525150
rect 679810 524211 679838 525141
rect 685474 524771 685502 525141
rect 685460 524762 685516 524771
rect 685460 524697 685516 524706
rect 679798 524205 679850 524211
rect 679798 524147 679850 524153
rect 679702 498305 679754 498311
rect 679702 498247 679754 498253
rect 679714 492211 679742 498247
rect 679700 492202 679756 492211
rect 679700 492137 679756 492146
rect 676724 490130 676780 490139
rect 676724 490065 676780 490074
rect 676642 489348 676766 489376
rect 676628 489242 676684 489251
rect 676628 489177 676684 489186
rect 676532 403994 676588 404003
rect 676532 403929 676588 403938
rect 673846 403289 673898 403295
rect 676054 403289 676106 403295
rect 673846 403231 673898 403237
rect 676052 403254 676054 403263
rect 676106 403254 676108 403263
rect 673750 395741 673802 395747
rect 673750 395683 673802 395689
rect 673654 394039 673706 394045
rect 673654 393981 673706 393987
rect 673666 376877 673694 393981
rect 673762 377247 673790 395683
rect 673750 377241 673802 377247
rect 673750 377183 673802 377189
rect 673654 376871 673706 376877
rect 673654 376813 673706 376819
rect 673858 358599 673886 403231
rect 676052 403189 676108 403198
rect 676052 402292 676108 402301
rect 676052 402227 676054 402236
rect 676106 402227 676108 402236
rect 676054 402195 676106 402201
rect 676642 402111 676670 489177
rect 676738 402967 676766 489348
rect 679988 481694 680044 481703
rect 679988 481629 680044 481638
rect 680002 481259 680030 481629
rect 679796 481250 679852 481259
rect 679796 481185 679852 481194
rect 679988 481250 680044 481259
rect 679988 481185 680044 481194
rect 679810 480815 679838 481185
rect 679796 480806 679852 480815
rect 679796 480741 679852 480750
rect 680002 479515 680030 481185
rect 679990 479509 680042 479515
rect 679990 479451 680042 479457
rect 676724 402958 676780 402967
rect 676724 402893 676780 402902
rect 676054 402105 676106 402111
rect 676054 402047 676106 402053
rect 676630 402105 676682 402111
rect 676630 402047 676682 402053
rect 676066 401783 676094 402047
rect 676052 401774 676108 401783
rect 676052 401709 676108 401718
rect 676066 401297 676094 401709
rect 676054 401291 676106 401297
rect 676054 401233 676106 401239
rect 676244 401034 676300 401043
rect 676244 400969 676246 400978
rect 676298 400969 676300 400978
rect 676246 400937 676298 400943
rect 676738 400409 676766 402893
rect 674326 400403 674378 400409
rect 674326 400345 674378 400351
rect 676726 400403 676778 400409
rect 676726 400345 676778 400351
rect 674338 385905 674366 400345
rect 676052 395780 676108 395789
rect 676052 395715 676054 395724
rect 676106 395715 676108 395724
rect 676054 395683 676106 395689
rect 676244 394078 676300 394087
rect 676244 394013 676246 394022
rect 676298 394013 676300 394022
rect 676246 393981 676298 393987
rect 679796 393486 679852 393495
rect 679796 393421 679852 393430
rect 679810 393051 679838 393421
rect 679796 393042 679852 393051
rect 679796 392977 679852 392986
rect 685556 393042 685612 393051
rect 685556 392977 685612 392986
rect 679810 391751 679838 392977
rect 685570 392607 685598 392977
rect 685556 392598 685612 392607
rect 685556 392533 685612 392542
rect 679798 391745 679850 391751
rect 679798 391687 679850 391693
rect 675764 385938 675820 385947
rect 674326 385899 674378 385905
rect 675764 385873 675820 385882
rect 674326 385841 674378 385847
rect 675778 385723 675806 385873
rect 675764 385642 675820 385651
rect 675764 385577 675820 385586
rect 675778 385096 675806 385577
rect 675764 384754 675820 384763
rect 675764 384689 675820 384698
rect 675778 384430 675806 384689
rect 675380 382978 675436 382987
rect 675380 382913 675436 382922
rect 675284 382830 675340 382839
rect 675284 382765 675340 382774
rect 675298 381410 675326 382765
rect 675394 382580 675422 382913
rect 675476 382238 675532 382247
rect 675476 382173 675532 382182
rect 675490 382062 675518 382173
rect 675298 381382 675408 381410
rect 675764 381202 675820 381211
rect 675764 381137 675820 381146
rect 675778 380730 675806 381137
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675764 377946 675820 377955
rect 675764 377881 675820 377890
rect 675778 377696 675806 377881
rect 675382 377241 675434 377247
rect 675382 377183 675434 377189
rect 675394 377075 675422 377183
rect 675286 376871 675338 376877
rect 675286 376813 675338 376819
rect 675298 376452 675326 376813
rect 675298 376424 675408 376452
rect 675764 375726 675820 375735
rect 675764 375661 675820 375670
rect 675778 375254 675806 375661
rect 675188 373802 675244 373811
rect 675188 373737 675244 373746
rect 675202 373418 675230 373737
rect 675202 373390 675408 373418
rect 675572 372026 675628 372035
rect 675572 371961 675628 371970
rect 675586 371554 675614 371961
rect 676054 360073 676106 360079
rect 676052 360038 676054 360047
rect 676106 360038 676108 360047
rect 676052 359973 676108 359982
rect 676246 359777 676298 359783
rect 676244 359742 676246 359751
rect 676298 359742 676300 359751
rect 676244 359677 676300 359686
rect 676054 359037 676106 359043
rect 676052 359002 676054 359011
rect 676106 359002 676108 359011
rect 676052 358937 676108 358946
rect 673846 358593 673898 358599
rect 676054 358593 676106 358599
rect 673846 358535 673898 358541
rect 676052 358558 676054 358567
rect 676106 358558 676108 358567
rect 676052 358493 676108 358502
rect 676246 357779 676298 357785
rect 676246 357721 676298 357727
rect 676258 357679 676286 357721
rect 676244 357670 676300 357679
rect 676244 357605 676300 357614
rect 676054 356595 676106 356601
rect 676052 356560 676054 356569
rect 676106 356560 676108 356569
rect 676052 356495 676108 356504
rect 675764 354562 675820 354571
rect 675764 354497 675820 354506
rect 675284 352638 675340 352647
rect 675284 352573 675340 352582
rect 674806 351415 674858 351421
rect 674806 351357 674858 351363
rect 673942 349935 673994 349941
rect 673942 349877 673994 349883
rect 673954 332255 673982 349877
rect 674038 349195 674090 349201
rect 674038 349137 674090 349143
rect 674050 332773 674078 349137
rect 674230 348603 674282 348609
rect 674230 348545 674282 348551
rect 674242 336103 674270 348545
rect 674710 348529 674762 348535
rect 674710 348471 674762 348477
rect 674230 336097 674282 336103
rect 674230 336039 674282 336045
rect 674038 332767 674090 332773
rect 674038 332709 674090 332715
rect 673942 332249 673994 332255
rect 673942 332191 673994 332197
rect 674722 331811 674750 348471
rect 674818 337953 674846 351357
rect 675298 339896 675326 352573
rect 675778 341209 675806 354497
rect 676052 354118 676108 354127
rect 676052 354053 676108 354062
rect 676066 351421 676094 354053
rect 676054 351415 676106 351421
rect 676054 351357 676106 351363
rect 676244 350418 676300 350427
rect 676244 350353 676300 350362
rect 676258 349941 676286 350353
rect 676246 349935 676298 349941
rect 676246 349877 676298 349883
rect 676244 349826 676300 349835
rect 676244 349761 676300 349770
rect 676052 349678 676108 349687
rect 676052 349613 676108 349622
rect 676066 349201 676094 349613
rect 676054 349195 676106 349201
rect 676054 349137 676106 349143
rect 676052 349086 676108 349095
rect 676052 349021 676108 349030
rect 676066 348535 676094 349021
rect 676258 348609 676286 349761
rect 676246 348603 676298 348609
rect 676246 348545 676298 348551
rect 676054 348529 676106 348535
rect 676054 348471 676106 348477
rect 679796 348346 679852 348355
rect 679796 348281 679852 348290
rect 679810 347763 679838 348281
rect 679796 347754 679852 347763
rect 679796 347689 679852 347698
rect 685460 347754 685516 347763
rect 685460 347689 685516 347698
rect 679810 345649 679838 347689
rect 685474 347319 685502 347689
rect 685460 347310 685516 347319
rect 685460 347245 685516 347254
rect 679798 345643 679850 345649
rect 679798 345585 679850 345591
rect 675766 341203 675818 341209
rect 675766 341145 675818 341151
rect 675766 340981 675818 340987
rect 675766 340923 675818 340929
rect 675778 340548 675806 340923
rect 675298 339868 675408 339896
rect 675764 339614 675820 339623
rect 675764 339549 675820 339558
rect 675778 339216 675806 339549
rect 674806 337947 674858 337953
rect 674806 337889 674858 337895
rect 675478 337947 675530 337953
rect 675478 337889 675530 337895
rect 675490 337395 675518 337889
rect 675476 337098 675532 337107
rect 675476 337033 675532 337042
rect 675490 336848 675518 337033
rect 675764 336506 675820 336515
rect 675764 336441 675820 336450
rect 675778 336182 675806 336441
rect 675382 336097 675434 336103
rect 675382 336039 675434 336045
rect 675394 335555 675422 336039
rect 675380 333546 675436 333555
rect 675380 333481 675436 333490
rect 675394 333074 675422 333481
rect 675382 332767 675434 332773
rect 675382 332709 675434 332715
rect 675394 332519 675422 332709
rect 675478 332249 675530 332255
rect 675478 332191 675530 332197
rect 675490 331890 675518 332191
rect 674710 331805 674762 331811
rect 674710 331747 674762 331753
rect 675382 331805 675434 331811
rect 675382 331747 675434 331753
rect 675394 331224 675422 331747
rect 675476 330586 675532 330595
rect 675476 330521 675532 330530
rect 675490 330040 675518 330521
rect 675380 328366 675436 328375
rect 675380 328301 675436 328310
rect 675394 328190 675422 328301
rect 675380 326886 675436 326895
rect 675380 326821 675436 326830
rect 675394 326340 675422 326821
rect 676054 315081 676106 315087
rect 676052 315046 676054 315055
rect 676106 315046 676108 315055
rect 676052 314981 676108 314990
rect 676246 314785 676298 314791
rect 676244 314750 676246 314759
rect 676298 314750 676300 314759
rect 676244 314685 676300 314694
rect 672598 314045 672650 314051
rect 676054 314045 676106 314051
rect 672598 313987 672650 313993
rect 676052 314010 676054 314019
rect 676106 314010 676108 314019
rect 676052 313945 676108 313954
rect 676052 310606 676108 310615
rect 676052 310541 676108 310550
rect 676066 309685 676094 310541
rect 674326 309679 674378 309685
rect 674326 309621 674378 309627
rect 676054 309679 676106 309685
rect 676054 309621 676106 309627
rect 674230 308199 674282 308205
rect 674230 308141 674282 308147
rect 674134 306423 674186 306429
rect 674134 306365 674186 306371
rect 674038 305387 674090 305393
rect 674038 305329 674090 305335
rect 673942 302501 673994 302507
rect 673942 302443 673994 302449
rect 673954 286597 673982 302443
rect 674050 291629 674078 305329
rect 674146 292073 674174 306365
rect 674242 295995 674270 308141
rect 674230 295989 674282 295995
rect 674230 295931 674282 295937
rect 674338 294589 674366 309621
rect 676052 309570 676108 309579
rect 676052 309505 676108 309514
rect 676066 308205 676094 309505
rect 676054 308199 676106 308205
rect 676054 308141 676106 308147
rect 676052 307646 676108 307655
rect 676052 307581 676108 307590
rect 676066 305319 676094 307581
rect 676244 306906 676300 306915
rect 676244 306841 676300 306850
rect 676258 306429 676286 306841
rect 676246 306423 676298 306429
rect 676246 306365 676298 306371
rect 676244 306314 676300 306323
rect 676244 306249 676300 306258
rect 676258 305393 676286 306249
rect 676246 305387 676298 305393
rect 676246 305329 676298 305335
rect 674518 305313 674570 305319
rect 674518 305255 674570 305261
rect 676054 305313 676106 305319
rect 676054 305255 676106 305261
rect 674422 302427 674474 302433
rect 674422 302369 674474 302375
rect 674326 294583 674378 294589
rect 674326 294525 674378 294531
rect 674134 292067 674186 292073
rect 674134 292009 674186 292015
rect 674038 291623 674090 291629
rect 674038 291565 674090 291571
rect 674434 291111 674462 302369
rect 674530 295403 674558 305255
rect 676244 304834 676300 304843
rect 676244 304769 676300 304778
rect 676052 304094 676108 304103
rect 676052 304029 676108 304038
rect 676066 302507 676094 304029
rect 676054 302501 676106 302507
rect 676054 302443 676106 302449
rect 676258 302433 676286 304769
rect 679892 303354 679948 303363
rect 679892 303289 679948 303298
rect 679906 302919 679934 303289
rect 679892 302910 679948 302919
rect 679892 302845 679948 302854
rect 679796 302762 679852 302771
rect 679796 302697 679852 302706
rect 676246 302427 676298 302433
rect 676246 302369 676298 302375
rect 679810 302327 679838 302697
rect 679906 302581 679934 302845
rect 679894 302575 679946 302581
rect 679894 302517 679946 302523
rect 679796 302318 679852 302327
rect 679796 302253 679852 302262
rect 675382 295989 675434 295995
rect 675382 295931 675434 295937
rect 675394 295523 675422 295931
rect 674518 295397 674570 295403
rect 674518 295339 674570 295345
rect 675478 295397 675530 295403
rect 675478 295339 675530 295345
rect 675490 294890 675518 295339
rect 675382 294583 675434 294589
rect 675382 294525 675434 294531
rect 675394 294224 675422 294525
rect 675380 292846 675436 292855
rect 675380 292781 675436 292790
rect 675394 292374 675422 292781
rect 675478 292067 675530 292073
rect 675478 292009 675530 292015
rect 675490 291856 675518 292009
rect 675382 291623 675434 291629
rect 675382 291565 675434 291571
rect 675394 291190 675422 291565
rect 674422 291105 674474 291111
rect 674422 291047 674474 291053
rect 675382 291105 675434 291111
rect 675382 291047 675434 291053
rect 675394 290555 675422 291047
rect 675476 288554 675532 288563
rect 675476 288489 675532 288498
rect 675490 288082 675518 288489
rect 675668 287814 675724 287823
rect 675668 287749 675724 287758
rect 675682 287519 675710 287749
rect 675476 287370 675532 287379
rect 675476 287305 675532 287314
rect 675490 286898 675518 287305
rect 673942 286591 673994 286597
rect 673942 286533 673994 286539
rect 675382 286591 675434 286597
rect 675382 286533 675434 286539
rect 675394 286232 675422 286533
rect 675476 285298 675532 285307
rect 675476 285233 675532 285242
rect 675490 285048 675518 285233
rect 675380 283670 675436 283679
rect 675380 283605 675436 283614
rect 675394 283198 675422 283605
rect 675380 281894 675436 281903
rect 675380 281829 675436 281838
rect 675394 281348 675422 281829
rect 672502 270089 672554 270095
rect 676054 270089 676106 270095
rect 672502 270031 672554 270037
rect 676052 270054 676054 270063
rect 676106 270054 676108 270063
rect 676052 269989 676108 269998
rect 676246 269793 676298 269799
rect 676244 269758 676246 269767
rect 676298 269758 676300 269767
rect 676244 269693 676300 269702
rect 676246 269201 676298 269207
rect 676244 269166 676246 269175
rect 676298 269166 676300 269175
rect 676244 269101 676300 269110
rect 675668 264578 675724 264587
rect 675668 264513 675724 264522
rect 674614 261431 674666 261437
rect 674614 261373 674666 261379
rect 674038 256473 674090 256479
rect 674038 256415 674090 256421
rect 674050 241827 674078 256415
rect 674626 247081 674654 261373
rect 674710 259359 674762 259365
rect 674710 259301 674762 259307
rect 674614 247075 674666 247081
rect 674614 247017 674666 247023
rect 674722 243011 674750 259301
rect 675682 251225 675710 264513
rect 675764 262654 675820 262663
rect 675764 262589 675820 262598
rect 675778 251225 675806 262589
rect 676244 261914 676300 261923
rect 676244 261849 676300 261858
rect 676258 261437 676286 261849
rect 676246 261431 676298 261437
rect 676246 261373 676298 261379
rect 676052 259620 676108 259629
rect 676052 259555 676108 259564
rect 676066 259365 676094 259555
rect 676054 259359 676106 259365
rect 676054 259301 676106 259307
rect 676052 259102 676108 259111
rect 676052 259037 676108 259046
rect 676066 256479 676094 259037
rect 679700 258362 679756 258371
rect 679700 258297 679756 258306
rect 679714 257779 679742 258297
rect 679700 257770 679756 257779
rect 679700 257705 679756 257714
rect 685460 257770 685516 257779
rect 685460 257705 685516 257714
rect 676054 256473 676106 256479
rect 676054 256415 676106 256421
rect 679714 256405 679742 257705
rect 685474 257335 685502 257705
rect 685460 257326 685516 257335
rect 685460 257261 685516 257270
rect 679702 256399 679754 256405
rect 679702 256341 679754 256347
rect 675670 251219 675722 251225
rect 675670 251161 675722 251167
rect 675766 251219 675818 251225
rect 675766 251161 675818 251167
rect 675670 250997 675722 251003
rect 675670 250939 675722 250945
rect 675682 250523 675710 250939
rect 675766 250257 675818 250263
rect 675766 250199 675818 250205
rect 675778 249898 675806 250199
rect 675764 249630 675820 249639
rect 675764 249565 675820 249574
rect 675778 249232 675806 249565
rect 675668 247558 675724 247567
rect 675668 247493 675724 247502
rect 675682 247382 675710 247493
rect 675478 247075 675530 247081
rect 675478 247017 675530 247023
rect 675490 246864 675518 247017
rect 675764 246670 675820 246679
rect 675764 246605 675820 246614
rect 675778 246198 675806 246605
rect 675764 245930 675820 245939
rect 675764 245865 675820 245874
rect 675778 245532 675806 245865
rect 675476 243562 675532 243571
rect 675476 243497 675532 243506
rect 675490 243090 675518 243497
rect 674710 243005 674762 243011
rect 674710 242947 674762 242953
rect 675382 243005 675434 243011
rect 675382 242947 675434 242953
rect 675394 242498 675422 242947
rect 675284 241934 675340 241943
rect 675340 241878 675408 241889
rect 675284 241869 675408 241878
rect 675298 241861 675408 241869
rect 674038 241821 674090 241827
rect 674038 241763 674090 241769
rect 675286 241821 675338 241827
rect 675286 241763 675338 241769
rect 675298 241254 675326 241763
rect 675298 241226 675408 241254
rect 675476 240602 675532 240611
rect 675476 240537 675532 240546
rect 675490 240056 675518 240537
rect 675284 238234 675340 238243
rect 675340 238192 675408 238220
rect 675284 238169 675340 238178
rect 675380 236902 675436 236911
rect 675380 236837 675436 236846
rect 675394 236356 675422 236837
rect 676246 225097 676298 225103
rect 676244 225062 676246 225071
rect 676298 225062 676300 225071
rect 676244 224997 676300 225006
rect 676054 224357 676106 224363
rect 676052 224322 676054 224331
rect 676106 224322 676108 224331
rect 676052 224257 676108 224266
rect 676054 223839 676106 223845
rect 676052 223804 676054 223813
rect 676106 223804 676108 223813
rect 676052 223739 676108 223748
rect 675764 219290 675820 219299
rect 675764 219225 675820 219234
rect 674806 216439 674858 216445
rect 674806 216381 674858 216387
rect 674422 214959 674474 214965
rect 674422 214901 674474 214907
rect 674434 197057 674462 214901
rect 674518 213331 674570 213337
rect 674518 213273 674570 213279
rect 674422 197051 674474 197057
rect 674422 196993 674474 196999
rect 674530 196613 674558 213273
rect 674614 213257 674666 213263
rect 674614 213199 674666 213205
rect 674626 197649 674654 213199
rect 674710 213183 674762 213189
rect 674710 213125 674762 213131
rect 674722 200905 674750 213125
rect 674818 202089 674846 216381
rect 675778 206011 675806 219225
rect 676052 216922 676108 216931
rect 676052 216857 676108 216866
rect 676066 216445 676094 216857
rect 676054 216439 676106 216445
rect 676054 216381 676106 216387
rect 676052 215368 676108 215377
rect 676052 215303 676108 215312
rect 676066 214965 676094 215303
rect 676054 214959 676106 214965
rect 676054 214901 676106 214907
rect 676052 214850 676108 214859
rect 676052 214785 676108 214794
rect 675956 213888 676012 213897
rect 675956 213823 676012 213832
rect 675970 213337 675998 213823
rect 675958 213331 676010 213337
rect 675958 213273 676010 213279
rect 676066 213189 676094 214785
rect 676244 214258 676300 214267
rect 676244 214193 676300 214202
rect 676258 213263 676286 214193
rect 679796 213518 679852 213527
rect 679796 213453 679852 213462
rect 676246 213257 676298 213263
rect 676246 213199 676298 213205
rect 676054 213183 676106 213189
rect 676054 213125 676106 213131
rect 679810 212639 679838 213453
rect 679796 212630 679852 212639
rect 679796 212565 679852 212574
rect 685460 212630 685516 212639
rect 685460 212565 685516 212574
rect 679810 210303 679838 212565
rect 685474 212195 685502 212565
rect 685460 212186 685516 212195
rect 685460 212121 685516 212130
rect 679798 210297 679850 210303
rect 679798 210239 679850 210245
rect 675766 206005 675818 206011
rect 675766 205947 675818 205953
rect 675766 205783 675818 205789
rect 675766 205725 675818 205731
rect 675778 205350 675806 205725
rect 675764 205082 675820 205091
rect 675764 205017 675820 205026
rect 675778 204684 675806 205017
rect 675476 204342 675532 204351
rect 675476 204277 675532 204286
rect 675490 204018 675518 204277
rect 675764 202714 675820 202723
rect 675764 202649 675820 202658
rect 675778 202168 675806 202649
rect 674806 202083 674858 202089
rect 674806 202025 674858 202031
rect 675478 202083 675530 202089
rect 675478 202025 675530 202031
rect 675490 201650 675518 202025
rect 675764 201382 675820 201391
rect 675764 201317 675820 201326
rect 675778 200984 675806 201317
rect 674710 200899 674762 200905
rect 674710 200841 674762 200847
rect 675382 200899 675434 200905
rect 675382 200841 675434 200847
rect 675394 200355 675422 200841
rect 675476 198422 675532 198431
rect 675476 198357 675532 198366
rect 675490 197876 675518 198357
rect 674614 197643 674666 197649
rect 674614 197585 674666 197591
rect 675382 197643 675434 197649
rect 675382 197585 675434 197591
rect 675394 197319 675422 197585
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 674518 196607 674570 196613
rect 674518 196549 674570 196555
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675476 195314 675532 195323
rect 675476 195249 675532 195258
rect 675490 194842 675518 195249
rect 675380 193538 675436 193547
rect 675380 193473 675436 193482
rect 675394 192992 675422 193473
rect 675380 191614 675436 191623
rect 675380 191549 675436 191558
rect 675394 191142 675422 191549
rect 676244 179626 676300 179635
rect 676244 179561 676300 179570
rect 676054 179365 676106 179371
rect 676052 179330 676054 179339
rect 676106 179330 676108 179339
rect 676052 179265 676108 179274
rect 676054 178847 676106 178853
rect 676052 178812 676054 178821
rect 676106 178812 676108 178821
rect 676052 178747 676108 178756
rect 676258 178705 676286 179561
rect 676246 178699 676298 178705
rect 676246 178641 676298 178647
rect 676052 175408 676108 175417
rect 676052 175343 676108 175352
rect 675380 174298 675436 174307
rect 675380 174233 675436 174242
rect 674518 172927 674570 172933
rect 674518 172869 674570 172875
rect 674530 159465 674558 172869
rect 674806 172853 674858 172859
rect 674806 172795 674858 172801
rect 674614 170041 674666 170047
rect 674614 169983 674666 169989
rect 674518 159459 674570 159465
rect 674518 159401 674570 159407
rect 674626 156357 674654 169983
rect 674710 169967 674762 169973
rect 674710 169909 674762 169915
rect 674722 156949 674750 169909
rect 674818 157763 674846 172795
rect 675190 167081 675242 167087
rect 675190 167023 675242 167029
rect 675202 158767 675230 167023
rect 675394 161019 675422 174233
rect 676066 172933 676094 175343
rect 676244 173706 676300 173715
rect 676244 173641 676300 173650
rect 676054 172927 676106 172933
rect 676054 172869 676106 172875
rect 676258 172859 676286 173641
rect 676246 172853 676298 172859
rect 676246 172795 676298 172801
rect 675476 172374 675532 172383
rect 675476 172309 675532 172318
rect 675490 167054 675518 172309
rect 676052 171930 676108 171939
rect 676052 171865 676108 171874
rect 675956 171338 676012 171347
rect 675956 171273 676012 171282
rect 675970 170047 675998 171273
rect 675958 170041 676010 170047
rect 675958 169983 676010 169989
rect 676066 169973 676094 171865
rect 676054 169967 676106 169973
rect 676054 169909 676106 169915
rect 676052 169858 676108 169867
rect 676052 169793 676108 169802
rect 676066 167087 676094 169793
rect 676244 168082 676300 168091
rect 676244 168017 676300 168026
rect 676148 167638 676204 167647
rect 676148 167573 676204 167582
rect 676162 167161 676190 167573
rect 676258 167383 676286 168017
rect 676246 167377 676298 167383
rect 676246 167319 676298 167325
rect 676246 167229 676298 167235
rect 676244 167194 676246 167203
rect 676298 167194 676300 167203
rect 676150 167155 676202 167161
rect 676244 167129 676300 167138
rect 676150 167097 676202 167103
rect 676054 167081 676106 167087
rect 675490 167026 675710 167054
rect 675682 161019 675710 167026
rect 676054 167023 676106 167029
rect 675382 161013 675434 161019
rect 675382 160955 675434 160961
rect 675670 161013 675722 161019
rect 675670 160955 675722 160961
rect 675382 160791 675434 160797
rect 675382 160733 675434 160739
rect 675394 160323 675422 160733
rect 675670 160051 675722 160057
rect 675670 159993 675722 159999
rect 675682 159692 675710 159993
rect 675382 159459 675434 159465
rect 675382 159401 675434 159407
rect 675394 159026 675422 159401
rect 675188 158758 675244 158767
rect 675188 158693 675244 158702
rect 675188 158462 675244 158471
rect 675188 158397 675244 158406
rect 674806 157757 674858 157763
rect 674806 157699 674858 157705
rect 674710 156943 674762 156949
rect 674710 156885 674762 156891
rect 674614 156351 674666 156357
rect 674614 156293 674666 156299
rect 675202 155913 675230 158397
rect 675478 157757 675530 157763
rect 675478 157699 675530 157705
rect 675490 157176 675518 157699
rect 675478 156943 675530 156949
rect 675478 156885 675530 156891
rect 675490 156658 675518 156885
rect 675382 156351 675434 156357
rect 675382 156293 675434 156299
rect 675394 155992 675422 156293
rect 675190 155907 675242 155913
rect 675190 155849 675242 155855
rect 675382 155907 675434 155913
rect 675382 155849 675434 155855
rect 675394 155355 675422 155849
rect 675476 153430 675532 153439
rect 675476 153365 675532 153374
rect 675490 152884 675518 153365
rect 675380 152542 675436 152551
rect 675380 152477 675436 152486
rect 675394 152292 675422 152477
rect 675476 151950 675532 151959
rect 675476 151885 675532 151894
rect 675490 151700 675518 151885
rect 675668 151358 675724 151367
rect 675668 151293 675724 151302
rect 675682 151034 675710 151293
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149850 675518 150257
rect 675476 148546 675532 148555
rect 675476 148481 675532 148490
rect 675490 148000 675518 148481
rect 675380 146622 675436 146631
rect 675380 146557 675436 146566
rect 675394 146150 675422 146557
rect 676148 134486 676204 134495
rect 676148 134421 676204 134430
rect 672406 134373 672458 134379
rect 672406 134315 672458 134321
rect 676052 132710 676108 132719
rect 676162 132677 676190 134421
rect 676246 134373 676298 134379
rect 676244 134338 676246 134347
rect 676298 134338 676300 134347
rect 676244 134273 676300 134282
rect 676244 133450 676300 133459
rect 676244 133385 676300 133394
rect 676258 132825 676286 133385
rect 676246 132819 676298 132825
rect 676246 132761 676298 132767
rect 676052 132645 676108 132654
rect 676150 132671 676202 132677
rect 676066 132529 676094 132645
rect 676150 132613 676202 132619
rect 676054 132523 676106 132529
rect 676054 132465 676106 132471
rect 676244 131378 676300 131387
rect 676244 131313 676300 131322
rect 676052 130638 676108 130647
rect 676052 130573 676108 130582
rect 676066 129865 676094 130573
rect 676054 129859 676106 129865
rect 676054 129801 676106 129807
rect 676258 129643 676286 131313
rect 676246 129637 676298 129643
rect 676246 129579 676298 129585
rect 675476 129158 675532 129167
rect 675476 129093 675532 129102
rect 674518 126751 674570 126757
rect 674518 126693 674570 126699
rect 674230 124753 674282 124759
rect 674230 124695 674282 124701
rect 674038 124013 674090 124019
rect 674038 123955 674090 123961
rect 674050 107369 674078 123955
rect 674134 123939 674186 123945
rect 674134 123881 674186 123887
rect 674146 110699 674174 123881
rect 674242 111217 674270 124695
rect 674422 124087 674474 124093
rect 674422 124029 674474 124035
rect 674434 111735 674462 124029
rect 674530 114843 674558 126693
rect 674614 121053 674666 121059
rect 674614 120995 674666 121001
rect 674518 114837 674570 114843
rect 674518 114779 674570 114785
rect 674422 111729 674474 111735
rect 674422 111671 674474 111677
rect 674230 111211 674282 111217
rect 674230 111153 674282 111159
rect 674134 110693 674186 110699
rect 674134 110635 674186 110641
rect 674038 107363 674090 107369
rect 674038 107305 674090 107311
rect 669524 106366 669580 106375
rect 669524 106301 669580 106310
rect 674626 106185 674654 120995
rect 675490 115805 675518 129093
rect 676052 127234 676108 127243
rect 676052 127169 676108 127178
rect 676066 126757 676094 127169
rect 676054 126751 676106 126757
rect 676054 126693 676106 126699
rect 676244 126494 676300 126503
rect 676244 126429 676300 126438
rect 676052 126124 676108 126133
rect 676052 126059 676108 126068
rect 676066 124759 676094 126059
rect 676054 124753 676106 124759
rect 676054 124695 676106 124701
rect 676052 124644 676108 124653
rect 676052 124579 676108 124588
rect 675956 124274 676012 124283
rect 675956 124209 676012 124218
rect 675970 124019 675998 124209
rect 675958 124013 676010 124019
rect 675958 123955 676010 123961
rect 676066 123945 676094 124579
rect 676258 124093 676286 126429
rect 676246 124087 676298 124093
rect 676246 124029 676298 124035
rect 676054 123939 676106 123945
rect 676054 123881 676106 123887
rect 676052 123682 676108 123691
rect 676052 123617 676108 123626
rect 676066 121059 676094 123617
rect 676340 122942 676396 122951
rect 676340 122877 676396 122886
rect 676148 122498 676204 122507
rect 676148 122433 676204 122442
rect 676162 121207 676190 122433
rect 676244 121906 676300 121915
rect 676244 121841 676300 121850
rect 676150 121201 676202 121207
rect 676150 121143 676202 121149
rect 676258 121133 676286 121841
rect 676354 121281 676382 122877
rect 676342 121275 676394 121281
rect 676342 121217 676394 121223
rect 676246 121127 676298 121133
rect 676246 121069 676298 121075
rect 676054 121053 676106 121059
rect 676054 120995 676106 121001
rect 675478 115799 675530 115805
rect 675478 115741 675530 115747
rect 675478 115577 675530 115583
rect 675478 115519 675530 115525
rect 675490 115144 675518 115519
rect 675382 114837 675434 114843
rect 675382 114779 675434 114785
rect 675394 114478 675422 114779
rect 675380 114358 675436 114367
rect 675380 114293 675436 114302
rect 675394 113812 675422 114293
rect 675380 112286 675436 112295
rect 675380 112221 675436 112230
rect 675394 111995 675422 112221
rect 675382 111729 675434 111735
rect 675382 111671 675434 111677
rect 675394 111444 675422 111671
rect 675382 111211 675434 111217
rect 675382 111153 675434 111159
rect 675394 110778 675422 111153
rect 675382 110693 675434 110699
rect 675382 110635 675434 110641
rect 675394 110155 675422 110635
rect 675476 108142 675532 108151
rect 675476 108077 675532 108086
rect 675490 107670 675518 108077
rect 675382 107363 675434 107369
rect 675382 107305 675434 107311
rect 675394 107119 675422 107305
rect 675394 106375 675422 106486
rect 675380 106366 675436 106375
rect 675380 106301 675436 106310
rect 674614 106179 674666 106185
rect 674614 106121 674666 106127
rect 675382 106179 675434 106185
rect 675382 106121 675434 106127
rect 675394 105820 675422 106121
rect 668180 105330 668236 105339
rect 668180 105265 668236 105274
rect 665300 105182 665356 105191
rect 665300 105117 665356 105126
rect 647924 104146 647980 104155
rect 647924 104081 647980 104090
rect 647938 103965 647966 104081
rect 647926 103959 647978 103965
rect 647926 103901 647978 103907
rect 661174 103959 661226 103965
rect 661174 103901 661226 103907
rect 657526 103737 657578 103743
rect 657526 103679 657578 103685
rect 652438 102109 652490 102115
rect 652438 102051 652490 102057
rect 647924 99706 647980 99715
rect 647924 99641 647980 99650
rect 647938 97971 647966 99641
rect 647926 97965 647978 97971
rect 647926 97907 647978 97913
rect 647732 94082 647788 94091
rect 647732 94017 647788 94026
rect 647158 92193 647210 92199
rect 647158 92135 647210 92141
rect 647062 87087 647114 87093
rect 647062 87029 647114 87035
rect 646966 77763 647018 77769
rect 646966 77705 647018 77711
rect 647062 74951 647114 74957
rect 647062 74893 647114 74899
rect 646868 68626 646924 68635
rect 646868 68561 646924 68570
rect 647074 60347 647102 74893
rect 647170 71891 647198 92135
rect 647746 81617 647774 94017
rect 649558 93599 649610 93605
rect 649558 93541 649610 93547
rect 647828 92750 647884 92759
rect 647828 92685 647884 92694
rect 647842 81839 647870 92685
rect 647926 87309 647978 87315
rect 647926 87251 647978 87257
rect 647938 87135 647966 87251
rect 647924 87126 647980 87135
rect 647924 87061 647980 87070
rect 649570 83689 649598 93541
rect 650902 87531 650954 87537
rect 650902 87473 650954 87479
rect 650914 86247 650942 87473
rect 650900 86238 650956 86247
rect 650900 86173 650956 86182
rect 652340 85350 652396 85359
rect 652340 85285 652396 85294
rect 651764 84314 651820 84323
rect 651764 84249 651820 84258
rect 649558 83683 649610 83689
rect 649558 83625 649610 83631
rect 651778 83615 651806 84249
rect 651766 83609 651818 83615
rect 651766 83551 651818 83557
rect 652244 83426 652300 83435
rect 652244 83361 652300 83370
rect 647924 82686 647980 82695
rect 647924 82621 647980 82630
rect 647938 81913 647966 82621
rect 647926 81907 647978 81913
rect 647926 81849 647978 81855
rect 647830 81833 647882 81839
rect 647830 81775 647882 81781
rect 647734 81611 647786 81617
rect 647734 81553 647786 81559
rect 647924 81058 647980 81067
rect 647924 80993 647980 81002
rect 647938 80803 647966 80993
rect 647926 80797 647978 80803
rect 647926 80739 647978 80745
rect 647926 77541 647978 77547
rect 647924 77506 647926 77515
rect 647978 77506 647980 77515
rect 647924 77441 647980 77450
rect 647924 73658 647980 73667
rect 647924 73593 647980 73602
rect 647938 72145 647966 73593
rect 647926 72139 647978 72145
rect 647926 72081 647978 72087
rect 647156 71882 647212 71891
rect 647156 71817 647212 71826
rect 647924 69662 647980 69671
rect 647924 69597 647926 69606
rect 647978 69597 647980 69606
rect 647926 69565 647978 69571
rect 647924 64186 647980 64195
rect 647924 64121 647980 64130
rect 647938 63635 647966 64121
rect 647926 63629 647978 63635
rect 647926 63571 647978 63577
rect 647924 62262 647980 62271
rect 647924 62197 647980 62206
rect 647938 61045 647966 62197
rect 647926 61039 647978 61045
rect 647926 60981 647978 60987
rect 647060 60338 647116 60347
rect 647060 60273 647116 60282
rect 652258 59121 652286 83361
rect 652354 66225 652382 85285
rect 652450 82695 652478 102051
rect 653686 95967 653738 95973
rect 653686 95909 653738 95915
rect 653698 86987 653726 95909
rect 657538 88000 657566 103679
rect 660694 92415 660746 92421
rect 660694 92357 660746 92363
rect 659830 92267 659882 92273
rect 659830 92209 659882 92215
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 657538 87972 657792 88000
rect 658882 87986 658910 92135
rect 659348 90826 659404 90835
rect 659348 90761 659404 90770
rect 659362 88000 659390 90761
rect 659842 88000 659870 92209
rect 659362 87972 659616 88000
rect 659842 87972 660144 88000
rect 660706 87986 660734 92357
rect 661186 88000 661214 103901
rect 662518 97965 662570 97971
rect 662518 97907 662570 97913
rect 661750 92341 661802 92347
rect 661750 92283 661802 92289
rect 661762 88000 661790 92283
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 97907
rect 668194 93605 668222 105265
rect 675380 105182 675436 105191
rect 675380 105117 675436 105126
rect 675394 104636 675422 105117
rect 675668 103258 675724 103267
rect 675668 103193 675724 103202
rect 675682 102786 675710 103193
rect 675380 101482 675436 101491
rect 675380 101417 675436 101426
rect 675394 100936 675422 101417
rect 668182 93599 668234 93605
rect 668182 93541 668234 93547
rect 663094 92711 663146 92717
rect 663094 92653 663146 92659
rect 663106 87986 663134 92653
rect 658006 87309 658058 87315
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 653684 86978 653740 86987
rect 653684 86913 653740 86922
rect 663298 86395 663326 87029
rect 663284 86386 663340 86395
rect 663284 86321 663340 86330
rect 663284 84758 663340 84767
rect 663202 84716 663284 84744
rect 657046 84201 657098 84207
rect 657046 84143 657098 84149
rect 652436 82686 652492 82695
rect 652436 82621 652492 82630
rect 657058 81691 657086 84143
rect 657046 81685 657098 81691
rect 657046 81627 657098 81633
rect 658582 81685 658634 81691
rect 662420 81650 662476 81659
rect 658634 81633 658896 81636
rect 658582 81627 658896 81633
rect 658594 81608 658896 81627
rect 662420 81585 662422 81594
rect 662474 81585 662476 81594
rect 662422 81553 662474 81559
rect 656962 81016 657216 81044
rect 657538 81016 657792 81044
rect 656962 77547 656990 81016
rect 656950 77541 657002 77547
rect 656950 77483 657002 77489
rect 657538 76141 657566 81016
rect 658306 77769 658334 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658294 77763 658346 77769
rect 658294 77705 658346 77711
rect 659458 77695 659486 80665
rect 659446 77689 659498 77695
rect 659446 77631 659498 77637
rect 657526 76135 657578 76141
rect 657526 76077 657578 76083
rect 660130 74957 660158 81030
rect 660118 74951 660170 74957
rect 660118 74893 660170 74899
rect 660706 72145 660734 81030
rect 661440 81016 661502 81044
rect 660694 72139 660746 72145
rect 660694 72081 660746 72087
rect 661474 69629 661502 81016
rect 661762 81016 662016 81044
rect 661762 77621 661790 81016
rect 662530 80803 662558 81030
rect 662518 80797 662570 80803
rect 662518 80739 662570 80745
rect 661750 77615 661802 77621
rect 661750 77557 661802 77563
rect 661462 69623 661514 69629
rect 661462 69565 661514 69571
rect 652342 66219 652394 66225
rect 652342 66161 652394 66167
rect 663202 63635 663230 84716
rect 663284 84693 663340 84702
rect 663476 84018 663532 84027
rect 663476 83953 663532 83962
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663190 63629 663242 63635
rect 663190 63571 663242 63577
rect 663490 61045 663518 83953
rect 663478 61039 663530 61045
rect 663478 60981 663530 60987
rect 652246 59115 652298 59121
rect 652246 59057 652298 59063
rect 646772 57082 646828 57091
rect 646772 57017 646828 57026
rect 646484 54714 646540 54723
rect 646484 54649 646540 54658
rect 633622 43279 633674 43285
rect 633622 43221 633674 43227
rect 640726 43279 640778 43285
rect 640726 43221 640778 43227
rect 545204 40654 545260 40663
rect 545204 40589 545260 40598
rect 633634 40515 633662 43221
rect 633620 40506 633676 40515
rect 633620 40441 633676 40450
rect 475606 37359 475658 37365
rect 475606 37301 475658 37307
rect 514006 37359 514058 37365
rect 514006 37301 514058 37307
<< via2 >>
rect 148532 1016214 148588 1016270
rect 250484 1016214 250540 1016270
rect 353396 1016214 353452 1016270
rect 146612 1007926 146668 1007982
rect 148532 1007926 148588 1007982
rect 102452 1006167 102508 1006206
rect 102452 1006150 102454 1006167
rect 102454 1006150 102506 1006167
rect 102506 1006150 102508 1006167
rect 85940 995790 85996 995846
rect 81620 995642 81676 995698
rect 81044 995494 81100 995550
rect 84500 994014 84556 994070
rect 92564 995790 92620 995846
rect 92660 995642 92716 995698
rect 101012 1005871 101068 1005910
rect 101012 1005854 101014 1005871
rect 101014 1005854 101066 1005871
rect 101066 1005854 101068 1005871
rect 109940 1005597 109942 1005614
rect 109942 1005597 109994 1005614
rect 109994 1005597 109996 1005614
rect 92852 995494 92908 995550
rect 88724 993866 88780 993922
rect 80180 993718 80236 993774
rect 42164 968706 42220 968762
rect 41780 967078 41836 967134
rect 41780 965006 41836 965062
rect 41780 963970 41836 964026
rect 41780 963378 41836 963434
rect 41780 962786 41836 962842
rect 41780 962194 41836 962250
rect 41780 959530 41836 959586
rect 41780 959086 41836 959142
rect 41876 957754 41932 957810
rect 42260 957458 42316 957514
rect 42260 956274 42316 956330
rect 34484 945026 34540 945082
rect 39764 943990 39820 944046
rect 41780 943807 41782 943824
rect 41782 943807 41834 943824
rect 41834 943807 41836 943824
rect 41780 943768 41836 943807
rect 41588 943585 41590 943602
rect 41590 943585 41642 943602
rect 41642 943585 41644 943602
rect 41588 943546 41644 943585
rect 40436 942658 40492 942714
rect 40244 941622 40300 941678
rect 40340 941030 40396 941086
rect 38804 937626 38860 937682
rect 28820 932594 28876 932650
rect 28820 932150 28876 932206
rect 39956 816266 40012 816322
rect 41684 942066 41740 942122
rect 41588 940586 41644 940642
rect 41588 932167 41644 932206
rect 41588 932150 41590 932167
rect 41590 932150 41642 932167
rect 41642 932150 41644 932167
rect 42260 939254 42316 939310
rect 41588 819265 41590 819282
rect 41590 819265 41642 819282
rect 41642 819265 41644 819282
rect 41588 819226 41644 819265
rect 41780 818525 41782 818542
rect 41782 818525 41834 818542
rect 41834 818525 41836 818542
rect 41780 818486 41836 818525
rect 41780 817894 41836 817950
rect 40436 817746 40492 817802
rect 41780 817023 41836 817062
rect 41780 817006 41782 817023
rect 41782 817006 41834 817023
rect 41834 817006 41836 817023
rect 40340 814786 40396 814842
rect 42068 814564 42124 814620
rect 41780 814046 41836 814102
rect 34388 813306 34444 813362
rect 23060 806794 23116 806850
rect 23060 806350 23116 806406
rect 41588 812862 41644 812918
rect 41876 811974 41932 812030
rect 34484 811382 34540 811438
rect 34388 802058 34444 802114
rect 41492 810642 41548 810698
rect 34484 801762 34540 801818
rect 41780 810050 41836 810106
rect 41684 809310 41740 809366
rect 41588 807830 41644 807886
rect 41588 806389 41590 806406
rect 41590 806389 41642 806406
rect 41642 806389 41644 806406
rect 41588 806350 41644 806389
rect 41684 800550 41740 800606
rect 41780 800282 41836 800338
rect 41972 811012 42028 811068
rect 42356 812566 42412 812622
rect 41972 808570 42028 808626
rect 41972 800282 42028 800338
rect 42164 809014 42220 809070
rect 42452 797470 42508 797526
rect 41780 796286 41836 796342
rect 41876 794214 41932 794270
rect 42740 790514 42796 790570
rect 42452 789182 42508 789238
rect 41588 776049 41590 776066
rect 41590 776049 41642 776066
rect 41642 776049 41644 776066
rect 41588 776010 41644 776049
rect 41780 775309 41782 775326
rect 41782 775309 41834 775326
rect 41834 775309 41836 775326
rect 41780 775270 41836 775309
rect 41780 774791 41782 774808
rect 41782 774791 41834 774808
rect 41834 774791 41836 774808
rect 41780 774752 41836 774791
rect 41588 774569 41590 774586
rect 41590 774569 41642 774586
rect 41642 774569 41644 774586
rect 41588 774530 41644 774569
rect 41588 773659 41644 773698
rect 41588 773642 41590 773659
rect 41590 773642 41642 773659
rect 41642 773642 41644 773659
rect 42164 773198 42220 773254
rect 42068 772310 42124 772366
rect 42068 771866 42124 771922
rect 41780 771348 41836 771404
rect 40436 770534 40492 770590
rect 33044 770090 33100 770146
rect 23060 763578 23116 763634
rect 23060 763134 23116 763190
rect 40340 768610 40396 768666
rect 33236 768166 33292 768222
rect 33236 758190 33292 758246
rect 33044 758042 33100 758098
rect 41780 769868 41836 769924
rect 41780 769350 41836 769406
rect 41684 766686 41740 766742
rect 41588 766111 41644 766150
rect 41588 766094 41590 766111
rect 41590 766094 41642 766111
rect 41642 766094 41644 766111
rect 41492 765206 41548 765262
rect 41588 763134 41644 763190
rect 41876 767870 41932 767926
rect 41972 767278 42028 767334
rect 41876 764836 41932 764892
rect 42164 765798 42220 765854
rect 42740 756474 42796 756530
rect 42932 757066 42988 757122
rect 42068 750998 42124 751054
rect 42644 748630 42700 748686
rect 42740 748482 42796 748538
rect 43028 749814 43084 749870
rect 41588 732833 41590 732850
rect 41590 732833 41642 732850
rect 41642 732833 41644 732850
rect 41588 732794 41644 732833
rect 41588 731797 41590 731814
rect 41590 731797 41642 731814
rect 41642 731797 41644 731814
rect 41588 731758 41644 731797
rect 41588 731353 41590 731370
rect 41590 731353 41642 731370
rect 41642 731353 41644 731370
rect 41588 731314 41644 731353
rect 41588 730443 41644 730482
rect 41588 730426 41590 730443
rect 41590 730426 41642 730443
rect 41642 730426 41644 730443
rect 41780 732093 41782 732110
rect 41782 732093 41834 732110
rect 41834 732093 41836 732110
rect 41780 732054 41836 732093
rect 42068 730056 42124 730112
rect 41684 729390 41740 729446
rect 41684 727910 41740 727966
rect 34388 726874 34444 726930
rect 23060 720362 23116 720418
rect 23060 719770 23116 719826
rect 41492 726430 41548 726486
rect 34484 724950 34540 725006
rect 34388 716958 34444 717014
rect 34484 716514 34540 716570
rect 41588 723914 41644 723970
rect 41588 721990 41644 722046
rect 41972 727614 42028 727670
rect 41876 725542 41932 725598
rect 41780 723618 41836 723674
rect 41780 723191 41836 723230
rect 41780 723174 41782 723191
rect 41782 723174 41834 723191
rect 41834 723174 41836 723191
rect 41780 721102 41836 721158
rect 41780 720179 41782 720196
rect 41782 720179 41834 720196
rect 41834 720179 41836 720196
rect 41780 720140 41836 720179
rect 41780 713998 41836 714054
rect 42068 726134 42124 726190
rect 41972 713850 42028 713906
rect 42164 724654 42220 724710
rect 42452 721546 42508 721602
rect 42164 713850 42220 713906
rect 42068 711630 42124 711686
rect 42452 706006 42508 706062
rect 42452 703638 42508 703694
rect 42932 709706 42988 709762
rect 43124 707190 43180 707246
rect 42836 703342 42892 703398
rect 41780 689469 41782 689486
rect 41782 689469 41834 689486
rect 41834 689469 41836 689486
rect 41780 689430 41836 689469
rect 41780 688877 41782 688894
rect 41782 688877 41834 688894
rect 41834 688877 41836 688894
rect 41780 688838 41836 688877
rect 41588 688581 41590 688598
rect 41590 688581 41642 688598
rect 41642 688581 41644 688598
rect 41588 688542 41644 688581
rect 41588 688137 41590 688154
rect 41590 688137 41642 688154
rect 41642 688137 41644 688154
rect 41588 688098 41644 688137
rect 41588 687227 41644 687266
rect 41588 687210 41590 687227
rect 41590 687210 41642 687227
rect 41642 687210 41644 687227
rect 41876 686914 41932 686970
rect 41780 685917 41782 685934
rect 41782 685917 41834 685934
rect 41834 685917 41836 685934
rect 41780 685878 41836 685917
rect 41780 684990 41836 685046
rect 41588 684250 41644 684306
rect 34388 683658 34444 683714
rect 23060 677146 23116 677202
rect 23060 676702 23116 676758
rect 41684 683214 41740 683270
rect 34484 681734 34540 681790
rect 34388 672558 34444 672614
rect 41588 680271 41644 680310
rect 41588 680254 41590 680271
rect 41590 680254 41642 680271
rect 41642 680254 41644 680271
rect 34484 672410 34540 672466
rect 41588 679235 41644 679274
rect 41588 679218 41590 679235
rect 41590 679218 41642 679235
rect 41642 679218 41644 679235
rect 42452 682918 42508 682974
rect 41876 682326 41932 682382
rect 41588 678774 41644 678830
rect 41780 678495 41836 678534
rect 41780 678478 41782 678495
rect 41782 678478 41834 678495
rect 41834 678478 41836 678495
rect 41780 677886 41836 677942
rect 41780 676941 41836 676980
rect 41780 676924 41782 676941
rect 41782 676924 41834 676941
rect 41834 676924 41836 676941
rect 41780 670634 41836 670690
rect 42164 681438 42220 681494
rect 42068 680846 42124 680902
rect 41972 679958 42028 680014
rect 42068 670634 42124 670690
rect 42452 670042 42508 670098
rect 42164 666638 42220 666694
rect 41780 663382 41836 663438
rect 42836 665158 42892 665214
rect 42836 660274 42892 660330
rect 43028 660866 43084 660922
rect 41780 646253 41782 646270
rect 41782 646253 41834 646270
rect 41834 646253 41836 646270
rect 41780 646214 41836 646253
rect 41780 645735 41782 645752
rect 41782 645735 41834 645752
rect 41834 645735 41836 645752
rect 41780 645696 41836 645735
rect 41588 645365 41590 645382
rect 41590 645365 41642 645382
rect 41642 645365 41644 645382
rect 41588 645326 41644 645365
rect 41780 644773 41782 644790
rect 41782 644773 41834 644790
rect 41834 644773 41836 644790
rect 41780 644734 41836 644773
rect 43796 644142 43852 644198
rect 43316 643698 43372 643754
rect 25844 642366 25900 642422
rect 23156 633930 23212 633986
rect 23156 633486 23212 633542
rect 41588 641478 41644 641534
rect 34388 640442 34444 640498
rect 41492 639998 41548 640054
rect 34484 638518 34540 638574
rect 34484 629046 34540 629102
rect 34388 627862 34444 627918
rect 41492 627862 41548 627918
rect 41780 641182 41836 641238
rect 41876 639702 41932 639758
rect 41780 639110 41836 639166
rect 41684 637055 41740 637094
rect 41684 637038 41686 637055
rect 41686 637038 41738 637055
rect 41738 637038 41740 637055
rect 41684 634983 41740 635022
rect 41684 634966 41686 634983
rect 41686 634966 41738 634983
rect 41738 634966 41740 634983
rect 41684 634522 41740 634578
rect 41684 633947 41740 633986
rect 41684 633930 41686 633947
rect 41686 633930 41738 633947
rect 41738 633930 41740 633947
rect 41588 627714 41644 627770
rect 42164 638222 42220 638278
rect 41972 637630 42028 637686
rect 42068 636150 42124 636206
rect 42932 636742 42988 636798
rect 42836 628010 42892 628066
rect 42164 627418 42220 627474
rect 42164 622090 42220 622146
rect 42836 621498 42892 621554
rect 41780 620906 41836 620962
rect 41780 616022 41836 616078
rect 42932 620166 42988 620222
rect 43028 618834 43084 618890
rect 42932 616466 42988 616522
rect 41780 603037 41782 603054
rect 41782 603037 41834 603054
rect 41834 603037 41836 603054
rect 41780 602998 41836 603037
rect 41588 602741 41590 602758
rect 41590 602741 41642 602758
rect 41642 602741 41644 602758
rect 41588 602702 41644 602741
rect 41588 602149 41590 602166
rect 41590 602149 41642 602166
rect 41642 602149 41644 602166
rect 41588 602110 41644 602149
rect 41780 601557 41782 601574
rect 41782 601557 41834 601574
rect 41834 601557 41836 601574
rect 41780 601518 41836 601557
rect 41780 601017 41836 601056
rect 41780 601000 41782 601017
rect 41782 601000 41834 601017
rect 41834 601000 41836 601017
rect 41588 599907 41644 599946
rect 41588 599890 41590 599907
rect 41590 599890 41642 599907
rect 41642 599890 41644 599907
rect 41780 599019 41836 599058
rect 41780 599002 41782 599019
rect 41782 599002 41834 599019
rect 41834 599002 41836 599019
rect 41492 598262 41548 598318
rect 34388 597226 34444 597282
rect 23060 590714 23116 590770
rect 23060 590270 23116 590326
rect 34484 595302 34540 595358
rect 34388 585526 34444 585582
rect 34484 585378 34540 585434
rect 41588 597818 41644 597874
rect 42068 597078 42124 597134
rect 41684 596338 41740 596394
rect 41588 591306 41644 591362
rect 41588 590731 41644 590770
rect 41588 590714 41590 590731
rect 41590 590714 41642 590731
rect 41642 590714 41644 590731
rect 41876 595968 41932 596024
rect 41780 594118 41836 594174
rect 41780 593543 41836 593582
rect 41780 593526 41782 593543
rect 41782 593526 41834 593543
rect 41834 593526 41836 593543
rect 41780 592581 41836 592620
rect 41780 592564 41782 592581
rect 41782 592564 41834 592581
rect 41834 592564 41836 592581
rect 41780 592046 41836 592102
rect 41492 584498 41548 584554
rect 41972 595006 42028 595062
rect 42164 594414 42220 594470
rect 42068 584202 42124 584258
rect 42452 592934 42508 592990
rect 42836 578726 42892 578782
rect 42356 574434 42412 574490
rect 42740 573990 42796 574046
rect 41780 559821 41782 559838
rect 41782 559821 41834 559838
rect 41834 559821 41836 559838
rect 41780 559782 41836 559821
rect 42932 577542 42988 577598
rect 42356 559338 42412 559394
rect 41780 558785 41782 558802
rect 41782 558785 41834 558802
rect 41834 558785 41836 558802
rect 41780 558746 41836 558785
rect 44372 619130 44428 619186
rect 41780 558341 41782 558358
rect 41782 558341 41834 558358
rect 41834 558341 41836 558358
rect 41780 558302 41836 558341
rect 41780 557875 41836 557914
rect 41780 557858 41782 557875
rect 41782 557858 41834 557875
rect 41834 557858 41836 557875
rect 42260 555342 42316 555398
rect 41588 554602 41644 554658
rect 34388 554010 34444 554066
rect 23060 547498 23116 547554
rect 23060 547054 23116 547110
rect 41684 554010 41740 554066
rect 34484 552086 34540 552142
rect 41492 551642 41548 551698
rect 41396 549126 41452 549182
rect 34484 541578 34540 541634
rect 34388 541430 34444 541486
rect 41588 550179 41644 550218
rect 41588 550162 41590 550179
rect 41590 550162 41642 550179
rect 41642 550162 41644 550179
rect 42164 553270 42220 553326
rect 41780 552826 41836 552882
rect 41684 541282 41740 541338
rect 41972 551272 42028 551328
rect 41876 550902 41932 550958
rect 41876 548847 41932 548886
rect 41876 548830 41878 548847
rect 41878 548830 41930 548847
rect 41930 548830 41932 548847
rect 41876 547367 41932 547406
rect 41876 547350 41878 547367
rect 41878 547350 41930 547367
rect 41930 547350 41932 547367
rect 42164 549718 42220 549774
rect 42740 541578 42796 541634
rect 41972 540986 42028 541042
rect 42164 540986 42220 541042
rect 42836 535658 42892 535714
rect 42164 535066 42220 535122
rect 42836 531366 42892 531422
rect 41972 530626 42028 530682
rect 41780 529590 41836 529646
rect 41780 526482 41836 526538
rect 41780 432245 41782 432262
rect 41782 432245 41834 432262
rect 41834 432245 41836 432262
rect 41780 432206 41836 432245
rect 41780 431727 41782 431744
rect 41782 431727 41834 431744
rect 41834 431727 41836 431744
rect 41780 431688 41836 431727
rect 41588 431357 41590 431374
rect 41590 431357 41642 431374
rect 41642 431357 41644 431374
rect 41588 431318 41644 431357
rect 41780 430765 41782 430782
rect 41782 430765 41834 430782
rect 41834 430765 41836 430782
rect 41780 430726 41836 430765
rect 41780 430225 41836 430264
rect 41780 430208 41782 430225
rect 41782 430208 41834 430225
rect 41834 430208 41836 430225
rect 40724 429838 40780 429894
rect 40724 428950 40780 429006
rect 28820 419922 28876 419978
rect 28820 419478 28876 419534
rect 41588 428523 41644 428562
rect 41588 428506 41590 428523
rect 41590 428506 41642 428523
rect 41642 428506 41644 428523
rect 41876 425176 41932 425232
rect 41780 423252 41836 423308
rect 41588 421550 41644 421606
rect 41588 420975 41644 421014
rect 41588 420958 41590 420975
rect 41590 420958 41642 420975
rect 41642 420958 41644 420975
rect 41780 419791 41836 419830
rect 41780 419774 41782 419791
rect 41782 419774 41834 419791
rect 41834 419774 41836 419791
rect 41972 422734 42028 422790
rect 41972 411190 42028 411246
rect 41780 406010 41836 406066
rect 41780 403790 41836 403846
rect 41780 403050 41836 403106
rect 41780 402458 41836 402514
rect 41780 401866 41836 401922
rect 41780 399942 41836 399998
rect 41780 399498 41836 399554
rect 41876 398906 41932 398962
rect 41876 390906 41932 390962
rect 41876 389286 41932 389342
rect 41780 389029 41782 389046
rect 41782 389029 41834 389046
rect 41834 389029 41836 389046
rect 41780 388990 41836 389029
rect 41588 388733 41590 388750
rect 41590 388733 41642 388750
rect 41642 388733 41644 388750
rect 41588 388694 41644 388733
rect 41780 387993 41782 388010
rect 41782 387993 41834 388010
rect 41834 387993 41836 388010
rect 41780 387954 41836 387993
rect 41780 387549 41782 387566
rect 41782 387549 41834 387566
rect 41834 387549 41836 387566
rect 41780 387510 41836 387549
rect 41780 387009 41836 387048
rect 41780 386992 41782 387009
rect 41782 386992 41834 387009
rect 41834 386992 41836 387009
rect 41876 386030 41932 386086
rect 34484 385142 34540 385198
rect 41588 385181 41590 385198
rect 41590 385181 41642 385198
rect 41642 385181 41644 385198
rect 41588 385142 41644 385181
rect 41876 381960 41932 382016
rect 41780 380127 41836 380166
rect 41780 380110 41782 380127
rect 41782 380110 41834 380127
rect 41834 380110 41836 380127
rect 41780 379518 41836 379574
rect 41588 378778 41644 378834
rect 41588 378334 41644 378390
rect 41780 378038 41836 378094
rect 40244 377298 40300 377354
rect 28820 376706 28876 376762
rect 41780 376575 41836 376614
rect 41780 376558 41782 376575
rect 41782 376558 41834 376575
rect 41834 376558 41836 376575
rect 28820 376262 28876 376318
rect 41972 368122 42028 368178
rect 41780 362794 41836 362850
rect 41780 359834 41836 359890
rect 41780 359390 41836 359446
rect 41780 358650 41836 358706
rect 41780 356874 41836 356930
rect 41780 356430 41836 356486
rect 41780 355542 41836 355598
rect 41780 345887 41782 345904
rect 41782 345887 41834 345904
rect 41834 345887 41836 345904
rect 41780 345848 41836 345887
rect 41588 345517 41590 345534
rect 41590 345517 41642 345534
rect 41642 345517 41644 345534
rect 41588 345478 41644 345517
rect 41780 344777 41782 344794
rect 41782 344777 41834 344794
rect 41834 344777 41836 344794
rect 41780 344738 41836 344777
rect 41780 344333 41782 344350
rect 41782 344333 41834 344350
rect 41834 344333 41836 344350
rect 41780 344294 41836 344333
rect 41780 343867 41836 343906
rect 41780 343850 41782 343867
rect 41782 343850 41834 343867
rect 41834 343850 41836 343867
rect 41780 343297 41782 343314
rect 41782 343297 41834 343314
rect 41834 343297 41836 343314
rect 41780 343258 41836 343297
rect 41780 342335 41782 342352
rect 41782 342335 41834 342352
rect 41834 342335 41836 342352
rect 41780 342296 41836 342335
rect 41588 341965 41590 341982
rect 41590 341965 41642 341982
rect 41642 341965 41644 341982
rect 41588 341926 41644 341965
rect 41876 338818 41932 338874
rect 41780 336894 41836 336950
rect 41588 336154 41644 336210
rect 41588 335118 41644 335174
rect 41780 334822 41836 334878
rect 28820 333490 28876 333546
rect 41780 333359 41836 333398
rect 41780 333342 41782 333359
rect 41782 333342 41834 333359
rect 41834 333342 41836 333359
rect 28820 333046 28876 333102
rect 42452 335710 42508 335766
rect 41780 324906 41836 324962
rect 41780 319726 41836 319782
rect 41780 316766 41836 316822
rect 41780 316026 41836 316082
rect 41780 315434 41836 315490
rect 41876 313658 41932 313714
rect 41780 313214 41836 313270
rect 41780 312326 41836 312382
rect 41780 302671 41782 302688
rect 41782 302671 41834 302688
rect 41834 302671 41836 302688
rect 41780 302632 41836 302671
rect 41588 302301 41590 302318
rect 41590 302301 41642 302318
rect 41642 302301 41644 302318
rect 41588 302262 41644 302301
rect 41780 301561 41782 301578
rect 41782 301561 41834 301578
rect 41834 301561 41836 301578
rect 41780 301522 41836 301561
rect 41780 301191 41782 301208
rect 41782 301191 41834 301208
rect 41834 301191 41836 301208
rect 41780 301152 41836 301191
rect 41780 300651 41836 300690
rect 41780 300634 41782 300651
rect 41782 300634 41834 300651
rect 41834 300634 41836 300651
rect 41780 300081 41782 300098
rect 41782 300081 41834 300098
rect 41834 300081 41836 300098
rect 41780 300042 41836 300081
rect 41780 299637 41782 299654
rect 41782 299637 41834 299654
rect 41834 299637 41836 299654
rect 41780 299598 41836 299637
rect 41588 299341 41590 299358
rect 41590 299341 41642 299358
rect 41642 299341 41644 299358
rect 41588 299302 41644 299341
rect 41780 298601 41782 298618
rect 41782 298601 41834 298618
rect 41834 298601 41836 298618
rect 41780 298562 41836 298601
rect 41972 295602 42028 295658
rect 41780 293678 41836 293734
rect 41588 292938 41644 292994
rect 41588 291458 41644 291514
rect 41876 292568 41932 292624
rect 41876 292198 41932 292254
rect 28820 290422 28876 290478
rect 41780 290143 41836 290182
rect 41780 290126 41782 290143
rect 41782 290126 41834 290143
rect 41834 290126 41836 290143
rect 28820 289830 28876 289886
rect 41780 281690 41836 281746
rect 41780 276510 41836 276566
rect 41780 273550 41836 273606
rect 41780 272810 41836 272866
rect 41780 272366 41836 272422
rect 41780 270442 41836 270498
rect 41780 269998 41836 270054
rect 41780 269110 41836 269166
rect 41588 259677 41590 259694
rect 41590 259677 41642 259694
rect 41642 259677 41644 259694
rect 41588 259638 41644 259677
rect 41780 258937 41782 258954
rect 41782 258937 41834 258954
rect 41834 258937 41836 258954
rect 41780 258898 41836 258937
rect 41780 258345 41782 258362
rect 41782 258345 41834 258362
rect 41834 258345 41836 258362
rect 41780 258306 41836 258345
rect 41780 257975 41782 257992
rect 41782 257975 41834 257992
rect 41834 257975 41836 257992
rect 41780 257936 41836 257975
rect 41780 257435 41836 257474
rect 41780 257418 41782 257435
rect 41782 257418 41834 257435
rect 41834 257418 41836 257435
rect 41780 256865 41782 256882
rect 41782 256865 41834 256882
rect 41834 256865 41836 256882
rect 41780 256826 41836 256865
rect 41780 256495 41782 256512
rect 41782 256495 41834 256512
rect 41834 256495 41836 256512
rect 41780 256456 41836 256495
rect 41780 255955 41836 255994
rect 41780 255938 41782 255955
rect 41782 255938 41834 255955
rect 41834 255938 41836 255955
rect 41780 255385 41782 255402
rect 41782 255385 41834 255402
rect 41834 255385 41836 255402
rect 41780 255346 41836 255385
rect 41876 252386 41932 252442
rect 41780 250462 41836 250518
rect 41588 249722 41644 249778
rect 41588 249130 41644 249186
rect 41588 248242 41644 248298
rect 41588 247689 41590 247706
rect 41590 247689 41642 247706
rect 41642 247689 41644 247706
rect 41588 247650 41644 247689
rect 41588 247206 41644 247262
rect 41684 246614 41740 246670
rect 41972 248982 42028 249038
rect 41780 238326 41836 238382
rect 41780 233294 41836 233350
rect 41780 230334 41836 230390
rect 41780 229742 41836 229798
rect 41780 229002 41836 229058
rect 41876 227374 41932 227430
rect 41780 226782 41836 226838
rect 41972 226190 42028 226246
rect 41588 216461 41590 216478
rect 41590 216461 41642 216478
rect 41642 216461 41644 216478
rect 41588 216422 41644 216461
rect 41780 215721 41782 215738
rect 41782 215721 41834 215738
rect 41834 215721 41836 215738
rect 41780 215682 41836 215721
rect 41780 215203 41782 215220
rect 41782 215203 41834 215220
rect 41834 215203 41836 215220
rect 41780 215164 41836 215203
rect 41588 214981 41590 214998
rect 41590 214981 41642 214998
rect 41642 214981 41644 214998
rect 41588 214942 41644 214981
rect 41780 214241 41782 214258
rect 41782 214241 41834 214258
rect 41834 214241 41836 214258
rect 41780 214202 41836 214241
rect 41780 213649 41782 213666
rect 41782 213649 41834 213666
rect 41834 213649 41836 213666
rect 41780 213610 41836 213649
rect 44468 558894 44524 558950
rect 44180 278434 44236 278490
rect 41780 213279 41782 213296
rect 41782 213279 41834 213296
rect 41834 213279 41836 213296
rect 41780 213240 41836 213279
rect 41588 212909 41590 212926
rect 41590 212909 41642 212926
rect 41642 212909 41644 212926
rect 41588 212870 41644 212909
rect 41780 212169 41782 212186
rect 41782 212169 41834 212186
rect 41834 212169 41836 212186
rect 41780 212130 41836 212169
rect 41972 209170 42028 209226
rect 41588 207098 41644 207154
rect 41780 206728 41836 206784
rect 41876 206227 41932 206266
rect 41876 206210 41878 206227
rect 41878 206210 41930 206227
rect 41930 206210 41932 206227
rect 41780 205766 41836 205822
rect 41588 205026 41644 205082
rect 41684 204917 41686 204934
rect 41686 204917 41738 204934
rect 41738 204917 41740 204934
rect 41684 204878 41740 204917
rect 41780 204325 41782 204342
rect 41782 204325 41834 204342
rect 41834 204325 41836 204342
rect 41780 204286 41836 204325
rect 41780 203733 41782 203750
rect 41782 203733 41834 203750
rect 41834 203733 41836 203750
rect 41780 203694 41836 203733
rect 41780 195110 41836 195166
rect 45716 772902 45772 772958
rect 59540 975958 59596 976014
rect 59540 962934 59596 962990
rect 59540 949910 59596 949966
rect 59540 936886 59596 936942
rect 58580 923714 58636 923770
rect 59540 910690 59596 910746
rect 59540 897814 59596 897870
rect 58004 884790 58060 884846
rect 59540 871618 59596 871674
rect 58388 858594 58444 858650
rect 59540 845570 59596 845626
rect 59540 832546 59596 832602
rect 59540 819374 59596 819430
rect 59540 806515 59596 806554
rect 59540 806498 59542 806515
rect 59542 806498 59594 806515
rect 59594 806498 59596 806515
rect 59540 793474 59596 793530
rect 59540 780450 59596 780506
rect 47444 607586 47500 607642
rect 59540 767426 59596 767482
rect 59540 754254 59596 754310
rect 58580 741230 58636 741286
rect 59156 728206 59212 728262
rect 59540 715330 59596 715386
rect 59540 702158 59596 702214
rect 59540 689134 59596 689190
rect 59060 676110 59116 676166
rect 58100 663086 58156 663142
rect 59540 650062 59596 650118
rect 59540 637038 59596 637094
rect 59540 624014 59596 624070
rect 59252 610990 59308 611046
rect 59348 597966 59404 598022
rect 59540 584794 59596 584850
rect 59540 571770 59596 571826
rect 59540 558763 59596 558802
rect 59540 558746 59542 558763
rect 59542 558746 59594 558763
rect 59594 558746 59596 558763
rect 59540 545870 59596 545926
rect 59540 532863 59596 532902
rect 59540 532846 59542 532863
rect 59542 532846 59594 532863
rect 59594 532846 59596 532863
rect 59540 519674 59596 519730
rect 59540 506650 59596 506706
rect 59540 493626 59596 493682
rect 59540 480602 59596 480658
rect 57812 467430 57868 467486
rect 59540 454554 59596 454610
rect 57812 441530 57868 441586
rect 59540 428506 59596 428562
rect 59540 415334 59596 415390
rect 59540 402310 59596 402366
rect 59540 389286 59596 389342
rect 109940 1005558 109996 1005597
rect 110516 1005575 110572 1005614
rect 110516 1005558 110518 1005575
rect 110518 1005558 110570 1005575
rect 110570 1005558 110572 1005575
rect 102068 1005449 102070 1005466
rect 102070 1005449 102122 1005466
rect 102122 1005449 102124 1005466
rect 102068 1005410 102124 1005449
rect 107060 1005301 107062 1005318
rect 107062 1005301 107114 1005318
rect 107114 1005301 107116 1005318
rect 107060 1005262 107116 1005301
rect 94964 1005114 95020 1005170
rect 97172 1005114 97228 1005170
rect 97940 1005114 97996 1005170
rect 105428 1005153 105430 1005170
rect 105430 1005153 105482 1005170
rect 105482 1005153 105484 1005170
rect 94964 995807 95020 995846
rect 94964 995790 94966 995807
rect 94966 995790 95018 995807
rect 95018 995790 95020 995807
rect 94964 995642 95020 995698
rect 105428 1005114 105484 1005153
rect 108020 1005153 108022 1005170
rect 108022 1005153 108074 1005170
rect 108074 1005153 108076 1005170
rect 108020 1005114 108076 1005153
rect 103028 1002467 103084 1002506
rect 103028 1002450 103030 1002467
rect 103030 1002450 103082 1002467
rect 103082 1002450 103084 1002467
rect 101492 1002341 101494 1002358
rect 101494 1002341 101546 1002358
rect 101546 1002341 101548 1002358
rect 101492 1002302 101548 1002341
rect 103604 1002319 103660 1002358
rect 103604 1002302 103606 1002319
rect 103606 1002302 103658 1002319
rect 103658 1002302 103660 1002319
rect 106004 997901 106006 997918
rect 106006 997901 106058 997918
rect 106058 997901 106060 997918
rect 106004 997862 106060 997901
rect 108500 996251 108556 996290
rect 108500 996234 108502 996251
rect 108502 996234 108554 996251
rect 108554 996234 108556 996251
rect 100532 996086 100588 996142
rect 103988 996086 104044 996142
rect 104468 996086 104524 996142
rect 108596 996086 108652 996142
rect 109556 996086 109612 996142
rect 103604 995938 103660 995994
rect 103988 994014 104044 994070
rect 104468 993718 104524 993774
rect 112340 995790 112396 995846
rect 110324 993866 110380 993922
rect 115220 995938 115276 995994
rect 133652 995790 133708 995846
rect 137972 995790 138028 995846
rect 137396 995642 137452 995698
rect 132404 995346 132460 995402
rect 132788 994162 132844 994218
rect 136724 995494 136780 995550
rect 136148 993866 136204 993922
rect 129716 993718 129772 993774
rect 158516 1005575 158572 1005614
rect 158516 1005558 158518 1005575
rect 158518 1005558 158570 1005575
rect 158570 1005558 158572 1005575
rect 161396 1005449 161398 1005466
rect 161398 1005449 161450 1005466
rect 161450 1005449 161452 1005466
rect 146708 995955 146764 995994
rect 146708 995938 146710 995955
rect 146710 995938 146762 995955
rect 146762 995938 146764 995955
rect 146804 995642 146860 995698
rect 146708 995346 146764 995402
rect 149684 994162 149740 994218
rect 161396 1005410 161452 1005449
rect 161876 1005427 161932 1005466
rect 161876 1005410 161878 1005427
rect 161878 1005410 161930 1005427
rect 161930 1005410 161932 1005427
rect 151988 996086 152044 996142
rect 152372 996086 152428 996142
rect 159476 1005301 159478 1005318
rect 159478 1005301 159530 1005318
rect 159530 1005301 159532 1005318
rect 159476 1005262 159532 1005301
rect 161492 1005279 161548 1005318
rect 161492 1005262 161494 1005279
rect 161494 1005262 161546 1005279
rect 161546 1005262 161548 1005279
rect 160916 1005153 160918 1005170
rect 160918 1005153 160970 1005170
rect 160970 1005153 160972 1005170
rect 160916 1005114 160972 1005153
rect 156980 1004835 157036 1004874
rect 156980 1004818 156982 1004835
rect 156982 1004818 157034 1004835
rect 157034 1004818 157036 1004835
rect 153044 1002319 153100 1002358
rect 153044 1002302 153046 1002319
rect 153046 1002302 153098 1002319
rect 153098 1002302 153100 1002319
rect 154964 999381 154966 999398
rect 154966 999381 155018 999398
rect 155018 999381 155020 999398
rect 154964 999342 155020 999381
rect 153428 996251 153484 996290
rect 153428 996234 153430 996251
rect 153430 996234 153482 996251
rect 153482 996234 153484 996251
rect 154388 996273 154390 996290
rect 154390 996273 154442 996290
rect 154442 996273 154444 996290
rect 154388 996234 154444 996273
rect 159956 996251 160012 996290
rect 159956 996234 159958 996251
rect 159958 996234 160010 996251
rect 160010 996234 160012 996251
rect 154004 996086 154060 996142
rect 156500 996086 156556 996142
rect 157364 996086 157420 996142
rect 158900 996103 158956 996142
rect 158900 996086 158902 996103
rect 158902 996086 158954 996103
rect 158954 996086 158956 996103
rect 156212 995938 156268 995994
rect 159668 995955 159724 995994
rect 159668 995938 159670 995955
rect 159670 995938 159722 995955
rect 159722 995938 159724 995955
rect 157364 993718 157420 993774
rect 207380 1005449 207382 1005466
rect 207382 1005449 207434 1005466
rect 207434 1005449 207436 1005466
rect 185108 995790 185164 995846
rect 184340 995642 184396 995698
rect 190580 995642 190636 995698
rect 183284 995494 183340 995550
rect 188084 995494 188140 995550
rect 187316 995198 187372 995254
rect 207380 1005410 207436 1005449
rect 210836 1005301 210838 1005318
rect 210838 1005301 210890 1005318
rect 210890 1005301 210892 1005318
rect 210836 1005262 210892 1005301
rect 212852 1005279 212908 1005318
rect 212852 1005262 212854 1005279
rect 212854 1005262 212906 1005279
rect 212906 1005262 212908 1005279
rect 198644 995938 198700 995994
rect 197204 995050 197260 995106
rect 191540 993718 191596 993774
rect 201524 995346 201580 995402
rect 209876 1005153 209878 1005170
rect 209878 1005153 209930 1005170
rect 209930 1005153 209932 1005170
rect 209876 1005114 209932 1005153
rect 208436 1000839 208492 1000878
rect 208436 1000822 208438 1000839
rect 208438 1000822 208490 1000839
rect 208490 1000822 208492 1000839
rect 206324 999381 206326 999398
rect 206326 999381 206378 999398
rect 206378 999381 206380 999398
rect 206324 999342 206380 999381
rect 204884 996251 204940 996290
rect 204884 996234 204886 996251
rect 204886 996234 204938 996251
rect 204938 996234 204940 996251
rect 202292 996086 202348 996142
rect 202868 996086 202924 996142
rect 203924 996086 203980 996142
rect 205268 996086 205324 996142
rect 205940 996086 205996 996142
rect 207860 996086 207916 996142
rect 210836 996103 210892 996142
rect 210836 996086 210838 996103
rect 210838 996086 210890 996103
rect 210890 996086 210892 996103
rect 202868 995494 202924 995550
rect 211412 996125 211414 996142
rect 211414 996125 211466 996142
rect 211466 996125 211468 996142
rect 211412 996086 211468 996125
rect 212756 996103 212812 996142
rect 212756 996086 212758 996103
rect 212758 996086 212810 996103
rect 212810 996086 212812 996103
rect 219092 996086 219148 996142
rect 210164 995938 210220 995994
rect 216020 995938 216076 995994
rect 209108 995494 209164 995550
rect 240212 995790 240268 995846
rect 241844 995790 241900 995846
rect 232148 995642 232204 995698
rect 231476 994014 231532 994070
rect 235220 995494 235276 995550
rect 246932 995938 246988 995994
rect 238676 994310 238732 994366
rect 234356 994162 234412 994218
rect 247028 995494 247084 995550
rect 243188 993866 243244 993922
rect 351284 1007926 351340 1007982
rect 353396 1007926 353452 1007982
rect 261332 1006463 261388 1006502
rect 261332 1006446 261334 1006463
rect 261334 1006446 261386 1006463
rect 261386 1006446 261388 1006463
rect 262292 1005871 262348 1005910
rect 262292 1005854 262294 1005871
rect 262294 1005854 262346 1005871
rect 262346 1005854 262348 1005871
rect 255284 1002467 255340 1002506
rect 255284 1002450 255286 1002467
rect 255286 1002450 255338 1002467
rect 255338 1002450 255340 1002467
rect 253652 1002341 253654 1002358
rect 253654 1002341 253706 1002358
rect 253706 1002341 253708 1002358
rect 253652 1002302 253708 1002341
rect 254228 1002319 254284 1002358
rect 254228 1002302 254230 1002319
rect 254230 1002302 254282 1002319
rect 254282 1002302 254284 1002319
rect 256628 999507 256684 999546
rect 256628 999490 256630 999507
rect 256630 999490 256682 999507
rect 256682 999490 256684 999507
rect 259796 999529 259798 999546
rect 259798 999529 259850 999546
rect 259850 999529 259852 999546
rect 259796 999490 259852 999529
rect 257780 999381 257782 999398
rect 257782 999381 257834 999398
rect 257834 999381 257836 999398
rect 257780 999342 257836 999381
rect 256244 996547 256300 996586
rect 256244 996530 256246 996547
rect 256246 996530 256298 996547
rect 256298 996530 256300 996547
rect 252308 996086 252364 996142
rect 252692 996086 252748 996142
rect 254804 996086 254860 996142
rect 258740 996086 258796 996142
rect 260372 996086 260428 996142
rect 262772 996125 262774 996142
rect 262774 996125 262826 996142
rect 262826 996125 262828 996142
rect 262772 996086 262828 996125
rect 263732 996103 263788 996142
rect 263732 996086 263734 996103
rect 263734 996086 263786 996103
rect 263786 996086 263788 996103
rect 258740 994162 258796 994218
rect 251828 993718 251884 993774
rect 270740 996086 270796 996142
rect 261524 995955 261580 995994
rect 261524 995938 261526 995955
rect 261526 995938 261578 995955
rect 261578 995938 261580 995955
rect 262484 995977 262486 995994
rect 262486 995977 262538 995994
rect 262538 995977 262540 995994
rect 262484 995938 262540 995977
rect 267860 995938 267916 995994
rect 267956 995790 268012 995846
rect 313844 1005279 313900 1005318
rect 313844 1005262 313846 1005279
rect 313846 1005262 313898 1005279
rect 313898 1005262 313900 1005279
rect 316436 1005301 316438 1005318
rect 316438 1005301 316490 1005318
rect 316490 1005301 316492 1005318
rect 316436 1005262 316492 1005301
rect 308276 1005153 308278 1005170
rect 308278 1005153 308330 1005170
rect 308330 1005153 308332 1005170
rect 286772 995790 286828 995846
rect 291764 995790 291820 995846
rect 293588 995642 293644 995698
rect 308276 1005114 308332 1005153
rect 312884 1005153 312886 1005170
rect 312886 1005153 312938 1005170
rect 312938 1005153 312940 1005170
rect 312884 1005114 312940 1005153
rect 306740 1002637 306742 1002654
rect 306742 1002637 306794 1002654
rect 306794 1002637 306796 1002654
rect 298484 995938 298540 995994
rect 306740 1002598 306796 1002637
rect 307316 1002615 307372 1002654
rect 307316 1002598 307318 1002615
rect 307318 1002598 307370 1002615
rect 307370 1002598 307372 1002615
rect 299540 995790 299596 995846
rect 299732 995642 299788 995698
rect 284372 995494 284428 995550
rect 287444 995346 287500 995402
rect 286004 994458 286060 994514
rect 283508 994162 283564 994218
rect 282836 994014 282892 994070
rect 305300 1002467 305356 1002506
rect 305300 1002450 305302 1002467
rect 305302 1002450 305354 1002467
rect 305354 1002450 305356 1002467
rect 307892 1002489 307894 1002506
rect 307894 1002489 307946 1002506
rect 307946 1002489 307948 1002506
rect 307892 1002450 307948 1002489
rect 305780 1002319 305836 1002358
rect 305780 1002302 305782 1002319
rect 305782 1002302 305834 1002319
rect 305834 1002302 305836 1002319
rect 306356 1002341 306358 1002358
rect 306358 1002341 306410 1002358
rect 306410 1002341 306412 1002358
rect 306356 1002302 306412 1002341
rect 311444 999529 311446 999546
rect 311446 999529 311498 999546
rect 311498 999529 311500 999546
rect 311444 999490 311500 999529
rect 309332 999381 309334 999398
rect 309334 999381 309386 999398
rect 309386 999381 309388 999398
rect 309332 999342 309388 999381
rect 309812 996547 309868 996586
rect 309812 996530 309814 996547
rect 309814 996530 309866 996547
rect 309866 996530 309868 996547
rect 304436 996086 304492 996142
rect 304916 996086 304972 996142
rect 305300 996086 305356 996142
rect 310868 996086 310924 996142
rect 314228 996125 314230 996142
rect 314230 996125 314282 996142
rect 314282 996125 314284 996142
rect 304820 995938 304876 995994
rect 303380 995790 303436 995846
rect 300116 995346 300172 995402
rect 303380 994458 303436 994514
rect 304820 994162 304876 994218
rect 294548 993718 294604 993774
rect 314228 996086 314284 996125
rect 319604 996086 319660 996142
rect 313076 995977 313078 995994
rect 313078 995977 313130 995994
rect 313130 995977 313132 995994
rect 313076 995938 313132 995977
rect 313844 995938 313900 995994
rect 310868 994014 310924 994070
rect 316724 993866 316780 993922
rect 319700 995938 319756 995994
rect 356372 1006041 356374 1006058
rect 356374 1006041 356426 1006058
rect 356426 1006041 356428 1006058
rect 356372 1006002 356428 1006041
rect 357908 1006019 357964 1006058
rect 558164 1006041 558166 1006058
rect 558166 1006041 558218 1006058
rect 558218 1006041 558220 1006058
rect 357908 1006002 357910 1006019
rect 357910 1006002 357962 1006019
rect 357962 1006002 357964 1006019
rect 358772 1005893 358774 1005910
rect 358774 1005893 358826 1005910
rect 358826 1005893 358828 1005910
rect 358772 1005854 358828 1005893
rect 359348 1005871 359404 1005910
rect 359348 1005854 359350 1005871
rect 359350 1005854 359402 1005871
rect 359402 1005854 359404 1005871
rect 361844 1005723 361900 1005762
rect 361844 1005706 361846 1005723
rect 361846 1005706 361898 1005723
rect 361898 1005706 361900 1005723
rect 356756 1005575 356812 1005614
rect 356756 1005558 356758 1005575
rect 356758 1005558 356810 1005575
rect 356810 1005558 356812 1005575
rect 357140 1005558 357196 1005614
rect 358292 1005597 358294 1005614
rect 358294 1005597 358346 1005614
rect 358346 1005597 358348 1005614
rect 358292 1005558 358348 1005597
rect 361268 1005427 361324 1005466
rect 361268 1005410 361270 1005427
rect 361270 1005410 361322 1005427
rect 361322 1005410 361324 1005427
rect 360884 1005301 360886 1005318
rect 360886 1005301 360938 1005318
rect 360938 1005301 360940 1005318
rect 360884 1005262 360940 1005301
rect 362324 1005279 362380 1005318
rect 362324 1005262 362326 1005279
rect 362326 1005262 362378 1005279
rect 362378 1005262 362380 1005279
rect 362804 1005153 362806 1005170
rect 362806 1005153 362858 1005170
rect 362858 1005153 362860 1005170
rect 362804 1005114 362860 1005153
rect 558164 1006002 558220 1006041
rect 359732 1000839 359788 1000878
rect 359732 1000822 359734 1000839
rect 359734 1000822 359786 1000839
rect 359786 1000822 359788 1000839
rect 363860 996086 363916 996142
rect 366260 996086 366316 996142
rect 366740 996103 366796 996142
rect 366740 996086 366742 996103
rect 366742 996086 366794 996103
rect 366794 996086 366796 996103
rect 360020 995642 360076 995698
rect 362900 995642 362956 995698
rect 363476 995642 363532 995698
rect 371540 996086 371596 996142
rect 364436 995642 364492 995698
rect 374420 995938 374476 995994
rect 374516 993866 374572 993922
rect 425684 1005893 425686 1005910
rect 425686 1005893 425738 1005910
rect 425738 1005893 425740 1005910
rect 425684 1005854 425740 1005893
rect 429716 1005871 429772 1005910
rect 429716 1005854 429718 1005871
rect 429718 1005854 429770 1005871
rect 429770 1005854 429772 1005871
rect 428276 1005745 428278 1005762
rect 428278 1005745 428330 1005762
rect 428330 1005745 428332 1005762
rect 428276 1005706 428332 1005745
rect 428660 1005723 428716 1005762
rect 428660 1005706 428662 1005723
rect 428662 1005706 428714 1005723
rect 428714 1005706 428716 1005723
rect 380180 995642 380236 995698
rect 382772 995790 382828 995846
rect 425300 1005575 425356 1005614
rect 425300 1005558 425302 1005575
rect 425302 1005558 425354 1005575
rect 425354 1005558 425356 1005575
rect 426740 1005597 426742 1005614
rect 426742 1005597 426794 1005614
rect 426794 1005597 426796 1005614
rect 426740 1005558 426796 1005597
rect 423764 1005449 423766 1005466
rect 423766 1005449 423818 1005466
rect 423818 1005449 423820 1005466
rect 423764 1005410 423820 1005449
rect 424724 1005427 424780 1005466
rect 424724 1005410 424726 1005427
rect 424726 1005410 424778 1005427
rect 424778 1005410 424780 1005427
rect 424148 1005301 424150 1005318
rect 424150 1005301 424202 1005318
rect 424202 1005301 424204 1005318
rect 424148 1005262 424204 1005301
rect 426164 1005279 426220 1005318
rect 426164 1005262 426166 1005279
rect 426166 1005262 426218 1005279
rect 426218 1005262 426220 1005279
rect 417524 1005114 417580 1005170
rect 420788 1005114 420844 1005170
rect 421556 1005114 421612 1005170
rect 388820 995790 388876 995846
rect 394868 995642 394924 995698
rect 392084 993866 392140 993922
rect 373940 993718 373996 993774
rect 374612 993718 374668 993774
rect 396980 993718 397036 993774
rect 430196 1000987 430252 1001026
rect 430196 1000970 430198 1000987
rect 430198 1000970 430250 1000987
rect 430250 1000970 430252 1000987
rect 427124 1000839 427180 1000878
rect 427124 1000822 427126 1000839
rect 427126 1000822 427178 1000839
rect 427178 1000822 427180 1000839
rect 429236 1000861 429238 1000878
rect 429238 1000861 429290 1000878
rect 429290 1000861 429292 1000878
rect 429236 1000822 429292 1000861
rect 430196 996086 430252 996142
rect 431252 996086 431308 996142
rect 432788 996125 432790 996142
rect 432790 996125 432842 996142
rect 432842 996125 432844 996142
rect 432788 996086 432844 996125
rect 433556 996086 433612 996142
rect 434132 996103 434188 996142
rect 434132 996086 434134 996103
rect 434134 996086 434186 996103
rect 434186 996086 434188 996103
rect 427412 995642 427468 995698
rect 430868 995494 430924 995550
rect 437972 996086 438028 996142
rect 431828 995494 431884 995550
rect 440660 995938 440716 995994
rect 551636 1005871 551692 1005910
rect 551636 1005854 551638 1005871
rect 551638 1005854 551690 1005871
rect 551690 1005854 551692 1005871
rect 501716 1005723 501772 1005762
rect 501716 1005706 501718 1005723
rect 501718 1005706 501770 1005723
rect 501770 1005706 501772 1005723
rect 502292 1005745 502294 1005762
rect 502294 1005745 502346 1005762
rect 502346 1005745 502348 1005762
rect 502292 1005706 502348 1005745
rect 553652 1005745 553654 1005762
rect 553654 1005745 553706 1005762
rect 553706 1005745 553708 1005762
rect 471860 995938 471916 995994
rect 502676 1005575 502732 1005614
rect 502676 1005558 502678 1005575
rect 502678 1005558 502730 1005575
rect 502730 1005558 502732 1005575
rect 500756 1005449 500758 1005466
rect 500758 1005449 500810 1005466
rect 500810 1005449 500812 1005466
rect 500756 1005410 500812 1005449
rect 503732 1005427 503788 1005466
rect 503732 1005410 503734 1005427
rect 503734 1005410 503786 1005427
rect 503786 1005410 503788 1005427
rect 503252 1005279 503308 1005318
rect 503252 1005262 503254 1005279
rect 503254 1005262 503306 1005279
rect 503306 1005262 503308 1005279
rect 505268 1005301 505270 1005318
rect 505270 1005301 505322 1005318
rect 505322 1005301 505324 1005318
rect 505268 1005262 505324 1005301
rect 501140 1005153 501142 1005170
rect 501142 1005153 501194 1005170
rect 501194 1005153 501196 1005170
rect 501140 1005114 501196 1005153
rect 506708 1005153 506710 1005170
rect 506710 1005153 506762 1005170
rect 506762 1005153 506764 1005170
rect 506708 1005114 506764 1005153
rect 505652 1002319 505708 1002358
rect 505652 1002302 505654 1002319
rect 505654 1002302 505706 1002319
rect 505706 1002302 505708 1002319
rect 472148 995790 472204 995846
rect 471956 995494 472012 995550
rect 507188 1000839 507244 1000878
rect 507188 1000822 507190 1000839
rect 507190 1000822 507242 1000839
rect 507242 1000822 507244 1000839
rect 506228 1000691 506284 1000730
rect 506228 1000674 506230 1000691
rect 506230 1000674 506282 1000691
rect 506282 1000674 506284 1000691
rect 504212 999507 504268 999546
rect 504212 999490 504214 999507
rect 504214 999490 504266 999507
rect 504266 999490 504268 999507
rect 499124 996086 499180 996142
rect 509780 996125 509782 996142
rect 509782 996125 509834 996142
rect 509834 996125 509836 996142
rect 509780 996086 509836 996125
rect 510740 996125 510742 996142
rect 510742 996125 510794 996142
rect 510794 996125 510796 996142
rect 510740 996086 510796 996125
rect 511124 996086 511180 996142
rect 515540 996086 515596 996142
rect 507860 995938 507916 995994
rect 508436 995938 508492 995994
rect 512660 995938 512716 995994
rect 478388 995790 478444 995846
rect 482036 995790 482092 995846
rect 495284 995790 495340 995846
rect 499124 995790 499180 995846
rect 481364 995494 481420 995550
rect 485588 995494 485644 995550
rect 471668 993866 471724 993922
rect 484148 993866 484204 993922
rect 466580 993718 466636 993774
rect 485972 993718 486028 993774
rect 491828 995494 491884 995550
rect 504404 995494 504460 995550
rect 507284 995494 507340 995550
rect 508820 995494 508876 995550
rect 517860 1000839 517916 1000878
rect 517860 1000822 517862 1000839
rect 517862 1000822 517914 1000839
rect 517914 1000822 517916 1000839
rect 518084 1000691 518140 1000730
rect 518084 1000674 518086 1000691
rect 518086 1000674 518138 1000691
rect 518138 1000674 518140 1000691
rect 518084 999342 518140 999398
rect 553652 1005706 553708 1005745
rect 554612 1005723 554668 1005762
rect 554612 1005706 554614 1005723
rect 554614 1005706 554666 1005723
rect 554666 1005706 554668 1005723
rect 520532 999638 520588 999694
rect 521300 999490 521356 999546
rect 521492 995938 521548 995994
rect 521396 995790 521452 995846
rect 554036 1005597 554038 1005614
rect 554038 1005597 554090 1005614
rect 554090 1005597 554092 1005614
rect 554036 1005558 554092 1005597
rect 555188 1005449 555190 1005466
rect 555190 1005449 555242 1005466
rect 555242 1005449 555244 1005466
rect 555188 1005410 555244 1005449
rect 552212 1005279 552268 1005318
rect 552212 1005262 552214 1005279
rect 552214 1005262 552266 1005279
rect 552266 1005262 552268 1005279
rect 552596 1005301 552598 1005318
rect 552598 1005301 552650 1005318
rect 552650 1005301 552652 1005318
rect 552596 1005262 552652 1005301
rect 552980 1005153 552982 1005170
rect 552982 1005153 553034 1005170
rect 553034 1005153 553036 1005170
rect 552980 1005114 553036 1005153
rect 558548 1002319 558604 1002358
rect 558548 1002302 558550 1002319
rect 558550 1002302 558602 1002319
rect 558602 1002302 558604 1002319
rect 523604 999638 523660 999694
rect 521588 995642 521644 995698
rect 523700 999490 523756 999546
rect 523892 1000822 523948 1000878
rect 523988 1000674 524044 1000730
rect 524084 999342 524140 999398
rect 527924 995790 527980 995846
rect 537236 995790 537292 995846
rect 555572 997605 555574 997622
rect 555574 997605 555626 997622
rect 555626 997605 555628 997622
rect 555572 997566 555628 997605
rect 557588 997457 557590 997474
rect 557590 997457 557642 997474
rect 557642 997457 557644 997474
rect 557588 997418 557644 997457
rect 555956 996086 556012 996142
rect 559124 996086 559180 996142
rect 561140 996103 561196 996142
rect 561140 996086 561142 996103
rect 561142 996086 561194 996103
rect 561194 996086 561196 996103
rect 532244 995642 532300 995698
rect 518516 995494 518572 995550
rect 518420 995346 518476 995402
rect 533396 995494 533452 995550
rect 535316 995346 535372 995402
rect 561908 996103 561964 996142
rect 561908 996086 561910 996103
rect 561910 996086 561962 996103
rect 561962 996086 561964 996103
rect 569876 996086 569932 996142
rect 560180 995938 560236 995994
rect 569780 995938 569836 995994
rect 567188 995790 567244 995846
rect 565844 995642 565900 995698
rect 561620 995198 561676 995254
rect 566036 995494 566092 995550
rect 567380 995346 567436 995402
rect 567380 994014 567436 994070
rect 573140 994458 573196 994514
rect 573044 994310 573100 994366
rect 573236 994162 573292 994218
rect 574676 993866 574732 993922
rect 572948 993718 573004 993774
rect 631796 994458 631852 994514
rect 630932 994310 630988 994366
rect 629972 994014 630028 994070
rect 636116 994162 636172 994218
rect 639188 993866 639244 993922
rect 637364 993718 637420 993774
rect 638516 993718 638572 993774
rect 641108 993718 641164 993774
rect 61940 384402 61996 384458
rect 59444 376262 59500 376318
rect 58388 363238 58444 363294
rect 59540 350214 59596 350270
rect 59540 337190 59596 337246
rect 59540 324166 59596 324222
rect 58580 311142 58636 311198
rect 59540 297970 59596 298026
rect 59540 285133 59542 285150
rect 59542 285133 59594 285150
rect 59594 285133 59596 285150
rect 59540 285094 59596 285133
rect 62228 389138 62284 389194
rect 62036 278286 62092 278342
rect 62228 278138 62284 278194
rect 63380 277990 63436 278046
rect 69428 272218 69484 272274
rect 67028 269406 67084 269462
rect 65876 269258 65932 269314
rect 71732 272070 71788 272126
rect 70580 269554 70636 269610
rect 130868 269850 130924 269906
rect 128564 269702 128620 269758
rect 41780 190078 41836 190134
rect 41780 187118 41836 187174
rect 41780 186674 41836 186730
rect 41780 185786 41836 185842
rect 41780 184010 41836 184066
rect 41780 183566 41836 183622
rect 41780 182974 41836 183030
rect 149396 244542 149452 244598
rect 148244 242026 148300 242082
rect 146900 229890 146956 229946
rect 146996 228114 147052 228170
rect 146900 165510 146956 165566
rect 148148 222638 148204 222694
rect 148052 221454 148108 221510
rect 147380 217754 147436 217810
rect 147284 216570 147340 216626
rect 147380 214794 147436 214850
rect 147092 212870 147148 212926
rect 147380 211686 147436 211742
rect 147284 209170 147340 209226
rect 147956 201622 148012 201678
rect 147860 198366 147916 198422
rect 147764 192150 147820 192206
rect 147572 190966 147628 191022
rect 147476 189782 147532 189838
rect 147188 177646 147244 177702
rect 147188 176462 147244 176518
rect 147092 175130 147148 175186
rect 146996 164326 147052 164382
rect 147380 178847 147436 178886
rect 147380 178830 147382 178847
rect 147382 178830 147434 178847
rect 147434 178830 147436 178847
rect 147380 173946 147436 174002
rect 147284 170246 147340 170302
rect 147092 129102 147148 129158
rect 146996 120518 147052 120574
rect 146900 111934 146956 111990
rect 147668 187414 147724 187470
rect 147572 183714 147628 183770
rect 148724 240842 148780 240898
rect 148532 238474 148588 238530
rect 148340 236698 148396 236754
rect 148436 233590 148492 233646
rect 148628 231074 148684 231130
rect 149396 239658 149452 239714
rect 149012 235958 149068 236014
rect 148820 226338 148876 226394
rect 148916 219678 148972 219734
rect 148916 184454 148972 184510
rect 148916 172762 148972 172818
rect 149396 234774 149452 234830
rect 149204 232258 149260 232314
rect 149108 225154 149164 225210
rect 148916 168026 148972 168082
rect 148340 159442 148396 159498
rect 148244 156926 148300 156982
rect 148052 148490 148108 148546
rect 148052 147306 148108 147362
rect 147956 146122 148012 146178
rect 147956 144363 148012 144402
rect 147956 144346 147958 144363
rect 147958 144346 148010 144363
rect 148010 144346 148012 144363
rect 147860 143606 147916 143662
rect 147860 142422 147916 142478
rect 147668 141255 147724 141294
rect 147668 141238 147670 141255
rect 147670 141238 147722 141255
rect 147722 141238 147724 141255
rect 147956 138722 148012 138778
rect 147860 135022 147916 135078
rect 147668 133838 147724 133894
rect 147572 130878 147628 130934
rect 147188 126586 147244 126642
rect 147284 125402 147340 125458
rect 147380 124218 147436 124274
rect 147476 122442 147532 122498
rect 147764 130286 147820 130342
rect 147668 103498 147724 103554
rect 148052 137538 148108 137594
rect 148148 132654 148204 132710
rect 147956 106014 148012 106070
rect 147572 94914 147628 94970
rect 148052 104682 148108 104738
rect 148820 157666 148876 157722
rect 148436 155742 148492 155798
rect 148628 154558 148684 154614
rect 148532 150858 148588 150914
rect 148340 109418 148396 109474
rect 148244 99798 148300 99854
rect 148148 98614 148204 98670
rect 148724 152042 148780 152098
rect 149012 161810 149068 161866
rect 149396 227374 149452 227430
rect 149300 206358 149356 206414
rect 149300 199550 149356 199606
rect 149300 195889 149302 195906
rect 149302 195889 149354 195906
rect 149354 195889 149356 195906
rect 149300 195850 149356 195889
rect 149492 223822 149548 223878
rect 149588 218955 149644 218994
rect 149588 218938 149590 218955
rect 149590 218938 149642 218955
rect 149642 218938 149644 218955
rect 149492 214054 149548 214110
rect 149492 210354 149548 210410
rect 149492 207986 149548 208042
rect 149492 205618 149548 205674
rect 149492 203250 149548 203306
rect 149492 200734 149548 200790
rect 149204 166250 149260 166306
rect 149108 160626 149164 160682
rect 149396 194683 149452 194722
rect 149396 194666 149398 194683
rect 149398 194666 149450 194683
rect 149450 194666 149452 194683
rect 149396 193055 149452 193094
rect 149396 193038 149398 193055
rect 149398 193038 149450 193055
rect 149450 193038 149452 193055
rect 149396 188006 149452 188062
rect 149396 186230 149452 186286
rect 149396 182530 149452 182586
rect 149396 179587 149452 179626
rect 149396 179570 149398 179587
rect 149398 179570 149450 179587
rect 149450 179570 149452 179587
rect 149396 170986 149452 171042
rect 149396 169062 149452 169118
rect 149204 139906 149260 139962
rect 149204 135762 149260 135818
rect 149396 163142 149452 163198
rect 149300 127918 149356 127974
rect 149684 204434 149740 204490
rect 149684 197034 149740 197090
rect 149684 181346 149740 181402
rect 149588 149822 149644 149878
rect 149300 121702 149356 121758
rect 149204 119334 149260 119390
rect 148916 118150 148972 118206
rect 148820 110898 148876 110954
rect 148436 108382 148492 108438
rect 148628 107198 148684 107254
rect 148532 102314 148588 102370
rect 148724 97430 148780 97486
rect 148340 85294 148396 85350
rect 148532 84110 148588 84166
rect 148436 81594 148492 81650
rect 149108 116818 149164 116874
rect 149012 114450 149068 114506
rect 148916 92546 148972 92602
rect 148820 86478 148876 86534
rect 148724 80410 148780 80466
rect 148628 77894 148684 77950
rect 149588 115634 149644 115690
rect 149492 113118 149548 113174
rect 149204 93730 149260 93786
rect 149012 91362 149068 91418
rect 149108 90178 149164 90234
rect 149492 95654 149548 95710
rect 149300 88994 149356 89050
rect 149396 87218 149452 87274
rect 185300 221010 185356 221066
rect 184340 219530 184396 219586
rect 184340 199698 184396 199754
rect 184244 197626 184300 197682
rect 184340 196738 184396 196794
rect 193076 272218 193132 272274
rect 192596 269406 192652 269462
rect 192404 269258 192460 269314
rect 185492 220270 185548 220326
rect 185588 218790 185644 218846
rect 185396 198218 185452 198274
rect 184436 195998 184492 196054
rect 184340 195258 184396 195314
rect 184436 194370 184492 194426
rect 184532 193778 184588 193834
rect 184436 192890 184492 192946
rect 184340 192298 184396 192354
rect 184532 191410 184588 191466
rect 184628 190670 184684 190726
rect 184340 189930 184396 189986
rect 184436 189190 184492 189246
rect 184532 188450 184588 188506
rect 184628 187562 184684 187618
rect 184436 186822 184492 186878
rect 184340 186082 184396 186138
rect 184628 185342 184684 185398
rect 184532 184602 184588 184658
rect 184340 183862 184396 183918
rect 184532 183122 184588 183178
rect 184436 182382 184492 182438
rect 184628 181494 184684 181550
rect 184340 180754 184396 180810
rect 184436 180014 184492 180070
rect 184532 179274 184588 179330
rect 184628 178534 184684 178590
rect 184340 177646 184396 177702
rect 184436 177054 184492 177110
rect 184532 176166 184588 176222
rect 184340 175613 184342 175630
rect 184342 175613 184394 175630
rect 184394 175613 184396 175630
rect 184340 175574 184396 175613
rect 184436 173946 184492 174002
rect 184340 172466 184396 172522
rect 184436 170838 184492 170894
rect 184532 170246 184588 170302
rect 184340 169358 184396 169414
rect 184436 168618 184492 168674
rect 184532 167878 184588 167934
rect 184628 167138 184684 167194
rect 184340 166398 184396 166454
rect 184436 165658 184492 165714
rect 184532 164770 184588 164826
rect 184340 164069 184342 164086
rect 184342 164069 184394 164086
rect 184394 164069 184396 164086
rect 184340 164030 184396 164069
rect 184340 163290 184396 163346
rect 184436 162550 184492 162606
rect 184532 161810 184588 161866
rect 184340 160922 184396 160978
rect 184436 160330 184492 160386
rect 184532 159442 184588 159498
rect 184628 158850 184684 158906
rect 184436 157962 184492 158018
rect 184532 157370 184588 157426
rect 184340 156482 184396 156538
rect 184628 155594 184684 155650
rect 184340 155002 184396 155058
rect 184436 154114 184492 154170
rect 184724 153522 184780 153578
rect 184532 152634 184588 152690
rect 184340 151894 184396 151950
rect 184532 151154 184588 151210
rect 184436 150414 184492 150470
rect 184340 148934 184396 148990
rect 184628 149674 184684 149730
rect 184436 148046 184492 148102
rect 184532 147306 184588 147362
rect 184340 145826 184396 145882
rect 184532 145086 184588 145142
rect 184436 144346 184492 144402
rect 184436 143606 184492 143662
rect 184340 142718 184396 142774
rect 184532 142126 184588 142182
rect 184628 141238 184684 141294
rect 184340 140498 184396 140554
rect 184532 139758 184588 139814
rect 184436 138870 184492 138926
rect 185876 201326 185932 201382
rect 186164 207246 186220 207302
rect 186452 211982 186508 212038
rect 186836 218050 186892 218106
rect 187124 243358 187180 243414
rect 187028 216422 187084 216478
rect 186932 214942 186988 214998
rect 186740 213462 186796 213518
rect 186644 210502 186700 210558
rect 186548 209022 186604 209078
rect 186356 205174 186412 205230
rect 186260 204286 186316 204342
rect 186068 202806 186124 202862
rect 194228 272070 194284 272126
rect 193748 269554 193804 269610
rect 206996 267926 207052 267982
rect 210740 269850 210796 269906
rect 210260 269702 210316 269758
rect 211412 267926 211468 267982
rect 368948 276362 369004 276418
rect 368372 268814 368428 268870
rect 370100 271922 370156 271978
rect 371252 273550 371308 273606
rect 370292 269258 370348 269314
rect 372692 268962 372748 269018
rect 375572 269110 375628 269166
rect 377012 273402 377068 273458
rect 379892 273254 379948 273310
rect 378644 270590 378700 270646
rect 381812 276214 381868 276270
rect 381236 270442 381292 270498
rect 383636 276066 383692 276122
rect 384884 275918 384940 275974
rect 385556 273106 385612 273162
rect 387764 275770 387820 275826
rect 387284 270294 387340 270350
rect 390836 275622 390892 275678
rect 387956 266742 388012 266798
rect 390164 270146 390220 270202
rect 389684 266890 389740 266946
rect 391988 275474 392044 275530
rect 391508 272958 391564 273014
rect 393236 275326 393292 275382
rect 394388 272810 394444 272866
rect 396308 275030 396364 275086
rect 395636 269998 395692 270054
rect 397556 275178 397612 275234
rect 399956 272662 400012 272718
rect 401300 269850 401356 269906
rect 401780 266594 401836 266650
rect 403028 272514 403084 272570
rect 402836 269258 402892 269314
rect 404180 269702 404236 269758
rect 405620 272366 405676 272422
rect 407828 266298 407884 266354
rect 408500 272218 408556 272274
rect 409172 266446 409228 266502
rect 409940 269554 409996 269610
rect 410420 269406 410476 269462
rect 411764 272070 411820 272126
rect 411572 269258 411628 269314
rect 542228 276362 542284 276418
rect 544628 271922 544684 271978
rect 541076 268814 541132 268870
rect 548180 273550 548236 273606
rect 551732 268962 551788 269018
rect 558836 269110 558892 269166
rect 562388 273402 562444 273458
rect 565844 270590 565900 270646
rect 569492 273254 569548 273310
rect 574196 276214 574252 276270
rect 572948 270442 573004 270498
rect 578900 276066 578956 276122
rect 581300 275918 581356 275974
rect 583604 273106 583660 273162
rect 588308 275770 588364 275826
rect 587156 270294 587212 270350
rect 596660 275622 596716 275678
rect 599060 275474 599116 275530
rect 597812 272958 597868 273014
rect 594356 270146 594412 270202
rect 593108 266890 593164 266946
rect 589556 266742 589612 266798
rect 602516 275326 602572 275382
rect 604916 272810 604972 272866
rect 609716 275030 609772 275086
rect 613172 275178 613228 275234
rect 608468 269998 608524 270054
rect 619028 272662 619084 272718
rect 622676 269850 622732 269906
rect 626132 272514 626188 272570
rect 623828 266594 623884 266650
rect 633332 272366 633388 272422
rect 629780 269702 629836 269758
rect 640436 272218 640492 272274
rect 643892 269554 643948 269610
rect 645140 269406 645196 269462
rect 648692 272070 648748 272126
rect 647540 269258 647596 269314
rect 641588 266446 641644 266502
rect 638036 266298 638092 266354
rect 420404 262171 420460 262210
rect 420404 262154 420406 262171
rect 420406 262154 420458 262171
rect 420458 262154 420460 262171
rect 420404 259786 420460 259842
rect 190004 259342 190060 259398
rect 189908 251646 189964 251702
rect 420404 256974 420460 257030
rect 420404 255198 420460 255254
rect 420404 252830 420460 252886
rect 420308 250462 420364 250518
rect 420404 248094 420460 248150
rect 420404 245282 420460 245338
rect 420404 243506 420460 243562
rect 420404 241138 420460 241194
rect 302900 228410 302956 228466
rect 310676 228558 310732 228614
rect 314900 228706 314956 228762
rect 316724 231222 316780 231278
rect 319508 231370 319564 231426
rect 324020 231518 324076 231574
rect 324788 225450 324844 225506
rect 327092 231666 327148 231722
rect 328052 225598 328108 225654
rect 330836 225746 330892 225802
rect 332468 228871 332524 228910
rect 332468 228854 332470 228871
rect 332470 228854 332522 228871
rect 332522 228854 332524 228871
rect 332564 225894 332620 225950
rect 335348 227374 335404 227430
rect 336788 236106 336844 236162
rect 339380 233146 339436 233202
rect 338708 228871 338764 228910
rect 338708 228854 338710 228871
rect 338710 228854 338762 228871
rect 338762 228854 338764 228871
rect 338612 227226 338668 227282
rect 341588 226930 341644 226986
rect 342548 234626 342604 234682
rect 342164 232998 342220 233054
rect 344372 235958 344428 236014
rect 344756 233294 344812 233350
rect 348788 230334 348844 230390
rect 348692 227078 348748 227134
rect 353492 234922 353548 234978
rect 354068 222786 354124 222842
rect 355700 222934 355756 222990
rect 356276 230186 356332 230242
rect 356852 226782 356908 226838
rect 359444 235366 359500 235422
rect 359060 230038 359116 230094
rect 358964 224562 359020 224618
rect 359828 224414 359884 224470
rect 361748 229890 361804 229946
rect 362516 234478 362572 234534
rect 362804 233294 362860 233350
rect 368564 234034 368620 234090
rect 369140 224266 369196 224322
rect 372212 236254 372268 236310
rect 371156 229742 371212 229798
rect 370292 224118 370348 224174
rect 373460 236846 373516 236902
rect 374324 232702 374380 232758
rect 374036 232554 374092 232610
rect 376724 236402 376780 236458
rect 376340 235810 376396 235866
rect 374900 223970 374956 224026
rect 377972 236994 378028 237050
rect 379124 234330 379180 234386
rect 380852 236550 380908 236606
rect 380468 232406 380524 232462
rect 379892 231962 379948 232018
rect 379796 223822 379852 223878
rect 381236 236698 381292 236754
rect 381332 232110 381388 232166
rect 382100 234182 382156 234238
rect 381716 229446 381772 229502
rect 383540 232258 383596 232314
rect 383828 236846 383884 236902
rect 384020 236846 384076 236902
rect 383636 229298 383692 229354
rect 385748 235662 385804 235718
rect 384980 229150 385036 229206
rect 382868 223674 382924 223730
rect 382772 223526 382828 223582
rect 388628 236994 388684 237050
rect 388820 236550 388876 236606
rect 388532 236254 388588 236310
rect 388724 236254 388780 236310
rect 386708 223378 386764 223434
rect 389012 236589 389014 236606
rect 389014 236589 389066 236606
rect 389066 236589 389068 236606
rect 389012 236550 389068 236589
rect 390356 236715 390412 236754
rect 390356 236698 390358 236715
rect 390358 236698 390410 236715
rect 390410 236698 390412 236715
rect 391604 226486 391660 226542
rect 394100 235218 394156 235274
rect 394484 235958 394540 236014
rect 393428 226634 393484 226690
rect 395348 235514 395404 235570
rect 395924 229002 395980 229058
rect 396788 226338 396844 226394
rect 397364 234330 397420 234386
rect 397364 232850 397420 232906
rect 397172 223230 397228 223286
rect 399092 235958 399148 236014
rect 398900 231814 398956 231870
rect 398804 229594 398860 229650
rect 400628 234626 400684 234682
rect 402164 235070 402220 235126
rect 402740 234330 402796 234386
rect 403220 235366 403276 235422
rect 403220 234922 403276 234978
rect 404372 234774 404428 234830
rect 405428 234922 405484 234978
rect 404756 234478 404812 234534
rect 404948 234478 405004 234534
rect 403988 228854 404044 228910
rect 405908 234626 405964 234682
rect 404756 222638 404812 222694
rect 408116 226190 408172 226246
rect 408500 226042 408556 226098
rect 409172 223082 409228 223138
rect 411380 235366 411436 235422
rect 411668 234034 411724 234090
rect 411668 228262 411724 228318
rect 413396 238918 413452 238974
rect 413684 238622 413740 238678
rect 413972 238326 414028 238382
rect 415700 228410 415756 228466
rect 415412 228262 415468 228318
rect 416948 234182 417004 234238
rect 430868 228558 430924 228614
rect 442868 231222 442924 231278
rect 439988 228706 440044 228762
rect 448916 231370 448972 231426
rect 458036 231518 458092 231574
rect 457268 225450 457324 225506
rect 464084 231666 464140 231722
rect 463316 225598 463372 225654
rect 471284 236106 471340 236162
rect 469364 225746 469420 225802
rect 472340 225894 472396 225950
rect 478388 227374 478444 227430
rect 484436 227226 484492 227282
rect 488276 233146 488332 233202
rect 490484 226930 490540 226986
rect 494228 232998 494284 233054
rect 495764 227078 495820 227134
rect 501044 234330 501100 234386
rect 504020 230334 504076 230390
rect 516212 234478 516268 234534
rect 516980 222786 517036 222842
rect 519188 230186 519244 230242
rect 521492 222934 521548 222990
rect 522932 226782 522988 226838
rect 525236 230038 525292 230094
rect 527540 224562 527596 224618
rect 528980 224414 529036 224470
rect 533492 229890 533548 229946
rect 532820 222638 532876 222694
rect 555380 238918 555436 238974
rect 553940 238326 553996 238382
rect 547124 224266 547180 224322
rect 547892 224118 547948 224174
rect 549428 229742 549484 229798
rect 557012 238622 557068 238678
rect 556148 236254 556204 236310
rect 555476 232702 555532 232758
rect 559892 235810 559948 235866
rect 557684 232554 557740 232610
rect 559220 223970 559276 224026
rect 576020 236994 576076 237050
rect 570260 236846 570316 236902
rect 567380 236698 567436 236754
rect 565268 236550 565324 236606
rect 562196 236402 562252 236458
rect 564404 235958 564460 236014
rect 565940 232850 565996 232906
rect 567476 232406 567532 232462
rect 569780 231962 569836 232018
rect 568244 223822 568300 223878
rect 570452 229446 570508 229502
rect 573524 232258 573580 232314
rect 572756 232110 572812 232166
rect 575060 229298 575116 229354
rect 574292 223526 574348 223582
rect 575828 223674 575884 223730
rect 579572 235662 579628 235718
rect 578900 229594 578956 229650
rect 576596 229150 576652 229206
rect 581780 223378 581836 223434
rect 588980 235514 589036 235570
rect 591668 226486 591724 226542
rect 596276 235218 596332 235274
rect 595412 226634 595468 226690
rect 599924 229002 599980 229058
rect 602228 226338 602284 226394
rect 605972 231814 606028 231870
rect 602996 223230 603052 223286
rect 609140 235366 609196 235422
rect 612788 235070 612844 235126
rect 618836 234922 618892 234978
rect 617300 234774 617356 234830
rect 616628 228854 616684 228910
rect 620372 234626 620428 234682
rect 621044 223082 621100 223138
rect 624884 226190 624940 226246
rect 625556 226042 625612 226098
rect 645140 221158 645196 221214
rect 645044 215830 645100 215886
rect 645140 212909 645142 212926
rect 645142 212909 645194 212926
rect 645194 212909 645196 212926
rect 645140 212870 645196 212909
rect 645140 209614 645196 209670
rect 645140 205914 645196 205970
rect 645140 201513 645142 201530
rect 645142 201513 645194 201530
rect 645194 201513 645196 201530
rect 645140 201474 645196 201513
rect 187220 199106 187276 199162
rect 645140 198218 645196 198274
rect 645140 193965 645142 193982
rect 645142 193965 645194 193982
rect 645194 193965 645196 193982
rect 645140 193926 645196 193965
rect 645140 190078 645196 190134
rect 646196 184306 646252 184362
rect 645908 182974 645964 183030
rect 646004 179274 646060 179330
rect 645140 174873 645142 174890
rect 645142 174873 645194 174890
rect 645194 174873 645196 174890
rect 645140 174834 645196 174873
rect 186164 174686 186220 174742
rect 185780 173206 185836 173262
rect 645140 170986 645196 171042
rect 645140 167730 645196 167786
rect 645524 161366 645580 161422
rect 645524 157518 645580 157574
rect 645140 155446 645196 155502
rect 646004 152525 646006 152542
rect 646006 152525 646058 152542
rect 646058 152525 646060 152542
rect 646004 152486 646060 152525
rect 645140 148046 645196 148102
rect 185780 146566 185836 146622
rect 646484 144198 646540 144254
rect 646580 140942 646636 140998
rect 184628 138278 184684 138334
rect 184340 137390 184396 137446
rect 184532 136798 184588 136854
rect 184436 135910 184492 135966
rect 184340 135209 184342 135226
rect 184342 135209 184394 135226
rect 184394 135209 184396 135226
rect 184340 135170 184396 135209
rect 184436 134430 184492 134486
rect 184340 133690 184396 133746
rect 184532 132950 184588 133006
rect 184340 132227 184396 132266
rect 184340 132210 184342 132227
rect 184342 132210 184394 132227
rect 184394 132210 184396 132227
rect 184436 131470 184492 131526
rect 184532 130582 184588 130638
rect 184628 129842 184684 129898
rect 184340 129102 184396 129158
rect 184436 128362 184492 128418
rect 184532 127622 184588 127678
rect 646580 128954 646636 129010
rect 184724 126882 184780 126938
rect 184340 125994 184396 126050
rect 646868 134726 646924 134782
rect 647828 130878 647884 130934
rect 646772 127622 646828 127678
rect 646676 125698 646732 125754
rect 186836 125402 186892 125458
rect 184436 124514 184492 124570
rect 184340 123774 184396 123830
rect 184436 122146 184492 122202
rect 184628 123034 184684 123090
rect 647732 121998 647788 122054
rect 184532 121554 184588 121610
rect 184340 120666 184396 120722
rect 184532 120074 184588 120130
rect 184628 119186 184684 119242
rect 184436 118594 184492 118650
rect 184340 117706 184396 117762
rect 184436 116966 184492 117022
rect 652244 175870 652300 175926
rect 652628 277990 652684 278046
rect 652436 175722 652492 175778
rect 654452 909506 654508 909562
rect 654452 896186 654508 896242
rect 654452 869694 654508 869750
rect 654452 856374 654508 856430
rect 654452 842906 654508 842962
rect 654740 829734 654796 829790
rect 654452 803094 654508 803150
rect 654452 763299 654508 763338
rect 654452 763282 654454 763299
rect 654454 763282 654506 763299
rect 654506 763282 654508 763299
rect 654452 750110 654508 750166
rect 654452 736790 654508 736846
rect 654452 710315 654508 710354
rect 654452 710298 654454 710315
rect 654454 710298 654506 710315
rect 654506 710298 654508 710315
rect 654452 696995 654508 697034
rect 654452 696978 654454 696995
rect 654454 696978 654506 696995
rect 654506 696978 654508 696995
rect 654452 683510 654508 683566
rect 654452 657018 654508 657074
rect 654452 643698 654508 643754
rect 654452 630526 654508 630582
rect 654548 617206 654604 617262
rect 654452 603886 654508 603942
rect 654452 590714 654508 590770
rect 654452 577394 654508 577450
rect 654836 550902 654892 550958
rect 654452 537582 654508 537638
rect 654452 524279 654508 524318
rect 654452 524262 654454 524279
rect 654454 524262 654506 524279
rect 654506 524262 654508 524279
rect 654452 510942 654508 510998
rect 654452 497622 654508 497678
rect 654452 484302 654508 484358
rect 654452 471130 654508 471186
rect 654452 457810 654508 457866
rect 654452 444490 654508 444546
rect 654452 431318 654508 431374
rect 654452 417998 654508 418054
rect 654452 404678 654508 404734
rect 654836 391506 654892 391562
rect 654452 378186 654508 378242
rect 654452 364883 654508 364922
rect 654452 364866 654454 364883
rect 654454 364866 654506 364883
rect 654506 364866 654508 364883
rect 654452 351546 654508 351602
rect 654836 324906 654892 324962
rect 654452 311734 654508 311790
rect 655220 975810 655276 975866
rect 655220 776602 655276 776658
rect 655220 723470 655276 723526
rect 655124 311142 655180 311198
rect 655124 298414 655180 298470
rect 655508 962490 655564 962546
rect 655700 949318 655756 949374
rect 655604 936146 655660 936202
rect 656372 922678 656428 922734
rect 656564 882866 656620 882922
rect 655508 816414 655564 816470
rect 655604 789922 655660 789978
rect 655508 670338 655564 670394
rect 656564 564074 656620 564130
rect 655316 338226 655372 338282
rect 655412 285242 655468 285298
rect 658196 264966 658252 265022
rect 658100 221750 658156 221806
rect 658004 218938 658060 218994
rect 658388 265114 658444 265170
rect 661172 625050 661228 625106
rect 660980 310994 661036 311050
rect 667988 625050 668044 625106
rect 666836 624162 666892 624218
rect 647924 123774 647980 123830
rect 647924 119482 647980 119538
rect 646676 117558 646732 117614
rect 184628 116226 184684 116282
rect 647924 115634 647980 115690
rect 184532 115338 184588 115394
rect 184340 114746 184396 114802
rect 184436 113858 184492 113914
rect 184532 113118 184588 113174
rect 646580 113118 646636 113174
rect 184628 112378 184684 112434
rect 184436 111638 184492 111694
rect 184340 110898 184396 110954
rect 184532 110158 184588 110214
rect 184436 108678 184492 108734
rect 184340 107790 184396 107846
rect 184532 107050 184588 107106
rect 184436 106310 184492 106366
rect 184340 105570 184396 105626
rect 184532 104830 184588 104886
rect 645908 106014 645964 106070
rect 184628 103942 184684 103998
rect 184340 103389 184342 103406
rect 184342 103389 184394 103406
rect 184394 103389 184396 103406
rect 184340 103350 184396 103389
rect 184532 102462 184588 102518
rect 184436 101870 184492 101926
rect 645140 102166 645196 102222
rect 149684 100834 149740 100890
rect 184628 100982 184684 101038
rect 184340 100242 184396 100298
rect 184436 99502 184492 99558
rect 184532 98614 184588 98670
rect 184628 98022 184684 98078
rect 184340 97134 184396 97190
rect 184436 96394 184492 96450
rect 645428 95967 645484 96006
rect 645428 95950 645430 95967
rect 645430 95950 645482 95967
rect 645482 95950 645484 95967
rect 184532 95654 184588 95710
rect 184340 94931 184396 94970
rect 184340 94914 184342 94931
rect 184342 94914 184394 94931
rect 184394 94914 184396 94931
rect 184532 94174 184588 94230
rect 184436 93434 184492 93490
rect 184340 92694 184396 92750
rect 184340 91845 184342 91862
rect 184342 91845 184394 91862
rect 184394 91845 184396 91862
rect 184340 91806 184396 91845
rect 184436 91066 184492 91122
rect 184532 90326 184588 90382
rect 184628 89586 184684 89642
rect 184340 88846 184396 88902
rect 184532 88106 184588 88162
rect 184436 87218 184492 87274
rect 184628 86626 184684 86682
rect 184340 85738 184396 85794
rect 184436 85146 184492 85202
rect 184532 84258 184588 84314
rect 184340 83387 184396 83426
rect 184340 83370 184342 83387
rect 184342 83370 184394 83387
rect 184394 83370 184396 83387
rect 149588 82334 149644 82390
rect 149108 76710 149164 76766
rect 149012 73010 149068 73066
rect 149396 75526 149452 75582
rect 149204 71974 149260 72030
rect 149396 70790 149452 70846
rect 149300 69458 149356 69514
rect 184532 82778 184588 82834
rect 184436 81890 184492 81946
rect 184628 81298 184684 81354
rect 184340 80410 184396 80466
rect 184436 79818 184492 79874
rect 149684 79226 149740 79282
rect 149588 73750 149644 73806
rect 184628 78930 184684 78986
rect 184532 78190 184588 78246
rect 184436 77450 184492 77506
rect 184532 76710 184588 76766
rect 184340 75970 184396 76026
rect 184628 75082 184684 75138
rect 184340 74342 184396 74398
rect 184436 73602 184492 73658
rect 184532 72862 184588 72918
rect 184628 72122 184684 72178
rect 184340 71382 184396 71438
rect 184436 70494 184492 70550
rect 184532 69902 184588 69958
rect 184340 69053 184342 69070
rect 184342 69053 184394 69070
rect 184394 69053 184396 69070
rect 184340 69014 184396 69053
rect 184340 68422 184396 68478
rect 149588 68274 149644 68330
rect 149492 67090 149548 67146
rect 149396 64574 149452 64630
rect 149300 63390 149356 63446
rect 184532 67534 184588 67590
rect 184436 66794 184492 66850
rect 184340 66071 184396 66110
rect 184340 66054 184342 66071
rect 184342 66054 184394 66071
rect 184394 66054 184396 66071
rect 149684 65314 149740 65370
rect 184532 65166 184588 65222
rect 184628 64574 184684 64630
rect 184436 63686 184492 63742
rect 184340 63133 184342 63150
rect 184342 63133 184394 63150
rect 184394 63133 184396 63150
rect 184340 63094 184396 63133
rect 149396 62206 149452 62262
rect 184436 62206 184492 62262
rect 184628 61466 184684 61522
rect 184532 60726 184588 60782
rect 149492 60578 149548 60634
rect 184340 59986 184396 60042
rect 149396 59690 149452 59746
rect 184436 59246 184492 59302
rect 149396 58506 149452 58562
rect 184532 58358 184588 58414
rect 184340 57618 184396 57674
rect 149492 57322 149548 57378
rect 149396 56177 149398 56194
rect 149398 56177 149450 56194
rect 149450 56177 149452 56194
rect 149396 56138 149452 56177
rect 184340 56878 184396 56934
rect 184340 56155 184396 56194
rect 184340 56138 184342 56155
rect 184342 56138 184394 56155
rect 184394 56138 184396 56155
rect 184436 55398 184492 55454
rect 149684 54806 149740 54862
rect 184340 54675 184396 54714
rect 184340 54658 184342 54675
rect 184342 54658 184394 54675
rect 184394 54658 184396 54675
rect 184340 53918 184396 53974
rect 149396 53770 149452 53826
rect 187604 41782 187660 41838
rect 194324 41782 194380 41838
rect 302900 41782 302956 41838
rect 307220 41782 307276 41838
rect 357716 42078 357772 42134
rect 337460 40898 337516 40954
rect 331220 40746 331276 40802
rect 216404 40348 216460 40404
rect 142292 40154 142348 40210
rect 406772 47406 406828 47462
rect 419732 47554 419788 47610
rect 415508 41930 415564 41986
rect 434900 41930 434956 41986
rect 416852 41782 416908 41838
rect 420692 40598 420748 40654
rect 474452 47406 474508 47462
rect 470324 41782 470380 41838
rect 492980 47554 493036 47610
rect 493940 40746 493996 40802
rect 506804 40154 506860 40210
rect 518708 41782 518764 41838
rect 520340 41782 520396 41838
rect 562484 47406 562540 47462
rect 645908 88846 645964 88902
rect 645908 84406 645964 84462
rect 645524 79374 645580 79430
rect 646004 75526 646060 75582
rect 646004 66219 646060 66258
rect 646004 66202 646006 66219
rect 646006 66202 646058 66219
rect 646058 66202 646060 66219
rect 646004 58950 646060 59006
rect 647060 111342 647116 111398
rect 646676 109418 646732 109474
rect 646772 107938 646828 107994
rect 646964 98022 647020 98078
rect 669620 356134 669676 356190
rect 675380 966190 675436 966246
rect 675476 965746 675532 965802
rect 675476 965006 675532 965062
rect 675380 963378 675436 963434
rect 675476 962638 675532 962694
rect 675764 962194 675820 962250
rect 675476 959086 675532 959142
rect 675764 958346 675820 958402
rect 675380 957606 675436 957662
rect 675764 957014 675820 957070
rect 675572 955978 675628 956034
rect 675476 953906 675532 953962
rect 674708 953314 674764 953370
rect 675764 951982 675820 952038
rect 676148 941030 676204 941086
rect 676052 939737 676054 939754
rect 676054 939737 676106 939754
rect 676106 939737 676108 939754
rect 676052 939698 676108 939737
rect 676052 939254 676108 939310
rect 676340 940438 676396 940494
rect 676244 939994 676300 940050
rect 669812 357022 669868 357078
rect 676244 938849 676246 938866
rect 676246 938849 676298 938866
rect 676298 938849 676300 938866
rect 676244 938810 676300 938849
rect 676244 938087 676300 938126
rect 676244 938070 676246 938087
rect 676246 938070 676298 938087
rect 676298 938070 676300 938087
rect 676052 937739 676054 937756
rect 676054 937739 676106 937756
rect 676106 937739 676108 937756
rect 676052 937700 676108 937739
rect 676052 937199 676108 937238
rect 676052 937182 676054 937199
rect 676054 937182 676106 937199
rect 676106 937182 676108 937199
rect 679796 929486 679852 929542
rect 679796 928894 679852 928950
rect 685460 928894 685516 928950
rect 685460 928450 685516 928506
rect 672500 624162 672556 624218
rect 669908 278434 669964 278490
rect 669716 278138 669772 278194
rect 675284 876354 675340 876410
rect 675284 876206 675340 876262
rect 675476 873986 675532 874042
rect 675380 869842 675436 869898
rect 675764 864662 675820 864718
rect 675380 862886 675436 862942
rect 675380 787850 675436 787906
rect 675380 786666 675436 786722
rect 675476 784742 675532 784798
rect 674612 777490 674668 777546
rect 675764 780598 675820 780654
rect 675764 779118 675820 779174
rect 675764 777342 675820 777398
rect 675764 775418 675820 775474
rect 674228 774826 674284 774882
rect 675476 773642 675532 773698
rect 676052 762877 676054 762894
rect 676054 762877 676106 762894
rect 676106 762877 676108 762894
rect 676052 762838 676108 762877
rect 676052 762285 676054 762302
rect 676054 762285 676106 762302
rect 676106 762285 676108 762302
rect 676052 762246 676108 762285
rect 676244 761989 676246 762006
rect 676246 761989 676298 762006
rect 676298 761989 676300 762006
rect 676244 761950 676300 761989
rect 676244 761545 676246 761562
rect 676246 761545 676298 761562
rect 676298 761545 676300 761562
rect 676244 761506 676300 761545
rect 676244 760635 676300 760674
rect 676244 760618 676246 760635
rect 676246 760618 676298 760635
rect 676298 760618 676300 760635
rect 676052 760287 676054 760304
rect 676054 760287 676106 760304
rect 676106 760287 676108 760304
rect 676052 760248 676108 760287
rect 676052 759895 676108 759934
rect 676052 759878 676054 759895
rect 676054 759878 676106 759895
rect 676106 759878 676108 759895
rect 676052 759325 676054 759342
rect 676054 759325 676106 759342
rect 676106 759325 676108 759342
rect 676052 759286 676108 759325
rect 676052 758807 676054 758824
rect 676054 758807 676106 758824
rect 676106 758807 676108 758824
rect 676052 758768 676108 758807
rect 676052 755403 676054 755420
rect 676054 755403 676106 755420
rect 676106 755403 676108 755420
rect 676052 755364 676108 755403
rect 676244 755033 676246 755050
rect 676246 755033 676298 755050
rect 676298 755033 676300 755050
rect 676244 754994 676300 755033
rect 676052 754293 676054 754310
rect 676054 754293 676106 754310
rect 676106 754293 676108 754310
rect 676052 754254 676108 754293
rect 676052 752813 676054 752830
rect 676054 752813 676106 752830
rect 676106 752813 676108 752830
rect 676052 752774 676108 752813
rect 676052 752369 676054 752386
rect 676054 752369 676106 752386
rect 676106 752369 676108 752386
rect 676052 752330 676108 752369
rect 676052 751851 676054 751868
rect 676054 751851 676106 751868
rect 676106 751851 676108 751868
rect 676052 751812 676108 751851
rect 679796 751442 679852 751498
rect 679796 750554 679852 750610
rect 685460 750554 685516 750610
rect 685460 750110 685516 750166
rect 675380 743154 675436 743210
rect 675764 742118 675820 742174
rect 675380 741674 675436 741730
rect 675476 740342 675532 740398
rect 675668 735458 675724 735514
rect 675764 734422 675820 734478
rect 676244 718033 676246 718050
rect 676246 718033 676298 718050
rect 676298 718033 676300 718050
rect 676244 717994 676300 718033
rect 676052 717293 676054 717310
rect 676054 717293 676106 717310
rect 676106 717293 676108 717310
rect 676052 717254 676108 717293
rect 676244 716997 676246 717014
rect 676246 716997 676298 717014
rect 676298 716997 676300 717014
rect 676244 716958 676300 716997
rect 679700 716514 679756 716570
rect 679700 715478 679756 715534
rect 676052 715295 676054 715312
rect 676054 715295 676106 715312
rect 676106 715295 676108 715312
rect 676052 715256 676108 715295
rect 676052 714903 676108 714942
rect 676052 714886 676054 714903
rect 676054 714886 676106 714903
rect 676106 714886 676108 714903
rect 676052 714333 676054 714350
rect 676054 714333 676106 714350
rect 676106 714333 676108 714350
rect 676052 714294 676108 714333
rect 676052 713741 676054 713758
rect 676054 713741 676106 713758
rect 676106 713741 676108 713758
rect 676052 713702 676108 713741
rect 676052 710411 676054 710428
rect 676054 710411 676106 710428
rect 676106 710411 676108 710428
rect 676052 710372 676108 710411
rect 676244 710041 676246 710058
rect 676246 710041 676298 710058
rect 676298 710041 676300 710058
rect 676244 710002 676300 710041
rect 676052 709301 676054 709318
rect 676054 709301 676106 709318
rect 676106 709301 676108 709318
rect 676052 709262 676108 709301
rect 676244 707969 676246 707986
rect 676246 707969 676298 707986
rect 676298 707969 676300 707986
rect 676244 707930 676300 707969
rect 676052 707377 676054 707394
rect 676054 707377 676106 707394
rect 676106 707377 676108 707394
rect 676052 707338 676108 707377
rect 676052 706859 676054 706876
rect 676054 706859 676106 706876
rect 676106 706859 676108 706876
rect 676052 706820 676108 706859
rect 679988 706450 680044 706506
rect 679796 705562 679852 705618
rect 679988 705562 680044 705618
rect 679796 705118 679852 705174
rect 675380 697866 675436 697922
rect 675764 697274 675820 697330
rect 675572 696830 675628 696886
rect 675380 694758 675436 694814
rect 675764 694166 675820 694222
rect 675476 690466 675532 690522
rect 675764 687358 675820 687414
rect 676052 672671 676054 672688
rect 676054 672671 676106 672688
rect 676106 672671 676108 672688
rect 676052 672632 676108 672671
rect 676244 672301 676246 672318
rect 676246 672301 676298 672318
rect 676298 672301 676300 672318
rect 676244 672262 676300 672301
rect 676052 671561 676054 671578
rect 676054 671561 676106 671578
rect 676106 671561 676108 671578
rect 676052 671522 676108 671561
rect 676052 671191 676054 671208
rect 676054 671191 676106 671208
rect 676106 671191 676108 671208
rect 676052 671152 676108 671191
rect 676052 670651 676108 670690
rect 676052 670634 676054 670651
rect 676054 670634 676106 670651
rect 676106 670634 676108 670651
rect 676052 670081 676054 670098
rect 676054 670081 676106 670098
rect 676106 670081 676108 670098
rect 676052 670042 676108 670081
rect 676052 669615 676108 669654
rect 676052 669598 676054 669615
rect 676054 669598 676106 669615
rect 676106 669598 676108 669615
rect 676244 669341 676246 669358
rect 676246 669341 676298 669358
rect 676298 669341 676300 669358
rect 676244 669302 676300 669341
rect 679892 668858 679948 668914
rect 676052 667600 676108 667656
rect 676244 665750 676300 665806
rect 676052 664605 676054 664622
rect 676054 664605 676106 664622
rect 676106 664605 676108 664622
rect 676052 664566 676108 664605
rect 676244 664309 676246 664326
rect 676246 664309 676298 664326
rect 676298 664309 676300 664326
rect 676244 664270 676300 664309
rect 676244 663865 676246 663882
rect 676246 663865 676298 663882
rect 676298 663865 676300 663882
rect 676244 663826 676300 663865
rect 676052 662607 676054 662624
rect 676054 662607 676106 662624
rect 676106 662607 676108 662624
rect 676052 662568 676108 662607
rect 676052 662237 676054 662254
rect 676054 662237 676106 662254
rect 676106 662237 676108 662254
rect 676052 662198 676108 662237
rect 676052 661645 676054 661662
rect 676054 661645 676106 661662
rect 676106 661645 676108 661662
rect 676052 661606 676108 661645
rect 679796 660866 679852 660922
rect 679796 660422 679852 660478
rect 685556 660422 685612 660478
rect 685556 659830 685612 659886
rect 675380 652578 675436 652634
rect 675380 651542 675436 651598
rect 675668 649618 675724 649674
rect 675476 645326 675532 645382
rect 675764 640294 675820 640350
rect 675476 638518 675532 638574
rect 676052 627679 676054 627696
rect 676054 627679 676106 627696
rect 676106 627679 676108 627696
rect 676052 627640 676108 627679
rect 676244 627309 676246 627326
rect 676246 627309 676298 627326
rect 676298 627309 676300 627326
rect 676244 627270 676300 627309
rect 676052 626569 676054 626586
rect 676054 626569 676106 626586
rect 676106 626569 676108 626586
rect 676052 626530 676108 626569
rect 679700 626382 679756 626438
rect 676052 625659 676108 625698
rect 676052 625642 676054 625659
rect 676054 625642 676106 625659
rect 676106 625642 676108 625659
rect 675956 624645 675958 624662
rect 675958 624645 676010 624662
rect 676010 624645 676012 624662
rect 675956 624606 676012 624645
rect 675956 623587 676012 623626
rect 675956 623570 675958 623587
rect 675958 623570 676010 623587
rect 676010 623570 676012 623587
rect 676052 622608 676108 622664
rect 676244 620758 676300 620814
rect 676052 619169 676054 619186
rect 676054 619169 676106 619186
rect 676106 619169 676108 619186
rect 676052 619130 676108 619169
rect 676052 618133 676054 618150
rect 676054 618133 676106 618150
rect 676106 618133 676108 618150
rect 676052 618094 676108 618133
rect 676052 617615 676054 617632
rect 676054 617615 676106 617632
rect 676106 617615 676108 617632
rect 676052 617576 676108 617615
rect 676244 617393 676246 617410
rect 676246 617393 676298 617410
rect 676298 617393 676300 617410
rect 676244 617354 676300 617393
rect 676052 616653 676054 616670
rect 676054 616653 676106 616670
rect 676106 616653 676108 616670
rect 676052 616614 676108 616653
rect 679796 615874 679852 615930
rect 679796 615282 679852 615338
rect 685460 615282 685516 615338
rect 685460 614838 685516 614894
rect 675380 607734 675436 607790
rect 675380 606402 675436 606458
rect 675380 604774 675436 604830
rect 675476 600186 675532 600242
rect 675764 595302 675820 595358
rect 675476 593378 675532 593434
rect 676052 582465 676054 582482
rect 676054 582465 676106 582482
rect 676106 582465 676108 582482
rect 676052 582426 676108 582465
rect 676052 581947 676054 581964
rect 676054 581947 676106 581964
rect 676106 581947 676108 581964
rect 676052 581908 676108 581947
rect 676244 581577 676246 581594
rect 676246 581577 676298 581594
rect 676298 581577 676300 581594
rect 676244 581538 676300 581577
rect 676052 580985 676054 581002
rect 676054 580985 676106 581002
rect 676106 580985 676108 581002
rect 676052 580946 676108 580985
rect 676244 580223 676300 580262
rect 676244 580206 676246 580223
rect 676246 580206 676298 580223
rect 676298 580206 676300 580223
rect 676052 579949 676054 579966
rect 676054 579949 676106 579966
rect 676106 579949 676108 579966
rect 676052 579910 676108 579949
rect 676052 579483 676108 579522
rect 676052 579466 676054 579483
rect 676054 579466 676106 579483
rect 676106 579466 676108 579483
rect 676052 578913 676054 578930
rect 676054 578913 676106 578930
rect 676106 578913 676108 578930
rect 676052 578874 676108 578913
rect 676052 578395 676054 578412
rect 676054 578395 676106 578412
rect 676106 578395 676108 578412
rect 676052 578356 676108 578395
rect 676052 574991 676054 575008
rect 676054 574991 676106 575008
rect 676106 574991 676108 575008
rect 676052 574952 676108 574991
rect 676244 574621 676246 574638
rect 676246 574621 676298 574638
rect 676298 574621 676300 574638
rect 676244 574582 676300 574621
rect 676052 573881 676054 573898
rect 676054 573881 676106 573898
rect 676106 573881 676108 573898
rect 676052 573842 676108 573881
rect 676052 573511 676054 573528
rect 676054 573511 676106 573528
rect 676106 573511 676108 573528
rect 676052 573472 676108 573511
rect 676052 572993 676054 573010
rect 676054 572993 676106 573010
rect 676106 572993 676108 573010
rect 676052 572954 676108 572993
rect 676052 572401 676054 572418
rect 676054 572401 676106 572418
rect 676106 572401 676108 572418
rect 676052 572362 676108 572401
rect 676052 571957 676054 571974
rect 676054 571957 676106 571974
rect 676106 571957 676108 571974
rect 676052 571918 676108 571957
rect 676244 571661 676246 571678
rect 676246 571661 676298 571678
rect 676298 571661 676300 571678
rect 676244 571622 676300 571661
rect 679988 571178 680044 571234
rect 679796 570142 679852 570198
rect 679988 570142 680044 570198
rect 679796 569698 679852 569754
rect 675476 562594 675532 562650
rect 675476 561706 675532 561762
rect 675476 561410 675532 561466
rect 675764 557562 675820 557618
rect 676052 537473 676054 537490
rect 676054 537473 676106 537490
rect 676106 537473 676108 537490
rect 676052 537434 676108 537473
rect 676052 536881 676054 536898
rect 676054 536881 676106 536898
rect 676106 536881 676108 536898
rect 676052 536842 676108 536881
rect 676244 536585 676246 536602
rect 676246 536585 676298 536602
rect 676298 536585 676300 536602
rect 676244 536546 676300 536585
rect 676532 535214 676588 535270
rect 676052 534883 676054 534900
rect 676054 534883 676106 534900
rect 676106 534883 676108 534900
rect 676052 534844 676108 534883
rect 676052 533921 676054 533938
rect 676054 533921 676106 533938
rect 676106 533921 676108 533938
rect 676052 533882 676108 533921
rect 676052 529999 676054 530016
rect 676054 529999 676106 530016
rect 676106 529999 676108 530016
rect 676052 529960 676108 529999
rect 676244 529629 676246 529646
rect 676246 529629 676298 529646
rect 676298 529629 676300 529646
rect 676244 529590 676300 529629
rect 676052 528889 676054 528906
rect 676054 528889 676106 528906
rect 676106 528889 676108 528906
rect 676052 528850 676108 528889
rect 676052 528445 676054 528462
rect 676054 528445 676106 528462
rect 676106 528445 676108 528462
rect 676052 528406 676108 528445
rect 676244 528149 676246 528166
rect 676246 528149 676298 528166
rect 676298 528149 676300 528166
rect 676244 528110 676300 528149
rect 676052 527409 676054 527426
rect 676054 527409 676106 527426
rect 676106 527409 676108 527426
rect 676052 527370 676108 527409
rect 676052 526965 676054 526982
rect 676054 526965 676106 526982
rect 676106 526965 676108 526982
rect 676052 526926 676108 526965
rect 676244 526669 676246 526686
rect 676246 526669 676298 526686
rect 676298 526669 676300 526686
rect 676244 526630 676300 526669
rect 676628 534178 676684 534234
rect 676244 493665 676246 493682
rect 676246 493665 676298 493682
rect 676298 493665 676300 493682
rect 676244 493626 676300 493665
rect 676052 492925 676054 492942
rect 676054 492925 676106 492942
rect 676106 492925 676108 492942
rect 676052 492886 676108 492925
rect 676052 492333 676054 492350
rect 676054 492333 676106 492350
rect 676106 492333 676108 492350
rect 676052 492294 676108 492333
rect 676532 491554 676588 491610
rect 676148 488594 676204 488650
rect 676052 487410 676108 487466
rect 676244 487114 676300 487170
rect 676244 486561 676246 486578
rect 676246 486561 676298 486578
rect 676298 486561 676300 486578
rect 676244 486522 676300 486561
rect 676052 485412 676108 485468
rect 676244 485081 676246 485098
rect 676246 485081 676298 485098
rect 676298 485081 676300 485098
rect 676244 485042 676300 485081
rect 676052 484489 676054 484506
rect 676054 484489 676106 484506
rect 676106 484489 676108 484506
rect 676052 484450 676108 484489
rect 676052 483971 676054 483988
rect 676054 483971 676106 483988
rect 676106 483971 676108 483988
rect 676052 483932 676108 483971
rect 676052 483009 676054 483026
rect 676054 483009 676106 483026
rect 676106 483009 676108 483026
rect 676052 482970 676108 483009
rect 676052 482417 676054 482434
rect 676054 482417 676106 482434
rect 676106 482417 676108 482434
rect 676052 482378 676108 482417
rect 670292 278582 670348 278638
rect 670100 278286 670156 278342
rect 676244 405457 676246 405474
rect 676246 405457 676298 405474
rect 676298 405457 676300 405474
rect 676244 405418 676300 405457
rect 676052 404717 676054 404734
rect 676054 404717 676106 404734
rect 676106 404717 676108 404734
rect 676052 404678 676108 404717
rect 676052 404199 676054 404216
rect 676054 404199 676106 404216
rect 676106 404199 676108 404216
rect 676052 404160 676108 404199
rect 679700 536102 679756 536158
rect 676724 533142 676780 533198
rect 676628 491110 676684 491166
rect 676628 490222 676684 490278
rect 679796 526038 679852 526094
rect 679796 525150 679852 525206
rect 685460 525150 685516 525206
rect 685460 524706 685516 524762
rect 679700 492146 679756 492202
rect 676724 490074 676780 490130
rect 676628 489186 676684 489242
rect 676532 403938 676588 403994
rect 676052 403237 676054 403254
rect 676054 403237 676106 403254
rect 676106 403237 676108 403254
rect 676052 403198 676108 403237
rect 676052 402253 676108 402292
rect 676052 402236 676054 402253
rect 676054 402236 676106 402253
rect 676106 402236 676108 402253
rect 679988 481638 680044 481694
rect 679796 481194 679852 481250
rect 679988 481194 680044 481250
rect 679796 480750 679852 480806
rect 676724 402902 676780 402958
rect 676052 401718 676108 401774
rect 676244 400995 676300 401034
rect 676244 400978 676246 400995
rect 676246 400978 676298 400995
rect 676298 400978 676300 400995
rect 676052 395741 676108 395780
rect 676052 395724 676054 395741
rect 676054 395724 676106 395741
rect 676106 395724 676108 395741
rect 676244 394039 676300 394078
rect 676244 394022 676246 394039
rect 676246 394022 676298 394039
rect 676298 394022 676300 394039
rect 679796 393430 679852 393486
rect 679796 392986 679852 393042
rect 685556 392986 685612 393042
rect 685556 392542 685612 392598
rect 675764 385882 675820 385938
rect 675764 385586 675820 385642
rect 675764 384698 675820 384754
rect 675380 382922 675436 382978
rect 675284 382774 675340 382830
rect 675476 382182 675532 382238
rect 675764 381146 675820 381202
rect 675476 378778 675532 378834
rect 675764 377890 675820 377946
rect 675764 375670 675820 375726
rect 675188 373746 675244 373802
rect 675572 371970 675628 372026
rect 676052 360021 676054 360038
rect 676054 360021 676106 360038
rect 676106 360021 676108 360038
rect 676052 359982 676108 360021
rect 676244 359725 676246 359742
rect 676246 359725 676298 359742
rect 676298 359725 676300 359742
rect 676244 359686 676300 359725
rect 676052 358985 676054 359002
rect 676054 358985 676106 359002
rect 676106 358985 676108 359002
rect 676052 358946 676108 358985
rect 676052 358541 676054 358558
rect 676054 358541 676106 358558
rect 676106 358541 676108 358558
rect 676052 358502 676108 358541
rect 676244 357614 676300 357670
rect 676052 356543 676054 356560
rect 676054 356543 676106 356560
rect 676106 356543 676108 356560
rect 676052 356504 676108 356543
rect 675764 354506 675820 354562
rect 675284 352582 675340 352638
rect 676052 354062 676108 354118
rect 676244 350362 676300 350418
rect 676244 349770 676300 349826
rect 676052 349622 676108 349678
rect 676052 349030 676108 349086
rect 679796 348290 679852 348346
rect 679796 347698 679852 347754
rect 685460 347698 685516 347754
rect 685460 347254 685516 347310
rect 675764 339558 675820 339614
rect 675476 337042 675532 337098
rect 675764 336450 675820 336506
rect 675380 333490 675436 333546
rect 675476 330530 675532 330586
rect 675380 328310 675436 328366
rect 675380 326830 675436 326886
rect 676052 315029 676054 315046
rect 676054 315029 676106 315046
rect 676106 315029 676108 315046
rect 676052 314990 676108 315029
rect 676244 314733 676246 314750
rect 676246 314733 676298 314750
rect 676298 314733 676300 314750
rect 676244 314694 676300 314733
rect 676052 313993 676054 314010
rect 676054 313993 676106 314010
rect 676106 313993 676108 314010
rect 676052 313954 676108 313993
rect 676052 310550 676108 310606
rect 676052 309514 676108 309570
rect 676052 307590 676108 307646
rect 676244 306850 676300 306906
rect 676244 306258 676300 306314
rect 676244 304778 676300 304834
rect 676052 304038 676108 304094
rect 679892 303298 679948 303354
rect 679892 302854 679948 302910
rect 679796 302706 679852 302762
rect 679796 302262 679852 302318
rect 675380 292790 675436 292846
rect 675476 288498 675532 288554
rect 675668 287758 675724 287814
rect 675476 287314 675532 287370
rect 675476 285242 675532 285298
rect 675380 283614 675436 283670
rect 675380 281838 675436 281894
rect 676052 270037 676054 270054
rect 676054 270037 676106 270054
rect 676106 270037 676108 270054
rect 676052 269998 676108 270037
rect 676244 269741 676246 269758
rect 676246 269741 676298 269758
rect 676298 269741 676300 269758
rect 676244 269702 676300 269741
rect 676244 269149 676246 269166
rect 676246 269149 676298 269166
rect 676298 269149 676300 269166
rect 676244 269110 676300 269149
rect 675668 264522 675724 264578
rect 675764 262598 675820 262654
rect 676244 261858 676300 261914
rect 676052 259564 676108 259620
rect 676052 259046 676108 259102
rect 679700 258306 679756 258362
rect 679700 257714 679756 257770
rect 685460 257714 685516 257770
rect 685460 257270 685516 257326
rect 675764 249574 675820 249630
rect 675668 247502 675724 247558
rect 675764 246614 675820 246670
rect 675764 245874 675820 245930
rect 675476 243506 675532 243562
rect 675284 241878 675340 241934
rect 675476 240546 675532 240602
rect 675284 238178 675340 238234
rect 675380 236846 675436 236902
rect 676244 225045 676246 225062
rect 676246 225045 676298 225062
rect 676298 225045 676300 225062
rect 676244 225006 676300 225045
rect 676052 224305 676054 224322
rect 676054 224305 676106 224322
rect 676106 224305 676108 224322
rect 676052 224266 676108 224305
rect 676052 223787 676054 223804
rect 676054 223787 676106 223804
rect 676106 223787 676108 223804
rect 676052 223748 676108 223787
rect 675764 219234 675820 219290
rect 676052 216866 676108 216922
rect 676052 215312 676108 215368
rect 676052 214794 676108 214850
rect 675956 213832 676012 213888
rect 676244 214202 676300 214258
rect 679796 213462 679852 213518
rect 679796 212574 679852 212630
rect 685460 212574 685516 212630
rect 685460 212130 685516 212186
rect 675764 205026 675820 205082
rect 675476 204286 675532 204342
rect 675764 202658 675820 202714
rect 675764 201326 675820 201382
rect 675476 198366 675532 198422
rect 675476 195258 675532 195314
rect 675380 193482 675436 193538
rect 675380 191558 675436 191614
rect 676244 179570 676300 179626
rect 676052 179313 676054 179330
rect 676054 179313 676106 179330
rect 676106 179313 676108 179330
rect 676052 179274 676108 179313
rect 676052 178795 676054 178812
rect 676054 178795 676106 178812
rect 676106 178795 676108 178812
rect 676052 178756 676108 178795
rect 676052 175352 676108 175408
rect 675380 174242 675436 174298
rect 676244 173650 676300 173706
rect 675476 172318 675532 172374
rect 676052 171874 676108 171930
rect 675956 171282 676012 171338
rect 676052 169802 676108 169858
rect 676244 168026 676300 168082
rect 676148 167582 676204 167638
rect 676244 167177 676246 167194
rect 676246 167177 676298 167194
rect 676298 167177 676300 167194
rect 676244 167138 676300 167177
rect 675188 158702 675244 158758
rect 675188 158406 675244 158462
rect 675476 153374 675532 153430
rect 675380 152486 675436 152542
rect 675476 151894 675532 151950
rect 675668 151302 675724 151358
rect 675476 150266 675532 150322
rect 675476 148490 675532 148546
rect 675380 146566 675436 146622
rect 676148 134430 676204 134486
rect 676052 132654 676108 132710
rect 676244 134321 676246 134338
rect 676246 134321 676298 134338
rect 676298 134321 676300 134338
rect 676244 134282 676300 134321
rect 676244 133394 676300 133450
rect 676244 131322 676300 131378
rect 676052 130582 676108 130638
rect 675476 129102 675532 129158
rect 669524 106310 669580 106366
rect 676052 127178 676108 127234
rect 676244 126438 676300 126494
rect 676052 126068 676108 126124
rect 676052 124588 676108 124644
rect 675956 124218 676012 124274
rect 676052 123626 676108 123682
rect 676340 122886 676396 122942
rect 676148 122442 676204 122498
rect 676244 121850 676300 121906
rect 675380 114302 675436 114358
rect 675380 112230 675436 112286
rect 675476 108086 675532 108142
rect 675380 106310 675436 106366
rect 668180 105274 668236 105330
rect 665300 105126 665356 105182
rect 647924 104090 647980 104146
rect 647924 99650 647980 99706
rect 647732 94026 647788 94082
rect 646868 68570 646924 68626
rect 647828 92694 647884 92750
rect 647924 87070 647980 87126
rect 650900 86182 650956 86238
rect 652340 85294 652396 85350
rect 651764 84258 651820 84314
rect 652244 83370 652300 83426
rect 647924 82630 647980 82686
rect 647924 81002 647980 81058
rect 647924 77489 647926 77506
rect 647926 77489 647978 77506
rect 647978 77489 647980 77506
rect 647924 77450 647980 77489
rect 647924 73602 647980 73658
rect 647156 71826 647212 71882
rect 647924 69623 647980 69662
rect 647924 69606 647926 69623
rect 647926 69606 647978 69623
rect 647978 69606 647980 69623
rect 647924 64130 647980 64186
rect 647924 62206 647980 62262
rect 647060 60282 647116 60338
rect 659348 90770 659404 90826
rect 675380 105126 675436 105182
rect 675668 103202 675724 103258
rect 675380 101426 675436 101482
rect 653684 86922 653740 86978
rect 663284 86330 663340 86386
rect 652436 82630 652492 82686
rect 662420 81611 662476 81650
rect 662420 81594 662422 81611
rect 662422 81594 662474 81611
rect 662474 81594 662476 81611
rect 663284 84702 663340 84758
rect 663476 83962 663532 84018
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 646772 57026 646828 57082
rect 646484 54658 646540 54714
rect 545204 40598 545260 40654
rect 633620 40450 633676 40506
<< metal3 >>
rect 148527 1016272 148593 1016275
rect 250479 1016272 250545 1016275
rect 353391 1016272 353457 1016275
rect 98370 1016212 99390 1016272
rect 94959 1005172 95025 1005175
rect 97167 1005172 97233 1005175
rect 94959 1005170 97233 1005172
rect 94959 1005114 94964 1005170
rect 95020 1005114 97172 1005170
rect 97228 1005114 97233 1005170
rect 94959 1005112 97233 1005114
rect 94959 1005109 95025 1005112
rect 97167 1005109 97233 1005112
rect 97935 1005172 98001 1005175
rect 98370 1005172 98430 1016212
rect 99330 1015946 99390 1016212
rect 148527 1016270 150750 1016272
rect 148527 1016214 148532 1016270
rect 148588 1016214 150750 1016270
rect 148527 1016212 150750 1016214
rect 148527 1016209 148593 1016212
rect 149730 1015946 149790 1016212
rect 150690 1015946 150750 1016212
rect 200610 1016212 201726 1016272
rect 200610 1015946 200670 1016212
rect 201666 1015946 201726 1016212
rect 250479 1016270 253566 1016272
rect 250479 1016214 250484 1016270
rect 250540 1016214 253566 1016270
rect 250479 1016212 253566 1016214
rect 250479 1016209 250545 1016212
rect 252546 1015946 252606 1016212
rect 253506 1015946 253566 1016212
rect 353391 1016270 355518 1016272
rect 353391 1016214 353396 1016270
rect 353452 1016214 355518 1016270
rect 353391 1016212 355518 1016214
rect 353391 1016209 353457 1016212
rect 354498 1015946 354558 1016212
rect 355458 1015946 355518 1016212
rect 421890 1016212 422910 1016272
rect 146607 1007984 146673 1007987
rect 148527 1007984 148593 1007987
rect 146607 1007982 148593 1007984
rect 146607 1007926 146612 1007982
rect 146668 1007926 148532 1007982
rect 148588 1007926 148593 1007982
rect 146607 1007924 148593 1007926
rect 146607 1007921 146673 1007924
rect 148527 1007921 148593 1007924
rect 351279 1007984 351345 1007987
rect 353391 1007984 353457 1007987
rect 351279 1007982 353457 1007984
rect 351279 1007926 351284 1007982
rect 351340 1007926 353396 1007982
rect 353452 1007926 353457 1007982
rect 351279 1007924 353457 1007926
rect 351279 1007921 351345 1007924
rect 353391 1007921 353457 1007924
rect 261327 1006504 261393 1006507
rect 261024 1006502 261393 1006504
rect 261024 1006446 261332 1006502
rect 261388 1006446 261393 1006502
rect 261024 1006444 261393 1006446
rect 261327 1006441 261393 1006444
rect 102447 1006208 102513 1006211
rect 102447 1006206 102816 1006208
rect 102447 1006150 102452 1006206
rect 102508 1006150 102816 1006206
rect 102447 1006148 102816 1006150
rect 102447 1006145 102513 1006148
rect 356367 1006060 356433 1006063
rect 357903 1006060 357969 1006063
rect 356064 1006058 356433 1006060
rect 356064 1006002 356372 1006058
rect 356428 1006002 356433 1006058
rect 356064 1006000 356433 1006002
rect 357600 1006058 357969 1006060
rect 357600 1006002 357908 1006058
rect 357964 1006002 357969 1006058
rect 357600 1006000 357969 1006002
rect 356367 1005997 356433 1006000
rect 357903 1005997 357969 1006000
rect 101007 1005912 101073 1005915
rect 262287 1005912 262353 1005915
rect 358767 1005912 358833 1005915
rect 359343 1005912 359409 1005915
rect 101007 1005910 101376 1005912
rect 101007 1005854 101012 1005910
rect 101068 1005854 101376 1005910
rect 101007 1005852 101376 1005854
rect 262080 1005910 262353 1005912
rect 262080 1005854 262292 1005910
rect 262348 1005854 262353 1005910
rect 262080 1005852 262353 1005854
rect 358560 1005910 358833 1005912
rect 358560 1005854 358772 1005910
rect 358828 1005854 358833 1005910
rect 358560 1005852 358833 1005854
rect 359040 1005910 359409 1005912
rect 359040 1005854 359348 1005910
rect 359404 1005854 359409 1005910
rect 359040 1005852 359409 1005854
rect 101007 1005849 101073 1005852
rect 262287 1005849 262353 1005852
rect 358767 1005849 358833 1005852
rect 359343 1005849 359409 1005852
rect 361839 1005764 361905 1005767
rect 361440 1005762 361905 1005764
rect 361440 1005706 361844 1005762
rect 361900 1005706 361905 1005762
rect 361440 1005704 361905 1005706
rect 361839 1005701 361905 1005704
rect 109935 1005616 110001 1005619
rect 110511 1005616 110577 1005619
rect 158511 1005616 158577 1005619
rect 356751 1005616 356817 1005619
rect 357135 1005616 357201 1005619
rect 358287 1005616 358353 1005619
rect 109935 1005614 110304 1005616
rect 109935 1005558 109940 1005614
rect 109996 1005558 110304 1005614
rect 109935 1005556 110304 1005558
rect 110511 1005614 110880 1005616
rect 110511 1005558 110516 1005614
rect 110572 1005558 110880 1005614
rect 110511 1005556 110880 1005558
rect 158208 1005614 158577 1005616
rect 158208 1005558 158516 1005614
rect 158572 1005558 158577 1005614
rect 158208 1005556 158577 1005558
rect 356640 1005614 356817 1005616
rect 356640 1005558 356756 1005614
rect 356812 1005558 356817 1005614
rect 356640 1005556 356817 1005558
rect 357024 1005614 357201 1005616
rect 357024 1005558 357140 1005614
rect 357196 1005558 357201 1005614
rect 357024 1005556 357201 1005558
rect 358080 1005614 358353 1005616
rect 358080 1005558 358292 1005614
rect 358348 1005558 358353 1005614
rect 358080 1005556 358353 1005558
rect 109935 1005553 110001 1005556
rect 110511 1005553 110577 1005556
rect 158511 1005553 158577 1005556
rect 356751 1005553 356817 1005556
rect 357135 1005553 357201 1005556
rect 358287 1005553 358353 1005556
rect 102063 1005468 102129 1005471
rect 161391 1005468 161457 1005471
rect 161871 1005468 161937 1005471
rect 207375 1005468 207441 1005471
rect 361263 1005468 361329 1005471
rect 102063 1005466 102240 1005468
rect 102063 1005410 102068 1005466
rect 102124 1005410 102240 1005466
rect 102063 1005408 102240 1005410
rect 161391 1005466 161760 1005468
rect 161391 1005410 161396 1005466
rect 161452 1005410 161760 1005466
rect 161391 1005408 161760 1005410
rect 161871 1005466 162240 1005468
rect 161871 1005410 161876 1005466
rect 161932 1005410 162240 1005466
rect 161871 1005408 162240 1005410
rect 207375 1005466 207648 1005468
rect 207375 1005410 207380 1005466
rect 207436 1005410 207648 1005466
rect 207375 1005408 207648 1005410
rect 361056 1005466 361329 1005468
rect 361056 1005410 361268 1005466
rect 361324 1005410 361329 1005466
rect 361056 1005408 361329 1005410
rect 102063 1005405 102129 1005408
rect 161391 1005405 161457 1005408
rect 161871 1005405 161937 1005408
rect 207375 1005405 207441 1005408
rect 361263 1005405 361329 1005408
rect 107055 1005320 107121 1005323
rect 159471 1005320 159537 1005323
rect 161487 1005320 161553 1005323
rect 210831 1005320 210897 1005323
rect 106848 1005318 107121 1005320
rect 106848 1005262 107060 1005318
rect 107116 1005262 107121 1005318
rect 106848 1005260 107121 1005262
rect 159264 1005318 159537 1005320
rect 159264 1005262 159476 1005318
rect 159532 1005262 159537 1005318
rect 159264 1005260 159537 1005262
rect 161184 1005318 161553 1005320
rect 161184 1005262 161492 1005318
rect 161548 1005262 161553 1005318
rect 161184 1005260 161553 1005262
rect 210720 1005318 210897 1005320
rect 210720 1005262 210836 1005318
rect 210892 1005262 210897 1005318
rect 210720 1005260 210897 1005262
rect 107055 1005257 107121 1005260
rect 159471 1005257 159537 1005260
rect 161487 1005257 161553 1005260
rect 210831 1005257 210897 1005260
rect 212847 1005320 212913 1005323
rect 313839 1005320 313905 1005323
rect 316431 1005320 316497 1005323
rect 360879 1005320 360945 1005323
rect 362319 1005320 362385 1005323
rect 212847 1005318 213120 1005320
rect 212847 1005262 212852 1005318
rect 212908 1005262 213120 1005318
rect 212847 1005260 213120 1005262
rect 313632 1005318 313905 1005320
rect 313632 1005262 313844 1005318
rect 313900 1005262 313905 1005318
rect 313632 1005260 313905 1005262
rect 316128 1005318 316497 1005320
rect 316128 1005262 316436 1005318
rect 316492 1005262 316497 1005318
rect 316128 1005260 316497 1005262
rect 360480 1005318 360945 1005320
rect 360480 1005262 360884 1005318
rect 360940 1005262 360945 1005318
rect 360480 1005260 360945 1005262
rect 362016 1005318 362385 1005320
rect 362016 1005262 362324 1005318
rect 362380 1005262 362385 1005318
rect 362016 1005260 362385 1005262
rect 212847 1005257 212913 1005260
rect 313839 1005257 313905 1005260
rect 316431 1005257 316497 1005260
rect 360879 1005257 360945 1005260
rect 362319 1005257 362385 1005260
rect 97935 1005170 98430 1005172
rect 97935 1005114 97940 1005170
rect 97996 1005142 98430 1005170
rect 105423 1005172 105489 1005175
rect 108015 1005172 108081 1005175
rect 160911 1005172 160977 1005175
rect 209871 1005172 209937 1005175
rect 105423 1005170 105888 1005172
rect 97996 1005114 98400 1005142
rect 97935 1005112 98400 1005114
rect 105423 1005114 105428 1005170
rect 105484 1005114 105888 1005170
rect 105423 1005112 105888 1005114
rect 107904 1005170 108081 1005172
rect 107904 1005114 108020 1005170
rect 108076 1005114 108081 1005170
rect 107904 1005112 108081 1005114
rect 160800 1005170 160977 1005172
rect 160800 1005114 160916 1005170
rect 160972 1005114 160977 1005170
rect 160800 1005112 160977 1005114
rect 209568 1005170 209937 1005172
rect 209568 1005114 209876 1005170
rect 209932 1005114 209937 1005170
rect 209568 1005112 209937 1005114
rect 97935 1005109 98001 1005112
rect 105423 1005109 105489 1005112
rect 108015 1005109 108081 1005112
rect 160911 1005109 160977 1005112
rect 209871 1005109 209937 1005112
rect 308271 1005172 308337 1005175
rect 312879 1005172 312945 1005175
rect 362799 1005172 362865 1005175
rect 308271 1005170 308640 1005172
rect 308271 1005114 308276 1005170
rect 308332 1005114 308640 1005170
rect 308271 1005112 308640 1005114
rect 312576 1005170 312945 1005172
rect 312576 1005114 312884 1005170
rect 312940 1005114 312945 1005170
rect 312576 1005112 312945 1005114
rect 362592 1005170 362865 1005172
rect 362592 1005114 362804 1005170
rect 362860 1005114 362865 1005170
rect 362592 1005112 362865 1005114
rect 308271 1005109 308337 1005112
rect 312879 1005109 312945 1005112
rect 362799 1005109 362865 1005112
rect 417519 1005172 417585 1005175
rect 420783 1005172 420849 1005175
rect 417519 1005170 420849 1005172
rect 417519 1005114 417524 1005170
rect 417580 1005114 420788 1005170
rect 420844 1005114 420849 1005170
rect 417519 1005112 420849 1005114
rect 417519 1005109 417585 1005112
rect 420783 1005109 420849 1005112
rect 421551 1005172 421617 1005175
rect 421890 1005172 421950 1016212
rect 422850 1015946 422910 1016212
rect 550338 1016212 551358 1016272
rect 550338 1015946 550398 1016212
rect 425679 1005912 425745 1005915
rect 429711 1005912 429777 1005915
rect 425472 1005910 425745 1005912
rect 425472 1005854 425684 1005910
rect 425740 1005854 425745 1005910
rect 425472 1005852 425745 1005854
rect 429408 1005910 429777 1005912
rect 429408 1005854 429716 1005910
rect 429772 1005854 429777 1005910
rect 551298 1005912 551358 1016212
rect 558159 1006060 558225 1006063
rect 557856 1006058 558225 1006060
rect 557856 1006002 558164 1006058
rect 558220 1006002 558225 1006058
rect 557856 1006000 558225 1006002
rect 558159 1005997 558225 1006000
rect 551631 1005912 551697 1005915
rect 551298 1005910 551697 1005912
rect 551298 1005882 551636 1005910
rect 429408 1005852 429777 1005854
rect 551328 1005854 551636 1005882
rect 551692 1005854 551697 1005910
rect 551328 1005852 551697 1005854
rect 425679 1005849 425745 1005852
rect 429711 1005849 429777 1005852
rect 551631 1005849 551697 1005852
rect 428271 1005764 428337 1005767
rect 428655 1005764 428721 1005767
rect 501711 1005764 501777 1005767
rect 502287 1005764 502353 1005767
rect 553647 1005764 553713 1005767
rect 554607 1005764 554673 1005767
rect 427968 1005762 428337 1005764
rect 427968 1005706 428276 1005762
rect 428332 1005706 428337 1005762
rect 427968 1005704 428337 1005706
rect 428448 1005762 428721 1005764
rect 428448 1005706 428660 1005762
rect 428716 1005706 428721 1005762
rect 428448 1005704 428721 1005706
rect 501408 1005762 501777 1005764
rect 501408 1005706 501716 1005762
rect 501772 1005706 501777 1005762
rect 501408 1005704 501777 1005706
rect 501984 1005762 502353 1005764
rect 501984 1005706 502292 1005762
rect 502348 1005706 502353 1005762
rect 501984 1005704 502353 1005706
rect 553344 1005762 553713 1005764
rect 553344 1005706 553652 1005762
rect 553708 1005706 553713 1005762
rect 553344 1005704 553713 1005706
rect 554304 1005762 554673 1005764
rect 554304 1005706 554612 1005762
rect 554668 1005706 554673 1005762
rect 554304 1005704 554673 1005706
rect 428271 1005701 428337 1005704
rect 428655 1005701 428721 1005704
rect 501711 1005701 501777 1005704
rect 502287 1005701 502353 1005704
rect 553647 1005701 553713 1005704
rect 554607 1005701 554673 1005704
rect 425295 1005616 425361 1005619
rect 426735 1005616 426801 1005619
rect 502671 1005616 502737 1005619
rect 554031 1005616 554097 1005619
rect 424992 1005614 425361 1005616
rect 424992 1005558 425300 1005614
rect 425356 1005558 425361 1005614
rect 424992 1005556 425361 1005558
rect 426432 1005614 426801 1005616
rect 426432 1005558 426740 1005614
rect 426796 1005558 426801 1005614
rect 426432 1005556 426801 1005558
rect 502464 1005614 502737 1005616
rect 502464 1005558 502676 1005614
rect 502732 1005558 502737 1005614
rect 502464 1005556 502737 1005558
rect 553920 1005614 554097 1005616
rect 553920 1005558 554036 1005614
rect 554092 1005558 554097 1005614
rect 553920 1005556 554097 1005558
rect 425295 1005553 425361 1005556
rect 426735 1005553 426801 1005556
rect 502671 1005553 502737 1005556
rect 554031 1005553 554097 1005556
rect 423759 1005468 423825 1005471
rect 424719 1005468 424785 1005471
rect 500751 1005468 500817 1005471
rect 503727 1005468 503793 1005471
rect 555183 1005468 555249 1005471
rect 423456 1005466 423825 1005468
rect 423456 1005410 423764 1005466
rect 423820 1005410 423825 1005466
rect 423456 1005408 423825 1005410
rect 424416 1005466 424785 1005468
rect 424416 1005410 424724 1005466
rect 424780 1005410 424785 1005466
rect 424416 1005408 424785 1005410
rect 500448 1005466 500817 1005468
rect 500448 1005410 500756 1005466
rect 500812 1005410 500817 1005466
rect 500448 1005408 500817 1005410
rect 503424 1005466 503793 1005468
rect 503424 1005410 503732 1005466
rect 503788 1005410 503793 1005466
rect 503424 1005408 503793 1005410
rect 554784 1005466 555249 1005468
rect 554784 1005410 555188 1005466
rect 555244 1005410 555249 1005466
rect 554784 1005408 555249 1005410
rect 423759 1005405 423825 1005408
rect 424719 1005405 424785 1005408
rect 500751 1005405 500817 1005408
rect 503727 1005405 503793 1005408
rect 555183 1005405 555249 1005408
rect 424143 1005320 424209 1005323
rect 426159 1005320 426225 1005323
rect 503247 1005320 503313 1005323
rect 505263 1005320 505329 1005323
rect 552207 1005320 552273 1005323
rect 552591 1005320 552657 1005323
rect 424032 1005318 424209 1005320
rect 424032 1005262 424148 1005318
rect 424204 1005262 424209 1005318
rect 424032 1005260 424209 1005262
rect 425952 1005318 426225 1005320
rect 425952 1005262 426164 1005318
rect 426220 1005262 426225 1005318
rect 425952 1005260 426225 1005262
rect 502944 1005318 503313 1005320
rect 502944 1005262 503252 1005318
rect 503308 1005262 503313 1005318
rect 502944 1005260 503313 1005262
rect 504960 1005318 505329 1005320
rect 504960 1005262 505268 1005318
rect 505324 1005262 505329 1005318
rect 504960 1005260 505329 1005262
rect 551904 1005318 552273 1005320
rect 551904 1005262 552212 1005318
rect 552268 1005262 552273 1005318
rect 551904 1005260 552273 1005262
rect 552384 1005318 552657 1005320
rect 552384 1005262 552596 1005318
rect 552652 1005262 552657 1005318
rect 552384 1005260 552657 1005262
rect 424143 1005257 424209 1005260
rect 426159 1005257 426225 1005260
rect 503247 1005257 503313 1005260
rect 505263 1005257 505329 1005260
rect 552207 1005257 552273 1005260
rect 552591 1005257 552657 1005260
rect 501135 1005172 501201 1005175
rect 506703 1005172 506769 1005175
rect 552975 1005172 553041 1005175
rect 421551 1005170 421950 1005172
rect 421551 1005114 421556 1005170
rect 421612 1005142 421950 1005170
rect 501024 1005170 501201 1005172
rect 421612 1005114 421920 1005142
rect 421551 1005112 421920 1005114
rect 501024 1005114 501140 1005170
rect 501196 1005114 501201 1005170
rect 501024 1005112 501201 1005114
rect 506400 1005170 506769 1005172
rect 506400 1005114 506708 1005170
rect 506764 1005114 506769 1005170
rect 506400 1005112 506769 1005114
rect 552864 1005170 553041 1005172
rect 552864 1005114 552980 1005170
rect 553036 1005114 553041 1005170
rect 552864 1005112 553041 1005114
rect 421551 1005109 421617 1005112
rect 501135 1005109 501201 1005112
rect 506703 1005109 506769 1005112
rect 552975 1005109 553041 1005112
rect 156975 1004876 157041 1004879
rect 156975 1004874 157248 1004876
rect 156975 1004818 156980 1004874
rect 157036 1004818 157248 1004874
rect 156975 1004816 157248 1004818
rect 156975 1004813 157041 1004816
rect 306735 1002656 306801 1002659
rect 307311 1002656 307377 1002659
rect 306735 1002654 307104 1002656
rect 306735 1002598 306740 1002654
rect 306796 1002598 307104 1002654
rect 306735 1002596 307104 1002598
rect 307311 1002654 307680 1002656
rect 307311 1002598 307316 1002654
rect 307372 1002598 307680 1002654
rect 307311 1002596 307680 1002598
rect 306735 1002593 306801 1002596
rect 307311 1002593 307377 1002596
rect 103023 1002508 103089 1002511
rect 255279 1002508 255345 1002511
rect 305295 1002508 305361 1002511
rect 307887 1002508 307953 1002511
rect 103023 1002506 103392 1002508
rect 103023 1002450 103028 1002506
rect 103084 1002450 103392 1002506
rect 103023 1002448 103392 1002450
rect 255279 1002506 255552 1002508
rect 255279 1002450 255284 1002506
rect 255340 1002450 255552 1002506
rect 255279 1002448 255552 1002450
rect 305295 1002506 305664 1002508
rect 305295 1002450 305300 1002506
rect 305356 1002450 305664 1002506
rect 305295 1002448 305664 1002450
rect 307887 1002506 308064 1002508
rect 307887 1002450 307892 1002506
rect 307948 1002450 308064 1002506
rect 307887 1002448 308064 1002450
rect 103023 1002445 103089 1002448
rect 255279 1002445 255345 1002448
rect 305295 1002445 305361 1002448
rect 307887 1002445 307953 1002448
rect 101487 1002360 101553 1002363
rect 103599 1002360 103665 1002363
rect 153039 1002360 153105 1002363
rect 253647 1002360 253713 1002363
rect 254223 1002360 254289 1002363
rect 305775 1002360 305841 1002363
rect 306351 1002360 306417 1002363
rect 505647 1002360 505713 1002363
rect 558543 1002360 558609 1002363
rect 101487 1002358 101856 1002360
rect 101487 1002302 101492 1002358
rect 101548 1002302 101856 1002358
rect 101487 1002300 101856 1002302
rect 103599 1002358 103776 1002360
rect 103599 1002302 103604 1002358
rect 103660 1002302 103776 1002358
rect 103599 1002300 103776 1002302
rect 153039 1002358 153312 1002360
rect 153039 1002302 153044 1002358
rect 153100 1002302 153312 1002358
rect 153039 1002300 153312 1002302
rect 253647 1002358 254112 1002360
rect 253647 1002302 253652 1002358
rect 253708 1002302 254112 1002358
rect 253647 1002300 254112 1002302
rect 254223 1002358 254592 1002360
rect 254223 1002302 254228 1002358
rect 254284 1002302 254592 1002358
rect 254223 1002300 254592 1002302
rect 305775 1002358 306144 1002360
rect 305775 1002302 305780 1002358
rect 305836 1002302 306144 1002358
rect 305775 1002300 306144 1002302
rect 306351 1002358 306624 1002360
rect 306351 1002302 306356 1002358
rect 306412 1002302 306624 1002358
rect 306351 1002300 306624 1002302
rect 505440 1002358 505713 1002360
rect 505440 1002302 505652 1002358
rect 505708 1002302 505713 1002358
rect 505440 1002300 505713 1002302
rect 558432 1002358 558609 1002360
rect 558432 1002302 558548 1002358
rect 558604 1002302 558609 1002358
rect 558432 1002300 558609 1002302
rect 101487 1002297 101553 1002300
rect 103599 1002297 103665 1002300
rect 153039 1002297 153105 1002300
rect 253647 1002297 253713 1002300
rect 254223 1002297 254289 1002300
rect 305775 1002297 305841 1002300
rect 306351 1002297 306417 1002300
rect 505647 1002297 505713 1002300
rect 558543 1002297 558609 1002300
rect 430191 1001028 430257 1001031
rect 429984 1001026 430257 1001028
rect 429984 1000970 430196 1001026
rect 430252 1000970 430257 1001026
rect 429984 1000968 430257 1000970
rect 430191 1000965 430257 1000968
rect 208431 1000880 208497 1000883
rect 359727 1000880 359793 1000883
rect 427119 1000880 427185 1000883
rect 429231 1000880 429297 1000883
rect 507183 1000880 507249 1000883
rect 208431 1000878 208608 1000880
rect 208431 1000822 208436 1000878
rect 208492 1000822 208608 1000878
rect 208431 1000820 208608 1000822
rect 359616 1000878 359793 1000880
rect 359616 1000822 359732 1000878
rect 359788 1000822 359793 1000878
rect 359616 1000820 359793 1000822
rect 427008 1000878 427185 1000880
rect 427008 1000822 427124 1000878
rect 427180 1000822 427185 1000878
rect 427008 1000820 427185 1000822
rect 428832 1000878 429297 1000880
rect 428832 1000822 429236 1000878
rect 429292 1000822 429297 1000878
rect 428832 1000820 429297 1000822
rect 506976 1000878 507249 1000880
rect 506976 1000822 507188 1000878
rect 507244 1000822 507249 1000878
rect 506976 1000820 507249 1000822
rect 208431 1000817 208497 1000820
rect 359727 1000817 359793 1000820
rect 427119 1000817 427185 1000820
rect 429231 1000817 429297 1000820
rect 507183 1000817 507249 1000820
rect 517855 1000880 517921 1000883
rect 523887 1000880 523953 1000883
rect 517855 1000878 523953 1000880
rect 517855 1000822 517860 1000878
rect 517916 1000822 523892 1000878
rect 523948 1000822 523953 1000878
rect 517855 1000820 523953 1000822
rect 517855 1000817 517921 1000820
rect 523887 1000817 523953 1000820
rect 506223 1000732 506289 1000735
rect 505920 1000730 506289 1000732
rect 505920 1000674 506228 1000730
rect 506284 1000674 506289 1000730
rect 505920 1000672 506289 1000674
rect 506223 1000669 506289 1000672
rect 518079 1000732 518145 1000735
rect 523983 1000732 524049 1000735
rect 518079 1000730 524049 1000732
rect 518079 1000674 518084 1000730
rect 518140 1000674 523988 1000730
rect 524044 1000674 524049 1000730
rect 518079 1000672 524049 1000674
rect 518079 1000669 518145 1000672
rect 523983 1000669 524049 1000672
rect 520527 999696 520593 999699
rect 523599 999696 523665 999699
rect 520527 999694 523665 999696
rect 520527 999638 520532 999694
rect 520588 999638 523604 999694
rect 523660 999638 523665 999694
rect 520527 999636 523665 999638
rect 520527 999633 520593 999636
rect 523599 999633 523665 999636
rect 256623 999548 256689 999551
rect 259791 999548 259857 999551
rect 311439 999548 311505 999551
rect 504207 999548 504273 999551
rect 256623 999546 256992 999548
rect 256623 999490 256628 999546
rect 256684 999490 256992 999546
rect 256623 999488 256992 999490
rect 259791 999546 260064 999548
rect 259791 999490 259796 999546
rect 259852 999490 260064 999546
rect 259791 999488 260064 999490
rect 311439 999546 311616 999548
rect 311439 999490 311444 999546
rect 311500 999490 311616 999546
rect 311439 999488 311616 999490
rect 504000 999546 504273 999548
rect 504000 999490 504212 999546
rect 504268 999490 504273 999546
rect 504000 999488 504273 999490
rect 256623 999485 256689 999488
rect 259791 999485 259857 999488
rect 311439 999485 311505 999488
rect 504207 999485 504273 999488
rect 521295 999548 521361 999551
rect 523695 999548 523761 999551
rect 521295 999546 523761 999548
rect 521295 999490 521300 999546
rect 521356 999490 523700 999546
rect 523756 999490 523761 999546
rect 521295 999488 523761 999490
rect 521295 999485 521361 999488
rect 523695 999485 523761 999488
rect 154959 999400 155025 999403
rect 206319 999400 206385 999403
rect 257775 999400 257841 999403
rect 309327 999400 309393 999403
rect 518079 999400 518145 999403
rect 524079 999400 524145 999403
rect 154959 999398 155232 999400
rect 154959 999342 154964 999398
rect 155020 999342 155232 999398
rect 154959 999340 155232 999342
rect 206319 999398 206592 999400
rect 206319 999342 206324 999398
rect 206380 999342 206592 999398
rect 206319 999340 206592 999342
rect 257775 999398 257952 999400
rect 257775 999342 257780 999398
rect 257836 999342 257952 999398
rect 257775 999340 257952 999342
rect 309327 999398 309600 999400
rect 309327 999342 309332 999398
rect 309388 999342 309600 999398
rect 309327 999340 309600 999342
rect 518079 999398 524145 999400
rect 518079 999342 518084 999398
rect 518140 999342 524084 999398
rect 524140 999342 524145 999398
rect 518079 999340 524145 999342
rect 154959 999337 155025 999340
rect 206319 999337 206385 999340
rect 257775 999337 257841 999340
rect 309327 999337 309393 999340
rect 518079 999337 518145 999340
rect 524079 999337 524145 999340
rect 105999 997920 106065 997923
rect 105999 997918 106368 997920
rect 105999 997862 106004 997918
rect 106060 997862 106368 997918
rect 105999 997860 106368 997862
rect 105999 997857 106065 997860
rect 555567 997624 555633 997627
rect 555360 997622 555633 997624
rect 555360 997566 555572 997622
rect 555628 997566 555633 997622
rect 555360 997564 555633 997566
rect 555567 997561 555633 997564
rect 557583 997476 557649 997479
rect 557280 997474 557649 997476
rect 557280 997418 557588 997474
rect 557644 997418 557649 997474
rect 557280 997416 557649 997418
rect 557583 997413 557649 997416
rect 256239 996588 256305 996591
rect 309807 996588 309873 996591
rect 256239 996586 256512 996588
rect 256239 996530 256244 996586
rect 256300 996530 256512 996586
rect 256239 996528 256512 996530
rect 309807 996586 310176 996588
rect 309807 996530 309812 996586
rect 309868 996530 310176 996586
rect 309807 996528 310176 996530
rect 256239 996525 256305 996528
rect 309807 996525 309873 996528
rect 108495 996292 108561 996295
rect 108288 996290 108561 996292
rect 108288 996234 108500 996290
rect 108556 996234 108561 996290
rect 108288 996232 108561 996234
rect 108495 996229 108561 996232
rect 153423 996292 153489 996295
rect 154383 996292 154449 996295
rect 159951 996292 160017 996295
rect 204879 996292 204945 996295
rect 153423 996290 153696 996292
rect 153423 996234 153428 996290
rect 153484 996234 153696 996290
rect 153423 996232 153696 996234
rect 154383 996290 154848 996292
rect 154383 996234 154388 996290
rect 154444 996234 154848 996290
rect 154383 996232 154848 996234
rect 159951 996290 160224 996292
rect 159951 996234 159956 996290
rect 160012 996234 160224 996290
rect 159951 996232 160224 996234
rect 204879 996290 205152 996292
rect 204879 996234 204884 996290
rect 204940 996234 205152 996290
rect 204879 996232 205152 996234
rect 264480 996232 264894 996292
rect 153423 996229 153489 996232
rect 154383 996229 154449 996232
rect 159951 996229 160017 996232
rect 204879 996229 204945 996232
rect 100527 996144 100593 996147
rect 103983 996144 104049 996147
rect 104463 996144 104529 996147
rect 108591 996144 108657 996147
rect 109551 996144 109617 996147
rect 151983 996144 152049 996147
rect 152367 996144 152433 996147
rect 153999 996144 154065 996147
rect 156495 996144 156561 996147
rect 157359 996144 157425 996147
rect 158895 996144 158961 996147
rect 100527 996142 100800 996144
rect 97794 995996 97854 996114
rect 98850 995996 98910 996114
rect 97794 995936 98910 995996
rect 85935 995848 86001 995851
rect 92559 995848 92625 995851
rect 85935 995846 92625 995848
rect 85935 995790 85940 995846
rect 85996 995790 92564 995846
rect 92620 995790 92625 995846
rect 85935 995788 92625 995790
rect 85935 995785 86001 995788
rect 92559 995785 92625 995788
rect 94959 995848 95025 995851
rect 99810 995848 99870 996114
rect 94959 995846 99870 995848
rect 94959 995790 94964 995846
rect 95020 995790 99870 995846
rect 94959 995788 99870 995790
rect 94959 995785 95025 995788
rect 81615 995700 81681 995703
rect 92655 995700 92721 995703
rect 81615 995698 92721 995700
rect 81615 995642 81620 995698
rect 81676 995642 92660 995698
rect 92716 995642 92721 995698
rect 81615 995640 92721 995642
rect 81615 995637 81681 995640
rect 92655 995637 92721 995640
rect 94959 995700 95025 995703
rect 100386 995700 100446 996114
rect 100527 996086 100532 996142
rect 100588 996086 100800 996142
rect 100527 996084 100800 996086
rect 103983 996142 104352 996144
rect 103983 996086 103988 996142
rect 104044 996086 104352 996142
rect 103983 996084 104352 996086
rect 104463 996142 104928 996144
rect 104463 996086 104468 996142
rect 104524 996086 104928 996142
rect 108591 996142 108768 996144
rect 104463 996084 104928 996086
rect 100527 996081 100593 996084
rect 103983 996081 104049 996084
rect 104463 996081 104529 996084
rect 103599 995996 103665 995999
rect 105282 995996 105342 996114
rect 103599 995994 105342 995996
rect 103599 995938 103604 995994
rect 103660 995938 105342 995994
rect 103599 995936 105342 995938
rect 103599 995933 103665 995936
rect 107298 995848 107358 996114
rect 108591 996086 108596 996142
rect 108652 996086 108768 996142
rect 109551 996142 109728 996144
rect 108591 996084 108768 996086
rect 108591 996081 108657 996084
rect 109314 995996 109374 996114
rect 109551 996086 109556 996142
rect 109612 996086 109728 996142
rect 109551 996084 109728 996086
rect 109551 996081 109617 996084
rect 115215 995996 115281 995999
rect 146703 995996 146769 995999
rect 109314 995994 115281 995996
rect 109314 995938 115220 995994
rect 115276 995938 115281 995994
rect 109314 995936 115281 995938
rect 115215 995933 115281 995936
rect 137730 995994 146769 995996
rect 137730 995938 146708 995994
rect 146764 995938 146769 995994
rect 137730 995936 146769 995938
rect 149154 995996 149214 996114
rect 150018 996084 150240 996144
rect 150978 996084 151200 996144
rect 151983 996142 152160 996144
rect 150018 995996 150078 996084
rect 149154 995936 150078 995996
rect 112335 995848 112401 995851
rect 107298 995846 112401 995848
rect 107298 995790 112340 995846
rect 112396 995790 112401 995846
rect 107298 995788 112401 995790
rect 112335 995785 112401 995788
rect 133647 995848 133713 995851
rect 137730 995848 137790 995936
rect 146703 995933 146769 995936
rect 133647 995846 137790 995848
rect 133647 995790 133652 995846
rect 133708 995790 137790 995846
rect 133647 995788 137790 995790
rect 137967 995848 138033 995851
rect 150978 995848 151038 996084
rect 137967 995846 151038 995848
rect 137967 995790 137972 995846
rect 138028 995790 151038 995846
rect 137967 995788 151038 995790
rect 133647 995785 133713 995788
rect 137967 995785 138033 995788
rect 94959 995698 100446 995700
rect 94959 995642 94964 995698
rect 95020 995642 100446 995698
rect 94959 995640 100446 995642
rect 137391 995700 137457 995703
rect 146799 995700 146865 995703
rect 137391 995698 146865 995700
rect 137391 995642 137396 995698
rect 137452 995642 146804 995698
rect 146860 995642 146865 995698
rect 137391 995640 146865 995642
rect 94959 995637 95025 995640
rect 137391 995637 137457 995640
rect 146799 995637 146865 995640
rect 81039 995552 81105 995555
rect 92847 995552 92913 995555
rect 81039 995550 92913 995552
rect 81039 995494 81044 995550
rect 81100 995494 92852 995550
rect 92908 995494 92913 995550
rect 81039 995492 92913 995494
rect 81039 995489 81105 995492
rect 92847 995489 92913 995492
rect 136719 995552 136785 995555
rect 151746 995552 151806 996114
rect 151983 996086 151988 996142
rect 152044 996086 152160 996142
rect 151983 996084 152160 996086
rect 152367 996142 152736 996144
rect 152367 996086 152372 996142
rect 152428 996086 152736 996142
rect 152367 996084 152736 996086
rect 153999 996142 154272 996144
rect 153999 996086 154004 996142
rect 154060 996086 154272 996142
rect 156495 996142 156672 996144
rect 153999 996084 154272 996086
rect 151983 996081 152049 996084
rect 152367 996081 152433 996084
rect 153999 996081 154065 996084
rect 136719 995550 151806 995552
rect 136719 995494 136724 995550
rect 136780 995494 151806 995550
rect 136719 995492 151806 995494
rect 136719 995489 136785 995492
rect 132399 995404 132465 995407
rect 146703 995404 146769 995407
rect 132399 995402 146769 995404
rect 132399 995346 132404 995402
rect 132460 995346 146708 995402
rect 146764 995346 146769 995402
rect 132399 995344 146769 995346
rect 132399 995341 132465 995344
rect 146703 995341 146769 995344
rect 132783 994220 132849 994223
rect 149679 994220 149745 994223
rect 132783 994218 149745 994220
rect 132783 994162 132788 994218
rect 132844 994162 149684 994218
rect 149740 994162 149745 994218
rect 132783 994160 149745 994162
rect 132783 994157 132849 994160
rect 149679 994157 149745 994160
rect 84495 994072 84561 994075
rect 103983 994072 104049 994075
rect 84495 994070 104049 994072
rect 84495 994014 84500 994070
rect 84556 994014 103988 994070
rect 104044 994014 104049 994070
rect 84495 994012 104049 994014
rect 84495 994009 84561 994012
rect 103983 994009 104049 994012
rect 88719 993924 88785 993927
rect 110319 993924 110385 993927
rect 88719 993922 110385 993924
rect 88719 993866 88724 993922
rect 88780 993866 110324 993922
rect 110380 993866 110385 993922
rect 88719 993864 110385 993866
rect 88719 993861 88785 993864
rect 110319 993861 110385 993864
rect 136143 993924 136209 993927
rect 155682 993924 155742 996114
rect 156258 995999 156318 996114
rect 156495 996086 156500 996142
rect 156556 996086 156672 996142
rect 156495 996084 156672 996086
rect 157359 996142 157728 996144
rect 157359 996086 157364 996142
rect 157420 996086 157728 996142
rect 157359 996084 157728 996086
rect 158688 996142 158961 996144
rect 158688 996086 158900 996142
rect 158956 996086 158961 996142
rect 202287 996144 202353 996147
rect 202863 996144 202929 996147
rect 203919 996144 203985 996147
rect 205263 996144 205329 996147
rect 205935 996144 206001 996147
rect 207855 996144 207921 996147
rect 210831 996144 210897 996147
rect 211407 996144 211473 996147
rect 212751 996144 212817 996147
rect 219087 996144 219153 996147
rect 252303 996144 252369 996147
rect 202287 996142 202656 996144
rect 158688 996084 158961 996086
rect 156495 996081 156561 996084
rect 157359 996081 157425 996084
rect 158895 996081 158961 996084
rect 156207 995994 156318 995999
rect 156207 995938 156212 995994
rect 156268 995938 156318 995994
rect 156207 995936 156318 995938
rect 159618 995999 159678 996114
rect 159618 995994 159729 995999
rect 159618 995938 159668 995994
rect 159724 995938 159729 995994
rect 159618 995936 159729 995938
rect 156207 995933 156273 995936
rect 159663 995933 159729 995936
rect 198639 995996 198705 995999
rect 201090 995996 201150 996114
rect 202050 995996 202110 996114
rect 202287 996086 202292 996142
rect 202348 996086 202656 996142
rect 202287 996084 202656 996086
rect 202863 996142 203232 996144
rect 202863 996086 202868 996142
rect 202924 996086 203232 996142
rect 203919 996142 204192 996144
rect 202863 996084 203232 996086
rect 202287 996081 202353 996084
rect 202863 996081 202929 996084
rect 198639 995994 202110 995996
rect 198639 995938 198644 995994
rect 198700 995938 202110 995994
rect 198639 995936 202110 995938
rect 198639 995933 198705 995936
rect 185103 995848 185169 995851
rect 203586 995848 203646 996114
rect 203919 996086 203924 996142
rect 203980 996086 204192 996142
rect 205263 996142 205632 996144
rect 203919 996084 204192 996086
rect 203919 996081 203985 996084
rect 185103 995846 203646 995848
rect 185103 995790 185108 995846
rect 185164 995790 203646 995846
rect 185103 995788 203646 995790
rect 185103 995785 185169 995788
rect 184335 995700 184401 995703
rect 190575 995700 190641 995703
rect 204642 995700 204702 996114
rect 205263 996086 205268 996142
rect 205324 996086 205632 996142
rect 205263 996084 205632 996086
rect 205935 996142 206208 996144
rect 205935 996086 205940 996142
rect 205996 996086 206208 996142
rect 207855 996142 208032 996144
rect 205935 996084 206208 996086
rect 205263 996081 205329 996084
rect 205935 996081 206001 996084
rect 184335 995698 187902 995700
rect 184335 995642 184340 995698
rect 184396 995642 187902 995698
rect 184335 995640 187902 995642
rect 184335 995637 184401 995640
rect 183279 995552 183345 995555
rect 183279 995550 187230 995552
rect 183279 995494 183284 995550
rect 183340 995494 187230 995550
rect 183279 995492 187230 995494
rect 183279 995489 183345 995492
rect 187170 995108 187230 995492
rect 187842 995404 187902 995640
rect 190575 995698 204702 995700
rect 190575 995642 190580 995698
rect 190636 995642 204702 995698
rect 190575 995640 204702 995642
rect 190575 995637 190641 995640
rect 188079 995552 188145 995555
rect 202863 995552 202929 995555
rect 188079 995550 202929 995552
rect 188079 995494 188084 995550
rect 188140 995494 202868 995550
rect 202924 995494 202929 995550
rect 188079 995492 202929 995494
rect 188079 995489 188145 995492
rect 202863 995489 202929 995492
rect 201519 995404 201585 995407
rect 187842 995402 201585 995404
rect 187842 995346 201524 995402
rect 201580 995346 201585 995402
rect 187842 995344 201585 995346
rect 201519 995341 201585 995344
rect 187311 995256 187377 995259
rect 207138 995256 207198 996114
rect 207855 996086 207860 996142
rect 207916 996086 208032 996142
rect 210831 996142 211104 996144
rect 207855 996084 208032 996086
rect 207855 996081 207921 996084
rect 209154 995555 209214 996114
rect 210114 995999 210174 996114
rect 210831 996086 210836 996142
rect 210892 996086 211104 996142
rect 210831 996084 211104 996086
rect 211407 996142 211680 996144
rect 211407 996086 211412 996142
rect 211468 996086 211680 996142
rect 212640 996142 212817 996144
rect 211407 996084 211680 996086
rect 210831 996081 210897 996084
rect 211407 996081 211473 996084
rect 210114 995994 210225 995999
rect 210114 995938 210164 995994
rect 210220 995938 210225 995994
rect 210114 995936 210225 995938
rect 212130 995996 212190 996114
rect 212640 996086 212756 996142
rect 212812 996086 212817 996142
rect 212640 996084 212817 996086
rect 213696 996142 219153 996144
rect 213696 996086 219092 996142
rect 219148 996086 219153 996142
rect 213696 996084 219153 996086
rect 252000 996142 252369 996144
rect 252000 996086 252308 996142
rect 252364 996086 252369 996142
rect 252000 996084 252369 996086
rect 212751 996081 212817 996084
rect 219087 996081 219153 996084
rect 252303 996081 252369 996084
rect 252687 996144 252753 996147
rect 254799 996144 254865 996147
rect 258735 996144 258801 996147
rect 260367 996144 260433 996147
rect 262767 996144 262833 996147
rect 263727 996144 263793 996147
rect 252687 996142 253152 996144
rect 252687 996086 252692 996142
rect 252748 996086 253152 996142
rect 252687 996084 253152 996086
rect 254799 996142 254976 996144
rect 254799 996086 254804 996142
rect 254860 996086 254976 996142
rect 254799 996084 254976 996086
rect 255810 996084 256032 996144
rect 258735 996142 259104 996144
rect 252687 996081 252753 996084
rect 254799 996081 254865 996084
rect 216015 995996 216081 995999
rect 246927 995996 246993 995999
rect 255810 995996 255870 996084
rect 212130 995994 216081 995996
rect 212130 995938 216020 995994
rect 216076 995938 216081 995994
rect 212130 995936 216081 995938
rect 210159 995933 210225 995936
rect 216015 995933 216081 995936
rect 240258 995994 246993 995996
rect 240258 995938 246932 995994
rect 246988 995938 246993 995994
rect 240258 995936 246993 995938
rect 240258 995851 240318 995936
rect 246927 995933 246993 995936
rect 247650 995936 255870 995996
rect 240207 995846 240318 995851
rect 240207 995790 240212 995846
rect 240268 995790 240318 995846
rect 240207 995788 240318 995790
rect 241839 995848 241905 995851
rect 247650 995848 247710 995936
rect 241839 995846 247710 995848
rect 241839 995790 241844 995846
rect 241900 995790 247710 995846
rect 241839 995788 247710 995790
rect 240207 995785 240273 995788
rect 241839 995785 241905 995788
rect 232143 995700 232209 995703
rect 257538 995700 257598 996114
rect 232143 995698 257598 995700
rect 232143 995642 232148 995698
rect 232204 995642 257598 995698
rect 232143 995640 257598 995642
rect 232143 995637 232209 995640
rect 209103 995550 209214 995555
rect 209103 995494 209108 995550
rect 209164 995494 209214 995550
rect 209103 995492 209214 995494
rect 235215 995552 235281 995555
rect 247023 995552 247089 995555
rect 235215 995550 247089 995552
rect 235215 995494 235220 995550
rect 235276 995494 247028 995550
rect 247084 995494 247089 995550
rect 235215 995492 247089 995494
rect 209103 995489 209169 995492
rect 235215 995489 235281 995492
rect 247023 995489 247089 995492
rect 187311 995254 207198 995256
rect 187311 995198 187316 995254
rect 187372 995198 207198 995254
rect 187311 995196 207198 995198
rect 187311 995193 187377 995196
rect 197199 995108 197265 995111
rect 187170 995106 197265 995108
rect 187170 995050 197204 995106
rect 197260 995050 197265 995106
rect 187170 995048 197265 995050
rect 197199 995045 197265 995048
rect 238671 994368 238737 994371
rect 258498 994368 258558 996114
rect 258735 996086 258740 996142
rect 258796 996086 259104 996142
rect 260367 996142 260640 996144
rect 258735 996084 259104 996086
rect 258735 996081 258801 996084
rect 238671 994366 258558 994368
rect 238671 994310 238676 994366
rect 238732 994310 258558 994366
rect 238671 994308 258558 994310
rect 238671 994305 238737 994308
rect 234351 994220 234417 994223
rect 258735 994220 258801 994223
rect 234351 994218 258801 994220
rect 234351 994162 234356 994218
rect 234412 994162 258740 994218
rect 258796 994162 258801 994218
rect 234351 994160 258801 994162
rect 234351 994157 234417 994160
rect 258735 994157 258801 994160
rect 231471 994072 231537 994075
rect 259458 994072 259518 996114
rect 260367 996086 260372 996142
rect 260428 996086 260640 996142
rect 262767 996142 263040 996144
rect 260367 996084 260640 996086
rect 260367 996081 260433 996084
rect 261474 995999 261534 996114
rect 262434 995999 262494 996114
rect 262767 996086 262772 996142
rect 262828 996086 263040 996142
rect 262767 996084 263040 996086
rect 263520 996142 263793 996144
rect 263520 996086 263732 996142
rect 263788 996086 263793 996142
rect 263520 996084 263793 996086
rect 262767 996081 262833 996084
rect 263727 996081 263793 996084
rect 261474 995994 261585 995999
rect 261474 995938 261524 995994
rect 261580 995938 261585 995994
rect 261474 995936 261585 995938
rect 262434 995994 262545 995999
rect 262434 995938 262484 995994
rect 262540 995938 262545 995994
rect 262434 995936 262545 995938
rect 261519 995933 261585 995936
rect 262479 995933 262545 995936
rect 263970 995848 264030 996114
rect 264834 995996 264894 996232
rect 270735 996144 270801 996147
rect 304431 996144 304497 996147
rect 265056 996142 270801 996144
rect 265056 996086 270740 996142
rect 270796 996086 270801 996142
rect 304128 996142 304497 996144
rect 265056 996084 270801 996086
rect 270735 996081 270801 996084
rect 267855 995996 267921 995999
rect 298479 995996 298545 995999
rect 264834 995994 267921 995996
rect 264834 995938 267860 995994
rect 267916 995938 267921 995994
rect 264834 995936 267921 995938
rect 267855 995933 267921 995936
rect 291522 995994 298545 995996
rect 291522 995938 298484 995994
rect 298540 995938 298545 995994
rect 291522 995936 298545 995938
rect 303618 995996 303678 996114
rect 304128 996086 304436 996142
rect 304492 996086 304497 996142
rect 304911 996144 304977 996147
rect 305295 996144 305361 996147
rect 304911 996142 305361 996144
rect 304128 996084 304497 996086
rect 304431 996081 304497 996084
rect 304674 995996 304734 996114
rect 304911 996086 304916 996142
rect 304972 996086 305300 996142
rect 305356 996086 305361 996142
rect 310863 996144 310929 996147
rect 314223 996144 314289 996147
rect 319599 996144 319665 996147
rect 363855 996144 363921 996147
rect 366255 996144 366321 996147
rect 366735 996144 366801 996147
rect 371535 996144 371601 996147
rect 310863 996142 311136 996144
rect 304911 996084 305361 996086
rect 304911 996081 304977 996084
rect 305295 996081 305361 996084
rect 303618 995936 304734 995996
rect 304815 995996 304881 995999
rect 309186 995996 309246 996114
rect 304815 995994 309246 995996
rect 304815 995938 304820 995994
rect 304876 995938 309246 995994
rect 304815 995936 309246 995938
rect 267951 995848 268017 995851
rect 263970 995846 268017 995848
rect 263970 995790 267956 995846
rect 268012 995790 268017 995846
rect 263970 995788 268017 995790
rect 267951 995785 268017 995788
rect 286767 995848 286833 995851
rect 291522 995848 291582 995936
rect 298479 995933 298545 995936
rect 304815 995933 304881 995936
rect 286767 995846 291582 995848
rect 286767 995790 286772 995846
rect 286828 995790 291582 995846
rect 286767 995788 291582 995790
rect 291759 995848 291825 995851
rect 299535 995848 299601 995851
rect 291759 995846 299601 995848
rect 291759 995790 291764 995846
rect 291820 995790 299540 995846
rect 299596 995790 299601 995846
rect 291759 995788 299601 995790
rect 286767 995785 286833 995788
rect 291759 995785 291825 995788
rect 299535 995785 299601 995788
rect 303375 995848 303441 995851
rect 310626 995848 310686 996114
rect 310863 996086 310868 996142
rect 310924 996086 311136 996142
rect 314112 996142 314289 996144
rect 310863 996084 311136 996086
rect 310863 996081 310929 996084
rect 303375 995846 310686 995848
rect 303375 995790 303380 995846
rect 303436 995790 310686 995846
rect 303375 995788 310686 995790
rect 303375 995785 303441 995788
rect 293583 995700 293649 995703
rect 299727 995700 299793 995703
rect 293583 995698 299793 995700
rect 293583 995642 293588 995698
rect 293644 995642 299732 995698
rect 299788 995642 299793 995698
rect 293583 995640 299793 995642
rect 293583 995637 293649 995640
rect 299727 995637 299793 995640
rect 284367 995552 284433 995555
rect 312162 995552 312222 996114
rect 313122 995999 313182 996114
rect 314112 996086 314228 996142
rect 314284 996086 314289 996142
rect 316704 996142 319665 996144
rect 314112 996084 314289 996086
rect 314223 996081 314289 996084
rect 313071 995994 313182 995999
rect 313071 995938 313076 995994
rect 313132 995938 313182 995994
rect 313071 995936 313182 995938
rect 313839 995996 313905 995999
rect 314562 995996 314622 996114
rect 313839 995994 314622 995996
rect 313839 995938 313844 995994
rect 313900 995938 314622 995994
rect 313839 995936 314622 995938
rect 315522 995996 315582 996114
rect 316704 996086 319604 996142
rect 319660 996086 319665 996142
rect 316704 996084 319665 996086
rect 353952 996084 354366 996144
rect 363855 996142 364128 996144
rect 319599 996081 319665 996084
rect 319695 995996 319761 995999
rect 315522 995994 319761 995996
rect 315522 995938 319700 995994
rect 319756 995938 319761 995994
rect 315522 995936 319761 995938
rect 354306 995996 354366 996084
rect 355074 995996 355134 996114
rect 354306 995936 355134 995996
rect 313071 995933 313137 995936
rect 313839 995933 313905 995936
rect 319695 995933 319761 995936
rect 359970 995703 360030 996114
rect 362946 995703 363006 996114
rect 363522 995703 363582 996114
rect 363855 996086 363860 996142
rect 363916 996086 364128 996142
rect 363855 996084 364128 996086
rect 363855 996081 363921 996084
rect 364482 995703 364542 996114
rect 365088 996084 365310 996144
rect 365952 996142 366321 996144
rect 365952 996086 366260 996142
rect 366316 996086 366321 996142
rect 365952 996084 366321 996086
rect 366528 996142 366801 996144
rect 366528 996086 366740 996142
rect 366796 996086 366801 996142
rect 366528 996084 366801 996086
rect 367008 996142 371601 996144
rect 367008 996086 371540 996142
rect 371596 996086 371601 996142
rect 430191 996144 430257 996147
rect 431247 996144 431313 996147
rect 432783 996144 432849 996147
rect 433551 996144 433617 996147
rect 434127 996144 434193 996147
rect 437967 996144 438033 996147
rect 499119 996144 499185 996147
rect 509775 996144 509841 996147
rect 510735 996144 510801 996147
rect 511119 996144 511185 996147
rect 515535 996144 515601 996147
rect 555951 996144 556017 996147
rect 430191 996142 430368 996144
rect 367008 996084 371601 996086
rect 365250 995996 365310 996084
rect 366255 996081 366321 996084
rect 366735 996081 366801 996084
rect 371535 996081 371601 996084
rect 374415 995996 374481 995999
rect 365250 995994 374481 995996
rect 365250 995938 374420 995994
rect 374476 995938 374481 995994
rect 365250 995936 374481 995938
rect 421410 995996 421470 996114
rect 422466 995996 422526 996114
rect 421410 995936 422526 995996
rect 374415 995933 374481 995936
rect 382767 995848 382833 995851
rect 388815 995848 388881 995851
rect 382767 995846 388881 995848
rect 382767 995790 382772 995846
rect 382828 995790 388820 995846
rect 388876 995790 388881 995846
rect 382767 995788 388881 995790
rect 382767 995785 382833 995788
rect 388815 995785 388881 995788
rect 427362 995703 427422 996114
rect 430191 996086 430196 996142
rect 430252 996086 430368 996142
rect 431247 996142 431520 996144
rect 430191 996084 430368 996086
rect 430191 996081 430257 996084
rect 359970 995698 360081 995703
rect 359970 995642 360020 995698
rect 360076 995642 360081 995698
rect 359970 995640 360081 995642
rect 360015 995637 360081 995640
rect 362895 995698 363006 995703
rect 362895 995642 362900 995698
rect 362956 995642 363006 995698
rect 362895 995640 363006 995642
rect 363471 995698 363582 995703
rect 363471 995642 363476 995698
rect 363532 995642 363582 995698
rect 363471 995640 363582 995642
rect 364431 995698 364542 995703
rect 364431 995642 364436 995698
rect 364492 995642 364542 995698
rect 364431 995640 364542 995642
rect 380175 995700 380241 995703
rect 394863 995700 394929 995703
rect 380175 995698 394929 995700
rect 380175 995642 380180 995698
rect 380236 995642 394868 995698
rect 394924 995642 394929 995698
rect 380175 995640 394929 995642
rect 427362 995698 427473 995703
rect 427362 995642 427412 995698
rect 427468 995642 427473 995698
rect 427362 995640 427473 995642
rect 362895 995637 362961 995640
rect 363471 995637 363537 995640
rect 364431 995637 364497 995640
rect 380175 995637 380241 995640
rect 394863 995637 394929 995640
rect 427407 995637 427473 995640
rect 430914 995555 430974 996114
rect 431247 996086 431252 996142
rect 431308 996086 431520 996142
rect 431247 996084 431520 996086
rect 431247 996081 431313 996084
rect 431874 995555 431934 996114
rect 432480 996084 432702 996144
rect 432642 995996 432702 996084
rect 432783 996142 432960 996144
rect 432783 996086 432788 996142
rect 432844 996086 432960 996142
rect 432783 996084 432960 996086
rect 433440 996142 433617 996144
rect 433440 996086 433556 996142
rect 433612 996086 433617 996142
rect 433440 996084 433617 996086
rect 433920 996142 434193 996144
rect 433920 996086 434132 996142
rect 434188 996086 434193 996142
rect 433920 996084 434193 996086
rect 434496 996142 438033 996144
rect 434496 996086 437972 996142
rect 438028 996086 438033 996142
rect 498912 996142 499185 996144
rect 434496 996084 438033 996086
rect 432783 996081 432849 996084
rect 433551 996081 433617 996084
rect 434127 996081 434193 996084
rect 437967 996081 438033 996084
rect 440655 995996 440721 995999
rect 432642 995994 440721 995996
rect 432642 995938 440660 995994
rect 440716 995938 440721 995994
rect 432642 995936 440721 995938
rect 440655 995933 440721 995936
rect 471855 995996 471921 995999
rect 498402 995996 498462 996114
rect 498912 996086 499124 996142
rect 499180 996086 499185 996142
rect 498912 996084 499185 996086
rect 499119 996081 499185 996084
rect 499458 995996 499518 996114
rect 471855 995994 480318 995996
rect 471855 995938 471860 995994
rect 471916 995938 480318 995994
rect 471855 995936 480318 995938
rect 498402 995936 499518 995996
rect 471855 995933 471921 995936
rect 472143 995848 472209 995851
rect 478383 995848 478449 995851
rect 472143 995846 478449 995848
rect 472143 995790 472148 995846
rect 472204 995790 478388 995846
rect 478444 995790 478449 995846
rect 472143 995788 478449 995790
rect 480258 995848 480318 995936
rect 482031 995848 482097 995851
rect 480258 995846 482097 995848
rect 480258 995790 482036 995846
rect 482092 995790 482097 995846
rect 480258 995788 482097 995790
rect 472143 995785 472209 995788
rect 478383 995785 478449 995788
rect 482031 995785 482097 995788
rect 495279 995848 495345 995851
rect 499119 995848 499185 995851
rect 499842 995848 499902 996114
rect 495279 995846 499902 995848
rect 495279 995790 495284 995846
rect 495340 995790 499124 995846
rect 499180 995790 499902 995846
rect 495279 995788 499902 995790
rect 495279 995785 495345 995788
rect 499119 995785 499185 995788
rect 504354 995555 504414 996114
rect 507330 995555 507390 996114
rect 507906 995999 507966 996114
rect 508482 995999 508542 996114
rect 507855 995994 507966 995999
rect 507855 995938 507860 995994
rect 507916 995938 507966 995994
rect 507855 995936 507966 995938
rect 508431 995994 508542 995999
rect 508431 995938 508436 995994
rect 508492 995938 508542 995994
rect 508431 995936 508542 995938
rect 507855 995933 507921 995936
rect 508431 995933 508497 995936
rect 508866 995555 508926 996114
rect 509472 996084 509694 996144
rect 509634 995996 509694 996084
rect 509775 996142 509952 996144
rect 509775 996086 509780 996142
rect 509836 996086 509952 996142
rect 509775 996084 509952 996086
rect 510432 996142 510801 996144
rect 510432 996086 510740 996142
rect 510796 996086 510801 996142
rect 510432 996084 510801 996086
rect 510912 996142 511185 996144
rect 510912 996086 511124 996142
rect 511180 996086 511185 996142
rect 510912 996084 511185 996086
rect 511488 996142 515601 996144
rect 511488 996086 515540 996142
rect 515596 996086 515601 996142
rect 511488 996084 515601 996086
rect 509775 996081 509841 996084
rect 510735 996081 510801 996084
rect 511119 996081 511185 996084
rect 515535 996081 515601 996084
rect 512655 995996 512721 995999
rect 509634 995994 512721 995996
rect 509634 995938 512660 995994
rect 512716 995938 512721 995994
rect 509634 995936 512721 995938
rect 512655 995933 512721 995936
rect 521487 995996 521553 995999
rect 549762 995996 549822 996114
rect 550530 996084 550944 996144
rect 555744 996142 556017 996144
rect 555744 996086 555956 996142
rect 556012 996086 556017 996142
rect 559119 996144 559185 996147
rect 561135 996144 561201 996147
rect 561903 996144 561969 996147
rect 569871 996144 569937 996147
rect 559119 996142 559392 996144
rect 555744 996084 556017 996086
rect 550530 995996 550590 996084
rect 555951 996081 556017 996084
rect 521487 995994 529470 995996
rect 521487 995938 521492 995994
rect 521548 995938 529470 995994
rect 521487 995936 529470 995938
rect 549762 995936 550590 995996
rect 521487 995933 521553 995936
rect 521391 995848 521457 995851
rect 527919 995848 527985 995851
rect 521391 995846 527985 995848
rect 521391 995790 521396 995846
rect 521452 995790 527924 995846
rect 527980 995790 527985 995846
rect 521391 995788 527985 995790
rect 529410 995848 529470 995936
rect 537231 995848 537297 995851
rect 529410 995846 537297 995848
rect 529410 995790 537236 995846
rect 537292 995790 537297 995846
rect 529410 995788 537297 995790
rect 521391 995785 521457 995788
rect 527919 995785 527985 995788
rect 537231 995785 537297 995788
rect 521583 995700 521649 995703
rect 532239 995700 532305 995703
rect 521583 995698 532305 995700
rect 521583 995642 521588 995698
rect 521644 995642 532244 995698
rect 532300 995642 532305 995698
rect 521583 995640 532305 995642
rect 521583 995637 521649 995640
rect 532239 995637 532305 995640
rect 284367 995550 312222 995552
rect 284367 995494 284372 995550
rect 284428 995494 312222 995550
rect 284367 995492 312222 995494
rect 430863 995550 430974 995555
rect 430863 995494 430868 995550
rect 430924 995494 430974 995550
rect 430863 995492 430974 995494
rect 431823 995550 431934 995555
rect 431823 995494 431828 995550
rect 431884 995494 431934 995550
rect 431823 995492 431934 995494
rect 471951 995552 472017 995555
rect 481359 995552 481425 995555
rect 471951 995550 481425 995552
rect 471951 995494 471956 995550
rect 472012 995494 481364 995550
rect 481420 995494 481425 995550
rect 471951 995492 481425 995494
rect 284367 995489 284433 995492
rect 430863 995489 430929 995492
rect 431823 995489 431889 995492
rect 471951 995489 472017 995492
rect 481359 995489 481425 995492
rect 485583 995552 485649 995555
rect 491823 995552 491889 995555
rect 485583 995550 491889 995552
rect 485583 995494 485588 995550
rect 485644 995494 491828 995550
rect 491884 995494 491889 995550
rect 485583 995492 491889 995494
rect 504354 995550 504465 995555
rect 504354 995494 504404 995550
rect 504460 995494 504465 995550
rect 504354 995492 504465 995494
rect 485583 995489 485649 995492
rect 491823 995489 491889 995492
rect 504399 995489 504465 995492
rect 507279 995550 507390 995555
rect 507279 995494 507284 995550
rect 507340 995494 507390 995550
rect 507279 995492 507390 995494
rect 508815 995550 508926 995555
rect 508815 995494 508820 995550
rect 508876 995494 508926 995550
rect 508815 995492 508926 995494
rect 518511 995552 518577 995555
rect 533391 995552 533457 995555
rect 518511 995550 533457 995552
rect 518511 995494 518516 995550
rect 518572 995494 533396 995550
rect 533452 995494 533457 995550
rect 518511 995492 533457 995494
rect 507279 995489 507345 995492
rect 508815 995489 508881 995492
rect 518511 995489 518577 995492
rect 533391 995489 533457 995492
rect 287439 995404 287505 995407
rect 300111 995404 300177 995407
rect 287439 995402 300177 995404
rect 287439 995346 287444 995402
rect 287500 995346 300116 995402
rect 300172 995346 300177 995402
rect 287439 995344 300177 995346
rect 287439 995341 287505 995344
rect 300111 995341 300177 995344
rect 518415 995404 518481 995407
rect 535311 995404 535377 995407
rect 518415 995402 535377 995404
rect 518415 995346 518420 995402
rect 518476 995346 535316 995402
rect 535372 995346 535377 995402
rect 518415 995344 535377 995346
rect 518415 995341 518481 995344
rect 535311 995341 535377 995344
rect 556290 995256 556350 996114
rect 556866 995404 556926 996114
rect 558786 995552 558846 996114
rect 559119 996086 559124 996142
rect 559180 996086 559392 996142
rect 561135 996142 561312 996144
rect 559119 996084 559392 996086
rect 559119 996081 559185 996084
rect 559842 995700 559902 996114
rect 560226 995999 560286 996114
rect 560175 995994 560286 995999
rect 560175 995938 560180 995994
rect 560236 995938 560286 995994
rect 560175 995936 560286 995938
rect 560175 995933 560241 995936
rect 560802 995848 560862 996114
rect 561135 996086 561140 996142
rect 561196 996086 561312 996142
rect 561135 996084 561312 996086
rect 561792 996142 561969 996144
rect 561792 996086 561908 996142
rect 561964 996086 561969 996142
rect 561792 996084 561969 996086
rect 562272 996084 562686 996144
rect 562848 996142 569937 996144
rect 562848 996086 569876 996142
rect 569932 996086 569937 996142
rect 562848 996084 569937 996086
rect 561135 996081 561201 996084
rect 561903 996081 561969 996084
rect 562626 995996 562686 996084
rect 569871 996081 569937 996084
rect 569775 995996 569841 995999
rect 562626 995994 569841 995996
rect 562626 995938 569780 995994
rect 569836 995938 569841 995994
rect 562626 995936 569841 995938
rect 569775 995933 569841 995936
rect 567183 995848 567249 995851
rect 560802 995846 567249 995848
rect 560802 995790 567188 995846
rect 567244 995790 567249 995846
rect 560802 995788 567249 995790
rect 567183 995785 567249 995788
rect 565839 995700 565905 995703
rect 559842 995698 565905 995700
rect 559842 995642 565844 995698
rect 565900 995642 565905 995698
rect 559842 995640 565905 995642
rect 565839 995637 565905 995640
rect 566031 995552 566097 995555
rect 558786 995550 566097 995552
rect 558786 995494 566036 995550
rect 566092 995494 566097 995550
rect 558786 995492 566097 995494
rect 566031 995489 566097 995492
rect 567375 995404 567441 995407
rect 556866 995402 567441 995404
rect 556866 995346 567380 995402
rect 567436 995346 567441 995402
rect 556866 995344 567441 995346
rect 567375 995341 567441 995344
rect 561615 995256 561681 995259
rect 556290 995254 561681 995256
rect 556290 995198 561620 995254
rect 561676 995198 561681 995254
rect 556290 995196 561681 995198
rect 561615 995193 561681 995196
rect 285999 994516 286065 994519
rect 303375 994516 303441 994519
rect 285999 994514 303441 994516
rect 285999 994458 286004 994514
rect 286060 994458 303380 994514
rect 303436 994458 303441 994514
rect 285999 994456 303441 994458
rect 285999 994453 286065 994456
rect 303375 994453 303441 994456
rect 573135 994516 573201 994519
rect 631791 994516 631857 994519
rect 573135 994514 631857 994516
rect 573135 994458 573140 994514
rect 573196 994458 631796 994514
rect 631852 994458 631857 994514
rect 573135 994456 631857 994458
rect 573135 994453 573201 994456
rect 631791 994453 631857 994456
rect 573039 994368 573105 994371
rect 630927 994368 630993 994371
rect 573039 994366 630993 994368
rect 573039 994310 573044 994366
rect 573100 994310 630932 994366
rect 630988 994310 630993 994366
rect 573039 994308 630993 994310
rect 573039 994305 573105 994308
rect 630927 994305 630993 994308
rect 283503 994220 283569 994223
rect 304815 994220 304881 994223
rect 283503 994218 304881 994220
rect 283503 994162 283508 994218
rect 283564 994162 304820 994218
rect 304876 994162 304881 994218
rect 283503 994160 304881 994162
rect 283503 994157 283569 994160
rect 304815 994157 304881 994160
rect 573231 994220 573297 994223
rect 636111 994220 636177 994223
rect 573231 994218 636177 994220
rect 573231 994162 573236 994218
rect 573292 994162 636116 994218
rect 636172 994162 636177 994218
rect 573231 994160 636177 994162
rect 573231 994157 573297 994160
rect 636111 994157 636177 994160
rect 231471 994070 259518 994072
rect 231471 994014 231476 994070
rect 231532 994014 259518 994070
rect 231471 994012 259518 994014
rect 282831 994072 282897 994075
rect 310863 994072 310929 994075
rect 282831 994070 310929 994072
rect 282831 994014 282836 994070
rect 282892 994014 310868 994070
rect 310924 994014 310929 994070
rect 282831 994012 310929 994014
rect 231471 994009 231537 994012
rect 282831 994009 282897 994012
rect 310863 994009 310929 994012
rect 567375 994072 567441 994075
rect 629967 994072 630033 994075
rect 567375 994070 630033 994072
rect 567375 994014 567380 994070
rect 567436 994014 629972 994070
rect 630028 994014 630033 994070
rect 567375 994012 630033 994014
rect 567375 994009 567441 994012
rect 629967 994009 630033 994012
rect 136143 993922 155742 993924
rect 136143 993866 136148 993922
rect 136204 993866 155742 993922
rect 136143 993864 155742 993866
rect 243183 993924 243249 993927
rect 316719 993924 316785 993927
rect 243183 993922 316785 993924
rect 243183 993866 243188 993922
rect 243244 993866 316724 993922
rect 316780 993866 316785 993922
rect 243183 993864 316785 993866
rect 136143 993861 136209 993864
rect 243183 993861 243249 993864
rect 316719 993861 316785 993864
rect 374511 993924 374577 993927
rect 392079 993924 392145 993927
rect 374511 993922 392145 993924
rect 374511 993866 374516 993922
rect 374572 993866 392084 993922
rect 392140 993866 392145 993922
rect 374511 993864 392145 993866
rect 374511 993861 374577 993864
rect 392079 993861 392145 993864
rect 471663 993924 471729 993927
rect 484143 993924 484209 993927
rect 471663 993922 484209 993924
rect 471663 993866 471668 993922
rect 471724 993866 484148 993922
rect 484204 993866 484209 993922
rect 471663 993864 484209 993866
rect 471663 993861 471729 993864
rect 484143 993861 484209 993864
rect 574671 993924 574737 993927
rect 639183 993924 639249 993927
rect 574671 993922 639249 993924
rect 574671 993866 574676 993922
rect 574732 993866 639188 993922
rect 639244 993866 639249 993922
rect 574671 993864 639249 993866
rect 574671 993861 574737 993864
rect 639183 993861 639249 993864
rect 80175 993776 80241 993779
rect 104463 993776 104529 993779
rect 80175 993774 104529 993776
rect 80175 993718 80180 993774
rect 80236 993718 104468 993774
rect 104524 993718 104529 993774
rect 80175 993716 104529 993718
rect 80175 993713 80241 993716
rect 104463 993713 104529 993716
rect 129711 993776 129777 993779
rect 157359 993776 157425 993779
rect 129711 993774 157425 993776
rect 129711 993718 129716 993774
rect 129772 993718 157364 993774
rect 157420 993718 157425 993774
rect 129711 993716 157425 993718
rect 129711 993713 129777 993716
rect 157359 993713 157425 993716
rect 191535 993776 191601 993779
rect 251823 993776 251889 993779
rect 191535 993774 251889 993776
rect 191535 993718 191540 993774
rect 191596 993718 251828 993774
rect 251884 993718 251889 993774
rect 191535 993716 251889 993718
rect 191535 993713 191601 993716
rect 251823 993713 251889 993716
rect 294543 993776 294609 993779
rect 373935 993776 374001 993779
rect 294543 993774 374001 993776
rect 294543 993718 294548 993774
rect 294604 993718 373940 993774
rect 373996 993718 374001 993774
rect 294543 993716 374001 993718
rect 294543 993713 294609 993716
rect 373935 993713 374001 993716
rect 374607 993776 374673 993779
rect 396975 993776 397041 993779
rect 374607 993774 397041 993776
rect 374607 993718 374612 993774
rect 374668 993718 396980 993774
rect 397036 993718 397041 993774
rect 374607 993716 397041 993718
rect 374607 993713 374673 993716
rect 396975 993713 397041 993716
rect 466575 993776 466641 993779
rect 485967 993776 486033 993779
rect 466575 993774 486033 993776
rect 466575 993718 466580 993774
rect 466636 993718 485972 993774
rect 486028 993718 486033 993774
rect 466575 993716 486033 993718
rect 466575 993713 466641 993716
rect 485967 993713 486033 993716
rect 572943 993776 573009 993779
rect 637359 993776 637425 993779
rect 572943 993774 637425 993776
rect 572943 993718 572948 993774
rect 573004 993718 637364 993774
rect 637420 993718 637425 993774
rect 572943 993716 637425 993718
rect 572943 993713 573009 993716
rect 637359 993713 637425 993716
rect 638511 993776 638577 993779
rect 641103 993776 641169 993779
rect 638511 993774 641169 993776
rect 638511 993718 638516 993774
rect 638572 993718 641108 993774
rect 641164 993718 641169 993774
rect 638511 993716 641169 993718
rect 638511 993713 638577 993716
rect 641103 993713 641169 993716
rect 59535 976016 59601 976019
rect 59535 976014 64416 976016
rect 59535 975958 59540 976014
rect 59596 975958 64416 976014
rect 59535 975956 64416 975958
rect 59535 975953 59601 975956
rect 655215 975868 655281 975871
rect 650208 975866 655281 975868
rect 650208 975810 655220 975866
rect 655276 975810 655281 975866
rect 650208 975808 655281 975810
rect 655215 975805 655281 975808
rect 42159 968766 42225 968767
rect 42106 968764 42112 968766
rect 42068 968704 42112 968764
rect 42176 968762 42225 968766
rect 42220 968706 42225 968762
rect 42106 968702 42112 968704
rect 42176 968702 42225 968706
rect 42159 968701 42225 968702
rect 41775 967138 41841 967139
rect 41722 967136 41728 967138
rect 41684 967076 41728 967136
rect 41792 967134 41841 967138
rect 41836 967078 41841 967134
rect 41722 967074 41728 967076
rect 41792 967074 41841 967078
rect 41775 967073 41841 967074
rect 674362 966186 674368 966250
rect 674432 966248 674438 966250
rect 675375 966248 675441 966251
rect 674432 966246 675441 966248
rect 674432 966190 675380 966246
rect 675436 966190 675441 966246
rect 674432 966188 675441 966190
rect 674432 966186 674438 966188
rect 675375 966185 675441 966188
rect 674170 965742 674176 965806
rect 674240 965804 674246 965806
rect 675471 965804 675537 965807
rect 674240 965802 675537 965804
rect 674240 965746 675476 965802
rect 675532 965746 675537 965802
rect 674240 965744 675537 965746
rect 674240 965742 674246 965744
rect 675471 965741 675537 965744
rect 40570 965002 40576 965066
rect 40640 965064 40646 965066
rect 41775 965064 41841 965067
rect 40640 965062 41841 965064
rect 40640 965006 41780 965062
rect 41836 965006 41841 965062
rect 40640 965004 41841 965006
rect 40640 965002 40646 965004
rect 41775 965001 41841 965004
rect 674554 965002 674560 965066
rect 674624 965064 674630 965066
rect 675471 965064 675537 965067
rect 674624 965062 675537 965064
rect 674624 965006 675476 965062
rect 675532 965006 675537 965062
rect 674624 965004 675537 965006
rect 674624 965002 674630 965004
rect 675471 965001 675537 965004
rect 40762 963966 40768 964030
rect 40832 964028 40838 964030
rect 41775 964028 41841 964031
rect 40832 964026 41841 964028
rect 40832 963970 41780 964026
rect 41836 963970 41841 964026
rect 40832 963968 41841 963970
rect 40832 963966 40838 963968
rect 41775 963965 41841 963968
rect 40954 963374 40960 963438
rect 41024 963436 41030 963438
rect 41775 963436 41841 963439
rect 41024 963434 41841 963436
rect 41024 963378 41780 963434
rect 41836 963378 41841 963434
rect 41024 963376 41841 963378
rect 41024 963374 41030 963376
rect 41775 963373 41841 963376
rect 674746 963374 674752 963438
rect 674816 963436 674822 963438
rect 675375 963436 675441 963439
rect 674816 963434 675441 963436
rect 674816 963378 675380 963434
rect 675436 963378 675441 963434
rect 674816 963376 675441 963378
rect 674816 963374 674822 963376
rect 675375 963373 675441 963376
rect 59535 962992 59601 962995
rect 59535 962990 64416 962992
rect 59535 962934 59540 962990
rect 59596 962934 64416 962990
rect 59535 962932 64416 962934
rect 59535 962929 59601 962932
rect 41146 962782 41152 962846
rect 41216 962844 41222 962846
rect 41775 962844 41841 962847
rect 41216 962842 41841 962844
rect 41216 962786 41780 962842
rect 41836 962786 41841 962842
rect 41216 962784 41841 962786
rect 41216 962782 41222 962784
rect 41775 962781 41841 962784
rect 674938 962634 674944 962698
rect 675008 962696 675014 962698
rect 675471 962696 675537 962699
rect 675008 962694 675537 962696
rect 675008 962638 675476 962694
rect 675532 962638 675537 962694
rect 675008 962636 675537 962638
rect 675008 962634 675014 962636
rect 675471 962633 675537 962636
rect 655503 962548 655569 962551
rect 650208 962546 655569 962548
rect 650208 962490 655508 962546
rect 655564 962490 655569 962546
rect 650208 962488 655569 962490
rect 655503 962485 655569 962488
rect 41530 962190 41536 962254
rect 41600 962252 41606 962254
rect 41775 962252 41841 962255
rect 675759 962254 675825 962255
rect 675706 962252 675712 962254
rect 41600 962250 41841 962252
rect 41600 962194 41780 962250
rect 41836 962194 41841 962250
rect 41600 962192 41841 962194
rect 675668 962192 675712 962252
rect 675776 962250 675825 962254
rect 675820 962194 675825 962250
rect 41600 962190 41606 962192
rect 41775 962189 41841 962192
rect 675706 962190 675712 962192
rect 675776 962190 675825 962194
rect 675759 962189 675825 962190
rect 41338 959526 41344 959590
rect 41408 959588 41414 959590
rect 41775 959588 41841 959591
rect 41408 959586 41841 959588
rect 41408 959530 41780 959586
rect 41836 959530 41841 959586
rect 41408 959528 41841 959530
rect 41408 959526 41414 959528
rect 41775 959525 41841 959528
rect 40378 959082 40384 959146
rect 40448 959144 40454 959146
rect 41775 959144 41841 959147
rect 40448 959142 41841 959144
rect 40448 959086 41780 959142
rect 41836 959086 41841 959142
rect 40448 959084 41841 959086
rect 40448 959082 40454 959084
rect 41775 959081 41841 959084
rect 675130 959082 675136 959146
rect 675200 959144 675206 959146
rect 675471 959144 675537 959147
rect 675200 959142 675537 959144
rect 675200 959086 675476 959142
rect 675532 959086 675537 959142
rect 675200 959084 675537 959086
rect 675200 959082 675206 959084
rect 675471 959081 675537 959084
rect 675759 958404 675825 958407
rect 676858 958404 676864 958406
rect 675759 958402 676864 958404
rect 675759 958346 675764 958402
rect 675820 958346 676864 958402
rect 675759 958344 676864 958346
rect 675759 958341 675825 958344
rect 676858 958342 676864 958344
rect 676928 958342 676934 958406
rect 41871 957814 41937 957815
rect 41871 957810 41920 957814
rect 41984 957812 41990 957814
rect 41871 957754 41876 957810
rect 41871 957750 41920 957754
rect 41984 957752 42028 957812
rect 41984 957750 41990 957752
rect 41871 957749 41937 957750
rect 675375 957666 675441 957667
rect 675322 957664 675328 957666
rect 675284 957604 675328 957664
rect 675392 957662 675441 957666
rect 675436 957606 675441 957662
rect 675322 957602 675328 957604
rect 675392 957602 675441 957606
rect 675375 957601 675441 957602
rect 42255 957518 42321 957519
rect 42255 957516 42304 957518
rect 42212 957514 42304 957516
rect 42212 957458 42260 957514
rect 42212 957456 42304 957458
rect 42255 957454 42304 957456
rect 42368 957454 42374 957518
rect 42255 957453 42321 957454
rect 675759 957070 675825 957075
rect 675759 957014 675764 957070
rect 675820 957014 675825 957070
rect 675759 957009 675825 957014
rect 42255 956332 42321 956335
rect 42490 956332 42496 956334
rect 42255 956330 42496 956332
rect 42255 956274 42260 956330
rect 42316 956274 42496 956330
rect 42255 956272 42496 956274
rect 42255 956269 42321 956272
rect 42490 956270 42496 956272
rect 42560 956270 42566 956334
rect 675762 956184 675822 957009
rect 675762 956124 677118 956184
rect 675567 956038 675633 956039
rect 677058 956038 677118 956124
rect 675514 956036 675520 956038
rect 675476 955976 675520 956036
rect 675584 956034 675633 956038
rect 675628 955978 675633 956034
rect 675514 955974 675520 955976
rect 675584 955974 675633 955978
rect 677050 955974 677056 956038
rect 677120 955974 677126 956038
rect 675567 955973 675633 955974
rect 673978 953902 673984 953966
rect 674048 953964 674054 953966
rect 675471 953964 675537 953967
rect 674048 953962 675537 953964
rect 674048 953906 675476 953962
rect 675532 953906 675537 953962
rect 674048 953904 675537 953906
rect 674048 953902 674054 953904
rect 675471 953901 675537 953904
rect 674703 953372 674769 953375
rect 677050 953372 677056 953374
rect 674703 953370 677056 953372
rect 674703 953314 674708 953370
rect 674764 953314 677056 953370
rect 674703 953312 677056 953314
rect 674703 953309 674769 953312
rect 677050 953310 677056 953312
rect 677120 953310 677126 953374
rect 675759 952040 675825 952043
rect 675898 952040 675904 952042
rect 675759 952038 675904 952040
rect 675759 951982 675764 952038
rect 675820 951982 675904 952038
rect 675759 951980 675904 951982
rect 675759 951977 675825 951980
rect 675898 951978 675904 951980
rect 675968 951978 675974 952042
rect 59535 949968 59601 949971
rect 59535 949966 64416 949968
rect 59535 949910 59540 949966
rect 59596 949910 64416 949966
rect 59535 949908 64416 949910
rect 59535 949905 59601 949908
rect 655695 949376 655761 949379
rect 650208 949374 655761 949376
rect 650208 949318 655700 949374
rect 655756 949318 655761 949374
rect 650208 949316 655761 949318
rect 655695 949313 655761 949316
rect 34479 945084 34545 945087
rect 34434 945082 34545 945084
rect 34434 945026 34484 945082
rect 34540 945026 34545 945082
rect 34434 945021 34545 945026
rect 34434 944906 34494 945021
rect 39810 944051 39870 944314
rect 39759 944046 39870 944051
rect 39759 943990 39764 944046
rect 39820 943990 39870 944046
rect 39759 943988 39870 943990
rect 39759 943985 39825 943988
rect 41775 943826 41841 943829
rect 41568 943824 41841 943826
rect 41568 943768 41780 943824
rect 41836 943768 41841 943824
rect 41568 943766 41841 943768
rect 41775 943763 41841 943766
rect 41583 943604 41649 943607
rect 41538 943602 41649 943604
rect 41538 943546 41588 943602
rect 41644 943546 41649 943602
rect 41538 943541 41649 943546
rect 41538 943426 41598 943541
rect 40386 942719 40446 942834
rect 40386 942714 40497 942719
rect 40386 942658 40436 942714
rect 40492 942658 40497 942714
rect 40386 942656 40497 942658
rect 40431 942653 40497 942656
rect 41538 942124 41598 942316
rect 41679 942124 41745 942127
rect 41538 942122 41745 942124
rect 41538 942066 41684 942122
rect 41740 942066 41745 942122
rect 41538 942064 41745 942066
rect 41679 942061 41745 942064
rect 40194 941683 40254 941946
rect 40194 941678 40305 941683
rect 40194 941622 40244 941678
rect 40300 941622 40305 941678
rect 40194 941620 40305 941622
rect 40239 941617 40305 941620
rect 40386 941091 40446 941354
rect 40335 941086 40446 941091
rect 40335 941030 40340 941086
rect 40396 941030 40446 941086
rect 40335 941028 40446 941030
rect 676143 941088 676209 941091
rect 676290 941088 676350 941280
rect 676143 941086 676350 941088
rect 676143 941030 676148 941086
rect 676204 941030 676350 941086
rect 676143 941028 676350 941030
rect 40335 941025 40401 941028
rect 676143 941025 676209 941028
rect 41538 940647 41598 940762
rect 41538 940642 41649 940647
rect 41538 940586 41588 940642
rect 41644 940586 41649 940642
rect 41538 940584 41649 940586
rect 41583 940581 41649 940584
rect 676290 940499 676350 940762
rect 42490 940496 42496 940498
rect 41538 940436 42496 940496
rect 41538 940392 41598 940436
rect 42490 940434 42496 940436
rect 42560 940434 42566 940498
rect 676290 940494 676401 940499
rect 676290 940438 676340 940494
rect 676396 940438 676401 940494
rect 676290 940436 676401 940438
rect 676335 940433 676401 940436
rect 676290 940055 676350 940170
rect 676239 940050 676350 940055
rect 676239 939994 676244 940050
rect 676300 939994 676350 940050
rect 676239 939992 676350 939994
rect 676239 939989 676305 939992
rect 41722 939904 41728 939906
rect 41568 939844 41728 939904
rect 41722 939842 41728 939844
rect 41792 939842 41798 939906
rect 676047 939756 676113 939759
rect 676047 939754 676320 939756
rect 676047 939698 676052 939754
rect 676108 939698 676320 939754
rect 676047 939696 676320 939698
rect 676047 939693 676113 939696
rect 42255 939312 42321 939315
rect 41568 939310 42321 939312
rect 41568 939254 42260 939310
rect 42316 939254 42321 939310
rect 41568 939252 42321 939254
rect 42255 939249 42321 939252
rect 676047 939312 676113 939315
rect 676047 939310 676320 939312
rect 676047 939254 676052 939310
rect 676108 939254 676320 939310
rect 676047 939252 676320 939254
rect 676047 939249 676113 939252
rect 41914 938942 41920 938944
rect 41568 938882 41920 938942
rect 41914 938880 41920 938882
rect 41984 938880 41990 938944
rect 676239 938868 676305 938871
rect 676239 938866 676350 938868
rect 676239 938810 676244 938866
rect 676300 938810 676350 938866
rect 676239 938805 676350 938810
rect 41530 938658 41536 938722
rect 41600 938658 41606 938722
rect 676290 938690 676350 938805
rect 41538 938394 41598 938658
rect 676290 938131 676350 938246
rect 676239 938126 676350 938131
rect 676239 938070 676244 938126
rect 676300 938070 676350 938126
rect 676239 938068 676350 938070
rect 676239 938065 676305 938068
rect 42106 937832 42112 937834
rect 41568 937772 42112 937832
rect 42106 937770 42112 937772
rect 42176 937770 42182 937834
rect 676047 937758 676113 937761
rect 676047 937756 676320 937758
rect 676047 937700 676052 937756
rect 676108 937700 676320 937756
rect 676047 937698 676320 937700
rect 676047 937695 676113 937698
rect 38799 937684 38865 937687
rect 38799 937682 38910 937684
rect 38799 937626 38804 937682
rect 38860 937626 38910 937682
rect 38799 937621 38910 937626
rect 38850 937358 38910 937621
rect 676047 937240 676113 937243
rect 676047 937238 676320 937240
rect 676047 937182 676052 937238
rect 676108 937182 676320 937238
rect 676047 937180 676320 937182
rect 676047 937177 676113 937180
rect 42298 936944 42304 936946
rect 41568 936884 42304 936944
rect 42298 936882 42304 936884
rect 42368 936882 42374 936946
rect 59535 936944 59601 936947
rect 59535 936942 64416 936944
rect 59535 936886 59540 936942
rect 59596 936886 64416 936942
rect 59535 936884 64416 936886
rect 59535 936881 59601 936884
rect 674554 936734 674560 936798
rect 674624 936796 674630 936798
rect 674624 936736 676320 936796
rect 674624 936734 674630 936736
rect 40378 936586 40384 936650
rect 40448 936586 40454 936650
rect 673978 936586 673984 936650
rect 674048 936648 674054 936650
rect 674048 936588 676350 936648
rect 674048 936586 674054 936588
rect 40386 936322 40446 936586
rect 676290 936248 676350 936588
rect 655599 936204 655665 936207
rect 650208 936202 655665 936204
rect 650208 936146 655604 936202
rect 655660 936146 655665 936202
rect 650208 936144 655665 936146
rect 655599 936141 655665 936144
rect 40578 935762 40638 935878
rect 40570 935698 40576 935762
rect 40640 935698 40646 935762
rect 40954 935698 40960 935762
rect 41024 935698 41030 935762
rect 674362 935698 674368 935762
rect 674432 935760 674438 935762
rect 674432 935700 676320 935760
rect 674432 935698 674438 935700
rect 40962 935360 41022 935698
rect 674746 935254 674752 935318
rect 674816 935316 674822 935318
rect 674816 935256 676320 935316
rect 674816 935254 674822 935256
rect 41338 935106 41344 935170
rect 41408 935106 41414 935170
rect 41346 934842 41406 935106
rect 675130 934662 675136 934726
rect 675200 934724 675206 934726
rect 675200 934664 676320 934724
rect 675200 934662 675206 934664
rect 41154 934282 41214 934398
rect 40762 934218 40768 934282
rect 40832 934218 40838 934282
rect 41146 934218 41152 934282
rect 41216 934218 41222 934282
rect 675898 934218 675904 934282
rect 675968 934280 675974 934282
rect 675968 934220 676320 934280
rect 675968 934218 675974 934220
rect 40770 933880 40830 934218
rect 674170 933774 674176 933838
rect 674240 933836 674246 933838
rect 674240 933776 676320 933836
rect 674240 933774 674246 933776
rect 41568 933332 41790 933392
rect 28866 932655 28926 932918
rect 41730 932800 41790 933332
rect 674938 933182 674944 933246
rect 675008 933244 675014 933246
rect 675008 933184 676320 933244
rect 675008 933182 675014 933184
rect 28815 932650 28926 932655
rect 28815 932594 28820 932650
rect 28876 932594 28926 932650
rect 28815 932592 28926 932594
rect 41538 932740 41790 932800
rect 28815 932589 28881 932592
rect 41538 932211 41598 932740
rect 675706 932664 675712 932728
rect 675776 932726 675782 932728
rect 675776 932666 676320 932726
rect 675776 932664 675782 932666
rect 675514 932294 675520 932358
rect 675584 932356 675590 932358
rect 675584 932296 676320 932356
rect 675584 932294 675590 932296
rect 28815 932208 28881 932211
rect 28815 932206 28926 932208
rect 28815 932150 28820 932206
rect 28876 932150 28926 932206
rect 28815 932145 28926 932150
rect 41538 932206 41649 932211
rect 41538 932150 41588 932206
rect 41644 932150 41649 932206
rect 41538 932148 41649 932150
rect 41583 932145 41649 932148
rect 28866 931882 28926 932145
rect 675322 931702 675328 931766
rect 675392 931764 675398 931766
rect 675392 931704 676320 931764
rect 675392 931702 675398 931704
rect 677050 931554 677056 931618
rect 677120 931554 677126 931618
rect 677058 931216 677118 931554
rect 676858 930962 676864 931026
rect 676928 930962 676934 931026
rect 676866 930846 676926 930962
rect 677242 930518 677248 930582
rect 677312 930518 677318 930582
rect 677250 930254 677310 930518
rect 679746 929547 679806 929662
rect 679746 929542 679857 929547
rect 679746 929486 679796 929542
rect 679852 929486 679857 929542
rect 679746 929484 679857 929486
rect 679791 929481 679857 929484
rect 685506 928955 685566 929292
rect 679791 928952 679857 928955
rect 679746 928950 679857 928952
rect 679746 928894 679796 928950
rect 679852 928894 679857 928950
rect 679746 928889 679857 928894
rect 685455 928950 685566 928955
rect 685455 928894 685460 928950
rect 685516 928894 685566 928950
rect 685455 928892 685566 928894
rect 685455 928889 685521 928892
rect 679746 928774 679806 928889
rect 685455 928508 685521 928511
rect 685455 928506 685566 928508
rect 685455 928450 685460 928506
rect 685516 928450 685566 928506
rect 685455 928445 685566 928450
rect 685506 928182 685566 928445
rect 58575 923772 58641 923775
rect 58575 923770 64416 923772
rect 58575 923714 58580 923770
rect 58636 923714 64416 923770
rect 58575 923712 64416 923714
rect 58575 923709 58641 923712
rect 656367 922736 656433 922739
rect 650208 922734 656433 922736
rect 650208 922678 656372 922734
rect 656428 922678 656433 922734
rect 650208 922676 656433 922678
rect 656367 922673 656433 922676
rect 59535 910748 59601 910751
rect 59535 910746 64416 910748
rect 59535 910690 59540 910746
rect 59596 910690 64416 910746
rect 59535 910688 64416 910690
rect 59535 910685 59601 910688
rect 654447 909564 654513 909567
rect 650208 909562 654513 909564
rect 650208 909506 654452 909562
rect 654508 909506 654513 909562
rect 650208 909504 654513 909506
rect 654447 909501 654513 909504
rect 59535 897872 59601 897875
rect 59535 897870 64416 897872
rect 59535 897814 59540 897870
rect 59596 897814 64416 897870
rect 59535 897812 64416 897814
rect 59535 897809 59601 897812
rect 654447 896244 654513 896247
rect 650208 896242 654513 896244
rect 650208 896186 654452 896242
rect 654508 896186 654513 896242
rect 650208 896184 654513 896186
rect 654447 896181 654513 896184
rect 57999 884848 58065 884851
rect 57999 884846 64416 884848
rect 57999 884790 58004 884846
rect 58060 884790 64416 884846
rect 57999 884788 64416 884790
rect 57999 884785 58065 884788
rect 656559 882924 656625 882927
rect 650208 882922 656625 882924
rect 650208 882866 656564 882922
rect 656620 882866 656625 882922
rect 650208 882864 656625 882866
rect 656559 882861 656625 882864
rect 673978 876350 673984 876414
rect 674048 876412 674054 876414
rect 675279 876412 675345 876415
rect 674048 876410 675345 876412
rect 674048 876354 675284 876410
rect 675340 876354 675345 876410
rect 674048 876352 675345 876354
rect 674048 876350 674054 876352
rect 675279 876349 675345 876352
rect 674170 876202 674176 876266
rect 674240 876264 674246 876266
rect 675279 876264 675345 876267
rect 674240 876262 675345 876264
rect 674240 876206 675284 876262
rect 675340 876206 675345 876262
rect 674240 876204 675345 876206
rect 674240 876202 674246 876204
rect 675279 876201 675345 876204
rect 674362 873982 674368 874046
rect 674432 874044 674438 874046
rect 675471 874044 675537 874047
rect 674432 874042 675537 874044
rect 674432 873986 675476 874042
rect 675532 873986 675537 874042
rect 674432 873984 675537 873986
rect 674432 873982 674438 873984
rect 675471 873981 675537 873984
rect 59535 871676 59601 871679
rect 59535 871674 64416 871676
rect 59535 871618 59540 871674
rect 59596 871618 64416 871674
rect 59535 871616 64416 871618
rect 59535 871613 59601 871616
rect 674554 869838 674560 869902
rect 674624 869900 674630 869902
rect 675375 869900 675441 869903
rect 674624 869898 675441 869900
rect 674624 869842 675380 869898
rect 675436 869842 675441 869898
rect 674624 869840 675441 869842
rect 674624 869838 674630 869840
rect 675375 869837 675441 869840
rect 654447 869752 654513 869755
rect 650208 869750 654513 869752
rect 650208 869694 654452 869750
rect 654508 869694 654513 869750
rect 650208 869692 654513 869694
rect 654447 869689 654513 869692
rect 675759 864722 675825 864723
rect 675706 864720 675712 864722
rect 675668 864660 675712 864720
rect 675776 864718 675825 864722
rect 675820 864662 675825 864718
rect 675706 864658 675712 864660
rect 675776 864658 675825 864662
rect 675759 864657 675825 864658
rect 674938 862882 674944 862946
rect 675008 862944 675014 862946
rect 675375 862944 675441 862947
rect 675008 862942 675441 862944
rect 675008 862886 675380 862942
rect 675436 862886 675441 862942
rect 675008 862884 675441 862886
rect 675008 862882 675014 862884
rect 675375 862881 675441 862884
rect 58383 858652 58449 858655
rect 58383 858650 64416 858652
rect 58383 858594 58388 858650
rect 58444 858594 64416 858650
rect 58383 858592 64416 858594
rect 58383 858589 58449 858592
rect 654447 856432 654513 856435
rect 650208 856430 654513 856432
rect 650208 856374 654452 856430
rect 654508 856374 654513 856430
rect 650208 856372 654513 856374
rect 654447 856369 654513 856372
rect 59535 845628 59601 845631
rect 59535 845626 64416 845628
rect 59535 845570 59540 845626
rect 59596 845570 64416 845626
rect 59535 845568 64416 845570
rect 59535 845565 59601 845568
rect 654447 842964 654513 842967
rect 650208 842962 654513 842964
rect 650208 842906 654452 842962
rect 654508 842906 654513 842962
rect 650208 842904 654513 842906
rect 654447 842901 654513 842904
rect 59535 832604 59601 832607
rect 59535 832602 64416 832604
rect 59535 832546 59540 832602
rect 59596 832546 64416 832602
rect 59535 832544 64416 832546
rect 59535 832541 59601 832544
rect 654735 829792 654801 829795
rect 650208 829790 654801 829792
rect 650208 829734 654740 829790
rect 654796 829734 654801 829790
rect 650208 829732 654801 829734
rect 654735 829729 654801 829732
rect 59535 819432 59601 819435
rect 59535 819430 64416 819432
rect 59535 819374 59540 819430
rect 59596 819374 64416 819430
rect 59535 819372 64416 819374
rect 59535 819369 59601 819372
rect 41583 819284 41649 819287
rect 41538 819282 41649 819284
rect 41538 819226 41588 819282
rect 41644 819226 41649 819282
rect 41538 819221 41649 819226
rect 41538 819106 41598 819221
rect 41775 818544 41841 818547
rect 41568 818542 41841 818544
rect 41568 818486 41780 818542
rect 41836 818486 41841 818542
rect 41568 818484 41841 818486
rect 41775 818481 41841 818484
rect 41775 817952 41841 817955
rect 41568 817950 41841 817952
rect 41568 817894 41780 817950
rect 41836 817894 41841 817950
rect 41568 817892 41841 817894
rect 41775 817889 41841 817892
rect 40431 817804 40497 817807
rect 40386 817802 40497 817804
rect 40386 817746 40436 817802
rect 40492 817746 40497 817802
rect 40386 817741 40497 817746
rect 40386 817626 40446 817741
rect 41775 817064 41841 817067
rect 41568 817062 41841 817064
rect 41568 817006 41780 817062
rect 41836 817006 41841 817062
rect 41568 817004 41841 817006
rect 41775 817001 41841 817004
rect 655503 816472 655569 816475
rect 650208 816470 655569 816472
rect 39951 816324 40017 816327
rect 40770 816326 40830 816442
rect 650208 816414 655508 816470
rect 655564 816414 655569 816470
rect 650208 816412 655569 816414
rect 655503 816409 655569 816412
rect 39951 816322 40062 816324
rect 39951 816266 39956 816322
rect 40012 816266 40062 816322
rect 39951 816261 40062 816266
rect 40762 816262 40768 816326
rect 40832 816262 40838 816326
rect 40002 816072 40062 816261
rect 41154 815290 41214 815554
rect 41146 815226 41152 815290
rect 41216 815226 41222 815290
rect 42106 814992 42112 814994
rect 41568 814962 42112 814992
rect 41538 814932 42112 814962
rect 40335 814844 40401 814847
rect 41538 814844 41598 814932
rect 42106 814930 42112 814932
rect 42176 814930 42182 814994
rect 40335 814842 41598 814844
rect 40335 814786 40340 814842
rect 40396 814786 41598 814842
rect 40335 814784 41598 814786
rect 40335 814781 40401 814784
rect 42063 814622 42129 814625
rect 41568 814620 42129 814622
rect 41568 814564 42068 814620
rect 42124 814564 42129 814620
rect 41568 814562 42129 814564
rect 42063 814559 42129 814562
rect 41775 814104 41841 814107
rect 41568 814102 41841 814104
rect 41568 814046 41780 814102
rect 41836 814046 41841 814102
rect 41568 814044 41841 814046
rect 41775 814041 41841 814044
rect 34434 813367 34494 813482
rect 34383 813362 34494 813367
rect 34383 813306 34388 813362
rect 34444 813306 34494 813362
rect 34383 813304 34494 813306
rect 34383 813301 34449 813304
rect 41538 812923 41598 813038
rect 41538 812918 41649 812923
rect 41538 812862 41588 812918
rect 41644 812862 41649 812918
rect 41538 812860 41649 812862
rect 41583 812857 41649 812860
rect 42351 812624 42417 812627
rect 41568 812622 42417 812624
rect 41568 812566 42356 812622
rect 42412 812566 42417 812622
rect 41568 812564 42417 812566
rect 42351 812561 42417 812564
rect 41871 812032 41937 812035
rect 41568 812030 41937 812032
rect 41568 811974 41876 812030
rect 41932 811974 41937 812030
rect 41568 811972 41937 811974
rect 41871 811969 41937 811972
rect 34434 811443 34494 811558
rect 34434 811438 34545 811443
rect 34434 811382 34484 811438
rect 34540 811382 34545 811438
rect 34434 811380 34545 811382
rect 34479 811377 34545 811380
rect 41967 811070 42033 811073
rect 41568 811068 42033 811070
rect 41568 811012 41972 811068
rect 42028 811012 42033 811068
rect 41568 811010 42033 811012
rect 41967 811007 42033 811010
rect 41487 810700 41553 810703
rect 41487 810698 41598 810700
rect 41487 810642 41492 810698
rect 41548 810642 41598 810698
rect 41487 810637 41598 810642
rect 41538 810522 41598 810637
rect 41775 810108 41841 810111
rect 41568 810106 41841 810108
rect 41568 810050 41780 810106
rect 41836 810050 41841 810106
rect 41568 810048 41841 810050
rect 41775 810045 41841 810048
rect 41538 809368 41598 809560
rect 41679 809368 41745 809371
rect 41538 809366 41745 809368
rect 41538 809310 41684 809366
rect 41740 809310 41745 809366
rect 41538 809308 41745 809310
rect 41679 809305 41745 809308
rect 42159 809072 42225 809075
rect 41568 809070 42225 809072
rect 41568 809014 42164 809070
rect 42220 809014 42225 809070
rect 41568 809012 42225 809014
rect 42159 809009 42225 809012
rect 41967 808628 42033 808631
rect 41568 808626 42033 808628
rect 41568 808570 41972 808626
rect 42028 808570 42033 808626
rect 41568 808568 42033 808570
rect 41967 808565 42033 808568
rect 41538 807891 41598 808006
rect 41538 807886 41649 807891
rect 41538 807830 41588 807886
rect 41644 807830 41649 807886
rect 41538 807828 41649 807830
rect 41583 807825 41649 807828
rect 41538 807296 41598 807562
rect 41538 807236 41790 807296
rect 23106 806855 23166 807118
rect 23055 806850 23166 806855
rect 41730 806852 41790 807236
rect 23055 806794 23060 806850
rect 23116 806794 23166 806850
rect 23055 806792 23166 806794
rect 41538 806792 41790 806852
rect 23055 806789 23121 806792
rect 41538 806411 41598 806792
rect 59535 806556 59601 806559
rect 59535 806554 64416 806556
rect 59535 806498 59540 806554
rect 59596 806498 64416 806554
rect 59535 806496 64416 806498
rect 59535 806493 59601 806496
rect 23055 806408 23121 806411
rect 23055 806406 23166 806408
rect 23055 806350 23060 806406
rect 23116 806350 23166 806406
rect 23055 806345 23166 806350
rect 41538 806406 41649 806411
rect 41538 806350 41588 806406
rect 41644 806350 41649 806406
rect 41538 806348 41649 806350
rect 41583 806345 41649 806348
rect 23106 806008 23166 806345
rect 654447 803152 654513 803155
rect 650208 803150 654513 803152
rect 650208 803094 654452 803150
rect 654508 803094 654513 803150
rect 650208 803092 654513 803094
rect 654447 803089 654513 803092
rect 34383 802116 34449 802119
rect 41530 802116 41536 802118
rect 34383 802114 41536 802116
rect 34383 802058 34388 802114
rect 34444 802058 41536 802114
rect 34383 802056 41536 802058
rect 34383 802053 34449 802056
rect 41530 802054 41536 802056
rect 41600 802054 41606 802118
rect 34479 801820 34545 801823
rect 41338 801820 41344 801822
rect 34479 801818 41344 801820
rect 34479 801762 34484 801818
rect 34540 801762 41344 801818
rect 34479 801760 41344 801762
rect 34479 801757 34545 801760
rect 41338 801758 41344 801760
rect 41408 801758 41414 801822
rect 41679 800608 41745 800611
rect 41914 800608 41920 800610
rect 41679 800606 41920 800608
rect 41679 800550 41684 800606
rect 41740 800550 41920 800606
rect 41679 800548 41920 800550
rect 41679 800545 41745 800548
rect 41914 800546 41920 800548
rect 41984 800546 41990 800610
rect 41775 800342 41841 800343
rect 41722 800278 41728 800342
rect 41792 800340 41841 800342
rect 41967 800340 42033 800343
rect 42298 800340 42304 800342
rect 41792 800338 41884 800340
rect 41836 800282 41884 800338
rect 41792 800280 41884 800282
rect 41967 800338 42304 800340
rect 41967 800282 41972 800338
rect 42028 800282 42304 800338
rect 41967 800280 42304 800282
rect 41792 800278 41841 800280
rect 41775 800277 41841 800278
rect 41967 800277 42033 800280
rect 42298 800278 42304 800280
rect 42368 800278 42374 800342
rect 42298 797466 42304 797530
rect 42368 797528 42374 797530
rect 42447 797528 42513 797531
rect 42368 797526 42513 797528
rect 42368 797470 42452 797526
rect 42508 797470 42513 797526
rect 42368 797468 42513 797470
rect 42368 797466 42374 797468
rect 42447 797465 42513 797468
rect 41775 796346 41841 796347
rect 41722 796344 41728 796346
rect 41684 796284 41728 796344
rect 41792 796342 41841 796346
rect 41836 796286 41841 796342
rect 41722 796282 41728 796284
rect 41792 796282 41841 796286
rect 41775 796281 41841 796282
rect 41871 794274 41937 794275
rect 41871 794270 41920 794274
rect 41984 794272 41990 794274
rect 41871 794214 41876 794270
rect 41871 794210 41920 794214
rect 41984 794212 42028 794272
rect 41984 794210 41990 794212
rect 41871 794209 41937 794210
rect 59535 793532 59601 793535
rect 59535 793530 64416 793532
rect 59535 793474 59540 793530
rect 59596 793474 64416 793530
rect 59535 793472 64416 793474
rect 59535 793469 59601 793472
rect 41338 790510 41344 790574
rect 41408 790572 41414 790574
rect 42735 790572 42801 790575
rect 41408 790570 42801 790572
rect 41408 790514 42740 790570
rect 42796 790514 42801 790570
rect 41408 790512 42801 790514
rect 41408 790510 41414 790512
rect 42735 790509 42801 790512
rect 655599 789980 655665 789983
rect 650208 789978 655665 789980
rect 650208 789922 655604 789978
rect 655660 789922 655665 789978
rect 650208 789920 655665 789922
rect 655599 789917 655665 789920
rect 41530 789178 41536 789242
rect 41600 789240 41606 789242
rect 42447 789240 42513 789243
rect 41600 789238 42513 789240
rect 41600 789182 42452 789238
rect 42508 789182 42513 789238
rect 41600 789180 42513 789182
rect 41600 789178 41606 789180
rect 42447 789177 42513 789180
rect 675375 787910 675441 787911
rect 675322 787908 675328 787910
rect 675284 787848 675328 787908
rect 675392 787906 675441 787910
rect 675436 787850 675441 787906
rect 675322 787846 675328 787848
rect 675392 787846 675441 787850
rect 675375 787845 675441 787846
rect 675130 786662 675136 786726
rect 675200 786724 675206 786726
rect 675375 786724 675441 786727
rect 675200 786722 675441 786724
rect 675200 786666 675380 786722
rect 675436 786666 675441 786722
rect 675200 786664 675441 786666
rect 675200 786662 675206 786664
rect 675375 786661 675441 786664
rect 675471 784802 675537 784803
rect 675471 784798 675520 784802
rect 675584 784800 675590 784802
rect 675471 784742 675476 784798
rect 675471 784738 675520 784742
rect 675584 784740 675628 784800
rect 675584 784738 675590 784740
rect 675471 784737 675537 784738
rect 675759 780656 675825 780659
rect 676282 780656 676288 780658
rect 675759 780654 676288 780656
rect 675759 780598 675764 780654
rect 675820 780598 676288 780654
rect 675759 780596 676288 780598
rect 675759 780593 675825 780596
rect 676282 780594 676288 780596
rect 676352 780594 676358 780658
rect 59535 780508 59601 780511
rect 59535 780506 64416 780508
rect 59535 780450 59540 780506
rect 59596 780450 64416 780506
rect 59535 780448 64416 780450
rect 59535 780445 59601 780448
rect 675759 779176 675825 779179
rect 676858 779176 676864 779178
rect 675759 779174 676864 779176
rect 675759 779118 675764 779174
rect 675820 779118 676864 779174
rect 675759 779116 676864 779118
rect 675759 779113 675825 779116
rect 676858 779114 676864 779116
rect 676928 779114 676934 779178
rect 674607 777548 674673 777551
rect 677050 777548 677056 777550
rect 674607 777546 677056 777548
rect 674607 777490 674612 777546
rect 674668 777490 677056 777546
rect 674607 777488 677056 777490
rect 674607 777485 674673 777488
rect 677050 777486 677056 777488
rect 677120 777486 677126 777550
rect 675759 777400 675825 777403
rect 677050 777400 677056 777402
rect 675759 777398 677056 777400
rect 675759 777342 675764 777398
rect 675820 777342 677056 777398
rect 675759 777340 677056 777342
rect 675759 777337 675825 777340
rect 677050 777338 677056 777340
rect 677120 777338 677126 777402
rect 655215 776660 655281 776663
rect 650208 776658 655281 776660
rect 650208 776602 655220 776658
rect 655276 776602 655281 776658
rect 650208 776600 655281 776602
rect 655215 776597 655281 776600
rect 41583 776068 41649 776071
rect 41538 776066 41649 776068
rect 41538 776010 41588 776066
rect 41644 776010 41649 776066
rect 41538 776005 41649 776010
rect 41538 775890 41598 776005
rect 675759 775476 675825 775479
rect 675898 775476 675904 775478
rect 675759 775474 675904 775476
rect 675759 775418 675764 775474
rect 675820 775418 675904 775474
rect 675759 775416 675904 775418
rect 675759 775413 675825 775416
rect 675898 775414 675904 775416
rect 675968 775414 675974 775478
rect 41775 775328 41841 775331
rect 41568 775326 41841 775328
rect 41568 775270 41780 775326
rect 41836 775270 41841 775326
rect 41568 775268 41841 775270
rect 41775 775265 41841 775268
rect 674223 774884 674289 774887
rect 677050 774884 677056 774886
rect 674223 774882 677056 774884
rect 674223 774826 674228 774882
rect 674284 774826 677056 774882
rect 674223 774824 677056 774826
rect 674223 774821 674289 774824
rect 677050 774822 677056 774824
rect 677120 774822 677126 774886
rect 41775 774810 41841 774813
rect 41568 774808 41841 774810
rect 41568 774752 41780 774808
rect 41836 774752 41841 774808
rect 41568 774750 41841 774752
rect 41775 774747 41841 774750
rect 41583 774588 41649 774591
rect 41538 774586 41649 774588
rect 41538 774530 41588 774586
rect 41644 774530 41649 774586
rect 41538 774525 41649 774530
rect 41538 774410 41598 774525
rect 41538 773703 41598 773818
rect 41538 773698 41649 773703
rect 41538 773642 41588 773698
rect 41644 773642 41649 773698
rect 41538 773640 41649 773642
rect 41583 773637 41649 773640
rect 674746 773638 674752 773702
rect 674816 773700 674822 773702
rect 675471 773700 675537 773703
rect 674816 773698 675537 773700
rect 674816 773642 675476 773698
rect 675532 773642 675537 773698
rect 674816 773640 675537 773642
rect 674816 773638 674822 773640
rect 675471 773637 675537 773640
rect 42159 773256 42225 773259
rect 40800 773254 42225 773256
rect 40800 773226 42164 773254
rect 40770 773198 42164 773226
rect 42220 773198 42225 773254
rect 40770 773196 42225 773198
rect 40770 773110 40830 773196
rect 42159 773193 42225 773196
rect 40762 773046 40768 773110
rect 40832 773046 40838 773110
rect 40954 773046 40960 773110
rect 41024 773108 41030 773110
rect 41024 773048 41598 773108
rect 41024 773046 41030 773048
rect 41538 772960 41598 773048
rect 45711 772960 45777 772963
rect 41538 772958 45777 772960
rect 41538 772930 45716 772958
rect 41568 772902 45716 772930
rect 45772 772902 45777 772958
rect 41568 772900 45777 772902
rect 45711 772897 45777 772900
rect 42063 772368 42129 772371
rect 40608 772366 42129 772368
rect 40608 772338 42068 772366
rect 40578 772310 42068 772338
rect 42124 772310 42129 772366
rect 40578 772308 42129 772310
rect 40578 772074 40638 772308
rect 42063 772305 42129 772308
rect 40570 772010 40576 772074
rect 40640 772010 40646 772074
rect 41146 772010 41152 772074
rect 41216 772072 41222 772074
rect 41216 772012 41790 772072
rect 41216 772010 41222 772012
rect 41730 771924 41790 772012
rect 42063 771924 42129 771927
rect 41730 771922 42129 771924
rect 41730 771866 42068 771922
rect 42124 771866 42129 771922
rect 41730 771864 42129 771866
rect 41730 771776 41790 771864
rect 42063 771861 42129 771864
rect 41568 771716 41790 771776
rect 41775 771406 41841 771409
rect 41568 771404 41841 771406
rect 41568 771348 41780 771404
rect 41836 771348 41841 771404
rect 41568 771346 41841 771348
rect 41775 771343 41841 771346
rect 40386 770595 40446 770858
rect 40386 770590 40497 770595
rect 40386 770534 40436 770590
rect 40492 770534 40497 770590
rect 40386 770532 40497 770534
rect 40431 770529 40497 770532
rect 33090 770151 33150 770266
rect 33039 770146 33150 770151
rect 33039 770090 33044 770146
rect 33100 770090 33150 770146
rect 33039 770088 33150 770090
rect 33039 770085 33105 770088
rect 41775 769926 41841 769929
rect 41568 769924 41841 769926
rect 41568 769868 41780 769924
rect 41836 769868 41841 769924
rect 41568 769866 41841 769868
rect 41775 769863 41841 769866
rect 41775 769408 41841 769411
rect 41568 769406 41841 769408
rect 41568 769350 41780 769406
rect 41836 769350 41841 769406
rect 41568 769348 41841 769350
rect 41775 769345 41841 769348
rect 40386 768671 40446 768786
rect 40335 768666 40446 768671
rect 40335 768610 40340 768666
rect 40396 768610 40446 768666
rect 40335 768608 40446 768610
rect 40335 768605 40401 768608
rect 33282 768227 33342 768342
rect 33231 768222 33342 768227
rect 33231 768166 33236 768222
rect 33292 768166 33342 768222
rect 33231 768164 33342 768166
rect 33231 768161 33297 768164
rect 41871 767928 41937 767931
rect 41568 767926 41937 767928
rect 41568 767870 41876 767926
rect 41932 767870 41937 767926
rect 41568 767868 41937 767870
rect 41871 767865 41937 767868
rect 59535 767484 59601 767487
rect 59535 767482 64416 767484
rect 59535 767426 59540 767482
rect 59596 767426 64416 767482
rect 59535 767424 64416 767426
rect 59535 767421 59601 767424
rect 41967 767336 42033 767339
rect 41568 767334 42033 767336
rect 41568 767278 41972 767334
rect 42028 767278 42033 767334
rect 41568 767276 42033 767278
rect 41967 767273 42033 767276
rect 41538 766744 41598 766862
rect 41679 766744 41745 766747
rect 41538 766742 41745 766744
rect 41538 766686 41684 766742
rect 41740 766686 41745 766742
rect 41538 766684 41745 766686
rect 41679 766681 41745 766684
rect 41538 766155 41598 766344
rect 41538 766150 41649 766155
rect 41538 766094 41588 766150
rect 41644 766094 41649 766150
rect 41538 766092 41649 766094
rect 41583 766089 41649 766092
rect 42159 765856 42225 765859
rect 41568 765854 42225 765856
rect 41568 765798 42164 765854
rect 42220 765798 42225 765854
rect 41568 765796 42225 765798
rect 42159 765793 42225 765796
rect 41538 765267 41598 765382
rect 41487 765262 41598 765267
rect 41487 765206 41492 765262
rect 41548 765206 41598 765262
rect 41487 765204 41598 765206
rect 41487 765201 41553 765204
rect 41871 764894 41937 764897
rect 41568 764892 41937 764894
rect 41568 764836 41876 764892
rect 41932 764836 41937 764892
rect 41568 764834 41937 764836
rect 41871 764831 41937 764834
rect 41538 764080 41598 764346
rect 41538 764020 41790 764080
rect 23106 763639 23166 763902
rect 23055 763634 23166 763639
rect 41730 763636 41790 764020
rect 23055 763578 23060 763634
rect 23116 763578 23166 763634
rect 23055 763576 23166 763578
rect 41538 763576 41790 763636
rect 23055 763573 23121 763576
rect 41538 763195 41598 763576
rect 654447 763340 654513 763343
rect 650208 763338 654513 763340
rect 650208 763282 654452 763338
rect 654508 763282 654513 763338
rect 650208 763280 654513 763282
rect 654447 763277 654513 763280
rect 23055 763192 23121 763195
rect 23055 763190 23166 763192
rect 23055 763134 23060 763190
rect 23116 763134 23166 763190
rect 23055 763129 23166 763134
rect 41538 763190 41649 763195
rect 41538 763134 41588 763190
rect 41644 763134 41649 763190
rect 41538 763132 41649 763134
rect 41583 763129 41649 763132
rect 23106 762866 23166 763129
rect 676047 762896 676113 762899
rect 676047 762894 676320 762896
rect 676047 762838 676052 762894
rect 676108 762838 676320 762894
rect 676047 762836 676320 762838
rect 676047 762833 676113 762836
rect 676047 762304 676113 762307
rect 676047 762302 676320 762304
rect 676047 762246 676052 762302
rect 676108 762246 676320 762302
rect 676047 762244 676320 762246
rect 676047 762241 676113 762244
rect 676239 762008 676305 762011
rect 676239 762006 676350 762008
rect 676239 761950 676244 762006
rect 676300 761950 676350 762006
rect 676239 761945 676350 761950
rect 676290 761830 676350 761945
rect 676239 761564 676305 761567
rect 676239 761562 676350 761564
rect 676239 761506 676244 761562
rect 676300 761506 676350 761562
rect 676239 761501 676350 761506
rect 676290 761386 676350 761501
rect 676290 760679 676350 760794
rect 676239 760674 676350 760679
rect 676239 760618 676244 760674
rect 676300 760618 676350 760674
rect 676239 760616 676350 760618
rect 676239 760613 676305 760616
rect 676047 760306 676113 760309
rect 676047 760304 676320 760306
rect 676047 760248 676052 760304
rect 676108 760248 676320 760304
rect 676047 760246 676320 760248
rect 676047 760243 676113 760246
rect 676047 759936 676113 759939
rect 676047 759934 676320 759936
rect 676047 759878 676052 759934
rect 676108 759878 676320 759934
rect 676047 759876 676320 759878
rect 676047 759873 676113 759876
rect 676047 759344 676113 759347
rect 676047 759342 676320 759344
rect 676047 759286 676052 759342
rect 676108 759286 676320 759342
rect 676047 759284 676320 759286
rect 676047 759281 676113 759284
rect 676047 758826 676113 758829
rect 676047 758824 676320 758826
rect 676047 758768 676052 758824
rect 676108 758768 676320 758824
rect 676047 758766 676320 758768
rect 676047 758763 676113 758766
rect 674170 758394 674176 758458
rect 674240 758456 674246 758458
rect 674240 758396 676320 758456
rect 674240 758394 674246 758396
rect 33231 758248 33297 758251
rect 40378 758248 40384 758250
rect 33231 758246 40384 758248
rect 33231 758190 33236 758246
rect 33292 758190 40384 758246
rect 33231 758188 40384 758190
rect 33231 758185 33297 758188
rect 40378 758186 40384 758188
rect 40448 758186 40454 758250
rect 33039 758100 33105 758103
rect 40954 758100 40960 758102
rect 33039 758098 40960 758100
rect 33039 758042 33044 758098
rect 33100 758042 40960 758098
rect 33039 758040 40960 758042
rect 33039 758037 33105 758040
rect 40954 758038 40960 758040
rect 41024 758038 41030 758102
rect 675706 757802 675712 757866
rect 675776 757864 675782 757866
rect 675776 757804 676320 757864
rect 675776 757802 675782 757804
rect 673978 757210 673984 757274
rect 674048 757272 674054 757274
rect 674048 757212 676320 757272
rect 674048 757210 674054 757212
rect 42927 757126 42993 757127
rect 42874 757124 42880 757126
rect 42836 757064 42880 757124
rect 42944 757122 42993 757126
rect 42988 757066 42993 757122
rect 42874 757062 42880 757064
rect 42944 757062 42993 757066
rect 674362 757062 674368 757126
rect 674432 757124 674438 757126
rect 674432 757064 676350 757124
rect 674432 757062 674438 757064
rect 42927 757061 42993 757062
rect 676290 756872 676350 757064
rect 42490 756470 42496 756534
rect 42560 756532 42566 756534
rect 42735 756532 42801 756535
rect 42560 756530 42801 756532
rect 42560 756474 42740 756530
rect 42796 756474 42801 756530
rect 42560 756472 42801 756474
rect 42560 756470 42566 756472
rect 42735 756469 42801 756472
rect 674554 756322 674560 756386
rect 674624 756384 674630 756386
rect 674624 756324 676320 756384
rect 674624 756322 674630 756324
rect 674938 755730 674944 755794
rect 675008 755792 675014 755794
rect 675008 755732 676320 755792
rect 675008 755730 675014 755732
rect 676047 755422 676113 755425
rect 676047 755420 676320 755422
rect 676047 755364 676052 755420
rect 676108 755364 676320 755420
rect 676047 755362 676320 755364
rect 676047 755359 676113 755362
rect 676239 755052 676305 755055
rect 676239 755050 676350 755052
rect 676239 754994 676244 755050
rect 676300 754994 676350 755050
rect 676239 754989 676350 754994
rect 676290 754874 676350 754989
rect 59535 754312 59601 754315
rect 676047 754312 676113 754315
rect 59535 754310 64416 754312
rect 59535 754254 59540 754310
rect 59596 754254 64416 754310
rect 59535 754252 64416 754254
rect 676047 754310 676320 754312
rect 676047 754254 676052 754310
rect 676108 754254 676320 754310
rect 676047 754252 676320 754254
rect 59535 754249 59601 754252
rect 676047 754249 676113 754252
rect 677050 754102 677056 754166
rect 677120 754102 677126 754166
rect 677058 753838 677118 754102
rect 677434 753658 677440 753722
rect 677504 753658 677510 753722
rect 677442 753394 677502 753658
rect 676047 752832 676113 752835
rect 676047 752830 676320 752832
rect 676047 752774 676052 752830
rect 676108 752774 676320 752830
rect 676047 752772 676320 752774
rect 676047 752769 676113 752772
rect 676047 752388 676113 752391
rect 676047 752386 676320 752388
rect 676047 752330 676052 752386
rect 676108 752330 676320 752386
rect 676047 752328 676320 752330
rect 676047 752325 676113 752328
rect 676047 751870 676113 751873
rect 676047 751868 676320 751870
rect 676047 751812 676052 751868
rect 676108 751812 676320 751868
rect 676047 751810 676320 751812
rect 676047 751807 676113 751810
rect 679791 751500 679857 751503
rect 679746 751498 679857 751500
rect 679746 751442 679796 751498
rect 679852 751442 679857 751498
rect 679746 751437 679857 751442
rect 679746 751322 679806 751437
rect 42063 751056 42129 751059
rect 42490 751056 42496 751058
rect 42063 751054 42496 751056
rect 42063 750998 42068 751054
rect 42124 750998 42496 751054
rect 42063 750996 42496 750998
rect 42063 750993 42129 750996
rect 42490 750994 42496 750996
rect 42560 750994 42566 751058
rect 685506 750615 685566 750878
rect 679791 750612 679857 750615
rect 679746 750610 679857 750612
rect 679746 750554 679796 750610
rect 679852 750554 679857 750610
rect 679746 750549 679857 750554
rect 685455 750610 685566 750615
rect 685455 750554 685460 750610
rect 685516 750554 685566 750610
rect 685455 750552 685566 750554
rect 685455 750549 685521 750552
rect 679746 750360 679806 750549
rect 654447 750168 654513 750171
rect 650208 750166 654513 750168
rect 650208 750110 654452 750166
rect 654508 750110 654513 750166
rect 650208 750108 654513 750110
rect 654447 750105 654513 750108
rect 685455 750168 685521 750171
rect 685455 750166 685566 750168
rect 685455 750110 685460 750166
rect 685516 750110 685566 750166
rect 685455 750105 685566 750110
rect 42874 749810 42880 749874
rect 42944 749872 42950 749874
rect 43023 749872 43089 749875
rect 42944 749870 43089 749872
rect 42944 749814 43028 749870
rect 43084 749814 43089 749870
rect 685506 749842 685566 750105
rect 42944 749812 43089 749814
rect 42944 749810 42950 749812
rect 43023 749809 43089 749812
rect 40378 748626 40384 748690
rect 40448 748688 40454 748690
rect 42639 748688 42705 748691
rect 40448 748686 42705 748688
rect 40448 748630 42644 748686
rect 42700 748630 42705 748686
rect 40448 748628 42705 748630
rect 40448 748626 40454 748628
rect 42639 748625 42705 748628
rect 40954 748478 40960 748542
rect 41024 748540 41030 748542
rect 42735 748540 42801 748543
rect 41024 748538 42801 748540
rect 41024 748482 42740 748538
rect 42796 748482 42801 748538
rect 41024 748480 42801 748482
rect 41024 748478 41030 748480
rect 42735 748477 42801 748480
rect 674362 743150 674368 743214
rect 674432 743212 674438 743214
rect 675375 743212 675441 743215
rect 674432 743210 675441 743212
rect 674432 743154 675380 743210
rect 675436 743154 675441 743210
rect 674432 743152 675441 743154
rect 674432 743150 674438 743152
rect 675375 743149 675441 743152
rect 675759 742176 675825 742179
rect 676090 742176 676096 742178
rect 675759 742174 676096 742176
rect 675759 742118 675764 742174
rect 675820 742118 676096 742174
rect 675759 742116 676096 742118
rect 675759 742113 675825 742116
rect 676090 742114 676096 742116
rect 676160 742114 676166 742178
rect 674554 741670 674560 741734
rect 674624 741732 674630 741734
rect 675375 741732 675441 741735
rect 674624 741730 675441 741732
rect 674624 741674 675380 741730
rect 675436 741674 675441 741730
rect 674624 741672 675441 741674
rect 674624 741670 674630 741672
rect 675375 741669 675441 741672
rect 58575 741288 58641 741291
rect 58575 741286 64416 741288
rect 58575 741230 58580 741286
rect 58636 741230 64416 741286
rect 58575 741228 64416 741230
rect 58575 741225 58641 741228
rect 674938 740338 674944 740402
rect 675008 740400 675014 740402
rect 675471 740400 675537 740403
rect 675008 740398 675537 740400
rect 675008 740342 675476 740398
rect 675532 740342 675537 740398
rect 675008 740340 675537 740342
rect 675008 740338 675014 740340
rect 675471 740337 675537 740340
rect 654447 736848 654513 736851
rect 650208 736846 654513 736848
rect 650208 736790 654452 736846
rect 654508 736790 654513 736846
rect 650208 736788 654513 736790
rect 654447 736785 654513 736788
rect 675663 735518 675729 735519
rect 675663 735514 675712 735518
rect 675776 735516 675782 735518
rect 675663 735458 675668 735514
rect 675663 735454 675712 735458
rect 675776 735456 675820 735516
rect 675776 735454 675782 735456
rect 675663 735453 675729 735454
rect 675759 734480 675825 734483
rect 677050 734480 677056 734482
rect 675759 734478 677056 734480
rect 675759 734422 675764 734478
rect 675820 734422 677056 734478
rect 675759 734420 677056 734422
rect 675759 734417 675825 734420
rect 677050 734418 677056 734420
rect 677120 734418 677126 734482
rect 41583 732852 41649 732855
rect 41538 732850 41649 732852
rect 41538 732794 41588 732850
rect 41644 732794 41649 732850
rect 41538 732789 41649 732794
rect 41538 732674 41598 732789
rect 41775 732112 41841 732115
rect 41568 732110 41841 732112
rect 41568 732054 41780 732110
rect 41836 732054 41841 732110
rect 41568 732052 41841 732054
rect 41775 732049 41841 732052
rect 41583 731816 41649 731819
rect 41538 731814 41649 731816
rect 41538 731758 41588 731814
rect 41644 731758 41649 731814
rect 41538 731753 41649 731758
rect 41538 731638 41598 731753
rect 41583 731372 41649 731375
rect 41538 731370 41649 731372
rect 41538 731314 41588 731370
rect 41644 731314 41649 731370
rect 41538 731309 41649 731314
rect 41538 731194 41598 731309
rect 41538 730487 41598 730602
rect 41538 730482 41649 730487
rect 41538 730426 41588 730482
rect 41644 730426 41649 730482
rect 41538 730424 41649 730426
rect 41583 730421 41649 730424
rect 42063 730114 42129 730117
rect 40992 730112 42129 730114
rect 40992 730084 42068 730112
rect 40962 730056 42068 730084
rect 42124 730056 42129 730112
rect 40962 730054 42129 730056
rect 40962 729894 41022 730054
rect 42063 730051 42129 730054
rect 40762 729830 40768 729894
rect 40832 729830 40838 729894
rect 40954 729830 40960 729894
rect 41024 729830 41030 729894
rect 40770 729714 40830 729830
rect 41679 729448 41745 729451
rect 41346 729446 41745 729448
rect 41346 729390 41684 729446
rect 41740 729390 41745 729446
rect 41346 729388 41745 729390
rect 41346 729152 41406 729388
rect 41679 729385 41745 729388
rect 40416 729122 41406 729152
rect 40386 729092 41376 729122
rect 40386 728858 40446 729092
rect 40570 728942 40576 729006
rect 40640 728942 40646 729006
rect 40378 728794 40384 728858
rect 40448 728794 40454 728858
rect 40578 728530 40638 728942
rect 59151 728264 59217 728267
rect 59151 728262 64416 728264
rect 41538 727968 41598 728234
rect 59151 728206 59156 728262
rect 59212 728206 64416 728262
rect 59151 728204 64416 728206
rect 59151 728201 59217 728204
rect 41679 727968 41745 727971
rect 41538 727966 41745 727968
rect 41538 727910 41684 727966
rect 41740 727910 41745 727966
rect 41538 727908 41745 727910
rect 41679 727905 41745 727908
rect 41967 727672 42033 727675
rect 41568 727670 42033 727672
rect 41568 727614 41972 727670
rect 42028 727614 42033 727670
rect 41568 727612 42033 727614
rect 41967 727609 42033 727612
rect 34434 726935 34494 727050
rect 34383 726930 34494 726935
rect 34383 726874 34388 726930
rect 34444 726874 34494 726930
rect 34383 726872 34494 726874
rect 34383 726869 34449 726872
rect 41538 726491 41598 726680
rect 41487 726486 41598 726491
rect 41487 726430 41492 726486
rect 41548 726430 41598 726486
rect 41487 726428 41598 726430
rect 41487 726425 41553 726428
rect 42063 726192 42129 726195
rect 41568 726190 42129 726192
rect 41568 726134 42068 726190
rect 42124 726134 42129 726190
rect 41568 726132 42129 726134
rect 42063 726129 42129 726132
rect 41871 725600 41937 725603
rect 41568 725598 41937 725600
rect 41568 725542 41876 725598
rect 41932 725542 41937 725598
rect 41568 725540 41937 725542
rect 41871 725537 41937 725540
rect 34434 725011 34494 725200
rect 34434 725006 34545 725011
rect 34434 724950 34484 725006
rect 34540 724950 34545 725006
rect 34434 724948 34545 724950
rect 34479 724945 34545 724948
rect 42159 724712 42225 724715
rect 41568 724710 42225 724712
rect 41568 724654 42164 724710
rect 42220 724654 42225 724710
rect 41568 724652 42225 724654
rect 42159 724649 42225 724652
rect 41538 723975 41598 724090
rect 41538 723970 41649 723975
rect 41538 723914 41588 723970
rect 41644 723914 41649 723970
rect 41538 723912 41649 723914
rect 41583 723909 41649 723912
rect 41775 723676 41841 723679
rect 41568 723674 41841 723676
rect 41568 723618 41780 723674
rect 41836 723618 41841 723674
rect 41568 723616 41841 723618
rect 41775 723613 41841 723616
rect 655215 723528 655281 723531
rect 650208 723526 655281 723528
rect 650208 723470 655220 723526
rect 655276 723470 655281 723526
rect 650208 723468 655281 723470
rect 655215 723465 655281 723468
rect 41775 723232 41841 723235
rect 41568 723230 41841 723232
rect 41568 723174 41780 723230
rect 41836 723174 41841 723230
rect 41568 723172 41841 723174
rect 41775 723169 41841 723172
rect 41722 722640 41728 722642
rect 41568 722580 41728 722640
rect 41722 722578 41728 722580
rect 41792 722578 41798 722642
rect 41538 722051 41598 722166
rect 41538 722046 41649 722051
rect 41538 721990 41588 722046
rect 41644 721990 41649 722046
rect 41538 721988 41649 721990
rect 41583 721985 41649 721988
rect 41538 721604 41598 721648
rect 42447 721604 42513 721607
rect 41538 721602 42513 721604
rect 41538 721546 42452 721602
rect 42508 721546 42513 721602
rect 41538 721544 42513 721546
rect 42447 721541 42513 721544
rect 41775 721160 41841 721163
rect 41568 721158 41841 721160
rect 41568 721102 41780 721158
rect 41836 721102 41841 721158
rect 41568 721100 41841 721102
rect 41775 721097 41841 721100
rect 23106 720423 23166 720686
rect 23055 720418 23166 720423
rect 23055 720362 23060 720418
rect 23116 720362 23166 720418
rect 23055 720360 23166 720362
rect 23055 720357 23121 720360
rect 41775 720198 41841 720201
rect 41568 720196 41841 720198
rect 41568 720140 41780 720196
rect 41836 720140 41841 720196
rect 41568 720138 41841 720140
rect 41775 720135 41841 720138
rect 23055 719828 23121 719831
rect 23055 719826 23166 719828
rect 23055 719770 23060 719826
rect 23116 719770 23166 719826
rect 23055 719765 23166 719770
rect 23106 719650 23166 719765
rect 676239 718052 676305 718055
rect 676239 718050 676350 718052
rect 676239 717994 676244 718050
rect 676300 717994 676350 718050
rect 676239 717989 676350 717994
rect 676290 717874 676350 717989
rect 676047 717312 676113 717315
rect 676047 717310 676320 717312
rect 676047 717254 676052 717310
rect 676108 717254 676320 717310
rect 676047 717252 676320 717254
rect 676047 717249 676113 717252
rect 34383 717016 34449 717019
rect 40762 717016 40768 717018
rect 34383 717014 40768 717016
rect 34383 716958 34388 717014
rect 34444 716958 40768 717014
rect 34383 716956 40768 716958
rect 34383 716953 34449 716956
rect 40762 716954 40768 716956
rect 40832 716954 40838 717018
rect 676239 717016 676305 717019
rect 676239 717014 676350 717016
rect 676239 716958 676244 717014
rect 676300 716958 676350 717014
rect 676239 716953 676350 716958
rect 676290 716838 676350 716953
rect 34479 716572 34545 716575
rect 40378 716572 40384 716574
rect 34479 716570 40384 716572
rect 34479 716514 34484 716570
rect 34540 716514 40384 716570
rect 34479 716512 40384 716514
rect 34479 716509 34545 716512
rect 40378 716510 40384 716512
rect 40448 716510 40454 716574
rect 679695 716572 679761 716575
rect 679695 716570 679806 716572
rect 679695 716514 679700 716570
rect 679756 716514 679806 716570
rect 679695 716509 679806 716514
rect 679746 716394 679806 716509
rect 679746 715539 679806 715802
rect 679695 715534 679806 715539
rect 679695 715478 679700 715534
rect 679756 715478 679806 715534
rect 679695 715476 679806 715478
rect 679695 715473 679761 715476
rect 59535 715388 59601 715391
rect 59535 715386 64416 715388
rect 59535 715330 59540 715386
rect 59596 715330 64416 715386
rect 59535 715328 64416 715330
rect 59535 715325 59601 715328
rect 676047 715314 676113 715317
rect 676047 715312 676320 715314
rect 676047 715256 676052 715312
rect 676108 715256 676320 715312
rect 676047 715254 676320 715256
rect 676047 715251 676113 715254
rect 676047 714944 676113 714947
rect 676047 714942 676320 714944
rect 676047 714886 676052 714942
rect 676108 714886 676320 714942
rect 676047 714884 676320 714886
rect 676047 714881 676113 714884
rect 676047 714352 676113 714355
rect 676047 714350 676320 714352
rect 676047 714294 676052 714350
rect 676108 714294 676320 714350
rect 676047 714292 676320 714294
rect 676047 714289 676113 714292
rect 41775 714056 41841 714059
rect 43066 714056 43072 714058
rect 41775 714054 43072 714056
rect 41775 713998 41780 714054
rect 41836 713998 43072 714054
rect 41775 713996 43072 713998
rect 41775 713993 41841 713996
rect 43066 713994 43072 713996
rect 43136 713994 43142 714058
rect 41967 713910 42033 713911
rect 41914 713846 41920 713910
rect 41984 713908 42033 713910
rect 42159 713908 42225 713911
rect 42874 713908 42880 713910
rect 41984 713906 42076 713908
rect 42028 713850 42076 713906
rect 41984 713848 42076 713850
rect 42159 713906 42880 713908
rect 42159 713850 42164 713906
rect 42220 713850 42880 713906
rect 42159 713848 42880 713850
rect 41984 713846 42033 713848
rect 41967 713845 42033 713846
rect 42159 713845 42225 713848
rect 42874 713846 42880 713848
rect 42944 713846 42950 713910
rect 676047 713760 676113 713763
rect 676047 713758 676320 713760
rect 676047 713702 676052 713758
rect 676108 713702 676320 713758
rect 676047 713700 676320 713702
rect 676047 713697 676113 713700
rect 675130 713402 675136 713466
rect 675200 713464 675206 713466
rect 675200 713404 676320 713464
rect 675200 713402 675206 713404
rect 675898 712810 675904 712874
rect 675968 712872 675974 712874
rect 675968 712812 676320 712872
rect 675968 712810 675974 712812
rect 675322 712218 675328 712282
rect 675392 712280 675398 712282
rect 675392 712220 676320 712280
rect 675392 712218 675398 712220
rect 675514 712070 675520 712134
rect 675584 712132 675590 712134
rect 675584 712072 676350 712132
rect 675584 712070 675590 712072
rect 676290 711880 676350 712072
rect 41914 711626 41920 711690
rect 41984 711688 41990 711690
rect 42063 711688 42129 711691
rect 41984 711686 42129 711688
rect 41984 711630 42068 711686
rect 42124 711630 42129 711686
rect 41984 711628 42129 711630
rect 41984 711626 41990 711628
rect 42063 711625 42129 711628
rect 676282 711626 676288 711690
rect 676352 711626 676358 711690
rect 676290 711362 676350 711626
rect 674746 710738 674752 710802
rect 674816 710800 674822 710802
rect 674816 710740 676320 710800
rect 674816 710738 674822 710740
rect 676047 710430 676113 710433
rect 676047 710428 676320 710430
rect 676047 710372 676052 710428
rect 676108 710372 676320 710428
rect 676047 710370 676320 710372
rect 676047 710367 676113 710370
rect 654447 710356 654513 710359
rect 650208 710354 654513 710356
rect 650208 710298 654452 710354
rect 654508 710298 654513 710354
rect 650208 710296 654513 710298
rect 654447 710293 654513 710296
rect 676239 710060 676305 710063
rect 676239 710058 676350 710060
rect 676239 710002 676244 710058
rect 676300 710002 676350 710058
rect 676239 709997 676350 710002
rect 676290 709882 676350 709997
rect 42927 709766 42993 709767
rect 42874 709702 42880 709766
rect 42944 709764 42993 709766
rect 42944 709762 43036 709764
rect 42988 709706 43036 709762
rect 42944 709704 43036 709706
rect 42944 709702 42993 709704
rect 42927 709701 42993 709702
rect 676047 709320 676113 709323
rect 676047 709318 676320 709320
rect 676047 709262 676052 709318
rect 676108 709262 676320 709318
rect 676047 709260 676320 709262
rect 676047 709257 676113 709260
rect 677242 709110 677248 709174
rect 677312 709110 677318 709174
rect 677250 708846 677310 709110
rect 676858 708518 676864 708582
rect 676928 708518 676934 708582
rect 676866 708402 676926 708518
rect 676239 707988 676305 707991
rect 676239 707986 676350 707988
rect 676239 707930 676244 707986
rect 676300 707930 676350 707986
rect 676239 707925 676350 707930
rect 676290 707810 676350 707925
rect 676047 707396 676113 707399
rect 676047 707394 676320 707396
rect 676047 707338 676052 707394
rect 676108 707338 676320 707394
rect 676047 707336 676320 707338
rect 676047 707333 676113 707336
rect 43119 707250 43185 707251
rect 43066 707186 43072 707250
rect 43136 707248 43185 707250
rect 43136 707246 43228 707248
rect 43180 707190 43228 707246
rect 43136 707188 43228 707190
rect 43136 707186 43185 707188
rect 43119 707185 43185 707186
rect 676047 706878 676113 706881
rect 676047 706876 676320 706878
rect 676047 706820 676052 706876
rect 676108 706820 676320 706876
rect 676047 706818 676320 706820
rect 676047 706815 676113 706818
rect 679983 706508 680049 706511
rect 679938 706506 680049 706508
rect 679938 706450 679988 706506
rect 680044 706450 680049 706506
rect 679938 706445 680049 706450
rect 679938 706330 679998 706445
rect 41722 706002 41728 706066
rect 41792 706064 41798 706066
rect 42447 706064 42513 706067
rect 41792 706062 42513 706064
rect 41792 706006 42452 706062
rect 42508 706006 42513 706062
rect 41792 706004 42513 706006
rect 41792 706002 41798 706004
rect 42447 706001 42513 706004
rect 679746 705623 679806 705886
rect 679746 705618 679857 705623
rect 679983 705620 680049 705623
rect 679746 705562 679796 705618
rect 679852 705562 679857 705618
rect 679746 705560 679857 705562
rect 679791 705557 679857 705560
rect 679938 705618 680049 705620
rect 679938 705562 679988 705618
rect 680044 705562 680049 705618
rect 679938 705557 680049 705562
rect 679938 705368 679998 705557
rect 679791 705176 679857 705179
rect 679746 705174 679857 705176
rect 679746 705118 679796 705174
rect 679852 705118 679857 705174
rect 679746 705113 679857 705118
rect 679746 704850 679806 705113
rect 40762 703634 40768 703698
rect 40832 703696 40838 703698
rect 42447 703696 42513 703699
rect 40832 703694 42513 703696
rect 40832 703638 42452 703694
rect 42508 703638 42513 703694
rect 40832 703636 42513 703638
rect 40832 703634 40838 703636
rect 42447 703633 42513 703636
rect 40378 703338 40384 703402
rect 40448 703400 40454 703402
rect 42831 703400 42897 703403
rect 40448 703398 42897 703400
rect 40448 703342 42836 703398
rect 42892 703342 42897 703398
rect 40448 703340 42897 703342
rect 40448 703338 40454 703340
rect 42831 703337 42897 703340
rect 59535 702216 59601 702219
rect 59535 702214 64416 702216
rect 59535 702158 59540 702214
rect 59596 702158 64416 702214
rect 59535 702156 64416 702158
rect 59535 702153 59601 702156
rect 675375 697926 675441 697927
rect 675322 697924 675328 697926
rect 675284 697864 675328 697924
rect 675392 697922 675441 697926
rect 675436 697866 675441 697922
rect 675322 697862 675328 697864
rect 675392 697862 675441 697866
rect 675375 697861 675441 697862
rect 675759 697332 675825 697335
rect 676282 697332 676288 697334
rect 675759 697330 676288 697332
rect 675759 697274 675764 697330
rect 675820 697274 676288 697330
rect 675759 697272 676288 697274
rect 675759 697269 675825 697272
rect 676282 697270 676288 697272
rect 676352 697270 676358 697334
rect 654447 697036 654513 697039
rect 650208 697034 654513 697036
rect 650208 696978 654452 697034
rect 654508 696978 654513 697034
rect 650208 696976 654513 696978
rect 654447 696973 654513 696976
rect 675567 696890 675633 696891
rect 675514 696888 675520 696890
rect 675476 696828 675520 696888
rect 675584 696886 675633 696890
rect 675628 696830 675633 696886
rect 675514 696826 675520 696828
rect 675584 696826 675633 696830
rect 675567 696825 675633 696826
rect 675130 694754 675136 694818
rect 675200 694816 675206 694818
rect 675375 694816 675441 694819
rect 675200 694814 675441 694816
rect 675200 694758 675380 694814
rect 675436 694758 675441 694814
rect 675200 694756 675441 694758
rect 675200 694754 675206 694756
rect 675375 694753 675441 694756
rect 675759 694224 675825 694227
rect 676474 694224 676480 694226
rect 675759 694222 676480 694224
rect 675759 694166 675764 694222
rect 675820 694166 676480 694222
rect 675759 694164 676480 694166
rect 675759 694161 675825 694164
rect 676474 694162 676480 694164
rect 676544 694162 676550 694226
rect 673978 690462 673984 690526
rect 674048 690524 674054 690526
rect 675471 690524 675537 690527
rect 674048 690522 675537 690524
rect 674048 690466 675476 690522
rect 675532 690466 675537 690522
rect 674048 690464 675537 690466
rect 674048 690462 674054 690464
rect 675471 690461 675537 690464
rect 41775 689488 41841 689491
rect 41568 689486 41841 689488
rect 41568 689430 41780 689486
rect 41836 689430 41841 689486
rect 41568 689428 41841 689430
rect 41775 689425 41841 689428
rect 59535 689192 59601 689195
rect 59535 689190 64416 689192
rect 59535 689134 59540 689190
rect 59596 689134 64416 689190
rect 59535 689132 64416 689134
rect 59535 689129 59601 689132
rect 41775 688896 41841 688899
rect 41568 688894 41841 688896
rect 41568 688838 41780 688894
rect 41836 688838 41841 688894
rect 41568 688836 41841 688838
rect 41775 688833 41841 688836
rect 41583 688600 41649 688603
rect 41538 688598 41649 688600
rect 41538 688542 41588 688598
rect 41644 688542 41649 688598
rect 41538 688537 41649 688542
rect 41538 688422 41598 688537
rect 41583 688156 41649 688159
rect 41538 688154 41649 688156
rect 41538 688098 41588 688154
rect 41644 688098 41649 688154
rect 41538 688093 41649 688098
rect 41538 687978 41598 688093
rect 675759 687416 675825 687419
rect 676858 687416 676864 687418
rect 675759 687414 676864 687416
rect 41538 687271 41598 687386
rect 675759 687358 675764 687414
rect 675820 687358 676864 687414
rect 675759 687356 676864 687358
rect 675759 687353 675825 687356
rect 676858 687354 676864 687356
rect 676928 687354 676934 687418
rect 41538 687266 41649 687271
rect 41538 687210 41588 687266
rect 41644 687210 41649 687266
rect 41538 687208 41649 687210
rect 41583 687205 41649 687208
rect 41871 686972 41937 686975
rect 41568 686970 41937 686972
rect 41568 686942 41876 686970
rect 41538 686914 41876 686942
rect 41932 686914 41937 686970
rect 41538 686912 41937 686914
rect 40762 686614 40768 686678
rect 40832 686614 40838 686678
rect 40954 686614 40960 686678
rect 41024 686676 41030 686678
rect 41538 686676 41598 686912
rect 41871 686909 41937 686912
rect 41024 686616 41598 686676
rect 41024 686614 41030 686616
rect 40770 686498 40830 686614
rect 41775 685936 41841 685939
rect 41184 685934 41841 685936
rect 41184 685906 41780 685934
rect 41154 685878 41780 685906
rect 41836 685878 41841 685934
rect 41154 685876 41841 685878
rect 41154 685790 41214 685876
rect 41775 685873 41841 685876
rect 41146 685726 41152 685790
rect 41216 685726 41222 685790
rect 40570 685578 40576 685642
rect 40640 685578 40646 685642
rect 40578 685492 40638 685578
rect 34434 685432 40638 685492
rect 34434 685388 34494 685432
rect 41775 685048 41841 685051
rect 41568 685046 41841 685048
rect 41568 684990 41780 685046
rect 41836 684990 41841 685046
rect 41568 684988 41841 684990
rect 41775 684985 41841 684988
rect 41538 684311 41598 684426
rect 41538 684306 41649 684311
rect 41538 684250 41588 684306
rect 41644 684250 41649 684306
rect 41538 684248 41649 684250
rect 41583 684245 41649 684248
rect 34434 683719 34494 683834
rect 34383 683714 34494 683719
rect 34383 683658 34388 683714
rect 34444 683658 34494 683714
rect 34383 683656 34494 683658
rect 34383 683653 34449 683656
rect 654447 683568 654513 683571
rect 650208 683566 654513 683568
rect 41538 683272 41598 683538
rect 650208 683510 654452 683566
rect 654508 683510 654513 683566
rect 650208 683508 654513 683510
rect 654447 683505 654513 683508
rect 41679 683272 41745 683275
rect 41538 683270 41745 683272
rect 41538 683214 41684 683270
rect 41740 683214 41745 683270
rect 41538 683212 41745 683214
rect 41679 683209 41745 683212
rect 42447 682976 42513 682979
rect 41568 682974 42513 682976
rect 41568 682918 42452 682974
rect 42508 682918 42513 682974
rect 41568 682916 42513 682918
rect 42447 682913 42513 682916
rect 41871 682384 41937 682387
rect 41568 682382 41937 682384
rect 41568 682326 41876 682382
rect 41932 682326 41937 682382
rect 41568 682324 41937 682326
rect 41871 682321 41937 682324
rect 34434 681795 34494 681984
rect 34434 681790 34545 681795
rect 34434 681734 34484 681790
rect 34540 681734 34545 681790
rect 34434 681732 34545 681734
rect 34479 681729 34545 681732
rect 42159 681496 42225 681499
rect 41568 681494 42225 681496
rect 41568 681438 42164 681494
rect 42220 681438 42225 681494
rect 41568 681436 42225 681438
rect 42159 681433 42225 681436
rect 42063 680904 42129 680907
rect 41568 680902 42129 680904
rect 41568 680846 42068 680902
rect 42124 680846 42129 680902
rect 41568 680844 42129 680846
rect 42063 680841 42129 680844
rect 41538 680315 41598 680504
rect 41538 680310 41649 680315
rect 41538 680254 41588 680310
rect 41644 680254 41649 680310
rect 41538 680252 41649 680254
rect 41583 680249 41649 680252
rect 41967 680016 42033 680019
rect 41568 680014 42033 680016
rect 41568 679958 41972 680014
rect 42028 679958 42033 680014
rect 41568 679956 42033 679958
rect 41967 679953 42033 679956
rect 41538 679279 41598 679394
rect 41538 679274 41649 679279
rect 41538 679218 41588 679274
rect 41644 679218 41649 679274
rect 41538 679216 41649 679218
rect 41583 679213 41649 679216
rect 41538 678835 41598 678950
rect 41538 678830 41649 678835
rect 41538 678774 41588 678830
rect 41644 678774 41649 678830
rect 41538 678772 41649 678774
rect 41583 678769 41649 678772
rect 41775 678536 41841 678539
rect 41568 678534 41841 678536
rect 41568 678478 41780 678534
rect 41836 678478 41841 678534
rect 41568 678476 41841 678478
rect 41775 678473 41841 678476
rect 41775 677944 41841 677947
rect 41568 677942 41841 677944
rect 41568 677886 41780 677942
rect 41836 677886 41841 677942
rect 41568 677884 41841 677886
rect 41775 677881 41841 677884
rect 23106 677207 23166 677470
rect 23055 677202 23166 677207
rect 23055 677146 23060 677202
rect 23116 677146 23166 677202
rect 23055 677144 23166 677146
rect 23055 677141 23121 677144
rect 41775 676982 41841 676985
rect 41568 676980 41841 676982
rect 41568 676924 41780 676980
rect 41836 676924 41841 676980
rect 41568 676922 41841 676924
rect 41775 676919 41841 676922
rect 23055 676760 23121 676763
rect 23055 676758 23166 676760
rect 23055 676702 23060 676758
rect 23116 676702 23166 676758
rect 23055 676697 23166 676702
rect 23106 676434 23166 676697
rect 59055 676168 59121 676171
rect 59055 676166 64416 676168
rect 59055 676110 59060 676166
rect 59116 676110 64416 676166
rect 59055 676108 64416 676110
rect 59055 676105 59121 676108
rect 676047 672690 676113 672693
rect 676047 672688 676320 672690
rect 676047 672632 676052 672688
rect 676108 672632 676320 672688
rect 676047 672630 676320 672632
rect 676047 672627 676113 672630
rect 34383 672616 34449 672619
rect 40570 672616 40576 672618
rect 34383 672614 40576 672616
rect 34383 672558 34388 672614
rect 34444 672558 40576 672614
rect 34383 672556 40576 672558
rect 34383 672553 34449 672556
rect 40570 672554 40576 672556
rect 40640 672554 40646 672618
rect 34479 672468 34545 672471
rect 40378 672468 40384 672470
rect 34479 672466 40384 672468
rect 34479 672410 34484 672466
rect 34540 672410 40384 672466
rect 34479 672408 40384 672410
rect 34479 672405 34545 672408
rect 40378 672406 40384 672408
rect 40448 672406 40454 672470
rect 676239 672320 676305 672323
rect 676239 672318 676350 672320
rect 676239 672262 676244 672318
rect 676300 672262 676350 672318
rect 676239 672257 676350 672262
rect 676290 672142 676350 672257
rect 676047 671580 676113 671583
rect 676047 671578 676320 671580
rect 676047 671522 676052 671578
rect 676108 671522 676320 671578
rect 676047 671520 676320 671522
rect 676047 671517 676113 671520
rect 676047 671210 676113 671213
rect 676047 671208 676320 671210
rect 676047 671152 676052 671208
rect 676108 671152 676320 671208
rect 676047 671150 676320 671152
rect 676047 671147 676113 671150
rect 41775 670694 41841 670695
rect 41722 670692 41728 670694
rect 41684 670632 41728 670692
rect 41792 670690 41841 670694
rect 41836 670634 41841 670690
rect 41722 670630 41728 670632
rect 41792 670630 41841 670634
rect 41775 670629 41841 670630
rect 42063 670692 42129 670695
rect 42490 670692 42496 670694
rect 42063 670690 42496 670692
rect 42063 670634 42068 670690
rect 42124 670634 42496 670690
rect 42063 670632 42496 670634
rect 42063 670629 42129 670632
rect 42490 670630 42496 670632
rect 42560 670630 42566 670694
rect 676047 670692 676113 670695
rect 676047 670690 676320 670692
rect 676047 670634 676052 670690
rect 676108 670634 676320 670690
rect 676047 670632 676320 670634
rect 676047 670629 676113 670632
rect 655503 670396 655569 670399
rect 650208 670394 655569 670396
rect 650208 670338 655508 670394
rect 655564 670338 655569 670394
rect 650208 670336 655569 670338
rect 655503 670333 655569 670336
rect 42298 670038 42304 670102
rect 42368 670100 42374 670102
rect 42447 670100 42513 670103
rect 42368 670098 42513 670100
rect 42368 670042 42452 670098
rect 42508 670042 42513 670098
rect 42368 670040 42513 670042
rect 42368 670038 42374 670040
rect 42447 670037 42513 670040
rect 676047 670100 676113 670103
rect 676047 670098 676320 670100
rect 676047 670042 676052 670098
rect 676108 670042 676320 670098
rect 676047 670040 676320 670042
rect 676047 670037 676113 670040
rect 676047 669656 676113 669659
rect 676047 669654 676320 669656
rect 676047 669598 676052 669654
rect 676108 669598 676320 669654
rect 676047 669596 676320 669598
rect 676047 669593 676113 669596
rect 676239 669360 676305 669363
rect 676239 669358 676350 669360
rect 676239 669302 676244 669358
rect 676300 669302 676350 669358
rect 676239 669297 676350 669302
rect 676290 669182 676350 669297
rect 679887 668916 679953 668919
rect 679887 668914 679998 668916
rect 679887 668858 679892 668914
rect 679948 668858 679998 668914
rect 679887 668853 679998 668858
rect 679938 668590 679998 668853
rect 674554 668114 674560 668178
rect 674624 668176 674630 668178
rect 674624 668116 676320 668176
rect 674624 668114 674630 668116
rect 676047 667658 676113 667661
rect 676047 667656 676320 667658
rect 676047 667600 676052 667656
rect 676108 667600 676320 667656
rect 676047 667598 676320 667600
rect 676047 667595 676113 667598
rect 674362 667078 674368 667142
rect 674432 667140 674438 667142
rect 674432 667080 676320 667140
rect 674432 667078 674438 667080
rect 42159 666696 42225 666699
rect 42298 666696 42304 666698
rect 42159 666694 42304 666696
rect 42159 666638 42164 666694
rect 42220 666638 42304 666694
rect 42159 666636 42304 666638
rect 42159 666633 42225 666636
rect 42298 666634 42304 666636
rect 42368 666634 42374 666698
rect 674938 666634 674944 666698
rect 675008 666696 675014 666698
rect 675008 666636 676320 666696
rect 675008 666634 675014 666636
rect 675706 666116 675712 666180
rect 675776 666178 675782 666180
rect 675776 666118 676320 666178
rect 675776 666116 675782 666118
rect 676239 665808 676305 665811
rect 676239 665806 676350 665808
rect 676239 665750 676244 665806
rect 676300 665750 676350 665806
rect 676239 665745 676350 665750
rect 676290 665630 676350 665745
rect 42490 665154 42496 665218
rect 42560 665216 42566 665218
rect 42831 665216 42897 665219
rect 42560 665214 42897 665216
rect 42560 665158 42836 665214
rect 42892 665158 42897 665214
rect 42560 665156 42897 665158
rect 42560 665154 42566 665156
rect 42831 665153 42897 665156
rect 676090 665006 676096 665070
rect 676160 665068 676166 665070
rect 676290 665068 676350 665186
rect 676160 665008 676350 665068
rect 676160 665006 676166 665008
rect 676047 664624 676113 664627
rect 676047 664622 676320 664624
rect 676047 664566 676052 664622
rect 676108 664566 676320 664622
rect 676047 664564 676320 664566
rect 676047 664561 676113 664564
rect 676239 664328 676305 664331
rect 676239 664326 676350 664328
rect 676239 664270 676244 664326
rect 676300 664270 676350 664326
rect 676239 664265 676350 664270
rect 676290 664150 676350 664265
rect 676239 663884 676305 663887
rect 676239 663882 676350 663884
rect 676239 663826 676244 663882
rect 676300 663826 676350 663882
rect 676239 663821 676350 663826
rect 676290 663706 676350 663821
rect 41775 663442 41841 663443
rect 41722 663378 41728 663442
rect 41792 663440 41841 663442
rect 41792 663438 41884 663440
rect 41836 663382 41884 663438
rect 41792 663380 41884 663382
rect 41792 663378 41841 663380
rect 677050 663378 677056 663442
rect 677120 663378 677126 663442
rect 41775 663377 41841 663378
rect 58095 663144 58161 663147
rect 58095 663142 64416 663144
rect 58095 663086 58100 663142
rect 58156 663086 64416 663142
rect 677058 663114 677118 663378
rect 58095 663084 64416 663086
rect 58095 663081 58161 663084
rect 676047 662626 676113 662629
rect 676047 662624 676320 662626
rect 676047 662568 676052 662624
rect 676108 662568 676320 662624
rect 676047 662566 676320 662568
rect 676047 662563 676113 662566
rect 676047 662256 676113 662259
rect 676047 662254 676320 662256
rect 676047 662198 676052 662254
rect 676108 662198 676320 662254
rect 676047 662196 676320 662198
rect 676047 662193 676113 662196
rect 676047 661664 676113 661667
rect 676047 661662 676320 661664
rect 676047 661606 676052 661662
rect 676108 661606 676320 661662
rect 676047 661604 676320 661606
rect 676047 661601 676113 661604
rect 679746 660927 679806 661116
rect 40570 660862 40576 660926
rect 40640 660924 40646 660926
rect 43023 660924 43089 660927
rect 40640 660922 43089 660924
rect 40640 660866 43028 660922
rect 43084 660866 43089 660922
rect 40640 660864 43089 660866
rect 679746 660922 679857 660927
rect 679746 660866 679796 660922
rect 679852 660866 679857 660922
rect 679746 660864 679857 660866
rect 40640 660862 40646 660864
rect 43023 660861 43089 660864
rect 679791 660861 679857 660864
rect 685506 660483 685566 660746
rect 679791 660480 679857 660483
rect 679746 660478 679857 660480
rect 679746 660422 679796 660478
rect 679852 660422 679857 660478
rect 679746 660417 679857 660422
rect 685506 660478 685617 660483
rect 685506 660422 685556 660478
rect 685612 660422 685617 660478
rect 685506 660420 685617 660422
rect 685551 660417 685617 660420
rect 40378 660270 40384 660334
rect 40448 660332 40454 660334
rect 42831 660332 42897 660335
rect 40448 660330 42897 660332
rect 40448 660274 42836 660330
rect 42892 660274 42897 660330
rect 40448 660272 42897 660274
rect 40448 660270 40454 660272
rect 42831 660269 42897 660272
rect 679746 660154 679806 660417
rect 685551 659888 685617 659891
rect 685506 659886 685617 659888
rect 685506 659830 685556 659886
rect 685612 659830 685617 659886
rect 685506 659825 685617 659830
rect 685506 659562 685566 659825
rect 654447 657076 654513 657079
rect 650208 657074 654513 657076
rect 650208 657018 654452 657074
rect 654508 657018 654513 657074
rect 650208 657016 654513 657018
rect 654447 657013 654513 657016
rect 674938 652574 674944 652638
rect 675008 652636 675014 652638
rect 675375 652636 675441 652639
rect 675008 652634 675441 652636
rect 675008 652578 675380 652634
rect 675436 652578 675441 652634
rect 675008 652576 675441 652578
rect 675008 652574 675014 652576
rect 675375 652573 675441 652576
rect 674554 651538 674560 651602
rect 674624 651600 674630 651602
rect 675375 651600 675441 651603
rect 674624 651598 675441 651600
rect 674624 651542 675380 651598
rect 675436 651542 675441 651598
rect 674624 651540 675441 651542
rect 674624 651538 674630 651540
rect 675375 651537 675441 651540
rect 59535 650120 59601 650123
rect 59535 650118 64416 650120
rect 59535 650062 59540 650118
rect 59596 650062 64416 650118
rect 59535 650060 64416 650062
rect 59535 650057 59601 650060
rect 675663 649678 675729 649679
rect 675663 649674 675712 649678
rect 675776 649676 675782 649678
rect 675663 649618 675668 649674
rect 675663 649614 675712 649618
rect 675776 649616 675820 649676
rect 675776 649614 675782 649616
rect 675663 649613 675729 649614
rect 41775 646272 41841 646275
rect 41568 646270 41841 646272
rect 41568 646214 41780 646270
rect 41836 646214 41841 646270
rect 41568 646212 41841 646214
rect 41775 646209 41841 646212
rect 41775 645754 41841 645757
rect 41568 645752 41841 645754
rect 41568 645696 41780 645752
rect 41836 645696 41841 645752
rect 41568 645694 41841 645696
rect 41775 645691 41841 645694
rect 41583 645384 41649 645387
rect 41538 645382 41649 645384
rect 41538 645326 41588 645382
rect 41644 645326 41649 645382
rect 41538 645321 41649 645326
rect 674170 645322 674176 645386
rect 674240 645384 674246 645386
rect 675471 645384 675537 645387
rect 674240 645382 675537 645384
rect 674240 645326 675476 645382
rect 675532 645326 675537 645382
rect 674240 645324 675537 645326
rect 674240 645322 674246 645324
rect 675471 645321 675537 645324
rect 41538 645206 41598 645321
rect 41775 644792 41841 644795
rect 41568 644790 41841 644792
rect 41568 644734 41780 644790
rect 41836 644734 41841 644790
rect 41568 644732 41841 644734
rect 41775 644729 41841 644732
rect 43791 644200 43857 644203
rect 41568 644198 43857 644200
rect 41568 644142 43796 644198
rect 43852 644142 43857 644198
rect 41568 644140 43857 644142
rect 43791 644137 43857 644140
rect 43311 643756 43377 643759
rect 654447 643756 654513 643759
rect 41568 643754 43377 643756
rect 41568 643698 43316 643754
rect 43372 643698 43377 643754
rect 41568 643696 43377 643698
rect 650208 643754 654513 643756
rect 650208 643698 654452 643754
rect 654508 643698 654513 643754
rect 650208 643696 654513 643698
rect 43311 643693 43377 643696
rect 654447 643693 654513 643696
rect 40762 643398 40768 643462
rect 40832 643398 40838 643462
rect 40770 643282 40830 643398
rect 25794 642427 25854 642690
rect 25794 642422 25905 642427
rect 25794 642366 25844 642422
rect 25900 642366 25905 642422
rect 25794 642364 25905 642366
rect 25839 642361 25905 642364
rect 41146 642362 41152 642426
rect 41216 642362 41222 642426
rect 41154 642246 41214 642362
rect 41538 641539 41598 641802
rect 41538 641534 41649 641539
rect 41538 641478 41588 641534
rect 41644 641478 41649 641534
rect 41538 641476 41649 641478
rect 41583 641473 41649 641476
rect 41775 641240 41841 641243
rect 41568 641238 41841 641240
rect 41568 641182 41780 641238
rect 41836 641182 41841 641238
rect 41568 641180 41841 641182
rect 41775 641177 41841 641180
rect 34434 640503 34494 640692
rect 34383 640498 34494 640503
rect 34383 640442 34388 640498
rect 34444 640442 34494 640498
rect 34383 640440 34494 640442
rect 34383 640437 34449 640440
rect 675759 640352 675825 640355
rect 675898 640352 675904 640354
rect 675759 640350 675904 640352
rect 41538 640059 41598 640322
rect 675759 640294 675764 640350
rect 675820 640294 675904 640350
rect 675759 640292 675904 640294
rect 675759 640289 675825 640292
rect 675898 640290 675904 640292
rect 675968 640290 675974 640354
rect 41487 640054 41598 640059
rect 41487 639998 41492 640054
rect 41548 639998 41598 640054
rect 41487 639996 41598 639998
rect 41487 639993 41553 639996
rect 41871 639760 41937 639763
rect 41568 639758 41937 639760
rect 41568 639702 41876 639758
rect 41932 639702 41937 639758
rect 41568 639700 41937 639702
rect 41871 639697 41937 639700
rect 41775 639168 41841 639171
rect 41568 639166 41841 639168
rect 41568 639110 41780 639166
rect 41836 639110 41841 639166
rect 41568 639108 41841 639110
rect 41775 639105 41841 639108
rect 34434 638579 34494 638842
rect 34434 638574 34545 638579
rect 34434 638518 34484 638574
rect 34540 638518 34545 638574
rect 34434 638516 34545 638518
rect 34479 638513 34545 638516
rect 674746 638514 674752 638578
rect 674816 638576 674822 638578
rect 675471 638576 675537 638579
rect 674816 638574 675537 638576
rect 674816 638518 675476 638574
rect 675532 638518 675537 638574
rect 674816 638516 675537 638518
rect 674816 638514 674822 638516
rect 675471 638513 675537 638516
rect 42159 638280 42225 638283
rect 41568 638278 42225 638280
rect 41568 638222 42164 638278
rect 42220 638222 42225 638278
rect 41568 638220 42225 638222
rect 42159 638217 42225 638220
rect 41967 637688 42033 637691
rect 41568 637686 42033 637688
rect 41568 637630 41972 637686
rect 42028 637630 42033 637686
rect 41568 637628 42033 637630
rect 41967 637625 42033 637628
rect 41538 637096 41598 637288
rect 41679 637096 41745 637099
rect 41538 637094 41745 637096
rect 41538 637038 41684 637094
rect 41740 637038 41745 637094
rect 41538 637036 41745 637038
rect 41679 637033 41745 637036
rect 59535 637096 59601 637099
rect 59535 637094 64416 637096
rect 59535 637038 59540 637094
rect 59596 637038 64416 637094
rect 59535 637036 64416 637038
rect 59535 637033 59601 637036
rect 42927 636800 42993 636803
rect 41568 636798 42993 636800
rect 41568 636742 42932 636798
rect 42988 636742 42993 636798
rect 41568 636740 42993 636742
rect 42927 636737 42993 636740
rect 42063 636208 42129 636211
rect 41568 636206 42129 636208
rect 41568 636150 42068 636206
rect 42124 636150 42129 636206
rect 41568 636148 42129 636150
rect 42063 636145 42129 636148
rect 41722 635838 41728 635840
rect 41568 635778 41728 635838
rect 41722 635776 41728 635778
rect 41792 635776 41798 635840
rect 41538 635024 41598 635290
rect 41679 635024 41745 635027
rect 41538 635022 41745 635024
rect 41538 634966 41684 635022
rect 41740 634966 41745 635022
rect 41538 634964 41745 634966
rect 41679 634961 41745 634964
rect 41538 634580 41598 634698
rect 41679 634580 41745 634583
rect 41538 634578 41745 634580
rect 41538 634522 41684 634578
rect 41740 634522 41745 634578
rect 41538 634520 41745 634522
rect 41679 634517 41745 634520
rect 23106 633991 23166 634254
rect 23106 633986 23217 633991
rect 41679 633988 41745 633991
rect 23106 633930 23156 633986
rect 23212 633930 23217 633986
rect 23106 633928 23217 633930
rect 23151 633925 23217 633928
rect 41538 633986 41745 633988
rect 41538 633930 41684 633986
rect 41740 633930 41745 633986
rect 41538 633928 41745 633930
rect 41538 633810 41598 633928
rect 41679 633925 41745 633928
rect 23151 633544 23217 633547
rect 23106 633542 23217 633544
rect 23106 633486 23156 633542
rect 23212 633486 23217 633542
rect 23106 633481 23217 633486
rect 23106 633218 23166 633481
rect 654447 630584 654513 630587
rect 650208 630582 654513 630584
rect 650208 630526 654452 630582
rect 654508 630526 654513 630582
rect 650208 630524 654513 630526
rect 654447 630521 654513 630524
rect 34479 629104 34545 629107
rect 40378 629104 40384 629106
rect 34479 629102 40384 629104
rect 34479 629046 34484 629102
rect 34540 629046 40384 629102
rect 34479 629044 40384 629046
rect 34479 629041 34545 629044
rect 40378 629042 40384 629044
rect 40448 629042 40454 629106
rect 42490 628006 42496 628070
rect 42560 628068 42566 628070
rect 42831 628068 42897 628071
rect 42560 628066 42897 628068
rect 42560 628010 42836 628066
rect 42892 628010 42897 628066
rect 42560 628008 42897 628010
rect 42560 628006 42566 628008
rect 42831 628005 42897 628008
rect 34383 627920 34449 627923
rect 41487 627922 41553 627923
rect 40570 627920 40576 627922
rect 34383 627918 40576 627920
rect 34383 627862 34388 627918
rect 34444 627862 40576 627918
rect 34383 627860 40576 627862
rect 34383 627857 34449 627860
rect 40570 627858 40576 627860
rect 40640 627858 40646 627922
rect 41487 627920 41536 627922
rect 41444 627918 41536 627920
rect 41444 627862 41492 627918
rect 41444 627860 41536 627862
rect 41487 627858 41536 627860
rect 41600 627858 41606 627922
rect 41487 627857 41553 627858
rect 41583 627772 41649 627775
rect 42298 627772 42304 627774
rect 41583 627770 42304 627772
rect 41583 627714 41588 627770
rect 41644 627714 42304 627770
rect 41583 627712 42304 627714
rect 41583 627709 41649 627712
rect 42298 627710 42304 627712
rect 42368 627710 42374 627774
rect 676047 627698 676113 627701
rect 676047 627696 676320 627698
rect 676047 627640 676052 627696
rect 676108 627640 676320 627696
rect 676047 627638 676320 627640
rect 676047 627635 676113 627638
rect 42159 627476 42225 627479
rect 42874 627476 42880 627478
rect 42159 627474 42880 627476
rect 42159 627418 42164 627474
rect 42220 627418 42880 627474
rect 42159 627416 42880 627418
rect 42159 627413 42225 627416
rect 42874 627414 42880 627416
rect 42944 627414 42950 627478
rect 676239 627328 676305 627331
rect 676239 627326 676350 627328
rect 676239 627270 676244 627326
rect 676300 627270 676350 627326
rect 676239 627265 676350 627270
rect 676290 627150 676350 627265
rect 676047 626588 676113 626591
rect 676047 626586 676320 626588
rect 676047 626530 676052 626586
rect 676108 626530 676320 626586
rect 676047 626528 676320 626530
rect 676047 626525 676113 626528
rect 679695 626440 679761 626443
rect 679695 626438 679806 626440
rect 679695 626382 679700 626438
rect 679756 626382 679806 626438
rect 679695 626377 679806 626382
rect 679746 626114 679806 626377
rect 676047 625700 676113 625703
rect 676047 625698 676320 625700
rect 676047 625642 676052 625698
rect 676108 625642 676320 625698
rect 676047 625640 676320 625642
rect 676047 625637 676113 625640
rect 661167 625108 661233 625111
rect 667983 625108 668049 625111
rect 661167 625106 676320 625108
rect 661167 625050 661172 625106
rect 661228 625050 667988 625106
rect 668044 625050 676320 625106
rect 661167 625048 676320 625050
rect 661167 625045 661233 625048
rect 667983 625045 668049 625048
rect 675951 624664 676017 624667
rect 675951 624662 676320 624664
rect 675951 624606 675956 624662
rect 676012 624606 676320 624662
rect 675951 624604 676320 624606
rect 675951 624601 676017 624604
rect 666831 624220 666897 624223
rect 672495 624220 672561 624223
rect 666831 624218 676320 624220
rect 666831 624162 666836 624218
rect 666892 624162 672500 624218
rect 672556 624162 676320 624218
rect 666831 624160 676320 624162
rect 666831 624157 666897 624160
rect 672495 624157 672561 624160
rect 59535 624072 59601 624075
rect 59535 624070 64416 624072
rect 59535 624014 59540 624070
rect 59596 624014 64416 624070
rect 59535 624012 64416 624014
rect 59535 624009 59601 624012
rect 675951 623628 676017 623631
rect 675951 623626 676320 623628
rect 675951 623570 675956 623626
rect 676012 623570 676320 623626
rect 675951 623568 676320 623570
rect 675951 623565 676017 623568
rect 675514 623122 675520 623186
rect 675584 623184 675590 623186
rect 675584 623124 676320 623184
rect 675584 623122 675590 623124
rect 676047 622666 676113 622669
rect 676047 622664 676320 622666
rect 676047 622608 676052 622664
rect 676108 622608 676320 622664
rect 676047 622606 676320 622608
rect 676047 622603 676113 622606
rect 42159 622148 42225 622151
rect 42490 622148 42496 622150
rect 42159 622146 42496 622148
rect 42159 622090 42164 622146
rect 42220 622090 42496 622146
rect 42159 622088 42496 622090
rect 42159 622085 42225 622088
rect 42490 622086 42496 622088
rect 42560 622086 42566 622150
rect 675322 622086 675328 622150
rect 675392 622148 675398 622150
rect 675392 622088 676320 622148
rect 675392 622086 675398 622088
rect 675130 621642 675136 621706
rect 675200 621704 675206 621706
rect 675200 621644 676320 621704
rect 675200 621642 675206 621644
rect 42298 621494 42304 621558
rect 42368 621556 42374 621558
rect 42831 621556 42897 621559
rect 42368 621554 42897 621556
rect 42368 621498 42836 621554
rect 42892 621498 42897 621554
rect 42368 621496 42897 621498
rect 42368 621494 42374 621496
rect 42831 621493 42897 621496
rect 673978 621050 673984 621114
rect 674048 621112 674054 621114
rect 674048 621052 676320 621112
rect 674048 621050 674054 621052
rect 41775 620966 41841 620967
rect 41722 620964 41728 620966
rect 41684 620904 41728 620964
rect 41792 620962 41841 620966
rect 41836 620906 41841 620962
rect 41722 620902 41728 620904
rect 41792 620902 41841 620906
rect 41775 620901 41841 620902
rect 676239 620816 676305 620819
rect 676239 620814 676350 620816
rect 676239 620758 676244 620814
rect 676300 620758 676350 620814
rect 676239 620753 676350 620758
rect 676290 620638 676350 620753
rect 676282 620310 676288 620374
rect 676352 620310 676358 620374
rect 42927 620226 42993 620227
rect 42874 620162 42880 620226
rect 42944 620224 42993 620226
rect 42944 620222 43036 620224
rect 42988 620166 43036 620222
rect 676290 620194 676350 620310
rect 42944 620164 43036 620166
rect 42944 620162 42993 620164
rect 42927 620161 42993 620162
rect 676474 619866 676480 619930
rect 676544 619866 676550 619930
rect 676482 619602 676542 619866
rect 41722 619126 41728 619190
rect 41792 619188 41798 619190
rect 44367 619188 44433 619191
rect 41792 619186 44433 619188
rect 41792 619130 44372 619186
rect 44428 619130 44433 619186
rect 41792 619128 44433 619130
rect 41792 619126 41798 619128
rect 44367 619125 44433 619128
rect 676047 619188 676113 619191
rect 676047 619186 676320 619188
rect 676047 619130 676052 619186
rect 676108 619130 676320 619186
rect 676047 619128 676320 619130
rect 676047 619125 676113 619128
rect 40570 618830 40576 618894
rect 40640 618892 40646 618894
rect 43023 618892 43089 618895
rect 40640 618890 43089 618892
rect 40640 618834 43028 618890
rect 43084 618834 43089 618890
rect 40640 618832 43089 618834
rect 40640 618830 40646 618832
rect 43023 618829 43089 618832
rect 676858 618830 676864 618894
rect 676928 618830 676934 618894
rect 676866 618714 676926 618830
rect 676047 618152 676113 618155
rect 676047 618150 676320 618152
rect 676047 618094 676052 618150
rect 676108 618094 676320 618150
rect 676047 618092 676320 618094
rect 676047 618089 676113 618092
rect 676047 617634 676113 617637
rect 676047 617632 676320 617634
rect 676047 617576 676052 617632
rect 676108 617576 676320 617632
rect 676047 617574 676320 617576
rect 676047 617571 676113 617574
rect 676239 617412 676305 617415
rect 676239 617410 676350 617412
rect 676239 617354 676244 617410
rect 676300 617354 676350 617410
rect 676239 617349 676350 617354
rect 654543 617264 654609 617267
rect 650208 617262 654609 617264
rect 650208 617206 654548 617262
rect 654604 617206 654609 617262
rect 676290 617234 676350 617349
rect 650208 617204 654609 617206
rect 654543 617201 654609 617204
rect 676047 616672 676113 616675
rect 676047 616670 676320 616672
rect 676047 616614 676052 616670
rect 676108 616614 676320 616670
rect 676047 616612 676320 616614
rect 676047 616609 676113 616612
rect 40378 616462 40384 616526
rect 40448 616524 40454 616526
rect 42927 616524 42993 616527
rect 40448 616522 42993 616524
rect 40448 616466 42932 616522
rect 42988 616466 42993 616522
rect 40448 616464 42993 616466
rect 40448 616462 40454 616464
rect 42927 616461 42993 616464
rect 41530 616018 41536 616082
rect 41600 616080 41606 616082
rect 41775 616080 41841 616083
rect 41600 616078 41841 616080
rect 41600 616022 41780 616078
rect 41836 616022 41841 616078
rect 41600 616020 41841 616022
rect 41600 616018 41606 616020
rect 41775 616017 41841 616020
rect 679746 615935 679806 616050
rect 679746 615930 679857 615935
rect 679746 615874 679796 615930
rect 679852 615874 679857 615930
rect 679746 615872 679857 615874
rect 679791 615869 679857 615872
rect 685506 615343 685566 615754
rect 679791 615340 679857 615343
rect 679746 615338 679857 615340
rect 679746 615282 679796 615338
rect 679852 615282 679857 615338
rect 679746 615277 679857 615282
rect 685455 615338 685566 615343
rect 685455 615282 685460 615338
rect 685516 615282 685566 615338
rect 685455 615280 685566 615282
rect 685455 615277 685521 615280
rect 679746 615162 679806 615277
rect 685455 614896 685521 614899
rect 685455 614894 685566 614896
rect 685455 614838 685460 614894
rect 685516 614838 685566 614894
rect 685455 614833 685566 614838
rect 685506 614570 685566 614833
rect 59247 611048 59313 611051
rect 59247 611046 64416 611048
rect 59247 610990 59252 611046
rect 59308 610990 64416 611046
rect 59247 610988 64416 610990
rect 59247 610985 59313 610988
rect 673978 607730 673984 607794
rect 674048 607792 674054 607794
rect 675375 607792 675441 607795
rect 674048 607790 675441 607792
rect 674048 607734 675380 607790
rect 675436 607734 675441 607790
rect 674048 607732 675441 607734
rect 674048 607730 674054 607732
rect 675375 607729 675441 607732
rect 41530 607582 41536 607646
rect 41600 607644 41606 607646
rect 47439 607644 47505 607647
rect 41600 607642 47505 607644
rect 41600 607586 47444 607642
rect 47500 607586 47505 607642
rect 41600 607584 47505 607586
rect 41600 607582 41606 607584
rect 47439 607581 47505 607584
rect 675130 606398 675136 606462
rect 675200 606460 675206 606462
rect 675375 606460 675441 606463
rect 675200 606458 675441 606460
rect 675200 606402 675380 606458
rect 675436 606402 675441 606458
rect 675200 606400 675441 606402
rect 675200 606398 675206 606400
rect 675375 606397 675441 606400
rect 674362 604770 674368 604834
rect 674432 604832 674438 604834
rect 675375 604832 675441 604835
rect 674432 604830 675441 604832
rect 674432 604774 675380 604830
rect 675436 604774 675441 604830
rect 674432 604772 675441 604774
rect 674432 604770 674438 604772
rect 675375 604769 675441 604772
rect 654447 603944 654513 603947
rect 650208 603942 654513 603944
rect 650208 603886 654452 603942
rect 654508 603886 654513 603942
rect 650208 603884 654513 603886
rect 654447 603881 654513 603884
rect 41775 603056 41841 603059
rect 41568 603054 41841 603056
rect 41568 602998 41780 603054
rect 41836 602998 41841 603054
rect 41568 602996 41841 602998
rect 41775 602993 41841 602996
rect 41583 602760 41649 602763
rect 41538 602758 41649 602760
rect 41538 602702 41588 602758
rect 41644 602702 41649 602758
rect 41538 602697 41649 602702
rect 41538 602582 41598 602697
rect 41583 602168 41649 602171
rect 41538 602166 41649 602168
rect 41538 602110 41588 602166
rect 41644 602110 41649 602166
rect 41538 602105 41649 602110
rect 41538 601990 41598 602105
rect 41775 601576 41841 601579
rect 41568 601574 41841 601576
rect 41568 601518 41780 601574
rect 41836 601518 41841 601574
rect 41568 601516 41841 601518
rect 41775 601513 41841 601516
rect 41775 601058 41841 601061
rect 41568 601056 41841 601058
rect 41568 601000 41780 601056
rect 41836 601000 41841 601056
rect 41568 600998 41841 601000
rect 41775 600995 41841 600998
rect 40762 600626 40768 600690
rect 40832 600626 40838 600690
rect 40770 600540 40830 600626
rect 41722 600540 41728 600542
rect 40770 600510 41728 600540
rect 40800 600480 41728 600510
rect 41722 600478 41728 600480
rect 41792 600478 41798 600542
rect 675322 600182 675328 600246
rect 675392 600244 675398 600246
rect 675471 600244 675537 600247
rect 675392 600242 675537 600244
rect 675392 600186 675476 600242
rect 675532 600186 675537 600242
rect 675392 600184 675537 600186
rect 675392 600182 675398 600184
rect 675471 600181 675537 600184
rect 41538 599951 41598 600066
rect 41538 599946 41649 599951
rect 41538 599890 41588 599946
rect 41644 599890 41649 599946
rect 41538 599888 41649 599890
rect 41583 599885 41649 599888
rect 41530 599738 41536 599802
rect 41600 599738 41606 599802
rect 41538 599504 41598 599738
rect 40608 599474 41598 599504
rect 40578 599444 41568 599474
rect 40578 599358 40638 599444
rect 40570 599294 40576 599358
rect 40640 599294 40646 599358
rect 41775 599060 41841 599063
rect 41568 599058 41841 599060
rect 41568 599002 41780 599058
rect 41836 599002 41841 599058
rect 41568 599000 41841 599002
rect 41775 598997 41841 599000
rect 41538 598323 41598 598586
rect 41487 598318 41598 598323
rect 41487 598262 41492 598318
rect 41548 598262 41598 598318
rect 41487 598260 41598 598262
rect 41487 598257 41553 598260
rect 59343 598024 59409 598027
rect 59343 598022 64416 598024
rect 41538 597879 41598 597994
rect 59343 597966 59348 598022
rect 59404 597966 64416 598022
rect 59343 597964 64416 597966
rect 59343 597961 59409 597964
rect 41538 597874 41649 597879
rect 41538 597818 41588 597874
rect 41644 597818 41649 597874
rect 41538 597816 41649 597818
rect 41583 597813 41649 597816
rect 34434 597287 34494 597550
rect 34383 597282 34494 597287
rect 34383 597226 34388 597282
rect 34444 597226 34494 597282
rect 34383 597224 34494 597226
rect 34383 597221 34449 597224
rect 42063 597136 42129 597139
rect 41568 597134 42129 597136
rect 41568 597078 42068 597134
rect 42124 597078 42129 597134
rect 41568 597076 42129 597078
rect 42063 597073 42129 597076
rect 41538 596396 41598 596514
rect 41679 596396 41745 596399
rect 41538 596394 41745 596396
rect 41538 596338 41684 596394
rect 41740 596338 41745 596394
rect 41538 596336 41745 596338
rect 41679 596333 41745 596336
rect 41871 596026 41937 596029
rect 41568 596024 41937 596026
rect 41568 595968 41876 596024
rect 41932 595968 41937 596024
rect 41568 595966 41937 595968
rect 41871 595963 41937 595966
rect 34434 595363 34494 595626
rect 34434 595358 34545 595363
rect 34434 595302 34484 595358
rect 34540 595302 34545 595358
rect 34434 595300 34545 595302
rect 34479 595297 34545 595300
rect 675759 595360 675825 595363
rect 676090 595360 676096 595362
rect 675759 595358 676096 595360
rect 675759 595302 675764 595358
rect 675820 595302 676096 595358
rect 675759 595300 676096 595302
rect 675759 595297 675825 595300
rect 676090 595298 676096 595300
rect 676160 595298 676166 595362
rect 41967 595064 42033 595067
rect 41568 595062 42033 595064
rect 41568 595006 41972 595062
rect 42028 595006 42033 595062
rect 41568 595004 42033 595006
rect 41967 595001 42033 595004
rect 42159 594472 42225 594475
rect 41568 594470 42225 594472
rect 41568 594414 42164 594470
rect 42220 594414 42225 594470
rect 41568 594412 42225 594414
rect 42159 594409 42225 594412
rect 41775 594176 41841 594179
rect 41568 594174 41841 594176
rect 41568 594118 41780 594174
rect 41836 594118 41841 594174
rect 41568 594116 41841 594118
rect 41775 594113 41841 594116
rect 41775 593584 41841 593587
rect 41568 593582 41841 593584
rect 41568 593526 41780 593582
rect 41836 593526 41841 593582
rect 41568 593524 41841 593526
rect 41775 593521 41841 593524
rect 675471 593438 675537 593439
rect 675471 593434 675520 593438
rect 675584 593436 675590 593438
rect 675471 593378 675476 593434
rect 675471 593374 675520 593378
rect 675584 593376 675628 593436
rect 675584 593374 675590 593376
rect 675471 593373 675537 593374
rect 42447 592992 42513 592995
rect 41568 592990 42513 592992
rect 41568 592934 42452 592990
rect 42508 592934 42513 592990
rect 41568 592932 42513 592934
rect 42447 592929 42513 592932
rect 41775 592622 41841 592625
rect 41568 592620 41841 592622
rect 41568 592564 41780 592620
rect 41836 592564 41841 592620
rect 41568 592562 41841 592564
rect 41775 592559 41841 592562
rect 41775 592104 41841 592107
rect 41568 592102 41841 592104
rect 41568 592046 41780 592102
rect 41836 592046 41841 592102
rect 41568 592044 41841 592046
rect 41775 592041 41841 592044
rect 41538 591367 41598 591482
rect 41538 591362 41649 591367
rect 41538 591306 41588 591362
rect 41644 591306 41649 591362
rect 41538 591304 41649 591306
rect 41583 591301 41649 591304
rect 23106 590775 23166 591112
rect 23055 590770 23166 590775
rect 41583 590772 41649 590775
rect 654447 590772 654513 590775
rect 23055 590714 23060 590770
rect 23116 590714 23166 590770
rect 23055 590712 23166 590714
rect 41538 590770 41649 590772
rect 41538 590714 41588 590770
rect 41644 590714 41649 590770
rect 23055 590709 23121 590712
rect 41538 590709 41649 590714
rect 650208 590770 654513 590772
rect 650208 590714 654452 590770
rect 654508 590714 654513 590770
rect 650208 590712 654513 590714
rect 654447 590709 654513 590712
rect 41538 590594 41598 590709
rect 23055 590328 23121 590331
rect 23055 590326 23166 590328
rect 23055 590270 23060 590326
rect 23116 590270 23166 590326
rect 23055 590265 23166 590270
rect 23106 590002 23166 590265
rect 34383 585584 34449 585587
rect 40378 585584 40384 585586
rect 34383 585582 40384 585584
rect 34383 585526 34388 585582
rect 34444 585526 40384 585582
rect 34383 585524 40384 585526
rect 34383 585521 34449 585524
rect 40378 585522 40384 585524
rect 40448 585522 40454 585586
rect 34479 585436 34545 585439
rect 40954 585436 40960 585438
rect 34479 585434 40960 585436
rect 34479 585378 34484 585434
rect 34540 585378 40960 585434
rect 34479 585376 40960 585378
rect 34479 585373 34545 585376
rect 40954 585374 40960 585376
rect 41024 585374 41030 585438
rect 59535 584852 59601 584855
rect 59535 584850 64416 584852
rect 59535 584794 59540 584850
rect 59596 584794 64416 584850
rect 59535 584792 64416 584794
rect 59535 584789 59601 584792
rect 41487 584556 41553 584559
rect 43066 584556 43072 584558
rect 41487 584554 43072 584556
rect 41487 584498 41492 584554
rect 41548 584498 43072 584554
rect 41487 584496 43072 584498
rect 41487 584493 41553 584496
rect 43066 584494 43072 584496
rect 43136 584494 43142 584558
rect 42063 584260 42129 584263
rect 42874 584260 42880 584262
rect 42063 584258 42880 584260
rect 42063 584202 42068 584258
rect 42124 584202 42880 584258
rect 42063 584200 42880 584202
rect 42063 584197 42129 584200
rect 42874 584198 42880 584200
rect 42944 584198 42950 584262
rect 676047 582484 676113 582487
rect 676047 582482 676320 582484
rect 676047 582426 676052 582482
rect 676108 582426 676320 582482
rect 676047 582424 676320 582426
rect 676047 582421 676113 582424
rect 676047 581966 676113 581969
rect 676047 581964 676320 581966
rect 676047 581908 676052 581964
rect 676108 581908 676320 581964
rect 676047 581906 676320 581908
rect 676047 581903 676113 581906
rect 676239 581596 676305 581599
rect 676239 581594 676350 581596
rect 676239 581538 676244 581594
rect 676300 581538 676350 581594
rect 676239 581533 676350 581538
rect 676290 581418 676350 581533
rect 676047 581004 676113 581007
rect 676047 581002 676320 581004
rect 676047 580946 676052 581002
rect 676108 580946 676320 581002
rect 676047 580944 676320 580946
rect 676047 580941 676113 580944
rect 676290 580267 676350 580382
rect 676239 580262 676350 580267
rect 676239 580206 676244 580262
rect 676300 580206 676350 580262
rect 676239 580204 676350 580206
rect 676239 580201 676305 580204
rect 676047 579968 676113 579971
rect 676047 579966 676320 579968
rect 676047 579910 676052 579966
rect 676108 579910 676320 579966
rect 676047 579908 676320 579910
rect 676047 579905 676113 579908
rect 676047 579524 676113 579527
rect 676047 579522 676320 579524
rect 676047 579466 676052 579522
rect 676108 579466 676320 579522
rect 676047 579464 676320 579466
rect 676047 579461 676113 579464
rect 676047 578932 676113 578935
rect 676047 578930 676320 578932
rect 676047 578874 676052 578930
rect 676108 578874 676320 578930
rect 676047 578872 676320 578874
rect 676047 578869 676113 578872
rect 42831 578786 42897 578787
rect 42831 578784 42880 578786
rect 42788 578782 42880 578784
rect 42788 578726 42836 578782
rect 42788 578724 42880 578726
rect 42831 578722 42880 578724
rect 42944 578722 42950 578786
rect 42831 578721 42897 578722
rect 676047 578414 676113 578417
rect 676047 578412 676320 578414
rect 676047 578356 676052 578412
rect 676108 578356 676320 578412
rect 676047 578354 676320 578356
rect 676047 578351 676113 578354
rect 674554 577982 674560 578046
rect 674624 578044 674630 578046
rect 674624 577984 676320 578044
rect 674624 577982 674630 577984
rect 42927 577600 42993 577603
rect 43066 577600 43072 577602
rect 42927 577598 43072 577600
rect 42927 577542 42932 577598
rect 42988 577542 43072 577598
rect 42927 577540 43072 577542
rect 42927 577537 42993 577540
rect 43066 577538 43072 577540
rect 43136 577538 43142 577602
rect 654447 577452 654513 577455
rect 650208 577450 654513 577452
rect 650208 577394 654452 577450
rect 654508 577394 654513 577450
rect 650208 577392 654513 577394
rect 654447 577389 654513 577392
rect 675898 577390 675904 577454
rect 675968 577452 675974 577454
rect 675968 577392 676320 577452
rect 675968 577390 675974 577392
rect 674938 577242 674944 577306
rect 675008 577304 675014 577306
rect 675008 577244 676350 577304
rect 675008 577242 675014 577244
rect 676290 576904 676350 577244
rect 675706 576502 675712 576566
rect 675776 576564 675782 576566
rect 675776 576504 676320 576564
rect 675776 576502 675782 576504
rect 674170 575910 674176 575974
rect 674240 575972 674246 575974
rect 674240 575912 676320 575972
rect 674240 575910 674246 575912
rect 674746 575318 674752 575382
rect 674816 575380 674822 575382
rect 674816 575320 676320 575380
rect 674816 575318 674822 575320
rect 676047 575010 676113 575013
rect 676047 575008 676320 575010
rect 676047 574952 676052 575008
rect 676108 574952 676320 575008
rect 676047 574950 676320 574952
rect 676047 574947 676113 574950
rect 676239 574640 676305 574643
rect 676239 574638 676350 574640
rect 676239 574582 676244 574638
rect 676300 574582 676350 574638
rect 676239 574577 676350 574582
rect 40954 574430 40960 574494
rect 41024 574492 41030 574494
rect 42351 574492 42417 574495
rect 41024 574490 42417 574492
rect 41024 574434 42356 574490
rect 42412 574434 42417 574490
rect 676290 574462 676350 574577
rect 41024 574432 42417 574434
rect 41024 574430 41030 574432
rect 42351 574429 42417 574432
rect 40378 573986 40384 574050
rect 40448 574048 40454 574050
rect 42735 574048 42801 574051
rect 40448 574046 42801 574048
rect 40448 573990 42740 574046
rect 42796 573990 42801 574046
rect 40448 573988 42801 573990
rect 40448 573986 40454 573988
rect 42735 573985 42801 573988
rect 676047 573900 676113 573903
rect 676047 573898 676320 573900
rect 676047 573842 676052 573898
rect 676108 573842 676320 573898
rect 676047 573840 676320 573842
rect 676047 573837 676113 573840
rect 676047 573530 676113 573533
rect 676047 573528 676320 573530
rect 676047 573472 676052 573528
rect 676108 573472 676320 573528
rect 676047 573470 676320 573472
rect 676047 573467 676113 573470
rect 676047 573012 676113 573015
rect 676047 573010 676320 573012
rect 676047 572954 676052 573010
rect 676108 572954 676320 573010
rect 676047 572952 676320 572954
rect 676047 572949 676113 572952
rect 676047 572420 676113 572423
rect 676047 572418 676320 572420
rect 676047 572362 676052 572418
rect 676108 572362 676320 572418
rect 676047 572360 676320 572362
rect 676047 572357 676113 572360
rect 676047 571976 676113 571979
rect 676047 571974 676320 571976
rect 676047 571918 676052 571974
rect 676108 571918 676320 571974
rect 676047 571916 676320 571918
rect 676047 571913 676113 571916
rect 59535 571828 59601 571831
rect 59535 571826 64416 571828
rect 59535 571770 59540 571826
rect 59596 571770 64416 571826
rect 59535 571768 64416 571770
rect 59535 571765 59601 571768
rect 676239 571680 676305 571683
rect 676239 571678 676350 571680
rect 676239 571622 676244 571678
rect 676300 571622 676350 571678
rect 676239 571617 676350 571622
rect 676290 571502 676350 571617
rect 679983 571236 680049 571239
rect 679938 571234 680049 571236
rect 679938 571178 679988 571234
rect 680044 571178 680049 571234
rect 679938 571173 680049 571178
rect 679938 570910 679998 571173
rect 679746 570203 679806 570466
rect 679746 570198 679857 570203
rect 679983 570200 680049 570203
rect 679746 570142 679796 570198
rect 679852 570142 679857 570198
rect 679746 570140 679857 570142
rect 679791 570137 679857 570140
rect 679938 570198 680049 570200
rect 679938 570142 679988 570198
rect 680044 570142 680049 570198
rect 679938 570137 680049 570142
rect 679938 569948 679998 570137
rect 679791 569756 679857 569759
rect 679746 569754 679857 569756
rect 679746 569698 679796 569754
rect 679852 569698 679857 569754
rect 679746 569693 679857 569698
rect 679746 569430 679806 569693
rect 656559 564132 656625 564135
rect 650208 564130 656625 564132
rect 650208 564074 656564 564130
rect 656620 564074 656625 564130
rect 650208 564072 656625 564074
rect 656559 564069 656625 564072
rect 674554 562590 674560 562654
rect 674624 562652 674630 562654
rect 675471 562652 675537 562655
rect 674624 562650 675537 562652
rect 674624 562594 675476 562650
rect 675532 562594 675537 562650
rect 674624 562592 675537 562594
rect 674624 562590 674630 562592
rect 675471 562589 675537 562592
rect 674938 561702 674944 561766
rect 675008 561764 675014 561766
rect 675471 561764 675537 561767
rect 675008 561762 675537 561764
rect 675008 561706 675476 561762
rect 675532 561706 675537 561762
rect 675008 561704 675537 561706
rect 675008 561702 675014 561704
rect 675471 561701 675537 561704
rect 674746 561406 674752 561470
rect 674816 561468 674822 561470
rect 675471 561468 675537 561471
rect 674816 561466 675537 561468
rect 674816 561410 675476 561466
rect 675532 561410 675537 561466
rect 674816 561408 675537 561410
rect 674816 561406 674822 561408
rect 675471 561405 675537 561408
rect 41775 559840 41841 559843
rect 41568 559838 41841 559840
rect 41568 559782 41780 559838
rect 41836 559782 41841 559838
rect 41568 559780 41841 559782
rect 41775 559777 41841 559780
rect 42351 559396 42417 559399
rect 41568 559394 42417 559396
rect 41568 559338 42356 559394
rect 42412 559338 42417 559394
rect 41568 559336 42417 559338
rect 42351 559333 42417 559336
rect 41722 558890 41728 558954
rect 41792 558952 41798 558954
rect 44463 558952 44529 558955
rect 41792 558950 44529 558952
rect 41792 558894 44468 558950
rect 44524 558894 44529 558950
rect 41792 558892 44529 558894
rect 41792 558890 41798 558892
rect 44463 558889 44529 558892
rect 41775 558804 41841 558807
rect 41568 558802 41841 558804
rect 41568 558746 41780 558802
rect 41836 558746 41841 558802
rect 41568 558744 41841 558746
rect 41775 558741 41841 558744
rect 59535 558804 59601 558807
rect 59535 558802 64416 558804
rect 59535 558746 59540 558802
rect 59596 558746 64416 558802
rect 59535 558744 64416 558746
rect 59535 558741 59601 558744
rect 41775 558360 41841 558363
rect 41568 558358 41841 558360
rect 41568 558302 41780 558358
rect 41836 558302 41841 558358
rect 41568 558300 41841 558302
rect 41775 558297 41841 558300
rect 41775 557916 41841 557919
rect 41568 557914 41841 557916
rect 41568 557858 41780 557914
rect 41836 557858 41841 557914
rect 41568 557856 41841 557858
rect 41775 557853 41841 557856
rect 675759 557620 675825 557623
rect 676858 557620 676864 557622
rect 675759 557618 676864 557620
rect 675759 557562 675764 557618
rect 675820 557562 676864 557618
rect 675759 557560 676864 557562
rect 675759 557557 675825 557560
rect 676858 557558 676864 557560
rect 676928 557558 676934 557622
rect 40378 557410 40384 557474
rect 40448 557410 40454 557474
rect 40386 557294 40446 557410
rect 40770 556734 40830 556850
rect 40762 556670 40768 556734
rect 40832 556670 40838 556734
rect 41722 556362 41728 556364
rect 40800 556332 41728 556362
rect 40770 556302 41728 556332
rect 40770 556142 40830 556302
rect 41722 556300 41728 556302
rect 41792 556300 41798 556364
rect 40762 556078 40768 556142
rect 40832 556078 40838 556142
rect 40570 555930 40576 555994
rect 40640 555930 40646 555994
rect 40578 555814 40638 555930
rect 42255 555400 42321 555403
rect 41568 555398 42321 555400
rect 41568 555342 42260 555398
rect 42316 555342 42321 555398
rect 41568 555340 42321 555342
rect 42255 555337 42321 555340
rect 41538 554663 41598 554778
rect 41538 554658 41649 554663
rect 41538 554602 41588 554658
rect 41644 554602 41649 554658
rect 41538 554600 41649 554602
rect 41583 554597 41649 554600
rect 34434 554071 34494 554334
rect 34383 554066 34494 554071
rect 41679 554068 41745 554071
rect 34383 554010 34388 554066
rect 34444 554010 34494 554066
rect 34383 554008 34494 554010
rect 41538 554066 41745 554068
rect 41538 554010 41684 554066
rect 41740 554010 41745 554066
rect 41538 554008 41745 554010
rect 34383 554005 34449 554008
rect 41538 553890 41598 554008
rect 41679 554005 41745 554008
rect 42159 553328 42225 553331
rect 41568 553326 42225 553328
rect 41568 553270 42164 553326
rect 42220 553270 42225 553326
rect 41568 553268 42225 553270
rect 42159 553265 42225 553268
rect 41775 552884 41841 552887
rect 41568 552882 41841 552884
rect 41568 552826 41780 552882
rect 41836 552826 41841 552882
rect 41568 552824 41841 552826
rect 41775 552821 41841 552824
rect 34434 552147 34494 552410
rect 34434 552142 34545 552147
rect 34434 552086 34484 552142
rect 34540 552086 34545 552142
rect 34434 552084 34545 552086
rect 34479 552081 34545 552084
rect 41538 551703 41598 551818
rect 41487 551698 41598 551703
rect 41487 551642 41492 551698
rect 41548 551642 41598 551698
rect 41487 551640 41598 551642
rect 41487 551637 41553 551640
rect 41967 551330 42033 551333
rect 41568 551328 42033 551330
rect 41568 551272 41972 551328
rect 42028 551272 42033 551328
rect 41568 551270 42033 551272
rect 41967 551267 42033 551270
rect 41871 550960 41937 550963
rect 654831 550960 654897 550963
rect 41568 550958 41937 550960
rect 41568 550902 41876 550958
rect 41932 550902 41937 550958
rect 41568 550900 41937 550902
rect 650208 550958 654897 550960
rect 650208 550902 654836 550958
rect 654892 550902 654897 550958
rect 650208 550900 654897 550902
rect 41871 550897 41937 550900
rect 654831 550897 654897 550900
rect 41538 550223 41598 550338
rect 41538 550218 41649 550223
rect 41538 550162 41588 550218
rect 41644 550162 41649 550218
rect 41538 550160 41649 550162
rect 41583 550157 41649 550160
rect 42159 549776 42225 549779
rect 41568 549774 42225 549776
rect 41568 549718 42164 549774
rect 42220 549718 42225 549774
rect 41568 549716 42225 549718
rect 42159 549713 42225 549716
rect 41346 549187 41406 549450
rect 41346 549182 41457 549187
rect 41346 549126 41396 549182
rect 41452 549126 41457 549182
rect 41346 549124 41457 549126
rect 41391 549121 41457 549124
rect 41871 548888 41937 548891
rect 41568 548886 41937 548888
rect 41568 548830 41876 548886
rect 41932 548830 41937 548886
rect 41568 548828 41937 548830
rect 41871 548825 41937 548828
rect 41538 548148 41598 548266
rect 41538 548088 41790 548148
rect 23106 547559 23166 547896
rect 41730 547704 41790 548088
rect 23055 547554 23166 547559
rect 23055 547498 23060 547554
rect 23116 547498 23166 547554
rect 23055 547496 23166 547498
rect 41538 547644 41790 547704
rect 23055 547493 23121 547496
rect 41538 547408 41598 547644
rect 41871 547408 41937 547411
rect 41538 547406 41937 547408
rect 41538 547378 41876 547406
rect 41568 547350 41876 547378
rect 41932 547350 41937 547406
rect 41568 547348 41937 547350
rect 41871 547345 41937 547348
rect 23055 547112 23121 547115
rect 23055 547110 23166 547112
rect 23055 547054 23060 547110
rect 23116 547054 23166 547110
rect 23055 547049 23166 547054
rect 23106 546786 23166 547049
rect 59535 545928 59601 545931
rect 59535 545926 64416 545928
rect 59535 545870 59540 545926
rect 59596 545870 64416 545926
rect 59535 545868 64416 545870
rect 59535 545865 59601 545868
rect 34479 541636 34545 541639
rect 40954 541636 40960 541638
rect 34479 541634 40960 541636
rect 34479 541578 34484 541634
rect 34540 541578 40960 541634
rect 34479 541576 40960 541578
rect 34479 541573 34545 541576
rect 40954 541574 40960 541576
rect 41024 541574 41030 541638
rect 42490 541574 42496 541638
rect 42560 541636 42566 541638
rect 42735 541636 42801 541639
rect 42560 541634 42801 541636
rect 42560 541578 42740 541634
rect 42796 541578 42801 541634
rect 42560 541576 42801 541578
rect 42560 541574 42566 541576
rect 42735 541573 42801 541576
rect 34383 541488 34449 541491
rect 41146 541488 41152 541490
rect 34383 541486 41152 541488
rect 34383 541430 34388 541486
rect 34444 541430 41152 541486
rect 34383 541428 41152 541430
rect 34383 541425 34449 541428
rect 41146 541426 41152 541428
rect 41216 541426 41222 541490
rect 41679 541342 41745 541343
rect 41679 541340 41728 541342
rect 41636 541338 41728 541340
rect 41636 541282 41684 541338
rect 41636 541280 41728 541282
rect 41679 541278 41728 541280
rect 41792 541278 41798 541342
rect 41679 541277 41745 541278
rect 41967 541046 42033 541047
rect 41914 541044 41920 541046
rect 41876 540984 41920 541044
rect 41984 541042 42033 541046
rect 42028 540986 42033 541042
rect 41914 540982 41920 540984
rect 41984 540982 42033 540986
rect 41967 540981 42033 540982
rect 42159 541044 42225 541047
rect 42298 541044 42304 541046
rect 42159 541042 42304 541044
rect 42159 540986 42164 541042
rect 42220 540986 42304 541042
rect 42159 540984 42304 540986
rect 42159 540981 42225 540984
rect 42298 540982 42304 540984
rect 42368 540982 42374 541046
rect 654447 537640 654513 537643
rect 650208 537638 654513 537640
rect 650208 537582 654452 537638
rect 654508 537582 654513 537638
rect 650208 537580 654513 537582
rect 654447 537577 654513 537580
rect 676047 537492 676113 537495
rect 676047 537490 676320 537492
rect 676047 537434 676052 537490
rect 676108 537434 676320 537490
rect 676047 537432 676320 537434
rect 676047 537429 676113 537432
rect 676047 536900 676113 536903
rect 676047 536898 676320 536900
rect 676047 536842 676052 536898
rect 676108 536842 676320 536898
rect 676047 536840 676320 536842
rect 676047 536837 676113 536840
rect 676239 536604 676305 536607
rect 676239 536602 676350 536604
rect 676239 536546 676244 536602
rect 676300 536546 676350 536602
rect 676239 536541 676350 536546
rect 676290 536426 676350 536541
rect 679695 536160 679761 536163
rect 679695 536158 679806 536160
rect 679695 536102 679700 536158
rect 679756 536102 679806 536158
rect 679695 536097 679806 536102
rect 679746 535982 679806 536097
rect 42298 535654 42304 535718
rect 42368 535716 42374 535718
rect 42831 535716 42897 535719
rect 42368 535714 42897 535716
rect 42368 535658 42836 535714
rect 42892 535658 42897 535714
rect 42368 535656 42897 535658
rect 42368 535654 42374 535656
rect 42831 535653 42897 535656
rect 676482 535275 676542 535390
rect 676482 535270 676593 535275
rect 676482 535214 676532 535270
rect 676588 535214 676593 535270
rect 676482 535212 676593 535214
rect 676527 535209 676593 535212
rect 42159 535124 42225 535127
rect 42490 535124 42496 535126
rect 42159 535122 42496 535124
rect 42159 535066 42164 535122
rect 42220 535066 42496 535122
rect 42159 535064 42496 535066
rect 42159 535061 42225 535064
rect 42490 535062 42496 535064
rect 42560 535062 42566 535126
rect 676047 534902 676113 534905
rect 676047 534900 676320 534902
rect 676047 534844 676052 534900
rect 676108 534844 676320 534900
rect 676047 534842 676320 534844
rect 676047 534839 676113 534842
rect 676674 534239 676734 534502
rect 676623 534234 676734 534239
rect 676623 534178 676628 534234
rect 676684 534178 676734 534234
rect 676623 534176 676734 534178
rect 676623 534173 676689 534176
rect 676047 533940 676113 533943
rect 676047 533938 676320 533940
rect 676047 533882 676052 533938
rect 676108 533882 676320 533938
rect 676047 533880 676320 533882
rect 676047 533877 676113 533880
rect 676674 533203 676734 533392
rect 676674 533198 676785 533203
rect 676674 533142 676724 533198
rect 676780 533142 676785 533198
rect 676674 533140 676785 533142
rect 676719 533137 676785 533140
rect 675130 532990 675136 533054
rect 675200 533052 675206 533054
rect 675200 532992 676320 533052
rect 675200 532990 675206 532992
rect 59535 532904 59601 532907
rect 59535 532902 64416 532904
rect 59535 532846 59540 532902
rect 59596 532846 64416 532902
rect 59535 532844 64416 532846
rect 59535 532841 59601 532844
rect 676090 532694 676096 532758
rect 676160 532756 676166 532758
rect 676160 532696 676350 532756
rect 676160 532694 676166 532696
rect 676290 532430 676350 532696
rect 673978 531806 673984 531870
rect 674048 531868 674054 531870
rect 674048 531808 676320 531868
rect 674048 531806 674054 531808
rect 674362 531510 674368 531574
rect 674432 531572 674438 531574
rect 674432 531512 676320 531572
rect 674432 531510 674438 531512
rect 40954 531362 40960 531426
rect 41024 531424 41030 531426
rect 42831 531424 42897 531427
rect 41024 531422 42897 531424
rect 41024 531366 42836 531422
rect 42892 531366 42897 531422
rect 41024 531364 42897 531366
rect 41024 531362 41030 531364
rect 42831 531361 42897 531364
rect 675322 530918 675328 530982
rect 675392 530980 675398 530982
rect 675392 530920 676320 530980
rect 675392 530918 675398 530920
rect 41967 530686 42033 530687
rect 41914 530622 41920 530686
rect 41984 530684 42033 530686
rect 41984 530682 42076 530684
rect 42028 530626 42076 530682
rect 41984 530624 42076 530626
rect 41984 530622 42033 530624
rect 41967 530621 42033 530622
rect 675514 530326 675520 530390
rect 675584 530388 675590 530390
rect 675584 530328 676320 530388
rect 675584 530326 675590 530328
rect 676047 530018 676113 530021
rect 676047 530016 676320 530018
rect 676047 529960 676052 530016
rect 676108 529960 676320 530016
rect 676047 529958 676320 529960
rect 676047 529955 676113 529958
rect 41775 529650 41841 529651
rect 41722 529648 41728 529650
rect 41684 529588 41728 529648
rect 41792 529646 41841 529650
rect 41836 529590 41841 529646
rect 41722 529586 41728 529588
rect 41792 529586 41841 529590
rect 41775 529585 41841 529586
rect 676239 529648 676305 529651
rect 676239 529646 676350 529648
rect 676239 529590 676244 529646
rect 676300 529590 676350 529646
rect 676239 529585 676350 529590
rect 676290 529470 676350 529585
rect 676047 528908 676113 528911
rect 676047 528906 676320 528908
rect 676047 528850 676052 528906
rect 676108 528850 676320 528906
rect 676047 528848 676320 528850
rect 676047 528845 676113 528848
rect 676047 528464 676113 528467
rect 676047 528462 676320 528464
rect 676047 528406 676052 528462
rect 676108 528406 676320 528462
rect 676047 528404 676320 528406
rect 676047 528401 676113 528404
rect 676239 528168 676305 528171
rect 676239 528166 676350 528168
rect 676239 528110 676244 528166
rect 676300 528110 676350 528166
rect 676239 528105 676350 528110
rect 676290 527990 676350 528105
rect 676047 527428 676113 527431
rect 676047 527426 676320 527428
rect 676047 527370 676052 527426
rect 676108 527370 676320 527426
rect 676047 527368 676320 527370
rect 676047 527365 676113 527368
rect 676047 526984 676113 526987
rect 676047 526982 676320 526984
rect 676047 526926 676052 526982
rect 676108 526926 676320 526982
rect 676047 526924 676320 526926
rect 676047 526921 676113 526924
rect 676239 526688 676305 526691
rect 676239 526686 676350 526688
rect 676239 526630 676244 526686
rect 676300 526630 676350 526686
rect 676239 526625 676350 526630
rect 41146 526478 41152 526542
rect 41216 526540 41222 526542
rect 41775 526540 41841 526543
rect 41216 526538 41841 526540
rect 41216 526482 41780 526538
rect 41836 526482 41841 526538
rect 676290 526510 676350 526625
rect 41216 526480 41841 526482
rect 41216 526478 41222 526480
rect 41775 526477 41841 526480
rect 679791 526096 679857 526099
rect 679746 526094 679857 526096
rect 679746 526038 679796 526094
rect 679852 526038 679857 526094
rect 679746 526033 679857 526038
rect 679746 525918 679806 526033
rect 685506 525211 685566 525474
rect 679791 525208 679857 525211
rect 679746 525206 679857 525208
rect 679746 525150 679796 525206
rect 679852 525150 679857 525206
rect 679746 525145 679857 525150
rect 685455 525206 685566 525211
rect 685455 525150 685460 525206
rect 685516 525150 685566 525206
rect 685455 525148 685566 525150
rect 685455 525145 685521 525148
rect 679746 524956 679806 525145
rect 685455 524764 685521 524767
rect 685455 524762 685566 524764
rect 685455 524706 685460 524762
rect 685516 524706 685566 524762
rect 685455 524701 685566 524706
rect 685506 524438 685566 524701
rect 654447 524320 654513 524323
rect 650208 524318 654513 524320
rect 650208 524262 654452 524318
rect 654508 524262 654513 524318
rect 650208 524260 654513 524262
rect 654447 524257 654513 524260
rect 59535 519732 59601 519735
rect 59535 519730 64416 519732
rect 59535 519674 59540 519730
rect 59596 519674 64416 519730
rect 59535 519672 64416 519674
rect 59535 519669 59601 519672
rect 654447 511000 654513 511003
rect 650208 510998 654513 511000
rect 650208 510942 654452 510998
rect 654508 510942 654513 510998
rect 650208 510940 654513 510942
rect 654447 510937 654513 510940
rect 59535 506708 59601 506711
rect 59535 506706 64416 506708
rect 59535 506650 59540 506706
rect 59596 506650 64416 506706
rect 59535 506648 64416 506650
rect 59535 506645 59601 506648
rect 654447 497680 654513 497683
rect 650208 497678 654513 497680
rect 650208 497622 654452 497678
rect 654508 497622 654513 497678
rect 650208 497620 654513 497622
rect 654447 497617 654513 497620
rect 59535 493684 59601 493687
rect 676239 493684 676305 493687
rect 59535 493682 64416 493684
rect 59535 493626 59540 493682
rect 59596 493626 64416 493682
rect 59535 493624 64416 493626
rect 676239 493682 676350 493684
rect 676239 493626 676244 493682
rect 676300 493626 676350 493682
rect 59535 493621 59601 493624
rect 676239 493621 676350 493626
rect 676290 493506 676350 493621
rect 676047 492944 676113 492947
rect 676047 492942 676320 492944
rect 676047 492886 676052 492942
rect 676108 492886 676320 492942
rect 676047 492884 676320 492886
rect 676047 492881 676113 492884
rect 676047 492352 676113 492355
rect 676047 492350 676320 492352
rect 676047 492294 676052 492350
rect 676108 492294 676320 492350
rect 676047 492292 676320 492294
rect 676047 492289 676113 492292
rect 679695 492204 679761 492207
rect 679695 492202 679806 492204
rect 679695 492146 679700 492202
rect 679756 492146 679806 492202
rect 679695 492141 679806 492146
rect 679746 492026 679806 492141
rect 676527 491612 676593 491615
rect 676482 491610 676593 491612
rect 676482 491554 676532 491610
rect 676588 491554 676593 491610
rect 676482 491549 676593 491554
rect 676482 491434 676542 491549
rect 676623 491168 676689 491171
rect 676623 491166 676734 491168
rect 676623 491110 676628 491166
rect 676684 491110 676734 491166
rect 676623 491105 676734 491110
rect 676674 490842 676734 491105
rect 676674 490283 676734 490472
rect 676623 490278 676734 490283
rect 676623 490222 676628 490278
rect 676684 490222 676734 490278
rect 676623 490220 676734 490222
rect 676623 490217 676689 490220
rect 676719 490132 676785 490135
rect 676674 490130 676785 490132
rect 676674 490074 676724 490130
rect 676780 490074 676785 490130
rect 676674 490069 676785 490074
rect 676674 489954 676734 490069
rect 676674 489247 676734 489362
rect 674546 489182 674552 489246
rect 674616 489244 674622 489246
rect 674616 489184 676350 489244
rect 674616 489182 674622 489184
rect 676290 488992 676350 489184
rect 676623 489242 676734 489247
rect 676623 489186 676628 489242
rect 676684 489186 676734 489242
rect 676623 489184 676734 489186
rect 676623 489181 676689 489184
rect 676143 488652 676209 488655
rect 676143 488650 676350 488652
rect 676143 488594 676148 488650
rect 676204 488594 676350 488650
rect 676143 488592 676350 488594
rect 676143 488589 676209 488592
rect 676290 488474 676350 488592
rect 674354 487850 674360 487914
rect 674424 487912 674430 487914
rect 674424 487852 676320 487912
rect 674424 487850 674430 487852
rect 676047 487468 676113 487471
rect 676047 487466 676320 487468
rect 676047 487410 676052 487466
rect 676108 487410 676320 487466
rect 676047 487408 676320 487410
rect 676047 487405 676113 487408
rect 676239 487172 676305 487175
rect 676239 487170 676350 487172
rect 676239 487114 676244 487170
rect 676300 487114 676350 487170
rect 676239 487109 676350 487114
rect 676290 486994 676350 487109
rect 676239 486580 676305 486583
rect 676239 486578 676350 486580
rect 676239 486522 676244 486578
rect 676300 486522 676350 486578
rect 676239 486517 676350 486522
rect 676290 486402 676350 486517
rect 674738 485926 674744 485990
rect 674808 485988 674814 485990
rect 674808 485928 676320 485988
rect 674808 485926 674814 485928
rect 676047 485470 676113 485473
rect 676047 485468 676320 485470
rect 676047 485412 676052 485468
rect 676108 485412 676320 485468
rect 676047 485410 676320 485412
rect 676047 485407 676113 485410
rect 676239 485100 676305 485103
rect 676239 485098 676350 485100
rect 676239 485042 676244 485098
rect 676300 485042 676350 485098
rect 676239 485037 676350 485042
rect 676290 484922 676350 485037
rect 676047 484508 676113 484511
rect 676047 484506 676320 484508
rect 676047 484450 676052 484506
rect 676108 484450 676320 484506
rect 676047 484448 676320 484450
rect 676047 484445 676113 484448
rect 654447 484360 654513 484363
rect 650208 484358 654513 484360
rect 650208 484302 654452 484358
rect 654508 484302 654513 484358
rect 650208 484300 654513 484302
rect 654447 484297 654513 484300
rect 676047 483990 676113 483993
rect 676047 483988 676320 483990
rect 676047 483932 676052 483988
rect 676108 483932 676320 483988
rect 676047 483930 676320 483932
rect 676047 483927 676113 483930
rect 676858 483706 676864 483770
rect 676928 483706 676934 483770
rect 676866 483442 676926 483706
rect 676047 483028 676113 483031
rect 676047 483026 676320 483028
rect 676047 482970 676052 483026
rect 676108 482970 676320 483026
rect 676047 482968 676320 482970
rect 676047 482965 676113 482968
rect 676047 482436 676113 482439
rect 676047 482434 676320 482436
rect 676047 482378 676052 482434
rect 676108 482378 676320 482434
rect 676047 482376 676320 482378
rect 676047 482373 676113 482376
rect 679938 481699 679998 481962
rect 679938 481694 680049 481699
rect 679938 481638 679988 481694
rect 680044 481638 680049 481694
rect 679938 481636 680049 481638
rect 679983 481633 680049 481636
rect 679746 481255 679806 481518
rect 679746 481250 679857 481255
rect 679983 481252 680049 481255
rect 679746 481194 679796 481250
rect 679852 481194 679857 481250
rect 679746 481192 679857 481194
rect 679791 481189 679857 481192
rect 679938 481250 680049 481252
rect 679938 481194 679988 481250
rect 680044 481194 680049 481250
rect 679938 481189 680049 481194
rect 679938 480926 679998 481189
rect 679791 480808 679857 480811
rect 679746 480806 679857 480808
rect 679746 480750 679796 480806
rect 679852 480750 679857 480806
rect 679746 480745 679857 480750
rect 59535 480660 59601 480663
rect 59535 480658 64416 480660
rect 59535 480602 59540 480658
rect 59596 480602 64416 480658
rect 59535 480600 64416 480602
rect 59535 480597 59601 480600
rect 679746 480408 679806 480745
rect 654447 471188 654513 471191
rect 650208 471186 654513 471188
rect 650208 471130 654452 471186
rect 654508 471130 654513 471186
rect 650208 471128 654513 471130
rect 654447 471125 654513 471128
rect 57807 467488 57873 467491
rect 57807 467486 64416 467488
rect 57807 467430 57812 467486
rect 57868 467430 64416 467486
rect 57807 467428 64416 467430
rect 57807 467425 57873 467428
rect 654447 457868 654513 457871
rect 650208 457866 654513 457868
rect 650208 457810 654452 457866
rect 654508 457810 654513 457866
rect 650208 457808 654513 457810
rect 654447 457805 654513 457808
rect 59535 454612 59601 454615
rect 59535 454610 64416 454612
rect 59535 454554 59540 454610
rect 59596 454554 64416 454610
rect 59535 454552 64416 454554
rect 59535 454549 59601 454552
rect 654447 444548 654513 444551
rect 650208 444546 654513 444548
rect 650208 444490 654452 444546
rect 654508 444490 654513 444546
rect 650208 444488 654513 444490
rect 654447 444485 654513 444488
rect 57807 441588 57873 441591
rect 57807 441586 64416 441588
rect 57807 441530 57812 441586
rect 57868 441530 64416 441586
rect 57807 441528 64416 441530
rect 57807 441525 57873 441528
rect 41775 432264 41841 432267
rect 41568 432262 41841 432264
rect 41568 432206 41780 432262
rect 41836 432206 41841 432262
rect 41568 432204 41841 432206
rect 41775 432201 41841 432204
rect 41775 431746 41841 431749
rect 41568 431744 41841 431746
rect 41568 431688 41780 431744
rect 41836 431688 41841 431744
rect 41568 431686 41841 431688
rect 41775 431683 41841 431686
rect 41583 431376 41649 431379
rect 654447 431376 654513 431379
rect 41538 431374 41649 431376
rect 41538 431318 41588 431374
rect 41644 431318 41649 431374
rect 41538 431313 41649 431318
rect 650208 431374 654513 431376
rect 650208 431318 654452 431374
rect 654508 431318 654513 431374
rect 650208 431316 654513 431318
rect 654447 431313 654513 431316
rect 41538 431198 41598 431313
rect 41775 430784 41841 430787
rect 41568 430782 41841 430784
rect 41568 430726 41780 430782
rect 41836 430726 41841 430782
rect 41568 430724 41841 430726
rect 41775 430721 41841 430724
rect 41775 430266 41841 430269
rect 41568 430264 41841 430266
rect 41568 430208 41780 430264
rect 41836 430208 41841 430264
rect 41568 430206 41841 430208
rect 41775 430203 41841 430206
rect 40570 429834 40576 429898
rect 40640 429896 40646 429898
rect 40719 429896 40785 429899
rect 40640 429894 40785 429896
rect 40640 429838 40724 429894
rect 40780 429838 40785 429894
rect 40640 429836 40785 429838
rect 40640 429834 40646 429836
rect 40719 429833 40785 429836
rect 41722 429748 41728 429750
rect 41568 429688 41728 429748
rect 41722 429686 41728 429688
rect 41792 429686 41798 429750
rect 40770 429011 40830 429274
rect 40719 429006 40830 429011
rect 40719 428950 40724 429006
rect 40780 428950 40830 429006
rect 40719 428948 40830 428950
rect 40719 428945 40785 428948
rect 41538 428567 41598 428682
rect 40762 428502 40768 428566
rect 40832 428502 40838 428566
rect 41538 428562 41649 428567
rect 41538 428506 41588 428562
rect 41644 428506 41649 428562
rect 41538 428504 41649 428506
rect 40770 428238 40830 428502
rect 41583 428501 41649 428504
rect 59535 428564 59601 428567
rect 59535 428562 64416 428564
rect 59535 428506 59540 428562
rect 59596 428506 64416 428562
rect 59535 428504 64416 428506
rect 59535 428501 59601 428504
rect 40770 427530 40830 427794
rect 40762 427466 40768 427530
rect 40832 427466 40838 427530
rect 41914 427232 41920 427234
rect 41568 427172 41920 427232
rect 41914 427170 41920 427172
rect 41984 427170 41990 427234
rect 41538 426492 41598 426684
rect 42298 426492 42304 426494
rect 41538 426432 42304 426492
rect 42298 426430 42304 426432
rect 42368 426430 42374 426494
rect 40962 426050 41022 426314
rect 40954 425986 40960 426050
rect 41024 425986 41030 426050
rect 40386 425458 40446 425722
rect 40378 425394 40384 425458
rect 40448 425394 40454 425458
rect 41871 425234 41937 425237
rect 41568 425232 41937 425234
rect 41568 425176 41876 425232
rect 41932 425176 41937 425232
rect 41568 425174 41937 425176
rect 41871 425171 41937 425174
rect 41154 424570 41214 424834
rect 41146 424506 41152 424570
rect 41216 424506 41222 424570
rect 41346 423978 41406 424242
rect 41338 423914 41344 423978
rect 41408 423914 41414 423978
rect 41538 423534 41598 423650
rect 41530 423470 41536 423534
rect 41600 423470 41606 423534
rect 41775 423310 41841 423313
rect 41568 423308 41841 423310
rect 41568 423252 41780 423308
rect 41836 423252 41841 423308
rect 41568 423250 41841 423252
rect 41775 423247 41841 423250
rect 41967 422792 42033 422795
rect 41568 422790 42033 422792
rect 41568 422734 41972 422790
rect 42028 422734 42033 422790
rect 41568 422732 42033 422734
rect 41967 422729 42033 422732
rect 40578 422054 40638 422170
rect 40570 421990 40576 422054
rect 40640 421990 40646 422054
rect 41538 421611 41598 421800
rect 41538 421606 41649 421611
rect 41538 421550 41588 421606
rect 41644 421550 41649 421606
rect 41538 421548 41649 421550
rect 41583 421545 41649 421548
rect 41538 421019 41598 421282
rect 41538 421014 41649 421019
rect 41538 420958 41588 421014
rect 41644 420958 41649 421014
rect 41538 420956 41649 420958
rect 41583 420953 41649 420956
rect 41538 420572 41598 420690
rect 41538 420512 41790 420572
rect 28866 419983 28926 420246
rect 41730 420128 41790 420512
rect 28815 419978 28926 419983
rect 28815 419922 28820 419978
rect 28876 419922 28926 419978
rect 28815 419920 28926 419922
rect 41538 420068 41790 420128
rect 28815 419917 28881 419920
rect 41538 419832 41598 420068
rect 41775 419832 41841 419835
rect 41538 419830 41841 419832
rect 41538 419802 41780 419830
rect 41568 419774 41780 419802
rect 41836 419774 41841 419830
rect 41568 419772 41841 419774
rect 41775 419769 41841 419772
rect 28815 419536 28881 419539
rect 28815 419534 28926 419536
rect 28815 419478 28820 419534
rect 28876 419478 28926 419534
rect 28815 419473 28926 419478
rect 28866 419210 28926 419473
rect 654447 418056 654513 418059
rect 650208 418054 654513 418056
rect 650208 417998 654452 418054
rect 654508 417998 654513 418054
rect 650208 417996 654513 417998
rect 654447 417993 654513 417996
rect 59535 415392 59601 415395
rect 59535 415390 64416 415392
rect 59535 415334 59540 415390
rect 59596 415334 64416 415390
rect 59535 415332 64416 415334
rect 59535 415329 59601 415332
rect 41967 411250 42033 411251
rect 41914 411248 41920 411250
rect 41876 411188 41920 411248
rect 41984 411246 42033 411250
rect 42028 411190 42033 411246
rect 41914 411186 41920 411188
rect 41984 411186 42033 411190
rect 41967 411185 42033 411186
rect 40378 406006 40384 406070
rect 40448 406068 40454 406070
rect 41775 406068 41841 406071
rect 40448 406066 41841 406068
rect 40448 406010 41780 406066
rect 41836 406010 41841 406066
rect 40448 406008 41841 406010
rect 40448 406006 40454 406008
rect 41775 406005 41841 406008
rect 676239 405476 676305 405479
rect 676239 405474 676350 405476
rect 676239 405418 676244 405474
rect 676300 405418 676350 405474
rect 676239 405413 676350 405418
rect 676290 405298 676350 405413
rect 654447 404736 654513 404739
rect 650208 404734 654513 404736
rect 650208 404678 654452 404734
rect 654508 404678 654513 404734
rect 650208 404676 654513 404678
rect 654447 404673 654513 404676
rect 676047 404736 676113 404739
rect 676047 404734 676320 404736
rect 676047 404678 676052 404734
rect 676108 404678 676320 404734
rect 676047 404676 676320 404678
rect 676047 404673 676113 404676
rect 676047 404218 676113 404221
rect 676047 404216 676320 404218
rect 676047 404160 676052 404216
rect 676108 404160 676320 404216
rect 676047 404158 676320 404160
rect 676047 404155 676113 404158
rect 676527 403996 676593 403999
rect 676482 403994 676593 403996
rect 676482 403938 676532 403994
rect 676588 403938 676593 403994
rect 676482 403933 676593 403938
rect 40570 403786 40576 403850
rect 40640 403848 40646 403850
rect 41775 403848 41841 403851
rect 40640 403846 41841 403848
rect 40640 403790 41780 403846
rect 41836 403790 41841 403846
rect 676482 403818 676542 403933
rect 40640 403788 41841 403790
rect 40640 403786 40646 403788
rect 41775 403785 41841 403788
rect 676047 403256 676113 403259
rect 676047 403254 676320 403256
rect 676047 403198 676052 403254
rect 676108 403198 676320 403254
rect 676047 403196 676320 403198
rect 676047 403193 676113 403196
rect 41530 403046 41536 403110
rect 41600 403108 41606 403110
rect 41775 403108 41841 403111
rect 41600 403106 41841 403108
rect 41600 403050 41780 403106
rect 41836 403050 41841 403106
rect 41600 403048 41841 403050
rect 41600 403046 41606 403048
rect 41775 403045 41841 403048
rect 676719 402960 676785 402963
rect 676674 402958 676785 402960
rect 676674 402902 676724 402958
rect 676780 402902 676785 402958
rect 676674 402897 676785 402902
rect 676674 402634 676734 402897
rect 41338 402454 41344 402518
rect 41408 402516 41414 402518
rect 41775 402516 41841 402519
rect 41408 402514 41841 402516
rect 41408 402458 41780 402514
rect 41836 402458 41841 402514
rect 41408 402456 41841 402458
rect 41408 402454 41414 402456
rect 41775 402453 41841 402456
rect 59535 402368 59601 402371
rect 59535 402366 64416 402368
rect 59535 402310 59540 402366
rect 59596 402310 64416 402366
rect 59535 402308 64416 402310
rect 59535 402305 59601 402308
rect 676047 402294 676113 402297
rect 676047 402292 676320 402294
rect 676047 402236 676052 402292
rect 676108 402236 676320 402292
rect 676047 402234 676320 402236
rect 676047 402231 676113 402234
rect 40954 401862 40960 401926
rect 41024 401924 41030 401926
rect 41775 401924 41841 401927
rect 41024 401922 41841 401924
rect 41024 401866 41780 401922
rect 41836 401866 41841 401922
rect 41024 401864 41841 401866
rect 41024 401862 41030 401864
rect 41775 401861 41841 401864
rect 676047 401776 676113 401779
rect 676047 401774 676320 401776
rect 676047 401718 676052 401774
rect 676108 401718 676320 401774
rect 676047 401716 676320 401718
rect 676047 401713 676113 401716
rect 676290 401039 676350 401154
rect 676239 401034 676350 401039
rect 676239 400978 676244 401034
rect 676300 400978 676350 401034
rect 676239 400976 676350 400978
rect 676239 400973 676305 400976
rect 676674 400446 676734 400784
rect 676666 400382 676672 400446
rect 676736 400382 676742 400446
rect 674170 400234 674176 400298
rect 674240 400296 674246 400298
rect 674240 400236 676320 400296
rect 674240 400234 674246 400236
rect 40762 399938 40768 400002
rect 40832 400000 40838 400002
rect 41775 400000 41841 400003
rect 40832 399998 41841 400000
rect 40832 399942 41780 399998
rect 41836 399942 41841 399998
rect 40832 399940 41841 399942
rect 40832 399938 40838 399940
rect 41775 399937 41841 399940
rect 41146 399494 41152 399558
rect 41216 399556 41222 399558
rect 41775 399556 41841 399559
rect 676482 399558 676542 399674
rect 41216 399554 41841 399556
rect 41216 399498 41780 399554
rect 41836 399498 41841 399554
rect 41216 399496 41841 399498
rect 41216 399494 41222 399496
rect 41775 399493 41841 399496
rect 676474 399494 676480 399558
rect 676544 399494 676550 399558
rect 674938 399198 674944 399262
rect 675008 399260 675014 399262
rect 675008 399200 676320 399260
rect 675008 399198 675014 399200
rect 41871 398966 41937 398967
rect 41871 398962 41920 398966
rect 41984 398964 41990 398966
rect 41871 398906 41876 398962
rect 41871 398902 41920 398906
rect 41984 398904 42028 398964
rect 41984 398902 41990 398904
rect 41871 398901 41937 398902
rect 674362 398754 674368 398818
rect 674432 398816 674438 398818
rect 674432 398756 676320 398816
rect 674432 398754 674438 398756
rect 675514 398162 675520 398226
rect 675584 398224 675590 398226
rect 675584 398164 676320 398224
rect 675584 398162 675590 398164
rect 675898 397718 675904 397782
rect 675968 397780 675974 397782
rect 675968 397720 676320 397780
rect 675968 397718 675974 397720
rect 675322 396830 675328 396894
rect 675392 396892 675398 396894
rect 676290 396892 676350 397232
rect 675392 396832 676350 396892
rect 675392 396830 675398 396832
rect 675130 396682 675136 396746
rect 675200 396744 675206 396746
rect 675200 396684 676320 396744
rect 675200 396682 675206 396684
rect 676090 395942 676096 396006
rect 676160 396004 676166 396006
rect 676290 396004 676350 396270
rect 676160 395944 676350 396004
rect 676160 395942 676166 395944
rect 676047 395782 676113 395785
rect 676047 395780 676320 395782
rect 676047 395724 676052 395780
rect 676108 395724 676320 395780
rect 676047 395722 676320 395724
rect 676047 395719 676113 395722
rect 675706 395202 675712 395266
rect 675776 395264 675782 395266
rect 675776 395204 676320 395264
rect 675776 395202 675782 395204
rect 676290 394674 676350 394790
rect 676282 394610 676288 394674
rect 676352 394610 676358 394674
rect 676290 394083 676350 394198
rect 676239 394078 676350 394083
rect 676239 394022 676244 394078
rect 676300 394022 676350 394078
rect 676239 394020 676350 394022
rect 676239 394017 676305 394020
rect 679746 393491 679806 393754
rect 679746 393486 679857 393491
rect 679746 393430 679796 393486
rect 679852 393430 679857 393486
rect 679746 393428 679857 393430
rect 679791 393425 679857 393428
rect 685506 393047 685566 393310
rect 679791 393044 679857 393047
rect 679746 393042 679857 393044
rect 679746 392986 679796 393042
rect 679852 392986 679857 393042
rect 679746 392981 679857 392986
rect 685506 393042 685617 393047
rect 685506 392986 685556 393042
rect 685612 392986 685617 393042
rect 685506 392984 685617 392986
rect 685551 392981 685617 392984
rect 679746 392718 679806 392981
rect 685551 392600 685617 392603
rect 685506 392598 685617 392600
rect 685506 392542 685556 392598
rect 685612 392542 685617 392598
rect 685506 392537 685617 392542
rect 685506 392200 685566 392537
rect 654831 391564 654897 391567
rect 650208 391562 654897 391564
rect 650208 391506 654836 391562
rect 654892 391506 654897 391562
rect 650208 391504 654897 391506
rect 654831 391501 654897 391504
rect 41122 390902 41128 390966
rect 41192 390964 41198 390966
rect 41871 390964 41937 390967
rect 41192 390962 41937 390964
rect 41192 390906 41876 390962
rect 41932 390906 41937 390962
rect 41192 390904 41937 390906
rect 41192 390902 41198 390904
rect 41871 390901 41937 390904
rect 41871 389344 41937 389347
rect 59535 389344 59601 389347
rect 41871 389342 54750 389344
rect 41871 389286 41876 389342
rect 41932 389286 54750 389342
rect 41871 389284 54750 389286
rect 41871 389281 41937 389284
rect 54690 389196 54750 389284
rect 59535 389342 64416 389344
rect 59535 389286 59540 389342
rect 59596 389286 64416 389342
rect 59535 389284 64416 389286
rect 59535 389281 59601 389284
rect 62223 389196 62289 389199
rect 54690 389194 62289 389196
rect 54690 389138 62228 389194
rect 62284 389138 62289 389194
rect 54690 389136 62289 389138
rect 62223 389133 62289 389136
rect 41775 389048 41841 389051
rect 41568 389046 41841 389048
rect 41568 388990 41780 389046
rect 41836 388990 41841 389046
rect 41568 388988 41841 388990
rect 41775 388985 41841 388988
rect 41583 388752 41649 388755
rect 41538 388750 41649 388752
rect 41538 388694 41588 388750
rect 41644 388694 41649 388750
rect 41538 388689 41649 388694
rect 41538 388574 41598 388689
rect 41775 388012 41841 388015
rect 41568 388010 41841 388012
rect 41568 387954 41780 388010
rect 41836 387954 41841 388010
rect 41568 387952 41841 387954
rect 41775 387949 41841 387952
rect 41775 387568 41841 387571
rect 41568 387566 41841 387568
rect 41568 387510 41780 387566
rect 41836 387510 41841 387566
rect 41568 387508 41841 387510
rect 41775 387505 41841 387508
rect 41775 387050 41841 387053
rect 41568 387048 41841 387050
rect 41568 386992 41780 387048
rect 41836 386992 41841 387048
rect 41568 386990 41841 386992
rect 41775 386987 41841 386990
rect 41722 386532 41728 386534
rect 41568 386472 41728 386532
rect 41722 386470 41728 386472
rect 41792 386470 41798 386534
rect 41871 386088 41937 386091
rect 41568 386086 41937 386088
rect 41568 386030 41876 386086
rect 41932 386030 41937 386086
rect 41568 386028 41937 386030
rect 41871 386025 41937 386028
rect 675759 385940 675825 385943
rect 676474 385940 676480 385942
rect 675759 385938 676480 385940
rect 675759 385882 675764 385938
rect 675820 385882 676480 385938
rect 675759 385880 676480 385882
rect 675759 385877 675825 385880
rect 676474 385878 676480 385880
rect 676544 385878 676550 385942
rect 675759 385644 675825 385647
rect 675898 385644 675904 385646
rect 675759 385642 675904 385644
rect 675759 385586 675764 385642
rect 675820 385586 675904 385642
rect 675759 385584 675904 385586
rect 675759 385581 675825 385584
rect 675898 385582 675904 385584
rect 675968 385582 675974 385646
rect 34434 385203 34494 385540
rect 34434 385198 34545 385203
rect 41583 385200 41649 385203
rect 34434 385142 34484 385198
rect 34540 385142 34545 385198
rect 34434 385140 34545 385142
rect 34479 385137 34545 385140
rect 41538 385198 41649 385200
rect 41538 385142 41588 385198
rect 41644 385142 41649 385198
rect 41538 385137 41649 385142
rect 41538 385022 41598 385137
rect 675759 384756 675825 384759
rect 676666 384756 676672 384758
rect 675759 384754 676672 384756
rect 675759 384698 675764 384754
rect 675820 384698 676672 384754
rect 675759 384696 676672 384698
rect 675759 384693 675825 384696
rect 676666 384694 676672 384696
rect 676736 384694 676742 384758
rect 40770 384314 40830 384578
rect 41722 384398 41728 384462
rect 41792 384460 41798 384462
rect 61935 384460 62001 384463
rect 41792 384458 62001 384460
rect 41792 384402 61940 384458
rect 61996 384402 62001 384458
rect 41792 384400 62001 384402
rect 41792 384398 41798 384400
rect 61935 384397 62001 384400
rect 40762 384250 40768 384314
rect 40832 384250 40838 384314
rect 41914 384016 41920 384018
rect 41568 383956 41920 384016
rect 41914 383954 41920 383956
rect 41984 383954 41990 384018
rect 40962 383278 41022 383542
rect 40954 383214 40960 383278
rect 41024 383214 41030 383278
rect 41346 382834 41406 383098
rect 674938 382918 674944 382982
rect 675008 382980 675014 382982
rect 675375 382980 675441 382983
rect 675008 382978 675441 382980
rect 675008 382922 675380 382978
rect 675436 382922 675441 382978
rect 675008 382920 675441 382922
rect 675008 382918 675014 382920
rect 675375 382917 675441 382920
rect 41338 382770 41344 382834
rect 41408 382770 41414 382834
rect 675130 382770 675136 382834
rect 675200 382832 675206 382834
rect 675279 382832 675345 382835
rect 675200 382830 675345 382832
rect 675200 382774 675284 382830
rect 675340 382774 675345 382830
rect 675200 382772 675345 382774
rect 675200 382770 675206 382772
rect 675279 382769 675345 382772
rect 40386 382242 40446 382506
rect 40378 382178 40384 382242
rect 40448 382178 40454 382242
rect 675322 382178 675328 382242
rect 675392 382240 675398 382242
rect 675471 382240 675537 382243
rect 675392 382238 675537 382240
rect 675392 382182 675476 382238
rect 675532 382182 675537 382238
rect 675392 382180 675537 382182
rect 675392 382178 675398 382180
rect 675471 382177 675537 382180
rect 41871 382018 41937 382021
rect 41568 382016 41937 382018
rect 41568 381960 41876 382016
rect 41932 381960 41937 382016
rect 41568 381958 41937 381960
rect 41871 381955 41937 381958
rect 41154 381354 41214 381618
rect 41146 381290 41152 381354
rect 41216 381290 41222 381354
rect 675759 381206 675825 381207
rect 675706 381142 675712 381206
rect 675776 381204 675825 381206
rect 675776 381202 675868 381204
rect 675820 381146 675868 381202
rect 675776 381144 675868 381146
rect 675776 381142 675825 381144
rect 675759 381141 675825 381142
rect 41722 381056 41728 381058
rect 41568 380996 41728 381056
rect 41722 380994 41728 380996
rect 41792 380994 41798 381058
rect 41538 380318 41598 380508
rect 41530 380254 41536 380318
rect 41600 380254 41606 380318
rect 41775 380168 41841 380171
rect 41568 380166 41841 380168
rect 41568 380110 41780 380166
rect 41836 380110 41841 380166
rect 41568 380108 41841 380110
rect 41775 380105 41841 380108
rect 41775 379576 41841 379579
rect 41568 379574 41841 379576
rect 41568 379518 41780 379574
rect 41836 379518 41841 379574
rect 41568 379516 41841 379518
rect 41775 379513 41841 379516
rect 41538 378839 41598 378954
rect 41538 378834 41649 378839
rect 41538 378778 41588 378834
rect 41644 378778 41649 378834
rect 41538 378776 41649 378778
rect 41583 378773 41649 378776
rect 674362 378774 674368 378838
rect 674432 378836 674438 378838
rect 675471 378836 675537 378839
rect 674432 378834 675537 378836
rect 674432 378778 675476 378834
rect 675532 378778 675537 378834
rect 674432 378776 675537 378778
rect 674432 378774 674438 378776
rect 675471 378773 675537 378776
rect 41538 378395 41598 378584
rect 41538 378390 41649 378395
rect 41538 378334 41588 378390
rect 41644 378334 41649 378390
rect 41538 378332 41649 378334
rect 41583 378329 41649 378332
rect 654447 378244 654513 378247
rect 650208 378242 654513 378244
rect 650208 378186 654452 378242
rect 654508 378186 654513 378242
rect 650208 378184 654513 378186
rect 654447 378181 654513 378184
rect 41775 378096 41841 378099
rect 41568 378094 41841 378096
rect 41568 378038 41780 378094
rect 41836 378038 41841 378094
rect 41568 378036 41841 378038
rect 41775 378033 41841 378036
rect 675759 377948 675825 377951
rect 676282 377948 676288 377950
rect 675759 377946 676288 377948
rect 675759 377890 675764 377946
rect 675820 377890 676288 377946
rect 675759 377888 676288 377890
rect 675759 377885 675825 377888
rect 676282 377886 676288 377888
rect 676352 377886 676358 377950
rect 40194 377359 40254 377474
rect 40194 377354 40305 377359
rect 40194 377298 40244 377354
rect 40300 377298 40305 377354
rect 40194 377296 40305 377298
rect 40239 377293 40305 377296
rect 28866 376767 28926 377104
rect 28815 376762 28926 376767
rect 28815 376706 28820 376762
rect 28876 376706 28926 376762
rect 28815 376704 28926 376706
rect 28815 376701 28881 376704
rect 41775 376616 41841 376619
rect 41568 376614 41841 376616
rect 41568 376558 41780 376614
rect 41836 376558 41841 376614
rect 41568 376556 41841 376558
rect 41775 376553 41841 376556
rect 28815 376320 28881 376323
rect 59439 376320 59505 376323
rect 28815 376318 28926 376320
rect 28815 376262 28820 376318
rect 28876 376262 28926 376318
rect 28815 376257 28926 376262
rect 59439 376318 64416 376320
rect 59439 376262 59444 376318
rect 59500 376262 64416 376318
rect 59439 376260 64416 376262
rect 59439 376257 59505 376260
rect 28866 375994 28926 376257
rect 675759 375728 675825 375731
rect 676090 375728 676096 375730
rect 675759 375726 676096 375728
rect 675759 375670 675764 375726
rect 675820 375670 676096 375726
rect 675759 375668 676096 375670
rect 675759 375665 675825 375668
rect 676090 375666 676096 375668
rect 676160 375666 676166 375730
rect 674170 373742 674176 373806
rect 674240 373804 674246 373806
rect 675183 373804 675249 373807
rect 674240 373802 675249 373804
rect 674240 373746 675188 373802
rect 675244 373746 675249 373802
rect 674240 373744 675249 373746
rect 674240 373742 674246 373744
rect 675183 373741 675249 373744
rect 675567 372030 675633 372031
rect 675514 372028 675520 372030
rect 675476 371968 675520 372028
rect 675584 372026 675633 372030
rect 675628 371970 675633 372026
rect 675514 371966 675520 371968
rect 675584 371966 675633 371970
rect 675567 371965 675633 371966
rect 41967 368182 42033 368183
rect 41914 368180 41920 368182
rect 41876 368120 41920 368180
rect 41984 368178 42033 368182
rect 42028 368122 42033 368178
rect 41914 368118 41920 368120
rect 41984 368118 42033 368122
rect 41967 368117 42033 368118
rect 654447 364924 654513 364927
rect 650208 364922 654513 364924
rect 650208 364866 654452 364922
rect 654508 364866 654513 364922
rect 650208 364864 654513 364866
rect 654447 364861 654513 364864
rect 58383 363296 58449 363299
rect 58383 363294 64416 363296
rect 58383 363238 58388 363294
rect 58444 363238 64416 363294
rect 58383 363236 64416 363238
rect 58383 363233 58449 363236
rect 40378 362790 40384 362854
rect 40448 362852 40454 362854
rect 41775 362852 41841 362855
rect 40448 362850 41841 362852
rect 40448 362794 41780 362850
rect 41836 362794 41841 362850
rect 40448 362792 41841 362794
rect 40448 362790 40454 362792
rect 41775 362789 41841 362792
rect 676047 360040 676113 360043
rect 676047 360038 676320 360040
rect 676047 359982 676052 360038
rect 676108 359982 676320 360038
rect 676047 359980 676320 359982
rect 676047 359977 676113 359980
rect 41530 359830 41536 359894
rect 41600 359892 41606 359894
rect 41775 359892 41841 359895
rect 41600 359890 41841 359892
rect 41600 359834 41780 359890
rect 41836 359834 41841 359890
rect 41600 359832 41841 359834
rect 41600 359830 41606 359832
rect 41775 359829 41841 359832
rect 676239 359744 676305 359747
rect 676239 359742 676350 359744
rect 676239 359686 676244 359742
rect 676300 359686 676350 359742
rect 676239 359681 676350 359686
rect 676290 359566 676350 359681
rect 41775 359450 41841 359451
rect 41722 359448 41728 359450
rect 41684 359388 41728 359448
rect 41792 359446 41841 359450
rect 41836 359390 41841 359446
rect 41722 359386 41728 359388
rect 41792 359386 41841 359390
rect 41775 359385 41841 359386
rect 676047 359004 676113 359007
rect 676047 359002 676320 359004
rect 676047 358946 676052 359002
rect 676108 358946 676320 359002
rect 676047 358944 676320 358946
rect 676047 358941 676113 358944
rect 41338 358646 41344 358710
rect 41408 358708 41414 358710
rect 41775 358708 41841 358711
rect 41408 358706 41841 358708
rect 41408 358650 41780 358706
rect 41836 358650 41841 358706
rect 41408 358648 41841 358650
rect 41408 358646 41414 358648
rect 41775 358645 41841 358648
rect 676047 358560 676113 358563
rect 676047 358558 676320 358560
rect 676047 358502 676052 358558
rect 676108 358502 676320 358558
rect 676047 358500 676320 358502
rect 676047 358497 676113 358500
rect 673978 358054 673984 358118
rect 674048 358116 674054 358118
rect 674048 358056 676320 358116
rect 674048 358054 674054 358056
rect 676239 357672 676305 357675
rect 676239 357670 676350 357672
rect 676239 357614 676244 357670
rect 676300 357614 676350 357670
rect 676239 357609 676350 357614
rect 676290 357494 676350 357609
rect 669807 357080 669873 357083
rect 674170 357080 674176 357082
rect 669807 357078 674176 357080
rect 669807 357022 669812 357078
rect 669868 357022 674176 357078
rect 669807 357020 674176 357022
rect 669807 357017 669873 357020
rect 674170 357018 674176 357020
rect 674240 357080 674246 357082
rect 674240 357020 676320 357080
rect 674240 357018 674246 357020
rect 40762 356870 40768 356934
rect 40832 356932 40838 356934
rect 41775 356932 41841 356935
rect 40832 356930 41841 356932
rect 40832 356874 41780 356930
rect 41836 356874 41841 356930
rect 40832 356872 41841 356874
rect 40832 356870 40838 356872
rect 41775 356869 41841 356872
rect 676047 356562 676113 356565
rect 676047 356560 676320 356562
rect 676047 356504 676052 356560
rect 676108 356504 676320 356560
rect 676047 356502 676320 356504
rect 676047 356499 676113 356502
rect 41146 356426 41152 356490
rect 41216 356488 41222 356490
rect 41775 356488 41841 356491
rect 41216 356486 41841 356488
rect 41216 356430 41780 356486
rect 41836 356430 41841 356486
rect 41216 356428 41841 356430
rect 41216 356426 41222 356428
rect 41775 356425 41841 356428
rect 669615 356192 669681 356195
rect 676090 356192 676096 356194
rect 669615 356190 676096 356192
rect 669615 356134 669620 356190
rect 669676 356134 676096 356190
rect 669615 356132 676096 356134
rect 669615 356129 669681 356132
rect 676090 356130 676096 356132
rect 676160 356192 676166 356194
rect 676160 356132 676350 356192
rect 676160 356130 676166 356132
rect 676290 356014 676350 356132
rect 40954 355538 40960 355602
rect 41024 355600 41030 355602
rect 41775 355600 41841 355603
rect 41024 355598 41841 355600
rect 41024 355542 41780 355598
rect 41836 355542 41841 355598
rect 41024 355540 41841 355542
rect 41024 355538 41030 355540
rect 41775 355537 41841 355540
rect 675898 355538 675904 355602
rect 675968 355600 675974 355602
rect 675968 355540 676320 355600
rect 675968 355538 675974 355540
rect 674554 354946 674560 355010
rect 674624 355008 674630 355010
rect 674624 354948 676320 355008
rect 674624 354946 674630 354948
rect 675759 354564 675825 354567
rect 675759 354562 676320 354564
rect 675759 354506 675764 354562
rect 675820 354506 676320 354562
rect 675759 354504 676320 354506
rect 675759 354501 675825 354504
rect 676047 354120 676113 354123
rect 676047 354118 676320 354120
rect 676047 354062 676052 354118
rect 676108 354062 676320 354118
rect 676047 354060 676320 354062
rect 676047 354057 676113 354060
rect 674938 353466 674944 353530
rect 675008 353528 675014 353530
rect 675008 353468 676320 353528
rect 675008 353466 675014 353468
rect 674746 353022 674752 353086
rect 674816 353084 674822 353086
rect 674816 353024 676320 353084
rect 674816 353022 674822 353024
rect 675279 352640 675345 352643
rect 675279 352638 676320 352640
rect 675279 352582 675284 352638
rect 675340 352582 676320 352638
rect 675279 352580 676320 352582
rect 675279 352577 675345 352580
rect 675514 351986 675520 352050
rect 675584 352048 675590 352050
rect 675584 351988 676320 352048
rect 675584 351986 675590 351988
rect 654447 351604 654513 351607
rect 650208 351602 654513 351604
rect 650208 351546 654452 351602
rect 654508 351546 654513 351602
rect 650208 351544 654513 351546
rect 654447 351541 654513 351544
rect 675706 351468 675712 351532
rect 675776 351530 675782 351532
rect 675776 351470 676320 351530
rect 675776 351468 675782 351470
rect 675130 351098 675136 351162
rect 675200 351160 675206 351162
rect 675200 351100 676320 351160
rect 675200 351098 675206 351100
rect 676290 350423 676350 350538
rect 676239 350418 676350 350423
rect 676239 350362 676244 350418
rect 676300 350362 676350 350418
rect 676239 350360 676350 350362
rect 676239 350357 676305 350360
rect 59535 350272 59601 350275
rect 59535 350270 64416 350272
rect 59535 350214 59540 350270
rect 59596 350214 64416 350270
rect 59535 350212 64416 350214
rect 59535 350209 59601 350212
rect 676290 349831 676350 349946
rect 676239 349826 676350 349831
rect 676239 349770 676244 349826
rect 676300 349770 676350 349826
rect 676239 349768 676350 349770
rect 676239 349765 676305 349768
rect 676047 349680 676113 349683
rect 676047 349678 676320 349680
rect 676047 349622 676052 349678
rect 676108 349622 676320 349678
rect 676047 349620 676320 349622
rect 676047 349617 676113 349620
rect 676047 349088 676113 349091
rect 676047 349086 676320 349088
rect 676047 349030 676052 349086
rect 676108 349030 676320 349086
rect 676047 349028 676320 349030
rect 676047 349025 676113 349028
rect 679746 348351 679806 348466
rect 679746 348346 679857 348351
rect 679746 348290 679796 348346
rect 679852 348290 679857 348346
rect 679746 348288 679857 348290
rect 679791 348285 679857 348288
rect 685506 347759 685566 348096
rect 679791 347756 679857 347759
rect 679746 347754 679857 347756
rect 679746 347698 679796 347754
rect 679852 347698 679857 347754
rect 679746 347693 679857 347698
rect 685455 347754 685566 347759
rect 685455 347698 685460 347754
rect 685516 347698 685566 347754
rect 685455 347696 685566 347698
rect 685455 347693 685521 347696
rect 679746 347578 679806 347693
rect 685455 347312 685521 347315
rect 685455 347310 685566 347312
rect 685455 347254 685460 347310
rect 685516 347254 685566 347310
rect 685455 347249 685566 347254
rect 685506 346986 685566 347249
rect 41775 345906 41841 345909
rect 41568 345904 41841 345906
rect 41568 345848 41780 345904
rect 41836 345848 41841 345904
rect 41568 345846 41841 345848
rect 41775 345843 41841 345846
rect 41583 345536 41649 345539
rect 41538 345534 41649 345536
rect 41538 345478 41588 345534
rect 41644 345478 41649 345534
rect 41538 345473 41649 345478
rect 41538 345358 41598 345473
rect 41775 344796 41841 344799
rect 41568 344794 41841 344796
rect 41568 344738 41780 344794
rect 41836 344738 41841 344794
rect 41568 344736 41841 344738
rect 41775 344733 41841 344736
rect 41775 344352 41841 344355
rect 41568 344350 41841 344352
rect 41568 344294 41780 344350
rect 41836 344294 41841 344350
rect 41568 344292 41841 344294
rect 41775 344289 41841 344292
rect 41775 343908 41841 343911
rect 41568 343906 41841 343908
rect 41568 343850 41780 343906
rect 41836 343850 41841 343906
rect 41568 343848 41841 343850
rect 41775 343845 41841 343848
rect 41775 343316 41841 343319
rect 41568 343314 41841 343316
rect 41568 343258 41780 343314
rect 41836 343258 41841 343314
rect 41568 343256 41841 343258
rect 41775 343253 41841 343256
rect 40578 342726 40638 342842
rect 40570 342662 40576 342726
rect 40640 342662 40646 342726
rect 41775 342354 41841 342357
rect 41568 342352 41841 342354
rect 41568 342296 41780 342352
rect 41836 342296 41841 342352
rect 41568 342294 41841 342296
rect 41775 342291 41841 342294
rect 41583 341984 41649 341987
rect 41538 341982 41649 341984
rect 41538 341926 41588 341982
rect 41644 341926 41649 341982
rect 41538 341921 41649 341926
rect 41538 341806 41598 341921
rect 40770 341098 40830 341362
rect 40762 341034 40768 341098
rect 40832 341034 40838 341098
rect 41722 340874 41728 340876
rect 41568 340814 41728 340874
rect 41722 340812 41728 340814
rect 41792 340812 41798 340876
rect 40570 340442 40576 340506
rect 40640 340442 40646 340506
rect 40578 340326 40638 340442
rect 41154 339618 41214 339882
rect 41146 339554 41152 339618
rect 41216 339554 41222 339618
rect 675759 339616 675825 339619
rect 675898 339616 675904 339618
rect 675759 339614 675904 339616
rect 675759 339558 675764 339614
rect 675820 339558 675904 339614
rect 675759 339556 675904 339558
rect 675759 339553 675825 339556
rect 675898 339554 675904 339556
rect 675968 339554 675974 339618
rect 40386 339026 40446 339290
rect 40378 338962 40384 339026
rect 40448 338962 40454 339026
rect 41871 338876 41937 338879
rect 41568 338874 41937 338876
rect 41568 338818 41876 338874
rect 41932 338818 41937 338874
rect 41568 338816 41937 338818
rect 41871 338813 41937 338816
rect 40962 338138 41022 338402
rect 655311 338284 655377 338287
rect 650208 338282 655377 338284
rect 650208 338226 655316 338282
rect 655372 338226 655377 338282
rect 650208 338224 655377 338226
rect 655311 338221 655377 338224
rect 40954 338074 40960 338138
rect 41024 338074 41030 338138
rect 41346 337546 41406 337810
rect 41338 337482 41344 337546
rect 41408 337482 41414 337546
rect 41538 337102 41598 337292
rect 59535 337248 59601 337251
rect 59535 337246 64416 337248
rect 59535 337190 59540 337246
rect 59596 337190 64416 337246
rect 59535 337188 64416 337190
rect 59535 337185 59601 337188
rect 675471 337102 675537 337103
rect 41530 337038 41536 337102
rect 41600 337038 41606 337102
rect 675471 337100 675520 337102
rect 675428 337098 675520 337100
rect 675428 337042 675476 337098
rect 675428 337040 675520 337042
rect 675471 337038 675520 337040
rect 675584 337038 675590 337102
rect 675471 337037 675537 337038
rect 41775 336952 41841 336955
rect 41568 336950 41841 336952
rect 41568 336894 41780 336950
rect 41836 336894 41841 336950
rect 41568 336892 41841 336894
rect 41775 336889 41841 336892
rect 675759 336510 675825 336511
rect 675706 336508 675712 336510
rect 675668 336448 675712 336508
rect 675776 336506 675825 336510
rect 675820 336450 675825 336506
rect 675706 336446 675712 336448
rect 675776 336446 675825 336450
rect 675759 336445 675825 336446
rect 41538 336215 41598 336330
rect 41538 336210 41649 336215
rect 41538 336154 41588 336210
rect 41644 336154 41649 336210
rect 41538 336152 41649 336154
rect 41583 336149 41649 336152
rect 41538 335768 41598 335812
rect 42447 335768 42513 335771
rect 41538 335766 42513 335768
rect 41538 335710 42452 335766
rect 42508 335710 42513 335766
rect 41538 335708 42513 335710
rect 42447 335705 42513 335708
rect 41538 335179 41598 335442
rect 41538 335174 41649 335179
rect 41538 335118 41588 335174
rect 41644 335118 41649 335174
rect 41538 335116 41649 335118
rect 41583 335113 41649 335116
rect 41775 334880 41841 334883
rect 41568 334878 41841 334880
rect 41568 334822 41780 334878
rect 41836 334822 41841 334878
rect 41568 334820 41841 334822
rect 41775 334817 41841 334820
rect 41538 334140 41598 334258
rect 41538 334080 41790 334140
rect 28866 333551 28926 333888
rect 41730 333696 41790 334080
rect 28815 333546 28926 333551
rect 28815 333490 28820 333546
rect 28876 333490 28926 333546
rect 28815 333488 28926 333490
rect 41538 333636 41790 333696
rect 28815 333485 28881 333488
rect 41538 333400 41598 333636
rect 674938 333486 674944 333550
rect 675008 333548 675014 333550
rect 675375 333548 675441 333551
rect 675008 333546 675441 333548
rect 675008 333490 675380 333546
rect 675436 333490 675441 333546
rect 675008 333488 675441 333490
rect 675008 333486 675014 333488
rect 675375 333485 675441 333488
rect 41775 333400 41841 333403
rect 41538 333398 41841 333400
rect 41538 333370 41780 333398
rect 41568 333342 41780 333370
rect 41836 333342 41841 333398
rect 41568 333340 41841 333342
rect 41775 333337 41841 333340
rect 28815 333104 28881 333107
rect 28815 333102 28926 333104
rect 28815 333046 28820 333102
rect 28876 333046 28926 333102
rect 28815 333041 28926 333046
rect 28866 332778 28926 333041
rect 675130 330526 675136 330590
rect 675200 330588 675206 330590
rect 675471 330588 675537 330591
rect 675200 330586 675537 330588
rect 675200 330530 675476 330586
rect 675532 330530 675537 330586
rect 675200 330528 675537 330530
rect 675200 330526 675206 330528
rect 675471 330525 675537 330528
rect 674554 328306 674560 328370
rect 674624 328368 674630 328370
rect 675375 328368 675441 328371
rect 674624 328366 675441 328368
rect 674624 328310 675380 328366
rect 675436 328310 675441 328366
rect 674624 328308 675441 328310
rect 674624 328306 674630 328308
rect 675375 328305 675441 328308
rect 674746 326826 674752 326890
rect 674816 326888 674822 326890
rect 675375 326888 675441 326891
rect 674816 326886 675441 326888
rect 674816 326830 675380 326886
rect 675436 326830 675441 326886
rect 674816 326828 675441 326830
rect 674816 326826 674822 326828
rect 675375 326825 675441 326828
rect 41775 324966 41841 324967
rect 41722 324964 41728 324966
rect 41684 324904 41728 324964
rect 41792 324962 41841 324966
rect 654831 324964 654897 324967
rect 41836 324906 41841 324962
rect 41722 324902 41728 324904
rect 41792 324902 41841 324906
rect 650208 324962 654897 324964
rect 650208 324906 654836 324962
rect 654892 324906 654897 324962
rect 650208 324904 654897 324906
rect 41775 324901 41841 324902
rect 654831 324901 654897 324904
rect 59535 324224 59601 324227
rect 59535 324222 64416 324224
rect 59535 324166 59540 324222
rect 59596 324166 64416 324222
rect 59535 324164 64416 324166
rect 59535 324161 59601 324164
rect 40378 319722 40384 319786
rect 40448 319784 40454 319786
rect 41775 319784 41841 319787
rect 40448 319782 41841 319784
rect 40448 319726 41780 319782
rect 41836 319726 41841 319782
rect 40448 319724 41841 319726
rect 40448 319722 40454 319724
rect 41775 319721 41841 319724
rect 41530 316762 41536 316826
rect 41600 316824 41606 316826
rect 41775 316824 41841 316827
rect 41600 316822 41841 316824
rect 41600 316766 41780 316822
rect 41836 316766 41841 316822
rect 41600 316764 41841 316766
rect 41600 316762 41606 316764
rect 41775 316761 41841 316764
rect 41338 316022 41344 316086
rect 41408 316084 41414 316086
rect 41775 316084 41841 316087
rect 41408 316082 41841 316084
rect 41408 316026 41780 316082
rect 41836 316026 41841 316082
rect 41408 316024 41841 316026
rect 41408 316022 41414 316024
rect 41775 316021 41841 316024
rect 41146 315430 41152 315494
rect 41216 315492 41222 315494
rect 41775 315492 41841 315495
rect 41216 315490 41841 315492
rect 41216 315434 41780 315490
rect 41836 315434 41841 315490
rect 41216 315432 41841 315434
rect 41216 315430 41222 315432
rect 41775 315429 41841 315432
rect 676047 315048 676113 315051
rect 676047 315046 676320 315048
rect 676047 314990 676052 315046
rect 676108 314990 676320 315046
rect 676047 314988 676320 314990
rect 676047 314985 676113 314988
rect 676239 314752 676305 314755
rect 676239 314750 676350 314752
rect 676239 314694 676244 314750
rect 676300 314694 676350 314750
rect 676239 314689 676350 314694
rect 676290 314574 676350 314689
rect 676047 314012 676113 314015
rect 676047 314010 676320 314012
rect 676047 313954 676052 314010
rect 676108 313954 676320 314010
rect 676047 313952 676320 313954
rect 676047 313949 676113 313952
rect 40762 313654 40768 313718
rect 40832 313716 40838 313718
rect 41871 313716 41937 313719
rect 40832 313714 41937 313716
rect 40832 313658 41876 313714
rect 41932 313658 41937 313714
rect 40832 313656 41937 313658
rect 40832 313654 40838 313656
rect 41871 313653 41937 313656
rect 673978 313506 673984 313570
rect 674048 313568 674054 313570
rect 674048 313508 676320 313568
rect 674048 313506 674054 313508
rect 40954 313210 40960 313274
rect 41024 313272 41030 313274
rect 41775 313272 41841 313275
rect 41024 313270 41841 313272
rect 41024 313214 41780 313270
rect 41836 313214 41841 313270
rect 41024 313212 41841 313214
rect 41024 313210 41030 313212
rect 41775 313209 41841 313212
rect 674362 312618 674368 312682
rect 674432 312680 674438 312682
rect 676290 312680 676350 313020
rect 674432 312620 676350 312680
rect 674432 312618 674438 312620
rect 674170 312470 674176 312534
rect 674240 312532 674246 312534
rect 674240 312472 676320 312532
rect 674240 312470 674246 312472
rect 40570 312322 40576 312386
rect 40640 312384 40646 312386
rect 41775 312384 41841 312387
rect 40640 312382 41841 312384
rect 40640 312326 41780 312382
rect 41836 312326 41841 312382
rect 40640 312324 41841 312326
rect 40640 312322 40646 312324
rect 41775 312321 41841 312324
rect 654447 311792 654513 311795
rect 673978 311792 673984 311794
rect 650208 311790 654513 311792
rect 650208 311734 654452 311790
rect 654508 311734 654513 311790
rect 650208 311732 654513 311734
rect 654447 311729 654513 311732
rect 659490 311732 673984 311792
rect 58575 311200 58641 311203
rect 655119 311200 655185 311203
rect 659490 311200 659550 311732
rect 673978 311730 673984 311732
rect 674048 311792 674054 311794
rect 676290 311792 676350 312058
rect 674048 311732 676350 311792
rect 674048 311730 674054 311732
rect 675898 311508 675904 311572
rect 675968 311570 675974 311572
rect 675968 311510 676320 311570
rect 675968 311508 675974 311510
rect 58575 311198 64416 311200
rect 58575 311142 58580 311198
rect 58636 311142 64416 311198
rect 58575 311140 64416 311142
rect 655119 311198 659550 311200
rect 655119 311142 655124 311198
rect 655180 311142 659550 311198
rect 655119 311140 659550 311142
rect 58575 311137 58641 311140
rect 655119 311137 655185 311140
rect 660975 311052 661041 311055
rect 674170 311052 674176 311054
rect 660975 311050 674176 311052
rect 660975 310994 660980 311050
rect 661036 310994 674176 311050
rect 660975 310992 674176 310994
rect 660975 310989 661041 310992
rect 674170 310990 674176 310992
rect 674240 311052 674246 311054
rect 674240 310992 676320 311052
rect 674240 310990 674246 310992
rect 676047 310608 676113 310611
rect 676047 310606 676320 310608
rect 676047 310550 676052 310606
rect 676108 310550 676320 310606
rect 676047 310548 676320 310550
rect 676047 310545 676113 310548
rect 674554 309954 674560 310018
rect 674624 310016 674630 310018
rect 674624 309956 676320 310016
rect 674624 309954 674630 309956
rect 676047 309572 676113 309575
rect 676047 309570 676320 309572
rect 676047 309514 676052 309570
rect 676108 309514 676320 309570
rect 676047 309512 676320 309514
rect 676047 309509 676113 309512
rect 675322 309066 675328 309130
rect 675392 309128 675398 309130
rect 675392 309068 676320 309128
rect 675392 309066 675398 309068
rect 675130 308474 675136 308538
rect 675200 308536 675206 308538
rect 675200 308476 676320 308536
rect 675200 308474 675206 308476
rect 674746 307734 674752 307798
rect 674816 307796 674822 307798
rect 676290 307796 676350 307988
rect 674816 307736 676350 307796
rect 674816 307734 674822 307736
rect 676047 307648 676113 307651
rect 676047 307646 676320 307648
rect 676047 307590 676052 307646
rect 676108 307590 676320 307646
rect 676047 307588 676320 307590
rect 676047 307585 676113 307588
rect 676290 306911 676350 307026
rect 676239 306906 676350 306911
rect 676239 306850 676244 306906
rect 676300 306850 676350 306906
rect 676239 306848 676350 306850
rect 676239 306845 676305 306848
rect 676290 306319 676350 306508
rect 676239 306314 676350 306319
rect 676239 306258 676244 306314
rect 676300 306258 676350 306314
rect 676239 306256 676350 306258
rect 676239 306253 676305 306256
rect 674938 306106 674944 306170
rect 675008 306168 675014 306170
rect 675008 306108 676320 306168
rect 675008 306106 675014 306108
rect 675514 305514 675520 305578
rect 675584 305576 675590 305578
rect 675584 305516 676320 305576
rect 675584 305514 675590 305516
rect 676290 304839 676350 304954
rect 676239 304834 676350 304839
rect 676239 304778 676244 304834
rect 676300 304778 676350 304834
rect 676239 304776 676350 304778
rect 676239 304773 676305 304776
rect 675706 304552 675712 304616
rect 675776 304614 675782 304616
rect 675776 304554 676320 304614
rect 675776 304552 675782 304554
rect 676047 304096 676113 304099
rect 676047 304094 676320 304096
rect 676047 304038 676052 304094
rect 676108 304038 676320 304094
rect 676047 304036 676320 304038
rect 676047 304033 676113 304036
rect 679938 303359 679998 303474
rect 679887 303354 679998 303359
rect 679887 303298 679892 303354
rect 679948 303298 679998 303354
rect 679887 303296 679998 303298
rect 679887 303293 679953 303296
rect 679746 302767 679806 303104
rect 679887 302912 679953 302915
rect 679887 302910 679998 302912
rect 679887 302854 679892 302910
rect 679948 302854 679998 302910
rect 679887 302849 679998 302854
rect 679746 302762 679857 302767
rect 679746 302706 679796 302762
rect 679852 302706 679857 302762
rect 679746 302704 679857 302706
rect 679791 302701 679857 302704
rect 41775 302690 41841 302693
rect 41568 302688 41841 302690
rect 41568 302632 41780 302688
rect 41836 302632 41841 302688
rect 41568 302630 41841 302632
rect 41775 302627 41841 302630
rect 679938 302586 679998 302849
rect 41583 302320 41649 302323
rect 679791 302320 679857 302323
rect 41538 302318 41649 302320
rect 41538 302262 41588 302318
rect 41644 302262 41649 302318
rect 41538 302257 41649 302262
rect 679746 302318 679857 302320
rect 679746 302262 679796 302318
rect 679852 302262 679857 302318
rect 679746 302257 679857 302262
rect 41538 302142 41598 302257
rect 679746 301994 679806 302257
rect 41775 301580 41841 301583
rect 41568 301578 41841 301580
rect 41568 301522 41780 301578
rect 41836 301522 41841 301578
rect 41568 301520 41841 301522
rect 41775 301517 41841 301520
rect 41775 301210 41841 301213
rect 41568 301208 41841 301210
rect 41568 301152 41780 301208
rect 41836 301152 41841 301208
rect 41568 301150 41841 301152
rect 41775 301147 41841 301150
rect 41775 300692 41841 300695
rect 41568 300690 41841 300692
rect 41568 300634 41780 300690
rect 41836 300634 41841 300690
rect 41568 300632 41841 300634
rect 41775 300629 41841 300632
rect 41775 300100 41841 300103
rect 41568 300098 41841 300100
rect 41568 300042 41780 300098
rect 41836 300042 41841 300098
rect 41568 300040 41841 300042
rect 41775 300037 41841 300040
rect 41775 299656 41841 299659
rect 41568 299654 41841 299656
rect 41568 299598 41780 299654
rect 41836 299598 41841 299654
rect 41568 299596 41841 299598
rect 41775 299593 41841 299596
rect 41583 299360 41649 299363
rect 41538 299358 41649 299360
rect 41538 299302 41588 299358
rect 41644 299302 41649 299358
rect 41538 299297 41649 299302
rect 41538 299182 41598 299297
rect 41775 298620 41841 298623
rect 41568 298618 41841 298620
rect 41568 298562 41780 298618
rect 41836 298562 41841 298618
rect 41568 298560 41841 298562
rect 41775 298557 41841 298560
rect 655119 298472 655185 298475
rect 650208 298470 655185 298472
rect 650208 298414 655124 298470
rect 655180 298414 655185 298470
rect 650208 298412 655185 298414
rect 655119 298409 655185 298412
rect 40578 297882 40638 298146
rect 59535 298028 59601 298031
rect 59535 298026 64416 298028
rect 59535 297970 59540 298026
rect 59596 297970 64416 298026
rect 59535 297968 64416 297970
rect 59535 297965 59601 297968
rect 40570 297818 40576 297882
rect 40640 297818 40646 297882
rect 41722 297658 41728 297660
rect 41568 297598 41728 297658
rect 41722 297596 41728 297598
rect 41792 297596 41798 297660
rect 40762 297226 40768 297290
rect 40832 297226 40838 297290
rect 40770 297110 40830 297226
rect 41154 296550 41214 296670
rect 41146 296486 41152 296550
rect 41216 296486 41222 296550
rect 41538 295810 41598 296148
rect 41530 295746 41536 295810
rect 41600 295746 41606 295810
rect 41967 295660 42033 295663
rect 41568 295658 42033 295660
rect 41568 295602 41972 295658
rect 42028 295602 42033 295658
rect 41568 295600 42033 295602
rect 41967 295597 42033 295600
rect 40962 294922 41022 295186
rect 40954 294858 40960 294922
rect 41024 294858 41030 294922
rect 40386 294330 40446 294594
rect 40378 294266 40384 294330
rect 40448 294266 40454 294330
rect 41346 293886 41406 294150
rect 41338 293822 41344 293886
rect 41408 293822 41414 293886
rect 41775 293736 41841 293739
rect 41568 293734 41841 293736
rect 41568 293678 41780 293734
rect 41836 293678 41841 293734
rect 41568 293676 41841 293678
rect 41775 293673 41841 293676
rect 41538 292999 41598 293114
rect 41538 292994 41649 292999
rect 41538 292938 41588 292994
rect 41644 292938 41649 292994
rect 41538 292936 41649 292938
rect 41583 292933 41649 292936
rect 675375 292850 675441 292851
rect 675322 292848 675328 292850
rect 675284 292788 675328 292848
rect 675392 292846 675441 292850
rect 675436 292790 675441 292846
rect 675322 292786 675328 292788
rect 675392 292786 675441 292790
rect 675375 292785 675441 292786
rect 41871 292626 41937 292629
rect 41568 292624 41937 292626
rect 41568 292568 41876 292624
rect 41932 292568 41937 292624
rect 41568 292566 41937 292568
rect 41871 292563 41937 292566
rect 41871 292256 41937 292259
rect 41568 292254 41937 292256
rect 41568 292198 41876 292254
rect 41932 292198 41937 292254
rect 41568 292196 41937 292198
rect 41871 292193 41937 292196
rect 41538 291519 41598 291634
rect 41538 291514 41649 291519
rect 41538 291458 41588 291514
rect 41644 291458 41649 291514
rect 41538 291456 41649 291458
rect 41583 291453 41649 291456
rect 41538 290924 41598 291116
rect 41538 290864 41790 290924
rect 28866 290483 28926 290746
rect 28815 290478 28926 290483
rect 41730 290480 41790 290864
rect 28815 290422 28820 290478
rect 28876 290422 28926 290478
rect 28815 290420 28926 290422
rect 41538 290420 41790 290480
rect 28815 290417 28881 290420
rect 41538 290184 41598 290420
rect 41775 290184 41841 290187
rect 41538 290182 41841 290184
rect 41538 290154 41780 290182
rect 41568 290126 41780 290154
rect 41836 290126 41841 290182
rect 41568 290124 41841 290126
rect 41775 290121 41841 290124
rect 28815 289888 28881 289891
rect 28815 289886 28926 289888
rect 28815 289830 28820 289886
rect 28876 289830 28926 289886
rect 28815 289825 28926 289830
rect 28866 289562 28926 289825
rect 675130 288494 675136 288558
rect 675200 288556 675206 288558
rect 675471 288556 675537 288559
rect 675200 288554 675537 288556
rect 675200 288498 675476 288554
rect 675532 288498 675537 288554
rect 675200 288496 675537 288498
rect 675200 288494 675206 288496
rect 675471 288493 675537 288496
rect 675663 287818 675729 287819
rect 675663 287814 675712 287818
rect 675776 287816 675782 287818
rect 675663 287758 675668 287814
rect 675663 287754 675712 287758
rect 675776 287756 675820 287816
rect 675776 287754 675782 287756
rect 675663 287753 675729 287754
rect 675471 287374 675537 287375
rect 675471 287370 675520 287374
rect 675584 287372 675590 287374
rect 675471 287314 675476 287370
rect 675471 287310 675520 287314
rect 675584 287312 675628 287372
rect 675584 287310 675590 287312
rect 675471 287309 675537 287310
rect 655407 285300 655473 285303
rect 650208 285298 655473 285300
rect 650208 285242 655412 285298
rect 655468 285242 655473 285298
rect 650208 285240 655473 285242
rect 655407 285237 655473 285240
rect 674938 285238 674944 285302
rect 675008 285300 675014 285302
rect 675471 285300 675537 285303
rect 675008 285298 675537 285300
rect 675008 285242 675476 285298
rect 675532 285242 675537 285298
rect 675008 285240 675537 285242
rect 675008 285238 675014 285240
rect 675471 285237 675537 285240
rect 59535 285152 59601 285155
rect 59535 285150 64416 285152
rect 59535 285094 59540 285150
rect 59596 285094 64416 285150
rect 59535 285092 64416 285094
rect 59535 285089 59601 285092
rect 674554 283610 674560 283674
rect 674624 283672 674630 283674
rect 675375 283672 675441 283675
rect 674624 283670 675441 283672
rect 674624 283614 675380 283670
rect 675436 283614 675441 283670
rect 674624 283612 675441 283614
rect 674624 283610 674630 283612
rect 675375 283609 675441 283612
rect 674746 281834 674752 281898
rect 674816 281896 674822 281898
rect 675375 281896 675441 281899
rect 674816 281894 675441 281896
rect 674816 281838 675380 281894
rect 675436 281838 675441 281894
rect 674816 281836 675441 281838
rect 674816 281834 674822 281836
rect 675375 281833 675441 281836
rect 41775 281750 41841 281751
rect 41722 281748 41728 281750
rect 41684 281688 41728 281748
rect 41792 281746 41841 281750
rect 41836 281690 41841 281746
rect 41722 281686 41728 281688
rect 41792 281686 41841 281690
rect 41775 281685 41841 281686
rect 42106 278578 42112 278642
rect 42176 278640 42182 278642
rect 670287 278640 670353 278643
rect 42176 278638 670353 278640
rect 42176 278582 670292 278638
rect 670348 278582 670353 278638
rect 42176 278580 670353 278582
rect 42176 278578 42182 278580
rect 670287 278577 670353 278580
rect 44175 278492 44241 278495
rect 669903 278492 669969 278495
rect 44175 278490 669969 278492
rect 44175 278434 44180 278490
rect 44236 278434 669908 278490
rect 669964 278434 669969 278490
rect 44175 278432 669969 278434
rect 44175 278429 44241 278432
rect 669903 278429 669969 278432
rect 62031 278344 62097 278347
rect 670095 278344 670161 278347
rect 62031 278342 670161 278344
rect 62031 278286 62036 278342
rect 62092 278286 670100 278342
rect 670156 278286 670161 278342
rect 62031 278284 670161 278286
rect 62031 278281 62097 278284
rect 670095 278281 670161 278284
rect 62223 278196 62289 278199
rect 669711 278196 669777 278199
rect 62223 278194 669777 278196
rect 62223 278138 62228 278194
rect 62284 278138 669716 278194
rect 669772 278138 669777 278194
rect 62223 278136 669777 278138
rect 62223 278133 62289 278136
rect 669711 278133 669777 278136
rect 63375 278048 63441 278051
rect 652623 278048 652689 278051
rect 63375 278046 652689 278048
rect 63375 277990 63380 278046
rect 63436 277990 652628 278046
rect 652684 277990 652689 278046
rect 63375 277988 652689 277990
rect 63375 277985 63441 277988
rect 652623 277985 652689 277988
rect 41530 276506 41536 276570
rect 41600 276568 41606 276570
rect 41775 276568 41841 276571
rect 41600 276566 41841 276568
rect 41600 276510 41780 276566
rect 41836 276510 41841 276566
rect 41600 276508 41841 276510
rect 41600 276506 41606 276508
rect 41775 276505 41841 276508
rect 368943 276420 369009 276423
rect 542223 276420 542289 276423
rect 368943 276418 542289 276420
rect 368943 276362 368948 276418
rect 369004 276362 542228 276418
rect 542284 276362 542289 276418
rect 368943 276360 542289 276362
rect 368943 276357 369009 276360
rect 542223 276357 542289 276360
rect 381807 276272 381873 276275
rect 574191 276272 574257 276275
rect 381807 276270 574257 276272
rect 381807 276214 381812 276270
rect 381868 276214 574196 276270
rect 574252 276214 574257 276270
rect 381807 276212 574257 276214
rect 381807 276209 381873 276212
rect 574191 276209 574257 276212
rect 383631 276124 383697 276127
rect 578895 276124 578961 276127
rect 383631 276122 578961 276124
rect 383631 276066 383636 276122
rect 383692 276066 578900 276122
rect 578956 276066 578961 276122
rect 383631 276064 578961 276066
rect 383631 276061 383697 276064
rect 578895 276061 578961 276064
rect 384879 275976 384945 275979
rect 581295 275976 581361 275979
rect 384879 275974 581361 275976
rect 384879 275918 384884 275974
rect 384940 275918 581300 275974
rect 581356 275918 581361 275974
rect 384879 275916 581361 275918
rect 384879 275913 384945 275916
rect 581295 275913 581361 275916
rect 387759 275828 387825 275831
rect 588303 275828 588369 275831
rect 387759 275826 588369 275828
rect 387759 275770 387764 275826
rect 387820 275770 588308 275826
rect 588364 275770 588369 275826
rect 387759 275768 588369 275770
rect 387759 275765 387825 275768
rect 588303 275765 588369 275768
rect 390831 275680 390897 275683
rect 596655 275680 596721 275683
rect 390831 275678 596721 275680
rect 390831 275622 390836 275678
rect 390892 275622 596660 275678
rect 596716 275622 596721 275678
rect 390831 275620 596721 275622
rect 390831 275617 390897 275620
rect 596655 275617 596721 275620
rect 391983 275532 392049 275535
rect 599055 275532 599121 275535
rect 391983 275530 599121 275532
rect 391983 275474 391988 275530
rect 392044 275474 599060 275530
rect 599116 275474 599121 275530
rect 391983 275472 599121 275474
rect 391983 275469 392049 275472
rect 599055 275469 599121 275472
rect 393231 275384 393297 275387
rect 602511 275384 602577 275387
rect 393231 275382 602577 275384
rect 393231 275326 393236 275382
rect 393292 275326 602516 275382
rect 602572 275326 602577 275382
rect 393231 275324 602577 275326
rect 393231 275321 393297 275324
rect 602511 275321 602577 275324
rect 397551 275236 397617 275239
rect 613167 275236 613233 275239
rect 397551 275234 613233 275236
rect 397551 275178 397556 275234
rect 397612 275178 613172 275234
rect 613228 275178 613233 275234
rect 397551 275176 613233 275178
rect 397551 275173 397617 275176
rect 613167 275173 613233 275176
rect 396303 275088 396369 275091
rect 609711 275088 609777 275091
rect 396303 275086 609777 275088
rect 396303 275030 396308 275086
rect 396364 275030 609716 275086
rect 609772 275030 609777 275086
rect 396303 275028 609777 275030
rect 396303 275025 396369 275028
rect 609711 275025 609777 275028
rect 41338 273546 41344 273610
rect 41408 273608 41414 273610
rect 41775 273608 41841 273611
rect 41408 273606 41841 273608
rect 41408 273550 41780 273606
rect 41836 273550 41841 273606
rect 41408 273548 41841 273550
rect 41408 273546 41414 273548
rect 41775 273545 41841 273548
rect 371247 273608 371313 273611
rect 548175 273608 548241 273611
rect 371247 273606 548241 273608
rect 371247 273550 371252 273606
rect 371308 273550 548180 273606
rect 548236 273550 548241 273606
rect 371247 273548 548241 273550
rect 371247 273545 371313 273548
rect 548175 273545 548241 273548
rect 377007 273460 377073 273463
rect 562383 273460 562449 273463
rect 377007 273458 562449 273460
rect 377007 273402 377012 273458
rect 377068 273402 562388 273458
rect 562444 273402 562449 273458
rect 377007 273400 562449 273402
rect 377007 273397 377073 273400
rect 562383 273397 562449 273400
rect 379887 273312 379953 273315
rect 569487 273312 569553 273315
rect 379887 273310 569553 273312
rect 379887 273254 379892 273310
rect 379948 273254 569492 273310
rect 569548 273254 569553 273310
rect 379887 273252 569553 273254
rect 379887 273249 379953 273252
rect 569487 273249 569553 273252
rect 385551 273164 385617 273167
rect 583599 273164 583665 273167
rect 385551 273162 583665 273164
rect 385551 273106 385556 273162
rect 385612 273106 583604 273162
rect 583660 273106 583665 273162
rect 385551 273104 583665 273106
rect 385551 273101 385617 273104
rect 583599 273101 583665 273104
rect 391503 273016 391569 273019
rect 597807 273016 597873 273019
rect 391503 273014 597873 273016
rect 391503 272958 391508 273014
rect 391564 272958 597812 273014
rect 597868 272958 597873 273014
rect 391503 272956 597873 272958
rect 391503 272953 391569 272956
rect 597807 272953 597873 272956
rect 40378 272806 40384 272870
rect 40448 272868 40454 272870
rect 41775 272868 41841 272871
rect 40448 272866 41841 272868
rect 40448 272810 41780 272866
rect 41836 272810 41841 272866
rect 40448 272808 41841 272810
rect 40448 272806 40454 272808
rect 41775 272805 41841 272808
rect 394383 272868 394449 272871
rect 604911 272868 604977 272871
rect 394383 272866 604977 272868
rect 394383 272810 394388 272866
rect 394444 272810 604916 272866
rect 604972 272810 604977 272866
rect 394383 272808 604977 272810
rect 394383 272805 394449 272808
rect 604911 272805 604977 272808
rect 399951 272720 400017 272723
rect 619023 272720 619089 272723
rect 399951 272718 619089 272720
rect 399951 272662 399956 272718
rect 400012 272662 619028 272718
rect 619084 272662 619089 272718
rect 399951 272660 619089 272662
rect 399951 272657 400017 272660
rect 619023 272657 619089 272660
rect 403023 272572 403089 272575
rect 626127 272572 626193 272575
rect 403023 272570 626193 272572
rect 403023 272514 403028 272570
rect 403084 272514 626132 272570
rect 626188 272514 626193 272570
rect 403023 272512 626193 272514
rect 403023 272509 403089 272512
rect 626127 272509 626193 272512
rect 41146 272362 41152 272426
rect 41216 272424 41222 272426
rect 41775 272424 41841 272427
rect 41216 272422 41841 272424
rect 41216 272366 41780 272422
rect 41836 272366 41841 272422
rect 41216 272364 41841 272366
rect 41216 272362 41222 272364
rect 41775 272361 41841 272364
rect 405615 272424 405681 272427
rect 633327 272424 633393 272427
rect 405615 272422 633393 272424
rect 405615 272366 405620 272422
rect 405676 272366 633332 272422
rect 633388 272366 633393 272422
rect 405615 272364 633393 272366
rect 405615 272361 405681 272364
rect 633327 272361 633393 272364
rect 69423 272276 69489 272279
rect 193071 272276 193137 272279
rect 69423 272274 193137 272276
rect 69423 272218 69428 272274
rect 69484 272218 193076 272274
rect 193132 272218 193137 272274
rect 69423 272216 193137 272218
rect 69423 272213 69489 272216
rect 193071 272213 193137 272216
rect 408495 272276 408561 272279
rect 640431 272276 640497 272279
rect 408495 272274 640497 272276
rect 408495 272218 408500 272274
rect 408556 272218 640436 272274
rect 640492 272218 640497 272274
rect 408495 272216 640497 272218
rect 408495 272213 408561 272216
rect 640431 272213 640497 272216
rect 71727 272128 71793 272131
rect 194223 272128 194289 272131
rect 71727 272126 194289 272128
rect 71727 272070 71732 272126
rect 71788 272070 194228 272126
rect 194284 272070 194289 272126
rect 71727 272068 194289 272070
rect 71727 272065 71793 272068
rect 194223 272065 194289 272068
rect 411759 272128 411825 272131
rect 648687 272128 648753 272131
rect 411759 272126 648753 272128
rect 411759 272070 411764 272126
rect 411820 272070 648692 272126
rect 648748 272070 648753 272126
rect 411759 272068 648753 272070
rect 411759 272065 411825 272068
rect 648687 272065 648753 272068
rect 370095 271980 370161 271983
rect 544623 271980 544689 271983
rect 370095 271978 544689 271980
rect 370095 271922 370100 271978
rect 370156 271922 544628 271978
rect 544684 271922 544689 271978
rect 370095 271920 544689 271922
rect 370095 271917 370161 271920
rect 544623 271917 544689 271920
rect 378639 270648 378705 270651
rect 565839 270648 565905 270651
rect 378639 270646 565905 270648
rect 378639 270590 378644 270646
rect 378700 270590 565844 270646
rect 565900 270590 565905 270646
rect 378639 270588 565905 270590
rect 378639 270585 378705 270588
rect 565839 270585 565905 270588
rect 40570 270438 40576 270502
rect 40640 270500 40646 270502
rect 41775 270500 41841 270503
rect 40640 270498 41841 270500
rect 40640 270442 41780 270498
rect 41836 270442 41841 270498
rect 40640 270440 41841 270442
rect 40640 270438 40646 270440
rect 41775 270437 41841 270440
rect 381231 270500 381297 270503
rect 572943 270500 573009 270503
rect 381231 270498 573009 270500
rect 381231 270442 381236 270498
rect 381292 270442 572948 270498
rect 573004 270442 573009 270498
rect 381231 270440 573009 270442
rect 381231 270437 381297 270440
rect 572943 270437 573009 270440
rect 387279 270352 387345 270355
rect 587151 270352 587217 270355
rect 387279 270350 587217 270352
rect 387279 270294 387284 270350
rect 387340 270294 587156 270350
rect 587212 270294 587217 270350
rect 387279 270292 587217 270294
rect 387279 270289 387345 270292
rect 587151 270289 587217 270292
rect 390159 270204 390225 270207
rect 594351 270204 594417 270207
rect 390159 270202 594417 270204
rect 390159 270146 390164 270202
rect 390220 270146 594356 270202
rect 594412 270146 594417 270202
rect 390159 270144 594417 270146
rect 390159 270141 390225 270144
rect 594351 270141 594417 270144
rect 40954 269994 40960 270058
rect 41024 270056 41030 270058
rect 41775 270056 41841 270059
rect 41024 270054 41841 270056
rect 41024 269998 41780 270054
rect 41836 269998 41841 270054
rect 41024 269996 41841 269998
rect 41024 269994 41030 269996
rect 41775 269993 41841 269996
rect 395631 270056 395697 270059
rect 608463 270056 608529 270059
rect 395631 270054 608529 270056
rect 395631 269998 395636 270054
rect 395692 269998 608468 270054
rect 608524 269998 608529 270054
rect 395631 269996 608529 269998
rect 395631 269993 395697 269996
rect 608463 269993 608529 269996
rect 676047 270056 676113 270059
rect 676047 270054 676320 270056
rect 676047 269998 676052 270054
rect 676108 269998 676320 270054
rect 676047 269996 676320 269998
rect 676047 269993 676113 269996
rect 130863 269908 130929 269911
rect 210735 269908 210801 269911
rect 130863 269906 210801 269908
rect 130863 269850 130868 269906
rect 130924 269850 210740 269906
rect 210796 269850 210801 269906
rect 130863 269848 210801 269850
rect 130863 269845 130929 269848
rect 210735 269845 210801 269848
rect 401295 269908 401361 269911
rect 622671 269908 622737 269911
rect 401295 269906 622737 269908
rect 401295 269850 401300 269906
rect 401356 269850 622676 269906
rect 622732 269850 622737 269906
rect 401295 269848 622737 269850
rect 401295 269845 401361 269848
rect 622671 269845 622737 269848
rect 128559 269760 128625 269763
rect 210255 269760 210321 269763
rect 128559 269758 210321 269760
rect 128559 269702 128564 269758
rect 128620 269702 210260 269758
rect 210316 269702 210321 269758
rect 128559 269700 210321 269702
rect 128559 269697 128625 269700
rect 210255 269697 210321 269700
rect 404175 269760 404241 269763
rect 629775 269760 629841 269763
rect 404175 269758 629841 269760
rect 404175 269702 404180 269758
rect 404236 269702 629780 269758
rect 629836 269702 629841 269758
rect 404175 269700 629841 269702
rect 404175 269697 404241 269700
rect 629775 269697 629841 269700
rect 676239 269760 676305 269763
rect 676239 269758 676350 269760
rect 676239 269702 676244 269758
rect 676300 269702 676350 269758
rect 676239 269697 676350 269702
rect 70575 269612 70641 269615
rect 193743 269612 193809 269615
rect 70575 269610 193809 269612
rect 70575 269554 70580 269610
rect 70636 269554 193748 269610
rect 193804 269554 193809 269610
rect 70575 269552 193809 269554
rect 70575 269549 70641 269552
rect 193743 269549 193809 269552
rect 409935 269612 410001 269615
rect 643887 269612 643953 269615
rect 409935 269610 643953 269612
rect 409935 269554 409940 269610
rect 409996 269554 643892 269610
rect 643948 269554 643953 269610
rect 676290 269582 676350 269697
rect 409935 269552 643953 269554
rect 409935 269549 410001 269552
rect 643887 269549 643953 269552
rect 67023 269464 67089 269467
rect 192591 269464 192657 269467
rect 67023 269462 192657 269464
rect 67023 269406 67028 269462
rect 67084 269406 192596 269462
rect 192652 269406 192657 269462
rect 67023 269404 192657 269406
rect 67023 269401 67089 269404
rect 192591 269401 192657 269404
rect 410415 269464 410481 269467
rect 645135 269464 645201 269467
rect 410415 269462 645201 269464
rect 410415 269406 410420 269462
rect 410476 269406 645140 269462
rect 645196 269406 645201 269462
rect 410415 269404 645201 269406
rect 410415 269401 410481 269404
rect 645135 269401 645201 269404
rect 65871 269316 65937 269319
rect 192399 269316 192465 269319
rect 65871 269314 192465 269316
rect 65871 269258 65876 269314
rect 65932 269258 192404 269314
rect 192460 269258 192465 269314
rect 65871 269256 192465 269258
rect 65871 269253 65937 269256
rect 192399 269253 192465 269256
rect 370287 269316 370353 269319
rect 402831 269316 402897 269319
rect 370287 269314 402897 269316
rect 370287 269258 370292 269314
rect 370348 269258 402836 269314
rect 402892 269258 402897 269314
rect 370287 269256 402897 269258
rect 370287 269253 370353 269256
rect 402831 269253 402897 269256
rect 411567 269316 411633 269319
rect 647535 269316 647601 269319
rect 411567 269314 647601 269316
rect 411567 269258 411572 269314
rect 411628 269258 647540 269314
rect 647596 269258 647601 269314
rect 411567 269256 647601 269258
rect 411567 269253 411633 269256
rect 647535 269253 647601 269256
rect 40762 269106 40768 269170
rect 40832 269168 40838 269170
rect 41775 269168 41841 269171
rect 40832 269166 41841 269168
rect 40832 269110 41780 269166
rect 41836 269110 41841 269166
rect 40832 269108 41841 269110
rect 40832 269106 40838 269108
rect 41775 269105 41841 269108
rect 375567 269168 375633 269171
rect 558831 269168 558897 269171
rect 375567 269166 558897 269168
rect 375567 269110 375572 269166
rect 375628 269110 558836 269166
rect 558892 269110 558897 269166
rect 375567 269108 558897 269110
rect 375567 269105 375633 269108
rect 558831 269105 558897 269108
rect 676239 269168 676305 269171
rect 676239 269166 676350 269168
rect 676239 269110 676244 269166
rect 676300 269110 676350 269166
rect 676239 269105 676350 269110
rect 372687 269020 372753 269023
rect 551727 269020 551793 269023
rect 372687 269018 551793 269020
rect 372687 268962 372692 269018
rect 372748 268962 551732 269018
rect 551788 268962 551793 269018
rect 676290 268990 676350 269105
rect 372687 268960 551793 268962
rect 372687 268957 372753 268960
rect 551727 268957 551793 268960
rect 368367 268872 368433 268875
rect 541071 268872 541137 268875
rect 368367 268870 541137 268872
rect 368367 268814 368372 268870
rect 368428 268814 541076 268870
rect 541132 268814 541137 268870
rect 368367 268812 541137 268814
rect 368367 268809 368433 268812
rect 541071 268809 541137 268812
rect 674362 268514 674368 268578
rect 674432 268576 674438 268578
rect 674432 268516 676320 268576
rect 674432 268514 674438 268516
rect 206991 267984 207057 267987
rect 211407 267984 211473 267987
rect 206991 267982 211473 267984
rect 206991 267926 206996 267982
rect 207052 267926 211412 267982
rect 211468 267926 211473 267982
rect 206991 267924 211473 267926
rect 206991 267921 207057 267924
rect 211407 267921 211473 267924
rect 675514 267922 675520 267986
rect 675584 267984 675590 267986
rect 676290 267984 676350 268028
rect 675584 267924 676350 267984
rect 675584 267922 675590 267924
rect 673978 267478 673984 267542
rect 674048 267540 674054 267542
rect 674048 267480 676320 267540
rect 674048 267478 674054 267480
rect 673978 267034 673984 267098
rect 674048 267096 674054 267098
rect 674048 267036 676320 267096
rect 674048 267034 674054 267036
rect 389679 266948 389745 266951
rect 593103 266948 593169 266951
rect 389679 266946 593169 266948
rect 389679 266890 389684 266946
rect 389740 266890 593108 266946
rect 593164 266890 593169 266946
rect 389679 266888 593169 266890
rect 389679 266885 389745 266888
rect 593103 266885 593169 266888
rect 387951 266800 388017 266803
rect 589551 266800 589617 266803
rect 387951 266798 589617 266800
rect 387951 266742 387956 266798
rect 388012 266742 589556 266798
rect 589612 266742 589617 266798
rect 387951 266740 589617 266742
rect 387951 266737 388017 266740
rect 589551 266737 589617 266740
rect 401775 266652 401841 266655
rect 623823 266652 623889 266655
rect 401775 266650 623889 266652
rect 401775 266594 401780 266650
rect 401836 266594 623828 266650
rect 623884 266594 623889 266650
rect 401775 266592 623889 266594
rect 401775 266589 401841 266592
rect 623823 266589 623889 266592
rect 409167 266504 409233 266507
rect 641583 266504 641649 266507
rect 409167 266502 641649 266504
rect 409167 266446 409172 266502
rect 409228 266446 641588 266502
rect 641644 266446 641649 266502
rect 409167 266444 641649 266446
rect 409167 266441 409233 266444
rect 641583 266441 641649 266444
rect 674170 266442 674176 266506
rect 674240 266504 674246 266506
rect 674240 266444 676320 266504
rect 674240 266442 674246 266444
rect 407823 266356 407889 266359
rect 638031 266356 638097 266359
rect 407823 266354 638097 266356
rect 407823 266298 407828 266354
rect 407884 266298 638036 266354
rect 638092 266298 638097 266354
rect 407823 266296 638097 266298
rect 407823 266293 407889 266296
rect 638031 266293 638097 266296
rect 674170 265764 674176 265766
rect 659490 265704 674176 265764
rect 658383 265172 658449 265175
rect 659490 265172 659550 265704
rect 674170 265702 674176 265704
rect 674240 265764 674246 265766
rect 676290 265764 676350 266030
rect 674240 265704 676350 265764
rect 674240 265702 674246 265704
rect 675898 265554 675904 265618
rect 675968 265616 675974 265618
rect 675968 265556 676320 265616
rect 675968 265554 675974 265556
rect 658383 265170 659550 265172
rect 658383 265114 658388 265170
rect 658444 265114 659550 265170
rect 658383 265112 659550 265114
rect 658383 265109 658449 265112
rect 658191 265024 658257 265027
rect 673978 265024 673984 265026
rect 658191 265022 673984 265024
rect 658191 264966 658196 265022
rect 658252 264966 673984 265022
rect 658191 264964 673984 264966
rect 658191 264961 658257 264964
rect 673978 264962 673984 264964
rect 674048 265024 674054 265026
rect 674362 265024 674368 265026
rect 674048 264964 674368 265024
rect 674048 264962 674054 264964
rect 674362 264962 674368 264964
rect 674432 264962 674438 265026
rect 674554 264962 674560 265026
rect 674624 265024 674630 265026
rect 674624 264964 676320 265024
rect 674624 264962 674630 264964
rect 675663 264580 675729 264583
rect 675663 264578 676320 264580
rect 675663 264522 675668 264578
rect 675724 264522 676320 264578
rect 675663 264520 676320 264522
rect 675663 264517 675729 264520
rect 675706 264074 675712 264138
rect 675776 264136 675782 264138
rect 675776 264076 676320 264136
rect 675776 264074 675782 264076
rect 673978 263482 673984 263546
rect 674048 263544 674054 263546
rect 674048 263484 676320 263544
rect 674048 263482 674054 263484
rect 674746 262742 674752 262806
rect 674816 262804 674822 262806
rect 676290 262804 676350 262996
rect 674816 262744 676350 262804
rect 674816 262742 674822 262744
rect 675759 262656 675825 262659
rect 675759 262654 676320 262656
rect 675759 262598 675764 262654
rect 675820 262598 676320 262654
rect 675759 262596 676320 262598
rect 675759 262593 675825 262596
rect 420399 262212 420465 262215
rect 412512 262210 420465 262212
rect 412512 262154 420404 262210
rect 420460 262154 420465 262210
rect 412512 262152 420465 262154
rect 420399 262149 420465 262152
rect 676290 261919 676350 262034
rect 676239 261914 676350 261919
rect 676239 261858 676244 261914
rect 676300 261858 676350 261914
rect 676239 261856 676350 261858
rect 676239 261853 676305 261856
rect 676290 261326 676350 261442
rect 676282 261262 676288 261326
rect 676352 261262 676358 261326
rect 674938 261114 674944 261178
rect 675008 261176 675014 261178
rect 675008 261116 676320 261176
rect 675008 261114 675014 261116
rect 675130 260522 675136 260586
rect 675200 260584 675206 260586
rect 675200 260524 676320 260584
rect 675200 260522 675206 260524
rect 420399 259844 420465 259847
rect 412512 259842 420465 259844
rect 412512 259786 420404 259842
rect 420460 259786 420465 259842
rect 412512 259784 420465 259786
rect 420399 259781 420465 259784
rect 676090 259782 676096 259846
rect 676160 259844 676166 259846
rect 676290 259844 676350 259962
rect 676160 259784 676350 259844
rect 676160 259782 676166 259784
rect 41583 259696 41649 259699
rect 41538 259694 41649 259696
rect 41538 259638 41588 259694
rect 41644 259638 41649 259694
rect 41538 259633 41649 259638
rect 41538 259518 41598 259633
rect 676047 259622 676113 259625
rect 676047 259620 676320 259622
rect 676047 259564 676052 259620
rect 676108 259564 676320 259620
rect 676047 259562 676320 259564
rect 676047 259559 676113 259562
rect 189999 259400 190065 259403
rect 189999 259398 191904 259400
rect 189999 259342 190004 259398
rect 190060 259342 191904 259398
rect 189999 259340 191904 259342
rect 189999 259337 190065 259340
rect 676047 259104 676113 259107
rect 676047 259102 676320 259104
rect 676047 259046 676052 259102
rect 676108 259046 676320 259102
rect 676047 259044 676320 259046
rect 676047 259041 676113 259044
rect 41775 258956 41841 258959
rect 41568 258954 41841 258956
rect 41568 258898 41780 258954
rect 41836 258898 41841 258954
rect 41568 258896 41841 258898
rect 41775 258893 41841 258896
rect 679746 258367 679806 258482
rect 41775 258364 41841 258367
rect 41568 258362 41841 258364
rect 41568 258306 41780 258362
rect 41836 258306 41841 258362
rect 41568 258304 41841 258306
rect 41775 258301 41841 258304
rect 679695 258362 679806 258367
rect 679695 258306 679700 258362
rect 679756 258306 679806 258362
rect 679695 258304 679806 258306
rect 679695 258301 679761 258304
rect 41775 257994 41841 257997
rect 41568 257992 41841 257994
rect 41568 257936 41780 257992
rect 41836 257936 41841 257992
rect 41568 257934 41841 257936
rect 41775 257931 41841 257934
rect 685506 257775 685566 258112
rect 679695 257772 679761 257775
rect 679695 257770 679806 257772
rect 679695 257714 679700 257770
rect 679756 257714 679806 257770
rect 679695 257709 679806 257714
rect 685455 257770 685566 257775
rect 685455 257714 685460 257770
rect 685516 257714 685566 257770
rect 685455 257712 685566 257714
rect 685455 257709 685521 257712
rect 679746 257594 679806 257709
rect 41775 257476 41841 257479
rect 41568 257474 41841 257476
rect 41568 257418 41780 257474
rect 41836 257418 41841 257474
rect 41568 257416 41841 257418
rect 41775 257413 41841 257416
rect 412482 257032 412542 257520
rect 685455 257328 685521 257331
rect 685455 257326 685566 257328
rect 685455 257270 685460 257326
rect 685516 257270 685566 257326
rect 685455 257265 685566 257270
rect 420399 257032 420465 257035
rect 412482 257030 420465 257032
rect 412482 256974 420404 257030
rect 420460 256974 420465 257030
rect 685506 257002 685566 257265
rect 412482 256972 420465 256974
rect 420399 256969 420465 256972
rect 41775 256884 41841 256887
rect 41568 256882 41841 256884
rect 41568 256826 41780 256882
rect 41836 256826 41841 256882
rect 41568 256824 41841 256826
rect 41775 256821 41841 256824
rect 41775 256514 41841 256517
rect 41568 256512 41841 256514
rect 41568 256456 41780 256512
rect 41836 256456 41841 256512
rect 41568 256454 41841 256456
rect 41775 256451 41841 256454
rect 41775 255996 41841 255999
rect 41568 255994 41841 255996
rect 41568 255938 41780 255994
rect 41836 255938 41841 255994
rect 41568 255936 41841 255938
rect 41775 255933 41841 255936
rect 41775 255404 41841 255407
rect 41568 255402 41841 255404
rect 41568 255346 41780 255402
rect 41836 255346 41841 255402
rect 41568 255344 41841 255346
rect 41775 255341 41841 255344
rect 420399 255256 420465 255259
rect 412512 255254 420465 255256
rect 412512 255198 420404 255254
rect 420460 255198 420465 255254
rect 412512 255196 420465 255198
rect 420399 255193 420465 255196
rect 40578 254666 40638 254930
rect 40570 254602 40576 254666
rect 40640 254602 40646 254666
rect 41722 254516 41728 254518
rect 41568 254456 41728 254516
rect 41722 254454 41728 254456
rect 41792 254454 41798 254518
rect 41914 253924 41920 253926
rect 41568 253864 41920 253924
rect 41914 253862 41920 253864
rect 41984 253862 41990 253926
rect 40962 253334 41022 253450
rect 40954 253270 40960 253334
rect 41024 253270 41030 253334
rect 41538 252594 41598 252932
rect 420399 252888 420465 252891
rect 412512 252886 420465 252888
rect 412512 252830 420404 252886
rect 420460 252830 420465 252886
rect 412512 252828 420465 252830
rect 420399 252825 420465 252828
rect 41530 252530 41536 252594
rect 41600 252530 41606 252594
rect 41871 252444 41937 252447
rect 41568 252442 41937 252444
rect 41568 252386 41876 252442
rect 41932 252386 41937 252442
rect 41568 252384 41937 252386
rect 41871 252381 41937 252384
rect 40770 251706 40830 251970
rect 40762 251642 40768 251706
rect 40832 251642 40838 251706
rect 189903 251704 189969 251707
rect 189903 251702 191904 251704
rect 189903 251646 189908 251702
rect 189964 251646 191904 251702
rect 189903 251644 191904 251646
rect 189903 251641 189969 251644
rect 41346 251114 41406 251452
rect 41146 251050 41152 251114
rect 41216 251050 41222 251114
rect 41338 251050 41344 251114
rect 41408 251050 41414 251114
rect 41154 250934 41214 251050
rect 41775 250520 41841 250523
rect 420303 250520 420369 250523
rect 41568 250518 41841 250520
rect 41568 250462 41780 250518
rect 41836 250462 41841 250518
rect 41568 250460 41841 250462
rect 412512 250518 420369 250520
rect 412512 250462 420308 250518
rect 420364 250462 420369 250518
rect 412512 250460 420369 250462
rect 41775 250457 41841 250460
rect 420303 250457 420369 250460
rect 41538 249783 41598 249898
rect 41538 249778 41649 249783
rect 41538 249722 41588 249778
rect 41644 249722 41649 249778
rect 41538 249720 41649 249722
rect 41583 249717 41649 249720
rect 675759 249632 675825 249635
rect 675898 249632 675904 249634
rect 675759 249630 675904 249632
rect 675759 249574 675764 249630
rect 675820 249574 675904 249630
rect 675759 249572 675904 249574
rect 675759 249569 675825 249572
rect 675898 249570 675904 249572
rect 675968 249570 675974 249634
rect 41538 249191 41598 249454
rect 41538 249186 41649 249191
rect 41538 249130 41588 249186
rect 41644 249130 41649 249186
rect 41538 249128 41649 249130
rect 41583 249125 41649 249128
rect 41967 249040 42033 249043
rect 41568 249038 42033 249040
rect 41568 248982 41972 249038
rect 42028 248982 42033 249038
rect 41568 248980 42033 248982
rect 41967 248977 42033 248980
rect 41538 248303 41598 248418
rect 41538 248298 41649 248303
rect 41538 248242 41588 248298
rect 41644 248242 41649 248298
rect 41538 248240 41649 248242
rect 41583 248237 41649 248240
rect 420399 248152 420465 248155
rect 412512 248150 420465 248152
rect 412512 248094 420404 248150
rect 420460 248094 420465 248150
rect 412512 248092 420465 248094
rect 420399 248089 420465 248092
rect 41538 247711 41598 247900
rect 41538 247706 41649 247711
rect 41538 247650 41588 247706
rect 41644 247650 41649 247706
rect 41538 247648 41649 247650
rect 41583 247645 41649 247648
rect 675663 247562 675729 247563
rect 675663 247558 675712 247562
rect 675776 247560 675782 247562
rect 41538 247267 41598 247530
rect 675663 247502 675668 247558
rect 675663 247498 675712 247502
rect 675776 247500 675820 247560
rect 675776 247498 675782 247500
rect 675663 247497 675729 247498
rect 41538 247262 41649 247267
rect 41538 247206 41588 247262
rect 41644 247206 41649 247262
rect 41538 247204 41649 247206
rect 41583 247201 41649 247204
rect 41538 246672 41598 246938
rect 41679 246672 41745 246675
rect 41538 246670 41745 246672
rect 41538 246614 41684 246670
rect 41740 246614 41745 246670
rect 41538 246612 41745 246614
rect 41679 246609 41745 246612
rect 675759 246672 675825 246675
rect 676282 246672 676288 246674
rect 675759 246670 676288 246672
rect 675759 246614 675764 246670
rect 675820 246614 676288 246670
rect 675759 246612 676288 246614
rect 675759 246609 675825 246612
rect 676282 246610 676288 246612
rect 676352 246610 676358 246674
rect 675759 245932 675825 245935
rect 676090 245932 676096 245934
rect 675759 245930 676096 245932
rect 675759 245874 675764 245930
rect 675820 245874 676096 245930
rect 675759 245872 676096 245874
rect 675759 245869 675825 245872
rect 676090 245870 676096 245872
rect 676160 245870 676166 245934
rect 412482 245340 412542 245828
rect 420399 245340 420465 245343
rect 412482 245338 420465 245340
rect 412482 245282 420404 245338
rect 420460 245282 420465 245338
rect 412482 245280 420465 245282
rect 420399 245277 420465 245280
rect 149391 244600 149457 244603
rect 143904 244598 149457 244600
rect 143904 244542 149396 244598
rect 149452 244542 149457 244598
rect 143904 244540 149457 244542
rect 149391 244537 149457 244540
rect 148324 243416 148330 243418
rect 143904 243356 148330 243416
rect 148324 243354 148330 243356
rect 148394 243354 148400 243418
rect 187119 243416 187185 243419
rect 191874 243416 191934 243904
rect 420399 243564 420465 243567
rect 412512 243562 420465 243564
rect 412512 243506 420404 243562
rect 420460 243506 420465 243562
rect 412512 243504 420465 243506
rect 420399 243501 420465 243504
rect 673978 243502 673984 243566
rect 674048 243564 674054 243566
rect 675471 243564 675537 243567
rect 674048 243562 675537 243564
rect 674048 243506 675476 243562
rect 675532 243506 675537 243562
rect 674048 243504 675537 243506
rect 674048 243502 674054 243504
rect 675471 243501 675537 243504
rect 187119 243414 191934 243416
rect 187119 243358 187124 243414
rect 187180 243358 191934 243414
rect 187119 243356 191934 243358
rect 187119 243353 187185 243356
rect 143874 242084 143934 242128
rect 148239 242084 148305 242087
rect 143874 242082 148305 242084
rect 143874 242026 148244 242082
rect 148300 242026 148305 242082
rect 143874 242024 148305 242026
rect 148239 242021 148305 242024
rect 675130 241874 675136 241938
rect 675200 241936 675206 241938
rect 675279 241936 675345 241939
rect 675200 241934 675345 241936
rect 675200 241878 675284 241934
rect 675340 241878 675345 241934
rect 675200 241876 675345 241878
rect 675200 241874 675206 241876
rect 675279 241873 675345 241876
rect 420399 241196 420465 241199
rect 412512 241194 420465 241196
rect 412512 241138 420404 241194
rect 420460 241138 420465 241194
rect 412512 241136 420465 241138
rect 420399 241133 420465 241136
rect 148719 240900 148785 240903
rect 143904 240898 148785 240900
rect 143904 240842 148724 240898
rect 148780 240842 148785 240898
rect 143904 240840 148785 240842
rect 148719 240837 148785 240840
rect 674938 240542 674944 240606
rect 675008 240604 675014 240606
rect 675471 240604 675537 240607
rect 675008 240602 675537 240604
rect 675008 240546 675476 240602
rect 675532 240546 675537 240602
rect 675008 240544 675537 240546
rect 675008 240542 675014 240544
rect 675471 240541 675537 240544
rect 149391 239716 149457 239719
rect 143904 239714 149457 239716
rect 143904 239658 149396 239714
rect 149452 239658 149457 239714
rect 143904 239656 149457 239658
rect 149391 239653 149457 239656
rect 413391 238976 413457 238979
rect 555375 238976 555441 238979
rect 413391 238974 555441 238976
rect 413391 238918 413396 238974
rect 413452 238918 555380 238974
rect 555436 238918 555441 238974
rect 413391 238916 555441 238918
rect 413391 238913 413457 238916
rect 555375 238913 555441 238916
rect 413679 238680 413745 238683
rect 557007 238680 557073 238683
rect 413679 238678 557073 238680
rect 413679 238622 413684 238678
rect 413740 238622 557012 238678
rect 557068 238622 557073 238678
rect 413679 238620 557073 238622
rect 413679 238617 413745 238620
rect 557007 238617 557073 238620
rect 148527 238532 148593 238535
rect 143904 238530 148593 238532
rect 143904 238474 148532 238530
rect 148588 238474 148593 238530
rect 143904 238472 148593 238474
rect 148527 238469 148593 238472
rect 41775 238386 41841 238387
rect 41722 238384 41728 238386
rect 41684 238324 41728 238384
rect 41792 238382 41841 238386
rect 41836 238326 41841 238382
rect 41722 238322 41728 238324
rect 41792 238322 41841 238326
rect 41775 238321 41841 238322
rect 413967 238384 414033 238387
rect 553935 238384 554001 238387
rect 413967 238382 554001 238384
rect 413967 238326 413972 238382
rect 414028 238326 553940 238382
rect 553996 238326 554001 238382
rect 413967 238324 554001 238326
rect 413967 238321 414033 238324
rect 553935 238321 554001 238324
rect 674554 238174 674560 238238
rect 674624 238236 674630 238238
rect 675279 238236 675345 238239
rect 674624 238234 675345 238236
rect 674624 238178 675284 238234
rect 675340 238178 675345 238234
rect 674624 238176 675345 238178
rect 674624 238174 674630 238176
rect 675279 238173 675345 238176
rect 143874 236756 143934 237244
rect 377967 237052 378033 237055
rect 388623 237052 388689 237055
rect 576015 237052 576081 237055
rect 377967 237050 388689 237052
rect 377967 236994 377972 237050
rect 378028 236994 388628 237050
rect 388684 236994 388689 237050
rect 377967 236992 388689 236994
rect 377967 236989 378033 236992
rect 388623 236989 388689 236992
rect 390018 237050 576081 237052
rect 390018 236994 576020 237050
rect 576076 236994 576081 237050
rect 390018 236992 576081 236994
rect 373455 236904 373521 236907
rect 383823 236904 383889 236907
rect 373455 236902 383889 236904
rect 373455 236846 373460 236902
rect 373516 236846 383828 236902
rect 383884 236846 383889 236902
rect 373455 236844 383889 236846
rect 373455 236841 373521 236844
rect 383823 236841 383889 236844
rect 384015 236904 384081 236907
rect 390018 236904 390078 236992
rect 576015 236989 576081 236992
rect 570255 236904 570321 236907
rect 384015 236902 390078 236904
rect 384015 236846 384020 236902
rect 384076 236846 390078 236902
rect 384015 236844 390078 236846
rect 390210 236902 570321 236904
rect 390210 236846 570260 236902
rect 570316 236846 570321 236902
rect 390210 236844 570321 236846
rect 384015 236841 384081 236844
rect 148335 236756 148401 236759
rect 143874 236754 148401 236756
rect 143874 236698 148340 236754
rect 148396 236698 148401 236754
rect 143874 236696 148401 236698
rect 148335 236693 148401 236696
rect 381231 236756 381297 236759
rect 390210 236756 390270 236844
rect 570255 236841 570321 236844
rect 674746 236842 674752 236906
rect 674816 236904 674822 236906
rect 675375 236904 675441 236907
rect 674816 236902 675441 236904
rect 674816 236846 675380 236902
rect 675436 236846 675441 236902
rect 674816 236844 675441 236846
rect 674816 236842 674822 236844
rect 675375 236841 675441 236844
rect 381231 236754 390270 236756
rect 381231 236698 381236 236754
rect 381292 236698 390270 236754
rect 381231 236696 390270 236698
rect 390351 236756 390417 236759
rect 567375 236756 567441 236759
rect 390351 236754 567441 236756
rect 390351 236698 390356 236754
rect 390412 236698 567380 236754
rect 567436 236698 567441 236754
rect 390351 236696 567441 236698
rect 381231 236693 381297 236696
rect 390351 236693 390417 236696
rect 567375 236693 567441 236696
rect 380847 236608 380913 236611
rect 388815 236608 388881 236611
rect 380847 236606 388881 236608
rect 380847 236550 380852 236606
rect 380908 236550 388820 236606
rect 388876 236550 388881 236606
rect 380847 236548 388881 236550
rect 380847 236545 380913 236548
rect 388815 236545 388881 236548
rect 389007 236608 389073 236611
rect 565263 236608 565329 236611
rect 389007 236606 565329 236608
rect 389007 236550 389012 236606
rect 389068 236550 565268 236606
rect 565324 236550 565329 236606
rect 389007 236548 565329 236550
rect 389007 236545 389073 236548
rect 565263 236545 565329 236548
rect 376719 236460 376785 236463
rect 562191 236460 562257 236463
rect 376719 236458 562257 236460
rect 376719 236402 376724 236458
rect 376780 236402 562196 236458
rect 562252 236402 562257 236458
rect 376719 236400 562257 236402
rect 376719 236397 376785 236400
rect 562191 236397 562257 236400
rect 372207 236312 372273 236315
rect 388527 236312 388593 236315
rect 372207 236310 388593 236312
rect 372207 236254 372212 236310
rect 372268 236254 388532 236310
rect 388588 236254 388593 236310
rect 372207 236252 388593 236254
rect 372207 236249 372273 236252
rect 388527 236249 388593 236252
rect 388719 236312 388785 236315
rect 556143 236312 556209 236315
rect 388719 236310 556209 236312
rect 388719 236254 388724 236310
rect 388780 236254 556148 236310
rect 556204 236254 556209 236310
rect 388719 236252 556209 236254
rect 388719 236249 388785 236252
rect 556143 236249 556209 236252
rect 336783 236164 336849 236167
rect 471279 236164 471345 236167
rect 336783 236162 471345 236164
rect 336783 236106 336788 236162
rect 336844 236106 471284 236162
rect 471340 236106 471345 236162
rect 336783 236104 471345 236106
rect 336783 236101 336849 236104
rect 471279 236101 471345 236104
rect 149007 236016 149073 236019
rect 143904 236014 149073 236016
rect 143904 235958 149012 236014
rect 149068 235958 149073 236014
rect 143904 235956 149073 235958
rect 149007 235953 149073 235956
rect 344367 236016 344433 236019
rect 394479 236016 394545 236019
rect 344367 236014 394545 236016
rect 344367 235958 344372 236014
rect 344428 235958 394484 236014
rect 394540 235958 394545 236014
rect 344367 235956 394545 235958
rect 344367 235953 344433 235956
rect 394479 235953 394545 235956
rect 399087 236016 399153 236019
rect 564399 236016 564465 236019
rect 399087 236014 564465 236016
rect 399087 235958 399092 236014
rect 399148 235958 564404 236014
rect 564460 235958 564465 236014
rect 399087 235956 564465 235958
rect 399087 235953 399153 235956
rect 564399 235953 564465 235956
rect 376335 235868 376401 235871
rect 559887 235868 559953 235871
rect 376335 235866 559953 235868
rect 376335 235810 376340 235866
rect 376396 235810 559892 235866
rect 559948 235810 559953 235866
rect 376335 235808 559953 235810
rect 376335 235805 376401 235808
rect 559887 235805 559953 235808
rect 385743 235720 385809 235723
rect 579567 235720 579633 235723
rect 385743 235718 579633 235720
rect 385743 235662 385748 235718
rect 385804 235662 579572 235718
rect 579628 235662 579633 235718
rect 385743 235660 579633 235662
rect 385743 235657 385809 235660
rect 579567 235657 579633 235660
rect 395343 235572 395409 235575
rect 588975 235572 589041 235575
rect 395343 235570 589041 235572
rect 395343 235514 395348 235570
rect 395404 235514 588980 235570
rect 589036 235514 589041 235570
rect 395343 235512 589041 235514
rect 395343 235509 395409 235512
rect 588975 235509 589041 235512
rect 359439 235424 359505 235427
rect 403215 235424 403281 235427
rect 359439 235422 403281 235424
rect 359439 235366 359444 235422
rect 359500 235366 403220 235422
rect 403276 235366 403281 235422
rect 359439 235364 403281 235366
rect 359439 235361 359505 235364
rect 403215 235361 403281 235364
rect 411375 235424 411441 235427
rect 609135 235424 609201 235427
rect 411375 235422 609201 235424
rect 411375 235366 411380 235422
rect 411436 235366 609140 235422
rect 609196 235366 609201 235422
rect 411375 235364 609201 235366
rect 411375 235361 411441 235364
rect 609135 235361 609201 235364
rect 394095 235276 394161 235279
rect 596271 235276 596337 235279
rect 394095 235274 596337 235276
rect 394095 235218 394100 235274
rect 394156 235218 596276 235274
rect 596332 235218 596337 235274
rect 394095 235216 596337 235218
rect 394095 235213 394161 235216
rect 596271 235213 596337 235216
rect 402159 235128 402225 235131
rect 612783 235128 612849 235131
rect 402159 235126 612849 235128
rect 402159 235070 402164 235126
rect 402220 235070 612788 235126
rect 612844 235070 612849 235126
rect 402159 235068 612849 235070
rect 402159 235065 402225 235068
rect 612783 235065 612849 235068
rect 353487 234980 353553 234983
rect 403215 234980 403281 234983
rect 353487 234978 403281 234980
rect 353487 234922 353492 234978
rect 353548 234922 403220 234978
rect 403276 234922 403281 234978
rect 353487 234920 403281 234922
rect 353487 234917 353553 234920
rect 403215 234917 403281 234920
rect 405423 234980 405489 234983
rect 618831 234980 618897 234983
rect 405423 234978 618897 234980
rect 405423 234922 405428 234978
rect 405484 234922 618836 234978
rect 618892 234922 618897 234978
rect 405423 234920 618897 234922
rect 405423 234917 405489 234920
rect 618831 234917 618897 234920
rect 149391 234832 149457 234835
rect 143904 234830 149457 234832
rect 143904 234774 149396 234830
rect 149452 234774 149457 234830
rect 143904 234772 149457 234774
rect 149391 234769 149457 234772
rect 404367 234832 404433 234835
rect 617295 234832 617361 234835
rect 404367 234830 617361 234832
rect 404367 234774 404372 234830
rect 404428 234774 617300 234830
rect 617356 234774 617361 234830
rect 404367 234772 617361 234774
rect 404367 234769 404433 234772
rect 617295 234769 617361 234772
rect 342543 234684 342609 234687
rect 400623 234684 400689 234687
rect 342543 234682 400689 234684
rect 342543 234626 342548 234682
rect 342604 234626 400628 234682
rect 400684 234626 400689 234682
rect 342543 234624 400689 234626
rect 342543 234621 342609 234624
rect 400623 234621 400689 234624
rect 405903 234684 405969 234687
rect 620367 234684 620433 234687
rect 405903 234682 620433 234684
rect 405903 234626 405908 234682
rect 405964 234626 620372 234682
rect 620428 234626 620433 234682
rect 405903 234624 620433 234626
rect 405903 234621 405969 234624
rect 620367 234621 620433 234624
rect 362511 234536 362577 234539
rect 404751 234536 404817 234539
rect 362511 234534 404817 234536
rect 362511 234478 362516 234534
rect 362572 234478 404756 234534
rect 404812 234478 404817 234534
rect 362511 234476 404817 234478
rect 362511 234473 362577 234476
rect 404751 234473 404817 234476
rect 404943 234536 405009 234539
rect 516207 234536 516273 234539
rect 404943 234534 516273 234536
rect 404943 234478 404948 234534
rect 405004 234478 516212 234534
rect 516268 234478 516273 234534
rect 404943 234476 516273 234478
rect 404943 234473 405009 234476
rect 516207 234473 516273 234476
rect 379119 234388 379185 234391
rect 397359 234388 397425 234391
rect 379119 234386 397425 234388
rect 379119 234330 379124 234386
rect 379180 234330 397364 234386
rect 397420 234330 397425 234386
rect 379119 234328 397425 234330
rect 379119 234325 379185 234328
rect 397359 234325 397425 234328
rect 402735 234388 402801 234391
rect 501039 234388 501105 234391
rect 402735 234386 501105 234388
rect 402735 234330 402740 234386
rect 402796 234330 501044 234386
rect 501100 234330 501105 234386
rect 402735 234328 501105 234330
rect 402735 234325 402801 234328
rect 501039 234325 501105 234328
rect 382095 234240 382161 234243
rect 416943 234240 417009 234243
rect 382095 234238 417009 234240
rect 382095 234182 382100 234238
rect 382156 234182 416948 234238
rect 417004 234182 417009 234238
rect 382095 234180 417009 234182
rect 382095 234177 382161 234180
rect 416943 234177 417009 234180
rect 368559 234092 368625 234095
rect 411663 234092 411729 234095
rect 368559 234090 411729 234092
rect 368559 234034 368564 234090
rect 368620 234034 411668 234090
rect 411724 234034 411729 234090
rect 368559 234032 411729 234034
rect 368559 234029 368625 234032
rect 411663 234029 411729 234032
rect 148431 233648 148497 233651
rect 143904 233646 148497 233648
rect 143904 233590 148436 233646
rect 148492 233590 148497 233646
rect 143904 233588 148497 233590
rect 148431 233585 148497 233588
rect 41530 233290 41536 233354
rect 41600 233352 41606 233354
rect 41775 233352 41841 233355
rect 41600 233350 41841 233352
rect 41600 233294 41780 233350
rect 41836 233294 41841 233350
rect 41600 233292 41841 233294
rect 41600 233290 41606 233292
rect 41775 233289 41841 233292
rect 344751 233352 344817 233355
rect 362799 233352 362865 233355
rect 344751 233350 362865 233352
rect 344751 233294 344756 233350
rect 344812 233294 362804 233350
rect 362860 233294 362865 233350
rect 344751 233292 362865 233294
rect 344751 233289 344817 233292
rect 362799 233289 362865 233292
rect 339375 233204 339441 233207
rect 488271 233204 488337 233207
rect 339375 233202 488337 233204
rect 339375 233146 339380 233202
rect 339436 233146 488276 233202
rect 488332 233146 488337 233202
rect 339375 233144 488337 233146
rect 339375 233141 339441 233144
rect 488271 233141 488337 233144
rect 342159 233056 342225 233059
rect 494223 233056 494289 233059
rect 342159 233054 494289 233056
rect 342159 232998 342164 233054
rect 342220 232998 494228 233054
rect 494284 232998 494289 233054
rect 342159 232996 494289 232998
rect 342159 232993 342225 232996
rect 494223 232993 494289 232996
rect 397359 232908 397425 232911
rect 565935 232908 566001 232911
rect 397359 232906 566001 232908
rect 397359 232850 397364 232906
rect 397420 232850 565940 232906
rect 565996 232850 566001 232906
rect 397359 232848 566001 232850
rect 397359 232845 397425 232848
rect 565935 232845 566001 232848
rect 374319 232760 374385 232763
rect 555471 232760 555537 232763
rect 374319 232758 555537 232760
rect 374319 232702 374324 232758
rect 374380 232702 555476 232758
rect 555532 232702 555537 232758
rect 374319 232700 555537 232702
rect 374319 232697 374385 232700
rect 555471 232697 555537 232700
rect 374031 232612 374097 232615
rect 557679 232612 557745 232615
rect 374031 232610 557745 232612
rect 374031 232554 374036 232610
rect 374092 232554 557684 232610
rect 557740 232554 557745 232610
rect 374031 232552 557745 232554
rect 374031 232549 374097 232552
rect 557679 232549 557745 232552
rect 380463 232464 380529 232467
rect 567471 232464 567537 232467
rect 380463 232462 567537 232464
rect 380463 232406 380468 232462
rect 380524 232406 567476 232462
rect 567532 232406 567537 232462
rect 380463 232404 567537 232406
rect 380463 232401 380529 232404
rect 567471 232401 567537 232404
rect 149199 232316 149265 232319
rect 143904 232314 149265 232316
rect 143904 232258 149204 232314
rect 149260 232258 149265 232314
rect 143904 232256 149265 232258
rect 149199 232253 149265 232256
rect 383535 232316 383601 232319
rect 573519 232316 573585 232319
rect 383535 232314 573585 232316
rect 383535 232258 383540 232314
rect 383596 232258 573524 232314
rect 573580 232258 573585 232314
rect 383535 232256 573585 232258
rect 383535 232253 383601 232256
rect 573519 232253 573585 232256
rect 381327 232168 381393 232171
rect 572751 232168 572817 232171
rect 381327 232166 572817 232168
rect 381327 232110 381332 232166
rect 381388 232110 572756 232166
rect 572812 232110 572817 232166
rect 381327 232108 572817 232110
rect 381327 232105 381393 232108
rect 572751 232105 572817 232108
rect 379887 232020 379953 232023
rect 569775 232020 569841 232023
rect 379887 232018 569841 232020
rect 379887 231962 379892 232018
rect 379948 231962 569780 232018
rect 569836 231962 569841 232018
rect 379887 231960 569841 231962
rect 379887 231957 379953 231960
rect 569775 231957 569841 231960
rect 398895 231872 398961 231875
rect 605967 231872 606033 231875
rect 398895 231870 606033 231872
rect 398895 231814 398900 231870
rect 398956 231814 605972 231870
rect 606028 231814 606033 231870
rect 398895 231812 606033 231814
rect 398895 231809 398961 231812
rect 605967 231809 606033 231812
rect 327087 231724 327153 231727
rect 464079 231724 464145 231727
rect 327087 231722 464145 231724
rect 327087 231666 327092 231722
rect 327148 231666 464084 231722
rect 464140 231666 464145 231722
rect 327087 231664 464145 231666
rect 327087 231661 327153 231664
rect 464079 231661 464145 231664
rect 324015 231576 324081 231579
rect 458031 231576 458097 231579
rect 324015 231574 458097 231576
rect 324015 231518 324020 231574
rect 324076 231518 458036 231574
rect 458092 231518 458097 231574
rect 324015 231516 458097 231518
rect 324015 231513 324081 231516
rect 458031 231513 458097 231516
rect 319503 231428 319569 231431
rect 448911 231428 448977 231431
rect 319503 231426 448977 231428
rect 319503 231370 319508 231426
rect 319564 231370 448916 231426
rect 448972 231370 448977 231426
rect 319503 231368 448977 231370
rect 319503 231365 319569 231368
rect 448911 231365 448977 231368
rect 316719 231280 316785 231283
rect 442863 231280 442929 231283
rect 316719 231278 442929 231280
rect 316719 231222 316724 231278
rect 316780 231222 442868 231278
rect 442924 231222 442929 231278
rect 316719 231220 442929 231222
rect 316719 231217 316785 231220
rect 442863 231217 442929 231220
rect 148623 231132 148689 231135
rect 143904 231130 148689 231132
rect 143904 231074 148628 231130
rect 148684 231074 148689 231130
rect 143904 231072 148689 231074
rect 148623 231069 148689 231072
rect 41146 230330 41152 230394
rect 41216 230392 41222 230394
rect 41775 230392 41841 230395
rect 41216 230390 41841 230392
rect 41216 230334 41780 230390
rect 41836 230334 41841 230390
rect 41216 230332 41841 230334
rect 41216 230330 41222 230332
rect 41775 230329 41841 230332
rect 348783 230392 348849 230395
rect 504015 230392 504081 230395
rect 348783 230390 504081 230392
rect 348783 230334 348788 230390
rect 348844 230334 504020 230390
rect 504076 230334 504081 230390
rect 348783 230332 504081 230334
rect 348783 230329 348849 230332
rect 504015 230329 504081 230332
rect 356271 230244 356337 230247
rect 519183 230244 519249 230247
rect 356271 230242 519249 230244
rect 356271 230186 356276 230242
rect 356332 230186 519188 230242
rect 519244 230186 519249 230242
rect 356271 230184 519249 230186
rect 356271 230181 356337 230184
rect 519183 230181 519249 230184
rect 359055 230096 359121 230099
rect 525231 230096 525297 230099
rect 359055 230094 525297 230096
rect 359055 230038 359060 230094
rect 359116 230038 525236 230094
rect 525292 230038 525297 230094
rect 359055 230036 525297 230038
rect 359055 230033 359121 230036
rect 525231 230033 525297 230036
rect 146895 229948 146961 229951
rect 143904 229946 146961 229948
rect 143904 229890 146900 229946
rect 146956 229890 146961 229946
rect 143904 229888 146961 229890
rect 146895 229885 146961 229888
rect 361743 229948 361809 229951
rect 533487 229948 533553 229951
rect 361743 229946 533553 229948
rect 361743 229890 361748 229946
rect 361804 229890 533492 229946
rect 533548 229890 533553 229946
rect 361743 229888 533553 229890
rect 361743 229885 361809 229888
rect 533487 229885 533553 229888
rect 41338 229738 41344 229802
rect 41408 229800 41414 229802
rect 41775 229800 41841 229803
rect 41408 229798 41841 229800
rect 41408 229742 41780 229798
rect 41836 229742 41841 229798
rect 41408 229740 41841 229742
rect 41408 229738 41414 229740
rect 41775 229737 41841 229740
rect 371151 229800 371217 229803
rect 549423 229800 549489 229803
rect 371151 229798 549489 229800
rect 371151 229742 371156 229798
rect 371212 229742 549428 229798
rect 549484 229742 549489 229798
rect 371151 229740 549489 229742
rect 371151 229737 371217 229740
rect 549423 229737 549489 229740
rect 398799 229652 398865 229655
rect 578895 229652 578961 229655
rect 398799 229650 578961 229652
rect 398799 229594 398804 229650
rect 398860 229594 578900 229650
rect 578956 229594 578961 229650
rect 398799 229592 578961 229594
rect 398799 229589 398865 229592
rect 578895 229589 578961 229592
rect 381711 229504 381777 229507
rect 570447 229504 570513 229507
rect 381711 229502 570513 229504
rect 381711 229446 381716 229502
rect 381772 229446 570452 229502
rect 570508 229446 570513 229502
rect 381711 229444 570513 229446
rect 381711 229441 381777 229444
rect 570447 229441 570513 229444
rect 383631 229356 383697 229359
rect 575055 229356 575121 229359
rect 383631 229354 575121 229356
rect 383631 229298 383636 229354
rect 383692 229298 575060 229354
rect 575116 229298 575121 229354
rect 383631 229296 575121 229298
rect 383631 229293 383697 229296
rect 575055 229293 575121 229296
rect 384975 229208 385041 229211
rect 576591 229208 576657 229211
rect 384975 229206 576657 229208
rect 384975 229150 384980 229206
rect 385036 229150 576596 229206
rect 576652 229150 576657 229206
rect 384975 229148 576657 229150
rect 384975 229145 385041 229148
rect 576591 229145 576657 229148
rect 40954 228998 40960 229062
rect 41024 229060 41030 229062
rect 41775 229060 41841 229063
rect 41024 229058 41841 229060
rect 41024 229002 41780 229058
rect 41836 229002 41841 229058
rect 41024 229000 41841 229002
rect 41024 228998 41030 229000
rect 41775 228997 41841 229000
rect 395919 229060 395985 229063
rect 599919 229060 599985 229063
rect 395919 229058 599985 229060
rect 395919 229002 395924 229058
rect 395980 229002 599924 229058
rect 599980 229002 599985 229058
rect 395919 229000 599985 229002
rect 395919 228997 395985 229000
rect 599919 228997 599985 229000
rect 332463 228912 332529 228915
rect 338703 228912 338769 228915
rect 332463 228910 338769 228912
rect 332463 228854 332468 228910
rect 332524 228854 338708 228910
rect 338764 228854 338769 228910
rect 332463 228852 338769 228854
rect 332463 228849 332529 228852
rect 338703 228849 338769 228852
rect 403983 228912 404049 228915
rect 616623 228912 616689 228915
rect 403983 228910 616689 228912
rect 403983 228854 403988 228910
rect 404044 228854 616628 228910
rect 616684 228854 616689 228910
rect 403983 228852 616689 228854
rect 403983 228849 404049 228852
rect 616623 228849 616689 228852
rect 314895 228764 314961 228767
rect 439983 228764 440049 228767
rect 314895 228762 440049 228764
rect 314895 228706 314900 228762
rect 314956 228706 439988 228762
rect 440044 228706 440049 228762
rect 314895 228704 440049 228706
rect 314895 228701 314961 228704
rect 439983 228701 440049 228704
rect 143874 228172 143934 228660
rect 310671 228616 310737 228619
rect 430863 228616 430929 228619
rect 310671 228614 430929 228616
rect 310671 228558 310676 228614
rect 310732 228558 430868 228614
rect 430924 228558 430929 228614
rect 310671 228556 430929 228558
rect 310671 228553 310737 228556
rect 430863 228553 430929 228556
rect 302895 228468 302961 228471
rect 415695 228468 415761 228471
rect 302895 228466 415761 228468
rect 302895 228410 302900 228466
rect 302956 228410 415700 228466
rect 415756 228410 415761 228466
rect 302895 228408 415761 228410
rect 302895 228405 302961 228408
rect 415695 228405 415761 228408
rect 411663 228320 411729 228323
rect 415407 228320 415473 228323
rect 411663 228318 415473 228320
rect 411663 228262 411668 228318
rect 411724 228262 415412 228318
rect 415468 228262 415473 228318
rect 411663 228260 415473 228262
rect 411663 228257 411729 228260
rect 415407 228257 415473 228260
rect 146991 228172 147057 228175
rect 143874 228170 147057 228172
rect 143874 228114 146996 228170
rect 147052 228114 147057 228170
rect 143874 228112 147057 228114
rect 146991 228109 147057 228112
rect 40570 227370 40576 227434
rect 40640 227432 40646 227434
rect 41871 227432 41937 227435
rect 149391 227432 149457 227435
rect 40640 227430 41937 227432
rect 40640 227374 41876 227430
rect 41932 227374 41937 227430
rect 40640 227372 41937 227374
rect 143904 227430 149457 227432
rect 143904 227374 149396 227430
rect 149452 227374 149457 227430
rect 143904 227372 149457 227374
rect 40640 227370 40646 227372
rect 41871 227369 41937 227372
rect 149391 227369 149457 227372
rect 335343 227432 335409 227435
rect 478383 227432 478449 227435
rect 335343 227430 478449 227432
rect 335343 227374 335348 227430
rect 335404 227374 478388 227430
rect 478444 227374 478449 227430
rect 335343 227372 478449 227374
rect 335343 227369 335409 227372
rect 478383 227369 478449 227372
rect 338607 227284 338673 227287
rect 484431 227284 484497 227287
rect 338607 227282 484497 227284
rect 338607 227226 338612 227282
rect 338668 227226 484436 227282
rect 484492 227226 484497 227282
rect 338607 227224 484497 227226
rect 338607 227221 338673 227224
rect 484431 227221 484497 227224
rect 348687 227136 348753 227139
rect 495759 227136 495825 227139
rect 348687 227134 495825 227136
rect 348687 227078 348692 227134
rect 348748 227078 495764 227134
rect 495820 227078 495825 227134
rect 348687 227076 495825 227078
rect 348687 227073 348753 227076
rect 495759 227073 495825 227076
rect 341583 226988 341649 226991
rect 490479 226988 490545 226991
rect 341583 226986 490545 226988
rect 341583 226930 341588 226986
rect 341644 226930 490484 226986
rect 490540 226930 490545 226986
rect 341583 226928 490545 226930
rect 341583 226925 341649 226928
rect 490479 226925 490545 226928
rect 40762 226778 40768 226842
rect 40832 226840 40838 226842
rect 41775 226840 41841 226843
rect 40832 226838 41841 226840
rect 40832 226782 41780 226838
rect 41836 226782 41841 226838
rect 40832 226780 41841 226782
rect 40832 226778 40838 226780
rect 41775 226777 41841 226780
rect 356847 226840 356913 226843
rect 522927 226840 522993 226843
rect 356847 226838 522993 226840
rect 356847 226782 356852 226838
rect 356908 226782 522932 226838
rect 522988 226782 522993 226838
rect 356847 226780 522993 226782
rect 356847 226777 356913 226780
rect 522927 226777 522993 226780
rect 393423 226692 393489 226695
rect 595407 226692 595473 226695
rect 393423 226690 595473 226692
rect 393423 226634 393428 226690
rect 393484 226634 595412 226690
rect 595468 226634 595473 226690
rect 393423 226632 595473 226634
rect 393423 226629 393489 226632
rect 595407 226629 595473 226632
rect 391599 226544 391665 226547
rect 591663 226544 591729 226547
rect 391599 226542 591729 226544
rect 391599 226486 391604 226542
rect 391660 226486 591668 226542
rect 591724 226486 591729 226542
rect 391599 226484 591729 226486
rect 391599 226481 391665 226484
rect 591663 226481 591729 226484
rect 148815 226396 148881 226399
rect 143904 226394 148881 226396
rect 143904 226338 148820 226394
rect 148876 226338 148881 226394
rect 143904 226336 148881 226338
rect 148815 226333 148881 226336
rect 396783 226396 396849 226399
rect 602223 226396 602289 226399
rect 396783 226394 602289 226396
rect 396783 226338 396788 226394
rect 396844 226338 602228 226394
rect 602284 226338 602289 226394
rect 396783 226336 602289 226338
rect 396783 226333 396849 226336
rect 602223 226333 602289 226336
rect 41967 226250 42033 226251
rect 41914 226248 41920 226250
rect 41876 226188 41920 226248
rect 41984 226246 42033 226250
rect 42028 226190 42033 226246
rect 41914 226186 41920 226188
rect 41984 226186 42033 226190
rect 41967 226185 42033 226186
rect 408111 226248 408177 226251
rect 624879 226248 624945 226251
rect 408111 226246 624945 226248
rect 408111 226190 408116 226246
rect 408172 226190 624884 226246
rect 624940 226190 624945 226246
rect 408111 226188 624945 226190
rect 408111 226185 408177 226188
rect 624879 226185 624945 226188
rect 408495 226100 408561 226103
rect 625551 226100 625617 226103
rect 408495 226098 625617 226100
rect 408495 226042 408500 226098
rect 408556 226042 625556 226098
rect 625612 226042 625617 226098
rect 408495 226040 625617 226042
rect 408495 226037 408561 226040
rect 625551 226037 625617 226040
rect 332559 225952 332625 225955
rect 472335 225952 472401 225955
rect 332559 225950 472401 225952
rect 332559 225894 332564 225950
rect 332620 225894 472340 225950
rect 472396 225894 472401 225950
rect 332559 225892 472401 225894
rect 332559 225889 332625 225892
rect 472335 225889 472401 225892
rect 330831 225804 330897 225807
rect 469359 225804 469425 225807
rect 330831 225802 469425 225804
rect 330831 225746 330836 225802
rect 330892 225746 469364 225802
rect 469420 225746 469425 225802
rect 330831 225744 469425 225746
rect 330831 225741 330897 225744
rect 469359 225741 469425 225744
rect 328047 225656 328113 225659
rect 463311 225656 463377 225659
rect 328047 225654 463377 225656
rect 328047 225598 328052 225654
rect 328108 225598 463316 225654
rect 463372 225598 463377 225654
rect 328047 225596 463377 225598
rect 328047 225593 328113 225596
rect 463311 225593 463377 225596
rect 324783 225508 324849 225511
rect 457263 225508 457329 225511
rect 324783 225506 457329 225508
rect 324783 225450 324788 225506
rect 324844 225450 457268 225506
rect 457324 225450 457329 225506
rect 324783 225448 457329 225450
rect 324783 225445 324849 225448
rect 457263 225445 457329 225448
rect 149103 225212 149169 225215
rect 143904 225210 149169 225212
rect 143904 225154 149108 225210
rect 149164 225154 149169 225210
rect 143904 225152 149169 225154
rect 149103 225149 149169 225152
rect 676239 225064 676305 225067
rect 676239 225062 676350 225064
rect 676239 225006 676244 225062
rect 676300 225006 676350 225062
rect 676239 225001 676350 225006
rect 676290 224886 676350 225001
rect 358959 224620 359025 224623
rect 527535 224620 527601 224623
rect 358959 224618 527601 224620
rect 358959 224562 358964 224618
rect 359020 224562 527540 224618
rect 527596 224562 527601 224618
rect 358959 224560 527601 224562
rect 358959 224557 359025 224560
rect 527535 224557 527601 224560
rect 359823 224472 359889 224475
rect 528975 224472 529041 224475
rect 359823 224470 529041 224472
rect 359823 224414 359828 224470
rect 359884 224414 528980 224470
rect 529036 224414 529041 224470
rect 359823 224412 529041 224414
rect 359823 224409 359889 224412
rect 528975 224409 529041 224412
rect 369135 224324 369201 224327
rect 547119 224324 547185 224327
rect 369135 224322 547185 224324
rect 369135 224266 369140 224322
rect 369196 224266 547124 224322
rect 547180 224266 547185 224322
rect 369135 224264 547185 224266
rect 369135 224261 369201 224264
rect 547119 224261 547185 224264
rect 676047 224324 676113 224327
rect 676047 224322 676320 224324
rect 676047 224266 676052 224322
rect 676108 224266 676320 224322
rect 676047 224264 676320 224266
rect 676047 224261 676113 224264
rect 370287 224176 370353 224179
rect 547887 224176 547953 224179
rect 370287 224174 547953 224176
rect 370287 224118 370292 224174
rect 370348 224118 547892 224174
rect 547948 224118 547953 224174
rect 370287 224116 547953 224118
rect 370287 224113 370353 224116
rect 547887 224113 547953 224116
rect 374895 224028 374961 224031
rect 559215 224028 559281 224031
rect 374895 224026 559281 224028
rect 374895 223970 374900 224026
rect 374956 223970 559220 224026
rect 559276 223970 559281 224026
rect 374895 223968 559281 223970
rect 374895 223965 374961 223968
rect 559215 223965 559281 223968
rect 149487 223880 149553 223883
rect 143904 223878 149553 223880
rect 143904 223822 149492 223878
rect 149548 223822 149553 223878
rect 143904 223820 149553 223822
rect 149487 223817 149553 223820
rect 379791 223880 379857 223883
rect 568239 223880 568305 223883
rect 379791 223878 568305 223880
rect 379791 223822 379796 223878
rect 379852 223822 568244 223878
rect 568300 223822 568305 223878
rect 379791 223820 568305 223822
rect 379791 223817 379857 223820
rect 568239 223817 568305 223820
rect 676047 223806 676113 223809
rect 676047 223804 676320 223806
rect 676047 223748 676052 223804
rect 676108 223748 676320 223804
rect 676047 223746 676320 223748
rect 676047 223743 676113 223746
rect 382863 223732 382929 223735
rect 575823 223732 575889 223735
rect 382863 223730 575889 223732
rect 382863 223674 382868 223730
rect 382924 223674 575828 223730
rect 575884 223674 575889 223730
rect 382863 223672 575889 223674
rect 382863 223669 382929 223672
rect 575823 223669 575889 223672
rect 382767 223584 382833 223587
rect 574287 223584 574353 223587
rect 382767 223582 574353 223584
rect 382767 223526 382772 223582
rect 382828 223526 574292 223582
rect 574348 223526 574353 223582
rect 382767 223524 574353 223526
rect 382767 223521 382833 223524
rect 574287 223521 574353 223524
rect 386703 223436 386769 223439
rect 581775 223436 581841 223439
rect 386703 223434 581841 223436
rect 386703 223378 386708 223434
rect 386764 223378 581780 223434
rect 581836 223378 581841 223434
rect 386703 223376 581841 223378
rect 386703 223373 386769 223376
rect 581775 223373 581841 223376
rect 675514 223374 675520 223438
rect 675584 223436 675590 223438
rect 675584 223376 676320 223436
rect 675584 223374 675590 223376
rect 397167 223288 397233 223291
rect 602991 223288 603057 223291
rect 397167 223286 603057 223288
rect 397167 223230 397172 223286
rect 397228 223230 602996 223286
rect 603052 223230 603057 223286
rect 397167 223228 603057 223230
rect 397167 223225 397233 223228
rect 602991 223225 603057 223228
rect 409167 223140 409233 223143
rect 621039 223140 621105 223143
rect 409167 223138 621105 223140
rect 409167 223082 409172 223138
rect 409228 223082 621044 223138
rect 621100 223082 621105 223138
rect 409167 223080 621105 223082
rect 409167 223077 409233 223080
rect 621039 223077 621105 223080
rect 355695 222992 355761 222995
rect 521487 222992 521553 222995
rect 355695 222990 521553 222992
rect 355695 222934 355700 222990
rect 355756 222934 521492 222990
rect 521548 222934 521553 222990
rect 355695 222932 521553 222934
rect 355695 222929 355761 222932
rect 521487 222929 521553 222932
rect 354063 222844 354129 222847
rect 516975 222844 517041 222847
rect 354063 222842 517041 222844
rect 354063 222786 354068 222842
rect 354124 222786 516980 222842
rect 517036 222786 517041 222842
rect 354063 222784 517041 222786
rect 354063 222781 354129 222784
rect 516975 222781 517041 222784
rect 675898 222782 675904 222846
rect 675968 222844 675974 222846
rect 675968 222784 676320 222844
rect 675968 222782 675974 222784
rect 148143 222696 148209 222699
rect 143904 222694 148209 222696
rect 143904 222638 148148 222694
rect 148204 222638 148209 222694
rect 143904 222636 148209 222638
rect 148143 222633 148209 222636
rect 404751 222696 404817 222699
rect 532815 222696 532881 222699
rect 404751 222694 532881 222696
rect 404751 222638 404756 222694
rect 404812 222638 532820 222694
rect 532876 222638 532881 222694
rect 404751 222636 532881 222638
rect 404751 222633 404817 222636
rect 532815 222633 532881 222636
rect 674362 222634 674368 222698
rect 674432 222696 674438 222698
rect 674432 222636 676350 222696
rect 674432 222634 674438 222636
rect 676290 222296 676350 222636
rect 673978 221956 673984 221958
rect 659490 221896 673984 221956
rect 658095 221808 658161 221811
rect 659490 221808 659550 221896
rect 673978 221894 673984 221896
rect 674048 221956 674054 221958
rect 674048 221896 676320 221956
rect 674048 221894 674054 221896
rect 658095 221806 659550 221808
rect 658095 221750 658100 221806
rect 658156 221750 659550 221806
rect 658095 221748 659550 221750
rect 658095 221745 658161 221748
rect 148047 221512 148113 221515
rect 143904 221510 148113 221512
rect 143904 221454 148052 221510
rect 148108 221454 148113 221510
rect 143904 221452 148113 221454
rect 148047 221449 148113 221452
rect 674170 221302 674176 221366
rect 674240 221364 674246 221366
rect 674240 221304 676320 221364
rect 674240 221302 674246 221304
rect 645135 221216 645201 221219
rect 640194 221214 645201 221216
rect 640194 221158 645140 221214
rect 645196 221158 645201 221214
rect 640194 221156 645201 221158
rect 185295 221068 185361 221071
rect 185295 221066 190560 221068
rect 185295 221010 185300 221066
rect 185356 221010 190560 221066
rect 185295 221008 190560 221010
rect 185295 221005 185361 221008
rect 185487 220328 185553 220331
rect 185487 220326 190560 220328
rect 185487 220270 185492 220326
rect 185548 220270 190560 220326
rect 185487 220268 190560 220270
rect 185487 220265 185553 220268
rect 143874 219736 143934 220224
rect 148911 219736 148977 219739
rect 143874 219734 148977 219736
rect 143874 219678 148916 219734
rect 148972 219678 148977 219734
rect 143874 219676 148977 219678
rect 148911 219673 148977 219676
rect 184335 219588 184401 219591
rect 184335 219586 190560 219588
rect 184335 219530 184340 219586
rect 184396 219530 190560 219586
rect 184335 219528 190560 219530
rect 184335 219525 184401 219528
rect 149583 218996 149649 218999
rect 143904 218994 149649 218996
rect 143904 218938 149588 218994
rect 149644 218938 149649 218994
rect 143904 218936 149649 218938
rect 149583 218933 149649 218936
rect 185583 218848 185649 218851
rect 185583 218846 190560 218848
rect 185583 218790 185588 218846
rect 185644 218790 190560 218846
rect 185583 218788 190560 218790
rect 185583 218785 185649 218788
rect 640194 218670 640254 221156
rect 645135 221153 645201 221156
rect 674170 220710 674176 220774
rect 674240 220772 674246 220774
rect 674240 220712 676320 220772
rect 674240 220710 674246 220712
rect 675514 219970 675520 220034
rect 675584 220032 675590 220034
rect 676290 220032 676350 220372
rect 675584 219972 676350 220032
rect 675584 219970 675590 219972
rect 674746 219822 674752 219886
rect 674816 219884 674822 219886
rect 674816 219824 676320 219884
rect 674816 219822 674822 219824
rect 675759 219292 675825 219295
rect 675759 219290 676320 219292
rect 675759 219234 675764 219290
rect 675820 219234 676320 219290
rect 675759 219232 676320 219234
rect 675759 219229 675825 219232
rect 657999 218996 658065 218999
rect 674170 218996 674176 218998
rect 657999 218994 674176 218996
rect 657999 218938 658004 218994
rect 658060 218938 674176 218994
rect 657999 218936 674176 218938
rect 657999 218933 658065 218936
rect 674170 218934 674176 218936
rect 674240 218934 674246 218998
rect 676290 218702 676350 218892
rect 676282 218638 676288 218702
rect 676352 218638 676358 218702
rect 675130 218342 675136 218406
rect 675200 218404 675206 218406
rect 675200 218344 676320 218404
rect 675200 218342 675206 218344
rect 186831 218108 186897 218111
rect 186831 218106 190560 218108
rect 186831 218050 186836 218106
rect 186892 218050 190560 218106
rect 186831 218048 190560 218050
rect 186831 218045 186897 218048
rect 147375 217812 147441 217815
rect 143904 217810 147441 217812
rect 143904 217754 147380 217810
rect 147436 217754 147441 217810
rect 143904 217752 147441 217754
rect 147375 217749 147441 217752
rect 190146 217294 190206 218048
rect 674554 217750 674560 217814
rect 674624 217812 674630 217814
rect 674624 217752 676320 217812
rect 674624 217750 674630 217752
rect 190146 217234 190560 217294
rect 676090 217010 676096 217074
rect 676160 217072 676166 217074
rect 676290 217072 676350 217338
rect 676160 217012 676350 217072
rect 676160 217010 676166 217012
rect 676047 216924 676113 216927
rect 676047 216922 676320 216924
rect 676047 216866 676052 216922
rect 676108 216866 676320 216922
rect 676047 216864 676320 216866
rect 676047 216861 676113 216864
rect 147279 216628 147345 216631
rect 143904 216626 147345 216628
rect 143904 216570 147284 216626
rect 147340 216570 147345 216626
rect 143904 216568 147345 216570
rect 147279 216565 147345 216568
rect 41583 216480 41649 216483
rect 41538 216478 41649 216480
rect 41538 216422 41588 216478
rect 41644 216422 41649 216478
rect 41538 216417 41649 216422
rect 187023 216480 187089 216483
rect 187023 216478 190560 216480
rect 187023 216422 187028 216478
rect 187084 216422 190560 216478
rect 187023 216420 190560 216422
rect 187023 216417 187089 216420
rect 41538 216302 41598 216417
rect 190146 215814 190206 216420
rect 640386 215888 640446 216746
rect 675706 216270 675712 216334
rect 675776 216332 675782 216334
rect 675776 216272 676320 216332
rect 675776 216270 675782 216272
rect 645039 215888 645105 215891
rect 640386 215886 645105 215888
rect 640386 215830 645044 215886
rect 645100 215830 645105 215886
rect 640386 215828 645105 215830
rect 190146 215754 190560 215814
rect 41775 215740 41841 215743
rect 41568 215738 41841 215740
rect 41568 215682 41780 215738
rect 41836 215682 41841 215738
rect 41568 215680 41841 215682
rect 41775 215677 41841 215680
rect 41775 215222 41841 215225
rect 41568 215220 41841 215222
rect 41568 215164 41780 215220
rect 41836 215164 41841 215220
rect 41568 215162 41841 215164
rect 41775 215159 41841 215162
rect 41583 215000 41649 215003
rect 41538 214998 41649 215000
rect 41538 214942 41588 214998
rect 41644 214942 41649 214998
rect 41538 214937 41649 214942
rect 41538 214822 41598 214937
rect 143874 214852 143934 215340
rect 186927 215000 186993 215003
rect 186927 214998 190560 215000
rect 186927 214942 186932 214998
rect 186988 214942 190560 214998
rect 186927 214940 190560 214942
rect 186927 214937 186993 214940
rect 147375 214852 147441 214855
rect 143874 214850 147441 214852
rect 143874 214794 147380 214850
rect 147436 214794 147441 214850
rect 143874 214792 147441 214794
rect 147375 214789 147441 214792
rect 190146 214334 190206 214940
rect 640386 214822 640446 215828
rect 645039 215825 645105 215828
rect 674938 215826 674944 215890
rect 675008 215888 675014 215890
rect 675008 215828 676320 215888
rect 675008 215826 675014 215828
rect 676047 215370 676113 215373
rect 676047 215368 676320 215370
rect 676047 215312 676052 215368
rect 676108 215312 676320 215368
rect 676047 215310 676320 215312
rect 676047 215307 676113 215310
rect 676047 214852 676113 214855
rect 676047 214850 676320 214852
rect 676047 214794 676052 214850
rect 676108 214794 676320 214850
rect 676047 214792 676320 214794
rect 676047 214789 676113 214792
rect 190146 214274 190560 214334
rect 676290 214263 676350 214378
rect 41775 214260 41841 214263
rect 41568 214258 41841 214260
rect 41568 214202 41780 214258
rect 41836 214202 41841 214258
rect 41568 214200 41841 214202
rect 41775 214197 41841 214200
rect 676239 214258 676350 214263
rect 676239 214202 676244 214258
rect 676300 214202 676350 214258
rect 676239 214200 676350 214202
rect 676239 214197 676305 214200
rect 149487 214112 149553 214115
rect 143904 214110 149553 214112
rect 143904 214054 149492 214110
rect 149548 214054 149553 214110
rect 143904 214052 149553 214054
rect 149487 214049 149553 214052
rect 675951 213890 676017 213893
rect 675951 213888 676320 213890
rect 675951 213832 675956 213888
rect 676012 213832 676320 213888
rect 675951 213830 676320 213832
rect 675951 213827 676017 213830
rect 41775 213668 41841 213671
rect 41568 213666 41841 213668
rect 41568 213610 41780 213666
rect 41836 213610 41841 213666
rect 41568 213608 41841 213610
rect 41775 213605 41841 213608
rect 186735 213520 186801 213523
rect 679791 213520 679857 213523
rect 186735 213518 190560 213520
rect 186735 213462 186740 213518
rect 186796 213462 190560 213518
rect 186735 213460 190560 213462
rect 679746 213518 679857 213520
rect 679746 213462 679796 213518
rect 679852 213462 679857 213518
rect 186735 213457 186801 213460
rect 41775 213298 41841 213301
rect 41568 213296 41841 213298
rect 41568 213240 41780 213296
rect 41836 213240 41841 213296
rect 41568 213238 41841 213240
rect 41775 213235 41841 213238
rect 41583 212928 41649 212931
rect 147087 212928 147153 212931
rect 41538 212926 41649 212928
rect 41538 212870 41588 212926
rect 41644 212870 41649 212926
rect 41538 212865 41649 212870
rect 143904 212926 147153 212928
rect 143904 212870 147092 212926
rect 147148 212870 147153 212926
rect 143904 212868 147153 212870
rect 147087 212865 147153 212868
rect 41538 212750 41598 212865
rect 190146 212706 190206 213460
rect 679746 213457 679857 213462
rect 679746 213342 679806 213457
rect 645135 212928 645201 212931
rect 640224 212926 645201 212928
rect 640224 212898 645140 212926
rect 640194 212870 645140 212898
rect 645196 212870 645201 212926
rect 640194 212868 645201 212870
rect 190146 212646 190560 212706
rect 41775 212188 41841 212191
rect 41568 212186 41841 212188
rect 41568 212130 41780 212186
rect 41836 212130 41841 212186
rect 41568 212128 41841 212130
rect 41775 212125 41841 212128
rect 186447 212040 186513 212043
rect 186447 212038 190560 212040
rect 186447 211982 186452 212038
rect 186508 211982 190560 212038
rect 186447 211980 190560 211982
rect 186447 211977 186513 211980
rect 40578 211450 40638 211788
rect 147375 211744 147441 211747
rect 143904 211742 147441 211744
rect 143904 211686 147380 211742
rect 147436 211686 147441 211742
rect 143904 211684 147441 211686
rect 147375 211681 147441 211684
rect 40570 211386 40576 211450
rect 40640 211386 40646 211450
rect 40386 211006 40446 211270
rect 190146 211152 190206 211980
rect 190146 211092 190560 211152
rect 40378 210942 40384 211006
rect 40448 210942 40454 211006
rect 640194 210974 640254 212868
rect 645135 212865 645201 212868
rect 685506 212635 685566 212898
rect 679791 212632 679857 212635
rect 679746 212630 679857 212632
rect 679746 212574 679796 212630
rect 679852 212574 679857 212630
rect 679746 212569 679857 212574
rect 685455 212630 685566 212635
rect 685455 212574 685460 212630
rect 685516 212574 685566 212630
rect 685455 212572 685566 212574
rect 685455 212569 685521 212572
rect 679746 212306 679806 212569
rect 685455 212188 685521 212191
rect 685455 212186 685566 212188
rect 685455 212130 685460 212186
rect 685516 212130 685566 212186
rect 685455 212125 685566 212130
rect 685506 211862 685566 212125
rect 41722 210708 41728 210710
rect 41568 210648 41728 210708
rect 41722 210646 41728 210648
rect 41792 210646 41798 210710
rect 186639 210560 186705 210563
rect 186639 210558 190206 210560
rect 186639 210502 186644 210558
rect 186700 210502 190206 210558
rect 186639 210500 190206 210502
rect 186639 210497 186705 210500
rect 190146 210486 190206 210500
rect 190146 210426 190560 210486
rect 149487 210412 149553 210415
rect 143904 210410 149553 210412
rect 143904 210354 149492 210410
rect 149548 210354 149553 210410
rect 143904 210352 149553 210354
rect 149487 210349 149553 210352
rect 41154 209970 41214 210234
rect 41146 209906 41152 209970
rect 41216 209906 41222 209970
rect 41538 209526 41598 209790
rect 190146 209672 190206 210426
rect 645135 209672 645201 209675
rect 190146 209612 190560 209672
rect 640386 209670 645201 209672
rect 640386 209614 645140 209670
rect 645196 209614 645201 209670
rect 640386 209612 645201 209614
rect 41530 209462 41536 209526
rect 41600 209462 41606 209526
rect 41967 209228 42033 209231
rect 147279 209228 147345 209231
rect 41568 209226 42033 209228
rect 41568 209170 41972 209226
rect 42028 209170 42033 209226
rect 41568 209168 42033 209170
rect 143904 209226 147345 209228
rect 143904 209170 147284 209226
rect 147340 209170 147345 209226
rect 143904 209168 147345 209170
rect 41967 209165 42033 209168
rect 147279 209165 147345 209168
rect 186543 209080 186609 209083
rect 186543 209078 190206 209080
rect 186543 209022 186548 209078
rect 186604 209022 190206 209078
rect 186543 209020 190206 209022
rect 186543 209017 186609 209020
rect 190146 209006 190206 209020
rect 190146 208946 190560 209006
rect 40770 208490 40830 208754
rect 40762 208426 40768 208490
rect 40832 208426 40838 208490
rect 41346 207898 41406 208236
rect 190146 208192 190206 208946
rect 190146 208132 190560 208192
rect 149487 208044 149553 208047
rect 640386 208044 640446 209612
rect 645135 209609 645201 209612
rect 143904 208042 149553 208044
rect 143904 207986 149492 208042
rect 149548 207986 149553 208042
rect 143904 207984 149553 207986
rect 149487 207981 149553 207984
rect 640194 207984 640446 208044
rect 40954 207834 40960 207898
rect 41024 207834 41030 207898
rect 41338 207834 41344 207898
rect 41408 207834 41414 207898
rect 40962 207718 41022 207834
rect 190146 207318 190560 207378
rect 186159 207304 186225 207307
rect 190146 207304 190206 207318
rect 186159 207302 190206 207304
rect 41538 207159 41598 207274
rect 186159 207246 186164 207302
rect 186220 207246 190206 207302
rect 640194 207274 640254 207984
rect 186159 207244 190206 207246
rect 186159 207241 186225 207244
rect 41538 207154 41649 207159
rect 41538 207098 41588 207154
rect 41644 207098 41649 207154
rect 41538 207096 41649 207098
rect 41583 207093 41649 207096
rect 41775 206786 41841 206789
rect 41568 206784 41841 206786
rect 41568 206728 41780 206784
rect 41836 206728 41841 206784
rect 41568 206726 41841 206728
rect 41775 206723 41841 206726
rect 143874 206416 143934 206904
rect 190146 206712 190206 207244
rect 190146 206652 190560 206712
rect 149295 206416 149361 206419
rect 143874 206414 149361 206416
rect 143874 206358 149300 206414
rect 149356 206358 149361 206414
rect 143874 206356 149361 206358
rect 149295 206353 149361 206356
rect 41871 206268 41937 206271
rect 41568 206266 41937 206268
rect 41568 206210 41876 206266
rect 41932 206210 41937 206266
rect 41568 206208 41937 206210
rect 41871 206205 41937 206208
rect 645135 205972 645201 205975
rect 640194 205970 645201 205972
rect 640194 205914 645140 205970
rect 645196 205914 645201 205970
rect 640194 205912 645201 205914
rect 190146 205838 190560 205898
rect 41775 205824 41841 205827
rect 41568 205822 41841 205824
rect 41568 205766 41780 205822
rect 41836 205766 41841 205822
rect 41568 205764 41841 205766
rect 41775 205761 41841 205764
rect 149487 205676 149553 205679
rect 143904 205674 149553 205676
rect 143904 205618 149492 205674
rect 149548 205618 149553 205674
rect 143904 205616 149553 205618
rect 149487 205613 149553 205616
rect 186351 205232 186417 205235
rect 190146 205232 190206 205838
rect 186351 205230 190560 205232
rect 41538 205087 41598 205202
rect 186351 205174 186356 205230
rect 186412 205174 190560 205230
rect 186351 205172 190560 205174
rect 186351 205169 186417 205172
rect 41538 205082 41649 205087
rect 41538 205026 41588 205082
rect 41644 205026 41649 205082
rect 41538 205024 41649 205026
rect 41583 205021 41649 205024
rect 41679 204936 41745 204939
rect 41538 204934 41745 204936
rect 41538 204878 41684 204934
rect 41740 204878 41745 204934
rect 41538 204876 41745 204878
rect 41538 204758 41598 204876
rect 41679 204873 41745 204876
rect 149679 204492 149745 204495
rect 143904 204490 149745 204492
rect 143904 204434 149684 204490
rect 149740 204434 149745 204490
rect 143904 204432 149745 204434
rect 149679 204429 149745 204432
rect 41775 204344 41841 204347
rect 41568 204342 41841 204344
rect 41568 204286 41780 204342
rect 41836 204286 41841 204342
rect 41568 204284 41841 204286
rect 41775 204281 41841 204284
rect 186255 204344 186321 204347
rect 186255 204342 190560 204344
rect 186255 204286 186260 204342
rect 186316 204286 190560 204342
rect 186255 204284 190560 204286
rect 186255 204281 186321 204284
rect 41775 203752 41841 203755
rect 41568 203750 41841 203752
rect 41568 203694 41780 203750
rect 41836 203694 41841 203750
rect 41568 203692 41841 203694
rect 41775 203689 41841 203692
rect 190146 203604 190206 204284
rect 190146 203544 190560 203604
rect 640194 203426 640254 205912
rect 645135 205909 645201 205912
rect 675759 205084 675825 205087
rect 676090 205084 676096 205086
rect 675759 205082 676096 205084
rect 675759 205026 675764 205082
rect 675820 205026 676096 205082
rect 675759 205024 676096 205026
rect 675759 205021 675825 205024
rect 676090 205022 676096 205024
rect 676160 205022 676166 205086
rect 675471 204346 675537 204347
rect 675471 204342 675520 204346
rect 675584 204344 675590 204346
rect 675471 204286 675476 204342
rect 675471 204282 675520 204286
rect 675584 204284 675628 204344
rect 675584 204282 675590 204284
rect 675471 204281 675537 204282
rect 149487 203308 149553 203311
rect 143904 203306 149553 203308
rect 143904 203250 149492 203306
rect 149548 203250 149553 203306
rect 143904 203248 149553 203250
rect 149487 203245 149553 203248
rect 186063 202864 186129 202867
rect 186063 202862 190560 202864
rect 186063 202806 186068 202862
rect 186124 202806 190560 202862
rect 186063 202804 190560 202806
rect 186063 202801 186129 202804
rect 190146 202124 190206 202804
rect 675759 202716 675825 202719
rect 676282 202716 676288 202718
rect 675759 202714 676288 202716
rect 675759 202658 675764 202714
rect 675820 202658 676288 202714
rect 675759 202656 676288 202658
rect 675759 202653 675825 202656
rect 676282 202654 676288 202656
rect 676352 202654 676358 202718
rect 190146 202064 190560 202124
rect 143874 201680 143934 202020
rect 147951 201680 148017 201683
rect 143874 201678 148017 201680
rect 143874 201622 147956 201678
rect 148012 201622 148017 201678
rect 143874 201620 148017 201622
rect 147951 201617 148017 201620
rect 645135 201532 645201 201535
rect 640416 201530 645201 201532
rect 640416 201502 645140 201530
rect 640386 201474 645140 201502
rect 645196 201474 645201 201530
rect 640386 201472 645201 201474
rect 185871 201384 185937 201387
rect 185871 201382 190560 201384
rect 185871 201326 185876 201382
rect 185932 201326 190560 201382
rect 185871 201324 190560 201326
rect 185871 201321 185937 201324
rect 149487 200792 149553 200795
rect 143904 200790 149553 200792
rect 143904 200734 149492 200790
rect 149548 200734 149553 200790
rect 143904 200732 149553 200734
rect 149487 200729 149553 200732
rect 190146 200570 190206 201324
rect 190146 200510 190560 200570
rect 184335 199756 184401 199759
rect 184335 199754 190560 199756
rect 184335 199698 184340 199754
rect 184396 199698 190560 199754
rect 184335 199696 190560 199698
rect 184335 199693 184401 199696
rect 149295 199608 149361 199611
rect 143904 199606 149361 199608
rect 143904 199550 149300 199606
rect 149356 199550 149361 199606
rect 640386 199578 640446 201472
rect 645135 201469 645201 201472
rect 675759 201386 675825 201387
rect 675706 201384 675712 201386
rect 675668 201324 675712 201384
rect 675776 201382 675825 201386
rect 675820 201326 675825 201382
rect 675706 201322 675712 201324
rect 675776 201322 675825 201326
rect 675759 201321 675825 201322
rect 143904 199548 149361 199550
rect 149295 199545 149361 199548
rect 187215 199164 187281 199167
rect 187215 199162 190014 199164
rect 187215 199106 187220 199162
rect 187276 199106 190014 199162
rect 187215 199104 190014 199106
rect 187215 199101 187281 199104
rect 189954 199090 190014 199104
rect 189954 199030 190560 199090
rect 147855 198424 147921 198427
rect 143904 198422 147921 198424
rect 143904 198366 147860 198422
rect 147916 198366 147921 198422
rect 143904 198364 147921 198366
rect 147855 198361 147921 198364
rect 675130 198362 675136 198426
rect 675200 198424 675206 198426
rect 675471 198424 675537 198427
rect 675200 198422 675537 198424
rect 675200 198366 675476 198422
rect 675532 198366 675537 198422
rect 675200 198364 675537 198366
rect 675200 198362 675206 198364
rect 675471 198361 675537 198364
rect 185391 198276 185457 198279
rect 645135 198276 645201 198279
rect 185391 198274 190560 198276
rect 185391 198218 185396 198274
rect 185452 198218 190560 198274
rect 185391 198216 190560 198218
rect 640386 198274 645201 198276
rect 640386 198218 645140 198274
rect 645196 198218 645201 198274
rect 640386 198216 645201 198218
rect 185391 198213 185457 198216
rect 184239 197684 184305 197687
rect 640386 197684 640446 198216
rect 645135 198213 645201 198216
rect 184239 197682 190014 197684
rect 184239 197626 184244 197682
rect 184300 197626 190014 197682
rect 640224 197654 640446 197684
rect 184239 197624 190014 197626
rect 184239 197621 184305 197624
rect 189954 197610 190014 197624
rect 640194 197624 640416 197654
rect 189954 197550 190560 197610
rect 149679 197092 149745 197095
rect 143904 197090 149745 197092
rect 143904 197034 149684 197090
rect 149740 197034 149745 197090
rect 143904 197032 149745 197034
rect 149679 197029 149745 197032
rect 184335 196796 184401 196799
rect 184335 196794 190560 196796
rect 184335 196738 184340 196794
rect 184396 196738 190560 196794
rect 184335 196736 190560 196738
rect 184335 196733 184401 196736
rect 184431 196056 184497 196059
rect 640194 196056 640254 197624
rect 184431 196054 190560 196056
rect 184431 195998 184436 196054
rect 184492 195998 190560 196054
rect 184431 195996 190560 195998
rect 640194 195996 640446 196056
rect 184431 195993 184497 195996
rect 149295 195908 149361 195911
rect 143904 195906 149361 195908
rect 143904 195850 149300 195906
rect 149356 195850 149361 195906
rect 143904 195848 149361 195850
rect 149295 195845 149361 195848
rect 640386 195730 640446 195996
rect 184335 195316 184401 195319
rect 184335 195314 190560 195316
rect 184335 195258 184340 195314
rect 184396 195258 190560 195314
rect 184335 195256 190560 195258
rect 184335 195253 184401 195256
rect 674938 195254 674944 195318
rect 675008 195316 675014 195318
rect 675471 195316 675537 195319
rect 675008 195314 675537 195316
rect 675008 195258 675476 195314
rect 675532 195258 675537 195314
rect 675008 195256 675537 195258
rect 675008 195254 675014 195256
rect 675471 195253 675537 195256
rect 40378 195106 40384 195170
rect 40448 195168 40454 195170
rect 41775 195168 41841 195171
rect 40448 195166 41841 195168
rect 40448 195110 41780 195166
rect 41836 195110 41841 195166
rect 40448 195108 41841 195110
rect 40448 195106 40454 195108
rect 41775 195105 41841 195108
rect 149391 194724 149457 194727
rect 143904 194722 149457 194724
rect 143904 194666 149396 194722
rect 149452 194666 149457 194722
rect 143904 194664 149457 194666
rect 149391 194661 149457 194664
rect 184431 194428 184497 194431
rect 184431 194426 190560 194428
rect 184431 194370 184436 194426
rect 184492 194370 190560 194426
rect 184431 194368 190560 194370
rect 184431 194365 184497 194368
rect 645135 193984 645201 193987
rect 640386 193982 645201 193984
rect 640386 193926 645140 193982
rect 645196 193926 645201 193982
rect 640386 193924 645201 193926
rect 184527 193836 184593 193839
rect 184527 193834 190014 193836
rect 184527 193778 184532 193834
rect 184588 193778 190014 193834
rect 184527 193776 190014 193778
rect 184527 193773 184593 193776
rect 189954 193762 190014 193776
rect 189954 193702 190560 193762
rect 143874 193096 143934 193436
rect 149391 193096 149457 193099
rect 143874 193094 149457 193096
rect 143874 193038 149396 193094
rect 149452 193038 149457 193094
rect 143874 193036 149457 193038
rect 149391 193033 149457 193036
rect 184431 192948 184497 192951
rect 184431 192946 190560 192948
rect 184431 192890 184436 192946
rect 184492 192890 190560 192946
rect 184431 192888 190560 192890
rect 184431 192885 184497 192888
rect 640386 192800 640446 193924
rect 645135 193921 645201 193924
rect 674746 193478 674752 193542
rect 674816 193540 674822 193542
rect 675375 193540 675441 193543
rect 674816 193538 675441 193540
rect 674816 193482 675380 193538
rect 675436 193482 675441 193538
rect 674816 193480 675441 193482
rect 674816 193478 674822 193480
rect 675375 193477 675441 193480
rect 640194 192740 640446 192800
rect 184335 192356 184401 192359
rect 184335 192354 190014 192356
rect 184335 192298 184340 192354
rect 184396 192298 190014 192354
rect 184335 192296 190014 192298
rect 184335 192293 184401 192296
rect 189954 192282 190014 192296
rect 189954 192222 190560 192282
rect 147759 192208 147825 192211
rect 143904 192206 147825 192208
rect 143904 192150 147764 192206
rect 147820 192150 147825 192206
rect 143904 192148 147825 192150
rect 147759 192145 147825 192148
rect 640194 192030 640254 192740
rect 674554 191554 674560 191618
rect 674624 191616 674630 191618
rect 675375 191616 675441 191619
rect 674624 191614 675441 191616
rect 674624 191558 675380 191614
rect 675436 191558 675441 191614
rect 674624 191556 675441 191558
rect 674624 191554 674630 191556
rect 675375 191553 675441 191556
rect 184527 191468 184593 191471
rect 184527 191466 190560 191468
rect 184527 191410 184532 191466
rect 184588 191410 190560 191466
rect 184527 191408 190560 191410
rect 184527 191405 184593 191408
rect 147567 191024 147633 191027
rect 143904 191022 147633 191024
rect 143904 190966 147572 191022
rect 147628 190966 147633 191022
rect 143904 190964 147633 190966
rect 147567 190961 147633 190964
rect 184623 190728 184689 190731
rect 184623 190726 190014 190728
rect 184623 190670 184628 190726
rect 184684 190670 190014 190726
rect 184623 190668 190014 190670
rect 184623 190665 184689 190668
rect 189954 190654 190014 190668
rect 189954 190594 190560 190654
rect 41530 190074 41536 190138
rect 41600 190136 41606 190138
rect 41775 190136 41841 190139
rect 645135 190136 645201 190139
rect 41600 190134 41841 190136
rect 41600 190078 41780 190134
rect 41836 190078 41841 190134
rect 640416 190134 645201 190136
rect 640416 190106 645140 190134
rect 41600 190076 41841 190078
rect 41600 190074 41606 190076
rect 41775 190073 41841 190076
rect 640386 190078 645140 190106
rect 645196 190078 645201 190134
rect 640386 190076 645201 190078
rect 184335 189988 184401 189991
rect 184335 189986 190560 189988
rect 184335 189930 184340 189986
rect 184396 189930 190560 189986
rect 184335 189928 190560 189930
rect 184335 189925 184401 189928
rect 147471 189840 147537 189843
rect 143904 189838 147537 189840
rect 143904 189782 147476 189838
rect 147532 189782 147537 189838
rect 143904 189780 147537 189782
rect 147471 189777 147537 189780
rect 184431 189248 184497 189251
rect 184431 189246 190014 189248
rect 184431 189190 184436 189246
rect 184492 189190 190014 189246
rect 184431 189188 190014 189190
rect 184431 189185 184497 189188
rect 189954 189174 190014 189188
rect 189954 189114 190560 189174
rect 143874 188064 143934 188552
rect 184527 188508 184593 188511
rect 184527 188506 190560 188508
rect 184527 188450 184532 188506
rect 184588 188450 190560 188506
rect 184527 188448 190560 188450
rect 184527 188445 184593 188448
rect 640386 188182 640446 190076
rect 645135 190073 645201 190076
rect 149391 188064 149457 188067
rect 143874 188062 149457 188064
rect 143874 188006 149396 188062
rect 149452 188006 149457 188062
rect 143874 188004 149457 188006
rect 149391 188001 149457 188004
rect 184623 187620 184689 187623
rect 184623 187618 190560 187620
rect 184623 187562 184628 187618
rect 184684 187562 190560 187618
rect 184623 187560 190560 187562
rect 184623 187557 184689 187560
rect 147663 187472 147729 187475
rect 143904 187470 147729 187472
rect 143904 187414 147668 187470
rect 147724 187414 147729 187470
rect 143904 187412 147729 187414
rect 147663 187409 147729 187412
rect 40954 187114 40960 187178
rect 41024 187176 41030 187178
rect 41775 187176 41841 187179
rect 41024 187174 41841 187176
rect 41024 187118 41780 187174
rect 41836 187118 41841 187174
rect 41024 187116 41841 187118
rect 41024 187114 41030 187116
rect 41775 187113 41841 187116
rect 184431 186880 184497 186883
rect 184431 186878 190560 186880
rect 184431 186822 184436 186878
rect 184492 186822 190560 186878
rect 184431 186820 190560 186822
rect 184431 186817 184497 186820
rect 41338 186670 41344 186734
rect 41408 186732 41414 186734
rect 41775 186732 41841 186735
rect 41408 186730 41841 186732
rect 41408 186674 41780 186730
rect 41836 186674 41841 186730
rect 41408 186672 41841 186674
rect 41408 186670 41414 186672
rect 41775 186669 41841 186672
rect 149391 186288 149457 186291
rect 143904 186286 149457 186288
rect 143904 186230 149396 186286
rect 149452 186230 149457 186286
rect 143904 186228 149457 186230
rect 149391 186225 149457 186228
rect 184335 186140 184401 186143
rect 184335 186138 190560 186140
rect 184335 186082 184340 186138
rect 184396 186082 190560 186138
rect 184335 186080 190560 186082
rect 184335 186077 184401 186080
rect 41146 185782 41152 185846
rect 41216 185844 41222 185846
rect 41775 185844 41841 185847
rect 41216 185842 41841 185844
rect 41216 185786 41780 185842
rect 41836 185786 41841 185842
rect 41216 185784 41841 185786
rect 41216 185782 41222 185784
rect 41775 185781 41841 185784
rect 184623 185400 184689 185403
rect 184623 185398 190014 185400
rect 184623 185342 184628 185398
rect 184684 185342 190014 185398
rect 184623 185340 190014 185342
rect 184623 185337 184689 185340
rect 189954 185326 190014 185340
rect 189954 185266 190560 185326
rect 143874 184512 143934 185000
rect 184527 184660 184593 184663
rect 184527 184658 190560 184660
rect 184527 184602 184532 184658
rect 184588 184602 190560 184658
rect 184527 184600 190560 184602
rect 184527 184597 184593 184600
rect 148911 184512 148977 184515
rect 143874 184510 148977 184512
rect 143874 184454 148916 184510
rect 148972 184454 148977 184510
rect 143874 184452 148977 184454
rect 148911 184449 148977 184452
rect 640386 184364 640446 186258
rect 646191 184364 646257 184367
rect 640386 184362 646257 184364
rect 640386 184334 646196 184362
rect 640416 184306 646196 184334
rect 646252 184306 646257 184362
rect 640416 184304 646257 184306
rect 646191 184301 646257 184304
rect 40570 184006 40576 184070
rect 40640 184068 40646 184070
rect 41775 184068 41841 184071
rect 40640 184066 41841 184068
rect 40640 184010 41780 184066
rect 41836 184010 41841 184066
rect 40640 184008 41841 184010
rect 40640 184006 40646 184008
rect 41775 184005 41841 184008
rect 184335 183920 184401 183923
rect 184335 183918 190014 183920
rect 184335 183862 184340 183918
rect 184396 183862 190014 183918
rect 184335 183860 190014 183862
rect 184335 183857 184401 183860
rect 189954 183846 190014 183860
rect 189954 183786 190560 183846
rect 147567 183772 147633 183775
rect 143904 183770 147633 183772
rect 143904 183714 147572 183770
rect 147628 183714 147633 183770
rect 143904 183712 147633 183714
rect 147567 183709 147633 183712
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 184527 183180 184593 183183
rect 184527 183178 190560 183180
rect 184527 183122 184532 183178
rect 184588 183122 190560 183178
rect 184527 183120 190560 183122
rect 184527 183117 184593 183120
rect 41775 183034 41841 183035
rect 41722 183032 41728 183034
rect 41684 182972 41728 183032
rect 41792 183030 41841 183034
rect 645903 183032 645969 183035
rect 41836 182974 41841 183030
rect 41722 182970 41728 182972
rect 41792 182970 41841 182974
rect 41775 182969 41841 182970
rect 640386 183030 645969 183032
rect 640386 182974 645908 183030
rect 645964 182974 645969 183030
rect 640386 182972 645969 182974
rect 149391 182588 149457 182591
rect 143904 182586 149457 182588
rect 143904 182530 149396 182586
rect 149452 182530 149457 182586
rect 143904 182528 149457 182530
rect 149391 182525 149457 182528
rect 184431 182440 184497 182443
rect 640386 182440 640446 182972
rect 645903 182969 645969 182972
rect 184431 182438 190014 182440
rect 184431 182382 184436 182438
rect 184492 182382 190014 182438
rect 640224 182410 640446 182440
rect 184431 182380 190014 182382
rect 184431 182377 184497 182380
rect 189954 182366 190014 182380
rect 640194 182380 640416 182410
rect 189954 182306 190560 182366
rect 184623 181552 184689 181555
rect 184623 181550 190560 181552
rect 184623 181494 184628 181550
rect 184684 181494 190560 181550
rect 184623 181492 190560 181494
rect 184623 181489 184689 181492
rect 149679 181404 149745 181407
rect 143904 181402 149745 181404
rect 143904 181346 149684 181402
rect 149740 181346 149745 181402
rect 143904 181344 149745 181346
rect 149679 181341 149745 181344
rect 184335 180812 184401 180815
rect 184335 180810 190560 180812
rect 184335 180754 184340 180810
rect 184396 180754 190560 180810
rect 184335 180752 190560 180754
rect 184335 180749 184401 180752
rect 640194 180560 640254 182380
rect 143874 179628 143934 180116
rect 184431 180072 184497 180075
rect 184431 180070 190560 180072
rect 184431 180014 184436 180070
rect 184492 180014 190560 180070
rect 184431 180012 190560 180014
rect 184431 180009 184497 180012
rect 676290 179631 676350 179894
rect 149391 179628 149457 179631
rect 143874 179626 149457 179628
rect 143874 179570 149396 179626
rect 149452 179570 149457 179626
rect 143874 179568 149457 179570
rect 149391 179565 149457 179568
rect 676239 179626 676350 179631
rect 676239 179570 676244 179626
rect 676300 179570 676350 179626
rect 676239 179568 676350 179570
rect 676239 179565 676305 179568
rect 184527 179332 184593 179335
rect 645999 179332 646065 179335
rect 184527 179330 190560 179332
rect 184527 179274 184532 179330
rect 184588 179274 190560 179330
rect 184527 179272 190560 179274
rect 640194 179330 646065 179332
rect 640194 179274 646004 179330
rect 646060 179274 646065 179330
rect 640194 179272 646065 179274
rect 184527 179269 184593 179272
rect 147375 178888 147441 178891
rect 143904 178886 147441 178888
rect 143904 178830 147380 178886
rect 147436 178830 147441 178886
rect 143904 178828 147441 178830
rect 147375 178825 147441 178828
rect 184623 178592 184689 178595
rect 184623 178590 190560 178592
rect 184623 178534 184628 178590
rect 184684 178534 190560 178590
rect 184623 178532 190560 178534
rect 184623 178529 184689 178532
rect 147183 177704 147249 177707
rect 143904 177702 147249 177704
rect 143904 177646 147188 177702
rect 147244 177646 147249 177702
rect 143904 177644 147249 177646
rect 147183 177641 147249 177644
rect 184335 177704 184401 177707
rect 184335 177702 190560 177704
rect 184335 177646 184340 177702
rect 184396 177646 190560 177702
rect 184335 177644 190560 177646
rect 184335 177641 184401 177644
rect 184431 177112 184497 177115
rect 184431 177110 190014 177112
rect 184431 177054 184436 177110
rect 184492 177054 190014 177110
rect 184431 177052 190014 177054
rect 184431 177049 184497 177052
rect 189954 177038 190014 177052
rect 189954 176978 190560 177038
rect 640194 176786 640254 179272
rect 645999 179269 646065 179272
rect 676047 179332 676113 179335
rect 676047 179330 676320 179332
rect 676047 179274 676052 179330
rect 676108 179274 676320 179330
rect 676047 179272 676320 179274
rect 676047 179269 676113 179272
rect 676047 178814 676113 178817
rect 676047 178812 676320 178814
rect 676047 178756 676052 178812
rect 676108 178756 676320 178812
rect 676047 178754 676320 178756
rect 676047 178751 676113 178754
rect 675898 178382 675904 178446
rect 675968 178444 675974 178446
rect 675968 178384 676320 178444
rect 675968 178382 675974 178384
rect 674362 177790 674368 177854
rect 674432 177852 674438 177854
rect 674432 177792 676320 177852
rect 674432 177790 674438 177792
rect 673978 177198 673984 177262
rect 674048 177260 674054 177262
rect 674048 177200 676320 177260
rect 674048 177198 674054 177200
rect 675514 176902 675520 176966
rect 675584 176964 675590 176966
rect 675584 176904 676320 176964
rect 675584 176902 675590 176904
rect 147183 176520 147249 176523
rect 143904 176518 147249 176520
rect 143904 176462 147188 176518
rect 147244 176462 147249 176518
rect 143904 176460 147249 176462
rect 147183 176457 147249 176460
rect 674170 176310 674176 176374
rect 674240 176372 674246 176374
rect 674240 176312 676320 176372
rect 674240 176310 674246 176312
rect 184527 176224 184593 176227
rect 184527 176222 190560 176224
rect 184527 176166 184532 176222
rect 184588 176166 190560 176222
rect 184527 176164 190560 176166
rect 184527 176161 184593 176164
rect 652239 175928 652305 175931
rect 675514 175928 675520 175930
rect 652239 175926 675520 175928
rect 652239 175870 652244 175926
rect 652300 175870 675520 175926
rect 652239 175868 675520 175870
rect 652239 175865 652305 175868
rect 675514 175866 675520 175868
rect 675584 175866 675590 175930
rect 652431 175780 652497 175783
rect 674170 175780 674176 175782
rect 652431 175778 674176 175780
rect 652431 175722 652436 175778
rect 652492 175722 674176 175778
rect 652431 175720 674176 175722
rect 652431 175717 652497 175720
rect 674170 175718 674176 175720
rect 674240 175780 674246 175782
rect 674240 175720 676320 175780
rect 674240 175718 674246 175720
rect 184335 175632 184401 175635
rect 184335 175630 190014 175632
rect 184335 175574 184340 175630
rect 184396 175574 190014 175630
rect 184335 175572 190014 175574
rect 184335 175569 184401 175572
rect 189954 175558 190014 175572
rect 189954 175498 190560 175558
rect 676047 175410 676113 175413
rect 676047 175408 676320 175410
rect 676047 175352 676052 175408
rect 676108 175352 676320 175408
rect 676047 175350 676320 175352
rect 676047 175347 676113 175350
rect 147087 175188 147153 175191
rect 143904 175186 147153 175188
rect 143904 175130 147092 175186
rect 147148 175130 147153 175186
rect 143904 175128 147153 175130
rect 147087 175125 147153 175128
rect 645135 174892 645201 174895
rect 640416 174890 645201 174892
rect 640416 174862 645140 174890
rect 640386 174834 645140 174862
rect 645196 174834 645201 174890
rect 640386 174832 645201 174834
rect 186159 174744 186225 174747
rect 186159 174742 190560 174744
rect 186159 174686 186164 174742
rect 186220 174686 190560 174742
rect 186159 174684 190560 174686
rect 186159 174681 186225 174684
rect 147375 174004 147441 174007
rect 143904 174002 147441 174004
rect 143904 173946 147380 174002
rect 147436 173946 147441 174002
rect 143904 173944 147441 173946
rect 147375 173941 147441 173944
rect 184431 174004 184497 174007
rect 184431 174002 190014 174004
rect 184431 173946 184436 174002
rect 184492 173946 190014 174002
rect 184431 173944 190014 173946
rect 184431 173941 184497 173944
rect 189954 173930 190014 173944
rect 189954 173870 190560 173930
rect 185775 173264 185841 173267
rect 185775 173262 190560 173264
rect 185775 173206 185780 173262
rect 185836 173206 190560 173262
rect 185775 173204 190560 173206
rect 185775 173201 185841 173204
rect 640386 172938 640446 174832
rect 645135 174829 645201 174832
rect 674746 174830 674752 174894
rect 674816 174892 674822 174894
rect 674816 174832 676320 174892
rect 674816 174830 674822 174832
rect 675375 174300 675441 174303
rect 675375 174298 676320 174300
rect 675375 174242 675380 174298
rect 675436 174242 676320 174298
rect 675375 174240 676320 174242
rect 675375 174237 675441 174240
rect 676290 173711 676350 173826
rect 676239 173706 676350 173711
rect 676239 173650 676244 173706
rect 676300 173650 676350 173706
rect 676239 173648 676350 173650
rect 676239 173645 676305 173648
rect 674938 173350 674944 173414
rect 675008 173412 675014 173414
rect 675008 173352 676320 173412
rect 675008 173350 675014 173352
rect 148911 172820 148977 172823
rect 143904 172818 148977 172820
rect 143904 172762 148916 172818
rect 148972 172762 148977 172818
rect 143904 172760 148977 172762
rect 148911 172757 148977 172760
rect 674554 172758 674560 172822
rect 674624 172820 674630 172822
rect 674624 172760 676320 172820
rect 674624 172758 674630 172760
rect 184335 172524 184401 172527
rect 184335 172522 190014 172524
rect 184335 172466 184340 172522
rect 184396 172466 190014 172522
rect 184335 172464 190014 172466
rect 184335 172461 184401 172464
rect 189954 172450 190014 172464
rect 189954 172390 190560 172450
rect 675471 172376 675537 172379
rect 675471 172374 676320 172376
rect 675471 172318 675476 172374
rect 675532 172318 676320 172374
rect 675471 172316 676320 172318
rect 675471 172313 675537 172316
rect 676047 171932 676113 171935
rect 676047 171930 676320 171932
rect 676047 171874 676052 171930
rect 676108 171874 676320 171930
rect 676047 171872 676320 171874
rect 676047 171869 676113 171872
rect 148324 171722 148330 171786
rect 148394 171784 148400 171786
rect 148394 171724 190560 171784
rect 148394 171722 148400 171724
rect 143874 171044 143934 171532
rect 675951 171340 676017 171343
rect 675951 171338 676320 171340
rect 675951 171282 675956 171338
rect 676012 171282 676320 171338
rect 675951 171280 676320 171282
rect 675951 171277 676017 171280
rect 149391 171044 149457 171047
rect 645135 171044 645201 171047
rect 143874 171042 149457 171044
rect 143874 170986 149396 171042
rect 149452 170986 149457 171042
rect 640416 171042 645201 171044
rect 640416 171014 645140 171042
rect 143874 170984 149457 170986
rect 149391 170981 149457 170984
rect 640386 170986 645140 171014
rect 645196 170986 645201 171042
rect 640386 170984 645201 170986
rect 184431 170896 184497 170899
rect 184431 170894 190560 170896
rect 184431 170838 184436 170894
rect 184492 170838 190560 170894
rect 184431 170836 190560 170838
rect 184431 170833 184497 170836
rect 147279 170304 147345 170307
rect 143904 170302 147345 170304
rect 143904 170246 147284 170302
rect 147340 170246 147345 170302
rect 143904 170244 147345 170246
rect 147279 170241 147345 170244
rect 184527 170304 184593 170307
rect 184527 170302 190014 170304
rect 184527 170246 184532 170302
rect 184588 170246 190014 170302
rect 184527 170244 190014 170246
rect 184527 170241 184593 170244
rect 189954 170230 190014 170244
rect 189954 170170 190560 170230
rect 184335 169416 184401 169419
rect 184335 169414 190560 169416
rect 184335 169358 184340 169414
rect 184396 169358 190560 169414
rect 184335 169356 190560 169358
rect 184335 169353 184401 169356
rect 149391 169120 149457 169123
rect 143904 169118 149457 169120
rect 143904 169062 149396 169118
rect 149452 169062 149457 169118
rect 640386 169090 640446 170984
rect 645135 170981 645201 170984
rect 673978 170834 673984 170898
rect 674048 170896 674054 170898
rect 674048 170836 676320 170896
rect 674048 170834 674054 170836
rect 675130 169946 675136 170010
rect 675200 170008 675206 170010
rect 676290 170008 676350 170348
rect 675200 169948 676350 170008
rect 675200 169946 675206 169948
rect 676047 169860 676113 169863
rect 676047 169858 676320 169860
rect 676047 169802 676052 169858
rect 676108 169802 676320 169858
rect 676047 169800 676320 169802
rect 676047 169797 676113 169800
rect 675322 169354 675328 169418
rect 675392 169416 675398 169418
rect 675392 169356 676320 169416
rect 675392 169354 675398 169356
rect 143904 169060 149457 169062
rect 149391 169057 149457 169060
rect 675706 168762 675712 168826
rect 675776 168824 675782 168826
rect 675776 168764 676320 168824
rect 675776 168762 675782 168764
rect 184431 168676 184497 168679
rect 184431 168674 190014 168676
rect 184431 168618 184436 168674
rect 184492 168618 190014 168674
rect 184431 168616 190014 168618
rect 184431 168613 184497 168616
rect 189954 168602 190014 168616
rect 189954 168542 190560 168602
rect 676290 168087 676350 168350
rect 148911 168084 148977 168087
rect 143904 168082 148977 168084
rect 143904 168026 148916 168082
rect 148972 168026 148977 168082
rect 143904 168024 148977 168026
rect 148911 168021 148977 168024
rect 676239 168082 676350 168087
rect 676239 168026 676244 168082
rect 676300 168026 676350 168082
rect 676239 168024 676350 168026
rect 676239 168021 676305 168024
rect 184527 167936 184593 167939
rect 184527 167934 190560 167936
rect 184527 167878 184532 167934
rect 184588 167878 190560 167934
rect 184527 167876 190560 167878
rect 184527 167873 184593 167876
rect 645135 167788 645201 167791
rect 640386 167786 645201 167788
rect 640386 167730 645140 167786
rect 645196 167730 645201 167786
rect 640386 167728 645201 167730
rect 184623 167196 184689 167199
rect 184623 167194 190014 167196
rect 184623 167138 184628 167194
rect 184684 167138 190014 167194
rect 184623 167136 190014 167138
rect 184623 167133 184689 167136
rect 189954 167122 190014 167136
rect 189954 167062 190560 167122
rect 143874 166308 143934 166796
rect 184335 166456 184401 166459
rect 184335 166454 190560 166456
rect 184335 166398 184340 166454
rect 184396 166398 190560 166454
rect 184335 166396 190560 166398
rect 184335 166393 184401 166396
rect 149199 166308 149265 166311
rect 143874 166306 149265 166308
rect 143874 166250 149204 166306
rect 149260 166250 149265 166306
rect 143874 166248 149265 166250
rect 149199 166245 149265 166248
rect 640386 166012 640446 167728
rect 645135 167725 645201 167728
rect 676143 167640 676209 167643
rect 676290 167640 676350 167906
rect 676143 167638 676350 167640
rect 676143 167582 676148 167638
rect 676204 167582 676350 167638
rect 676143 167580 676350 167582
rect 676143 167577 676209 167580
rect 676290 167199 676350 167314
rect 676239 167194 676350 167199
rect 676239 167138 676244 167194
rect 676300 167138 676350 167194
rect 676239 167136 676350 167138
rect 676239 167133 676305 167136
rect 640194 165952 640446 166012
rect 184431 165716 184497 165719
rect 184431 165714 190014 165716
rect 184431 165658 184436 165714
rect 184492 165658 190014 165714
rect 184431 165656 190014 165658
rect 184431 165653 184497 165656
rect 189954 165642 190014 165656
rect 189954 165582 190560 165642
rect 146895 165568 146961 165571
rect 143904 165566 146961 165568
rect 143904 165510 146900 165566
rect 146956 165510 146961 165566
rect 143904 165508 146961 165510
rect 146895 165505 146961 165508
rect 640194 165242 640254 165952
rect 184527 164828 184593 164831
rect 184527 164826 190560 164828
rect 184527 164770 184532 164826
rect 184588 164770 190560 164826
rect 184527 164768 190560 164770
rect 184527 164765 184593 164768
rect 146991 164384 147057 164387
rect 143904 164382 147057 164384
rect 143904 164326 146996 164382
rect 147052 164326 147057 164382
rect 143904 164324 147057 164326
rect 146991 164321 147057 164324
rect 184335 164088 184401 164091
rect 184335 164086 190560 164088
rect 184335 164030 184340 164086
rect 184396 164030 190560 164086
rect 184335 164028 190560 164030
rect 184335 164025 184401 164028
rect 184335 163348 184401 163351
rect 184335 163346 190560 163348
rect 184335 163290 184340 163346
rect 184396 163290 190560 163346
rect 184335 163288 190560 163290
rect 184335 163285 184401 163288
rect 149391 163200 149457 163203
rect 143904 163198 149457 163200
rect 143904 163142 149396 163198
rect 149452 163142 149457 163198
rect 143904 163140 149457 163142
rect 149391 163137 149457 163140
rect 184431 162608 184497 162611
rect 184431 162606 190560 162608
rect 184431 162550 184436 162606
rect 184492 162550 190560 162606
rect 184431 162548 190560 162550
rect 184431 162545 184497 162548
rect 149007 161868 149073 161871
rect 143904 161866 149073 161868
rect 143904 161810 149012 161866
rect 149068 161810 149073 161866
rect 143904 161808 149073 161810
rect 149007 161805 149073 161808
rect 184527 161868 184593 161871
rect 184527 161866 190560 161868
rect 184527 161810 184532 161866
rect 184588 161810 190560 161866
rect 184527 161808 190560 161810
rect 184527 161805 184593 161808
rect 640386 161424 640446 163318
rect 645519 161424 645585 161427
rect 640386 161422 645585 161424
rect 640386 161394 645524 161422
rect 640416 161366 645524 161394
rect 645580 161366 645585 161422
rect 640416 161364 645585 161366
rect 645519 161361 645585 161364
rect 184335 160980 184401 160983
rect 184335 160978 190560 160980
rect 184335 160922 184340 160978
rect 184396 160922 190560 160978
rect 184335 160920 190560 160922
rect 184335 160917 184401 160920
rect 149103 160684 149169 160687
rect 143904 160682 149169 160684
rect 143904 160626 149108 160682
rect 149164 160626 149169 160682
rect 143904 160624 149169 160626
rect 149103 160621 149169 160624
rect 184431 160388 184497 160391
rect 184431 160386 190014 160388
rect 184431 160330 184436 160386
rect 184492 160330 190014 160386
rect 184431 160328 190014 160330
rect 184431 160325 184497 160328
rect 189954 160314 190014 160328
rect 189954 160254 190560 160314
rect 148335 159500 148401 159503
rect 143904 159498 148401 159500
rect 143904 159442 148340 159498
rect 148396 159442 148401 159498
rect 143904 159440 148401 159442
rect 148335 159437 148401 159440
rect 184527 159500 184593 159503
rect 184527 159498 190560 159500
rect 184527 159442 184532 159498
rect 184588 159442 190560 159498
rect 184527 159440 190560 159442
rect 184527 159437 184593 159440
rect 184623 158908 184689 158911
rect 184623 158906 190014 158908
rect 184623 158850 184628 158906
rect 184684 158850 190014 158906
rect 184623 158848 190014 158850
rect 184623 158845 184689 158848
rect 189954 158834 190014 158848
rect 189954 158774 190560 158834
rect 143874 157724 143934 158212
rect 184431 158020 184497 158023
rect 184431 158018 190560 158020
rect 184431 157962 184436 158018
rect 184492 157962 190560 158018
rect 184431 157960 190560 157962
rect 184431 157957 184497 157960
rect 148815 157724 148881 157727
rect 143874 157722 148881 157724
rect 143874 157666 148820 157722
rect 148876 157666 148881 157722
rect 143874 157664 148881 157666
rect 148815 157661 148881 157664
rect 640386 157576 640446 159470
rect 675183 158760 675249 158763
rect 675138 158758 675249 158760
rect 675138 158702 675188 158758
rect 675244 158702 675249 158758
rect 675138 158697 675249 158702
rect 675138 158467 675198 158697
rect 675138 158462 675249 158467
rect 675138 158406 675188 158462
rect 675244 158406 675249 158462
rect 675138 158404 675249 158406
rect 675183 158401 675249 158404
rect 645519 157576 645585 157579
rect 640386 157574 645585 157576
rect 640386 157546 645524 157574
rect 640416 157518 645524 157546
rect 645580 157518 645585 157574
rect 640416 157516 645585 157518
rect 645519 157513 645585 157516
rect 184527 157428 184593 157431
rect 184527 157426 190014 157428
rect 184527 157370 184532 157426
rect 184588 157370 190014 157426
rect 184527 157368 190014 157370
rect 184527 157365 184593 157368
rect 189954 157354 190014 157368
rect 189954 157294 190560 157354
rect 148239 156984 148305 156987
rect 143904 156982 148305 156984
rect 143904 156926 148244 156982
rect 148300 156926 148305 156982
rect 143904 156924 148305 156926
rect 148239 156921 148305 156924
rect 184335 156540 184401 156543
rect 184335 156538 190560 156540
rect 184335 156482 184340 156538
rect 184396 156482 190560 156538
rect 184335 156480 190560 156482
rect 184335 156477 184401 156480
rect 148431 155800 148497 155803
rect 143904 155798 148497 155800
rect 143904 155742 148436 155798
rect 148492 155742 148497 155798
rect 143904 155740 148497 155742
rect 148431 155737 148497 155740
rect 184623 155652 184689 155655
rect 184623 155650 190560 155652
rect 184623 155594 184628 155650
rect 184684 155594 190560 155650
rect 184623 155592 190560 155594
rect 184623 155589 184689 155592
rect 640194 155504 640254 155622
rect 645135 155504 645201 155507
rect 640194 155502 645201 155504
rect 640194 155446 645140 155502
rect 645196 155446 645201 155502
rect 640194 155444 645201 155446
rect 184335 155060 184401 155063
rect 184335 155058 190560 155060
rect 184335 155002 184340 155058
rect 184396 155002 190560 155058
rect 184335 155000 190560 155002
rect 184335 154997 184401 155000
rect 148623 154616 148689 154619
rect 143904 154614 148689 154616
rect 143904 154558 148628 154614
rect 148684 154558 148689 154614
rect 143904 154556 148689 154558
rect 148623 154553 148689 154556
rect 184431 154172 184497 154175
rect 184431 154170 190560 154172
rect 184431 154114 184436 154170
rect 184492 154114 190560 154170
rect 184431 154112 190560 154114
rect 184431 154109 184497 154112
rect 640386 153772 640446 155444
rect 645135 155441 645201 155444
rect 184719 153580 184785 153583
rect 184719 153578 190014 153580
rect 184719 153522 184724 153578
rect 184780 153522 190014 153578
rect 184719 153520 190014 153522
rect 184719 153517 184785 153520
rect 189954 153506 190014 153520
rect 189954 153446 190560 153506
rect 674938 153370 674944 153434
rect 675008 153432 675014 153434
rect 675471 153432 675537 153435
rect 675008 153430 675537 153432
rect 675008 153374 675476 153430
rect 675532 153374 675537 153430
rect 675008 153372 675537 153374
rect 675008 153370 675014 153372
rect 675471 153369 675537 153372
rect 143874 152840 143934 153328
rect 148282 152840 148288 152842
rect 143874 152780 148288 152840
rect 148282 152778 148288 152780
rect 148352 152778 148358 152842
rect 184527 152692 184593 152695
rect 184527 152690 190560 152692
rect 184527 152634 184532 152690
rect 184588 152634 190560 152690
rect 184527 152632 190560 152634
rect 184527 152629 184593 152632
rect 645999 152544 646065 152547
rect 675375 152546 675441 152547
rect 675322 152544 675328 152546
rect 640194 152542 646065 152544
rect 640194 152486 646004 152542
rect 646060 152486 646065 152542
rect 640194 152484 646065 152486
rect 675284 152484 675328 152544
rect 675392 152542 675441 152546
rect 675436 152486 675441 152542
rect 148719 152100 148785 152103
rect 143904 152098 148785 152100
rect 143904 152042 148724 152098
rect 148780 152042 148785 152098
rect 143904 152040 148785 152042
rect 148719 152037 148785 152040
rect 184335 151952 184401 151955
rect 184335 151950 190014 151952
rect 184335 151894 184340 151950
rect 184396 151894 190014 151950
rect 184335 151892 190014 151894
rect 184335 151889 184401 151892
rect 189954 151878 190014 151892
rect 189954 151818 190560 151878
rect 184527 151212 184593 151215
rect 184527 151210 190560 151212
rect 184527 151154 184532 151210
rect 184588 151154 190560 151210
rect 184527 151152 190560 151154
rect 184527 151149 184593 151152
rect 148527 150916 148593 150919
rect 143904 150914 148593 150916
rect 143904 150858 148532 150914
rect 148588 150858 148593 150914
rect 143904 150856 148593 150858
rect 148527 150853 148593 150856
rect 184431 150472 184497 150475
rect 184431 150470 190014 150472
rect 184431 150414 184436 150470
rect 184492 150414 190014 150470
rect 184431 150412 190014 150414
rect 184431 150409 184497 150412
rect 189954 150398 190014 150412
rect 189954 150338 190560 150398
rect 640194 149998 640254 152484
rect 645999 152481 646065 152484
rect 675322 152482 675328 152484
rect 675392 152482 675441 152486
rect 675375 152481 675441 152482
rect 675130 151890 675136 151954
rect 675200 151952 675206 151954
rect 675471 151952 675537 151955
rect 675200 151950 675537 151952
rect 675200 151894 675476 151950
rect 675532 151894 675537 151950
rect 675200 151892 675537 151894
rect 675200 151890 675206 151892
rect 675471 151889 675537 151892
rect 675663 151362 675729 151363
rect 675663 151358 675712 151362
rect 675776 151360 675782 151362
rect 675663 151302 675668 151358
rect 675663 151298 675712 151302
rect 675776 151300 675820 151360
rect 675776 151298 675782 151300
rect 675663 151297 675729 151298
rect 673978 150262 673984 150326
rect 674048 150324 674054 150326
rect 675471 150324 675537 150327
rect 674048 150322 675537 150324
rect 674048 150266 675476 150322
rect 675532 150266 675537 150322
rect 674048 150264 675537 150266
rect 674048 150262 674054 150264
rect 675471 150261 675537 150264
rect 149583 149880 149649 149883
rect 143874 149878 149649 149880
rect 143874 149822 149588 149878
rect 149644 149822 149649 149878
rect 143874 149820 149649 149822
rect 143874 149776 143934 149820
rect 149583 149817 149649 149820
rect 184623 149732 184689 149735
rect 184623 149730 190560 149732
rect 184623 149674 184628 149730
rect 184684 149674 190560 149730
rect 184623 149672 190560 149674
rect 184623 149669 184689 149672
rect 184335 148992 184401 148995
rect 184335 148990 190014 148992
rect 184335 148934 184340 148990
rect 184396 148934 190014 148990
rect 184335 148932 190014 148934
rect 184335 148929 184401 148932
rect 189954 148918 190014 148932
rect 189954 148858 190560 148918
rect 148047 148548 148113 148551
rect 143904 148546 148113 148548
rect 143904 148490 148052 148546
rect 148108 148490 148113 148546
rect 143904 148488 148113 148490
rect 148047 148485 148113 148488
rect 674746 148486 674752 148550
rect 674816 148548 674822 148550
rect 675471 148548 675537 148551
rect 674816 148546 675537 148548
rect 674816 148490 675476 148546
rect 675532 148490 675537 148546
rect 674816 148488 675537 148490
rect 674816 148486 674822 148488
rect 675471 148485 675537 148488
rect 184431 148104 184497 148107
rect 645135 148104 645201 148107
rect 184431 148102 190560 148104
rect 184431 148046 184436 148102
rect 184492 148046 190560 148102
rect 640416 148102 645201 148104
rect 640416 148074 645140 148102
rect 184431 148044 190560 148046
rect 640386 148046 645140 148074
rect 645196 148046 645201 148102
rect 640386 148044 645201 148046
rect 184431 148041 184497 148044
rect 148047 147364 148113 147367
rect 143904 147362 148113 147364
rect 143904 147306 148052 147362
rect 148108 147306 148113 147362
rect 143904 147304 148113 147306
rect 148047 147301 148113 147304
rect 184527 147364 184593 147367
rect 184527 147362 190560 147364
rect 184527 147306 184532 147362
rect 184588 147306 190560 147362
rect 184527 147304 190560 147306
rect 184527 147301 184593 147304
rect 185775 146624 185841 146627
rect 185775 146622 190560 146624
rect 185775 146566 185780 146622
rect 185836 146566 190560 146622
rect 185775 146564 190560 146566
rect 185775 146561 185841 146564
rect 147951 146180 148017 146183
rect 143904 146178 148017 146180
rect 143904 146122 147956 146178
rect 148012 146122 148017 146178
rect 640386 146150 640446 148044
rect 645135 148041 645201 148044
rect 674554 146562 674560 146626
rect 674624 146624 674630 146626
rect 675375 146624 675441 146627
rect 674624 146622 675441 146624
rect 674624 146566 675380 146622
rect 675436 146566 675441 146622
rect 674624 146564 675441 146566
rect 674624 146562 674630 146564
rect 675375 146561 675441 146564
rect 143904 146120 148017 146122
rect 147951 146117 148017 146120
rect 184335 145884 184401 145887
rect 184335 145882 190560 145884
rect 184335 145826 184340 145882
rect 184396 145826 190560 145882
rect 184335 145824 190560 145826
rect 184335 145821 184401 145824
rect 184527 145144 184593 145147
rect 184527 145142 190014 145144
rect 184527 145086 184532 145142
rect 184588 145086 190014 145142
rect 184527 145084 190014 145086
rect 184527 145081 184593 145084
rect 189954 145070 190014 145084
rect 189954 145010 190560 145070
rect 143874 144404 143934 144892
rect 147951 144404 148017 144407
rect 143874 144402 148017 144404
rect 143874 144346 147956 144402
rect 148012 144346 148017 144402
rect 143874 144344 148017 144346
rect 147951 144341 148017 144344
rect 184431 144404 184497 144407
rect 184431 144402 190560 144404
rect 184431 144346 184436 144402
rect 184492 144346 190560 144402
rect 184431 144344 190560 144346
rect 184431 144341 184497 144344
rect 646479 144256 646545 144259
rect 640416 144254 646545 144256
rect 640416 144226 646484 144254
rect 640386 144198 646484 144226
rect 646540 144198 646545 144254
rect 640386 144196 646545 144198
rect 147855 143664 147921 143667
rect 143904 143662 147921 143664
rect 143904 143606 147860 143662
rect 147916 143606 147921 143662
rect 143904 143604 147921 143606
rect 147855 143601 147921 143604
rect 184431 143664 184497 143667
rect 184431 143662 190014 143664
rect 184431 143606 184436 143662
rect 184492 143606 190014 143662
rect 184431 143604 190014 143606
rect 184431 143601 184497 143604
rect 189954 143590 190014 143604
rect 189954 143530 190560 143590
rect 184335 142776 184401 142779
rect 184335 142774 190560 142776
rect 184335 142718 184340 142774
rect 184396 142718 190560 142774
rect 184335 142716 190560 142718
rect 184335 142713 184401 142716
rect 147855 142480 147921 142483
rect 143904 142478 147921 142480
rect 143904 142422 147860 142478
rect 147916 142422 147921 142478
rect 143904 142420 147921 142422
rect 147855 142417 147921 142420
rect 640386 142302 640446 144196
rect 646479 144193 646545 144196
rect 184527 142184 184593 142187
rect 184527 142182 190014 142184
rect 184527 142126 184532 142182
rect 184588 142126 190014 142182
rect 184527 142124 190014 142126
rect 184527 142121 184593 142124
rect 189954 142110 190014 142124
rect 189954 142050 190560 142110
rect 147663 141296 147729 141299
rect 143904 141294 147729 141296
rect 143904 141238 147668 141294
rect 147724 141238 147729 141294
rect 143904 141236 147729 141238
rect 147663 141233 147729 141236
rect 184623 141296 184689 141299
rect 184623 141294 190560 141296
rect 184623 141238 184628 141294
rect 184684 141238 190560 141294
rect 184623 141236 190560 141238
rect 184623 141233 184689 141236
rect 646575 141000 646641 141003
rect 640386 140998 646641 141000
rect 640386 140942 646580 140998
rect 646636 140942 646641 140998
rect 640386 140940 646641 140942
rect 184335 140556 184401 140559
rect 184335 140554 190560 140556
rect 184335 140498 184340 140554
rect 184396 140498 190560 140554
rect 184335 140496 190560 140498
rect 184335 140493 184401 140496
rect 640386 140408 640446 140940
rect 646575 140937 646641 140940
rect 640224 140378 640446 140408
rect 640194 140348 640416 140378
rect 149199 139964 149265 139967
rect 143904 139962 149265 139964
rect 143904 139906 149204 139962
rect 149260 139906 149265 139962
rect 143904 139904 149265 139906
rect 149199 139901 149265 139904
rect 184527 139816 184593 139819
rect 184527 139814 190560 139816
rect 184527 139758 184532 139814
rect 184588 139758 190560 139814
rect 184527 139756 190560 139758
rect 184527 139753 184593 139756
rect 184431 138928 184497 138931
rect 184431 138926 190560 138928
rect 184431 138870 184436 138926
rect 184492 138870 190560 138926
rect 184431 138868 190560 138870
rect 184431 138865 184497 138868
rect 147951 138780 148017 138783
rect 143904 138778 148017 138780
rect 143904 138722 147956 138778
rect 148012 138722 148017 138778
rect 143904 138720 148017 138722
rect 147951 138717 148017 138720
rect 640194 138528 640254 140348
rect 184623 138336 184689 138339
rect 184623 138334 190560 138336
rect 184623 138278 184628 138334
rect 184684 138278 190560 138334
rect 184623 138276 190560 138278
rect 184623 138273 184689 138276
rect 148047 137596 148113 137599
rect 143904 137594 148113 137596
rect 143904 137538 148052 137594
rect 148108 137538 148113 137594
rect 143904 137536 148113 137538
rect 148047 137533 148113 137536
rect 184335 137448 184401 137451
rect 184335 137446 190560 137448
rect 184335 137390 184340 137446
rect 184396 137390 190560 137446
rect 184335 137388 190560 137390
rect 184335 137385 184401 137388
rect 184527 136856 184593 136859
rect 184527 136854 190014 136856
rect 184527 136798 184532 136854
rect 184588 136798 190014 136854
rect 184527 136796 190014 136798
rect 184527 136793 184593 136796
rect 189954 136782 190014 136796
rect 189954 136722 190560 136782
rect 143874 135820 143934 136308
rect 184431 135968 184497 135971
rect 184431 135966 190560 135968
rect 184431 135910 184436 135966
rect 184492 135910 190560 135966
rect 184431 135908 190560 135910
rect 184431 135905 184497 135908
rect 149199 135820 149265 135823
rect 143874 135818 149265 135820
rect 143874 135762 149204 135818
rect 149260 135762 149265 135818
rect 143874 135760 149265 135762
rect 149199 135757 149265 135760
rect 184335 135228 184401 135231
rect 184335 135226 190014 135228
rect 184335 135170 184340 135226
rect 184396 135170 190014 135226
rect 184335 135168 190014 135170
rect 184335 135165 184401 135168
rect 189954 135154 190014 135168
rect 189954 135094 190560 135154
rect 147855 135080 147921 135083
rect 143904 135078 147921 135080
rect 143904 135022 147860 135078
rect 147916 135022 147921 135078
rect 143904 135020 147921 135022
rect 147855 135017 147921 135020
rect 646863 134784 646929 134787
rect 640416 134782 646929 134784
rect 640416 134726 646868 134782
rect 646924 134726 646929 134782
rect 640416 134724 646929 134726
rect 646863 134721 646929 134724
rect 184431 134488 184497 134491
rect 676143 134488 676209 134491
rect 676290 134488 676350 134680
rect 184431 134486 190560 134488
rect 184431 134430 184436 134486
rect 184492 134430 190560 134486
rect 184431 134428 190560 134430
rect 676143 134486 676350 134488
rect 676143 134430 676148 134486
rect 676204 134430 676350 134486
rect 676143 134428 676350 134430
rect 184431 134425 184497 134428
rect 676143 134425 676209 134428
rect 676239 134340 676305 134343
rect 676239 134338 676350 134340
rect 676239 134282 676244 134338
rect 676300 134282 676350 134338
rect 676239 134277 676350 134282
rect 676290 134162 676350 134277
rect 147663 133896 147729 133899
rect 143904 133894 147729 133896
rect 143904 133838 147668 133894
rect 147724 133838 147729 133894
rect 143904 133836 147729 133838
rect 147663 133833 147729 133836
rect 184335 133748 184401 133751
rect 184335 133746 190014 133748
rect 184335 133690 184340 133746
rect 184396 133690 190014 133746
rect 184335 133688 190014 133690
rect 184335 133685 184401 133688
rect 189954 133674 190014 133688
rect 189954 133614 190560 133674
rect 676290 133455 676350 133570
rect 676239 133450 676350 133455
rect 676239 133394 676244 133450
rect 676300 133394 676350 133450
rect 676239 133392 676350 133394
rect 676239 133389 676305 133392
rect 673362 133094 673368 133158
rect 673432 133156 673438 133158
rect 673432 133096 676320 133156
rect 673432 133094 673438 133096
rect 184527 133008 184593 133011
rect 184527 133006 190560 133008
rect 184527 132950 184532 133006
rect 184588 132950 190560 133006
rect 184527 132948 190560 132950
rect 184527 132945 184593 132948
rect 148143 132712 148209 132715
rect 143904 132710 148209 132712
rect 143904 132654 148148 132710
rect 148204 132654 148209 132710
rect 143904 132652 148209 132654
rect 148143 132649 148209 132652
rect 676047 132712 676113 132715
rect 676047 132710 676320 132712
rect 676047 132654 676052 132710
rect 676108 132654 676320 132710
rect 676047 132652 676320 132654
rect 676047 132649 676113 132652
rect 184335 132268 184401 132271
rect 184335 132266 190014 132268
rect 184335 132210 184340 132266
rect 184396 132210 190014 132266
rect 184335 132208 190014 132210
rect 184335 132205 184401 132208
rect 189954 132194 190014 132208
rect 189954 132134 190560 132194
rect 674514 132058 674520 132122
rect 674584 132120 674590 132122
rect 674584 132060 676320 132120
rect 674584 132058 674590 132060
rect 184431 131528 184497 131531
rect 184431 131526 190560 131528
rect 184431 131470 184436 131526
rect 184492 131470 190560 131526
rect 184431 131468 190560 131470
rect 184431 131465 184497 131468
rect 143874 130936 143934 131424
rect 676290 131383 676350 131646
rect 676239 131378 676350 131383
rect 676239 131322 676244 131378
rect 676300 131322 676350 131378
rect 676239 131320 676350 131322
rect 676239 131317 676305 131320
rect 673170 131170 673176 131234
rect 673240 131232 673246 131234
rect 673240 131172 676350 131232
rect 673240 131170 673246 131172
rect 676290 131128 676350 131172
rect 147567 130936 147633 130939
rect 647823 130936 647889 130939
rect 143874 130934 147633 130936
rect 143874 130878 147572 130934
rect 147628 130878 147633 130934
rect 143874 130876 147633 130878
rect 640416 130934 647889 130936
rect 640416 130878 647828 130934
rect 647884 130878 647889 130934
rect 640416 130876 647889 130878
rect 147567 130873 147633 130876
rect 647823 130873 647889 130876
rect 184527 130640 184593 130643
rect 676047 130640 676113 130643
rect 184527 130638 190560 130640
rect 184527 130582 184532 130638
rect 184588 130582 190560 130638
rect 184527 130580 190560 130582
rect 676047 130638 676320 130640
rect 676047 130582 676052 130638
rect 676108 130582 676320 130638
rect 676047 130580 676320 130582
rect 184527 130577 184593 130580
rect 676047 130577 676113 130580
rect 147759 130344 147825 130347
rect 143904 130342 147825 130344
rect 143904 130286 147764 130342
rect 147820 130286 147825 130342
rect 143904 130284 147825 130286
rect 147759 130281 147825 130284
rect 674938 130134 674944 130198
rect 675008 130196 675014 130198
rect 675008 130136 676320 130196
rect 675008 130134 675014 130136
rect 184623 129900 184689 129903
rect 184623 129898 190560 129900
rect 184623 129842 184628 129898
rect 184684 129842 190560 129898
rect 184623 129840 190560 129842
rect 184623 129837 184689 129840
rect 675706 129616 675712 129680
rect 675776 129678 675782 129680
rect 675776 129618 676320 129678
rect 675776 129616 675782 129618
rect 147087 129160 147153 129163
rect 143904 129158 147153 129160
rect 143904 129102 147092 129158
rect 147148 129102 147153 129158
rect 143904 129100 147153 129102
rect 147087 129097 147153 129100
rect 184335 129160 184401 129163
rect 675471 129160 675537 129163
rect 184335 129158 190560 129160
rect 184335 129102 184340 129158
rect 184396 129102 190560 129158
rect 184335 129100 190560 129102
rect 675471 129158 676320 129160
rect 675471 129102 675476 129158
rect 675532 129102 676320 129158
rect 675471 129100 676320 129102
rect 184335 129097 184401 129100
rect 675471 129097 675537 129100
rect 646575 129012 646641 129015
rect 640416 129010 646641 129012
rect 640416 128954 646580 129010
rect 646636 128954 646641 129010
rect 640416 128952 646641 128954
rect 646575 128949 646641 128952
rect 675130 128654 675136 128718
rect 675200 128716 675206 128718
rect 675200 128656 676320 128716
rect 675200 128654 675206 128656
rect 184431 128420 184497 128423
rect 184431 128418 190014 128420
rect 184431 128362 184436 128418
rect 184492 128362 190014 128418
rect 184431 128360 190014 128362
rect 184431 128357 184497 128360
rect 189954 128346 190014 128360
rect 189954 128286 190560 128346
rect 674362 128062 674368 128126
rect 674432 128124 674438 128126
rect 674432 128064 676320 128124
rect 674432 128062 674438 128064
rect 149295 127976 149361 127979
rect 143904 127974 149361 127976
rect 143904 127918 149300 127974
rect 149356 127918 149361 127974
rect 143904 127916 149361 127918
rect 149295 127913 149361 127916
rect 184527 127680 184593 127683
rect 646767 127680 646833 127683
rect 184527 127678 190560 127680
rect 184527 127622 184532 127678
rect 184588 127622 190560 127678
rect 184527 127620 190560 127622
rect 640386 127678 646833 127680
rect 640386 127622 646772 127678
rect 646828 127622 646833 127678
rect 640386 127620 646833 127622
rect 184527 127617 184593 127620
rect 640386 127058 640446 127620
rect 646767 127617 646833 127620
rect 675322 127618 675328 127682
rect 675392 127680 675398 127682
rect 675392 127620 676320 127680
rect 675392 127618 675398 127620
rect 676047 127236 676113 127239
rect 676047 127234 676320 127236
rect 676047 127178 676052 127234
rect 676108 127178 676320 127234
rect 676047 127176 676320 127178
rect 676047 127173 676113 127176
rect 184719 126940 184785 126943
rect 184719 126938 190014 126940
rect 184719 126882 184724 126938
rect 184780 126882 190014 126938
rect 184719 126880 190014 126882
rect 184719 126877 184785 126880
rect 189954 126866 190014 126880
rect 189954 126806 190560 126866
rect 147183 126644 147249 126647
rect 143904 126642 147249 126644
rect 143904 126586 147188 126642
rect 147244 126586 147249 126642
rect 143904 126584 147249 126586
rect 147183 126581 147249 126584
rect 676290 126499 676350 126614
rect 676239 126494 676350 126499
rect 676239 126438 676244 126494
rect 676300 126438 676350 126494
rect 676239 126436 676350 126438
rect 676239 126433 676305 126436
rect 676047 126126 676113 126129
rect 676047 126124 676320 126126
rect 676047 126068 676052 126124
rect 676108 126068 676320 126124
rect 676047 126066 676320 126068
rect 676047 126063 676113 126066
rect 184335 126052 184401 126055
rect 184335 126050 190560 126052
rect 184335 125994 184340 126050
rect 184396 125994 190560 126050
rect 184335 125992 190560 125994
rect 184335 125989 184401 125992
rect 646671 125756 646737 125759
rect 640386 125754 646737 125756
rect 640386 125698 646676 125754
rect 646732 125698 646737 125754
rect 640386 125696 646737 125698
rect 147279 125460 147345 125463
rect 143904 125458 147345 125460
rect 143904 125402 147284 125458
rect 147340 125402 147345 125458
rect 143904 125400 147345 125402
rect 147279 125397 147345 125400
rect 186831 125460 186897 125463
rect 186831 125458 190014 125460
rect 186831 125402 186836 125458
rect 186892 125402 190014 125458
rect 186831 125400 190014 125402
rect 186831 125397 186897 125400
rect 189954 125386 190014 125400
rect 189954 125326 190560 125386
rect 640386 125208 640446 125696
rect 646671 125693 646737 125696
rect 674554 125694 674560 125758
rect 674624 125756 674630 125758
rect 674624 125696 676320 125756
rect 674624 125694 674630 125696
rect 674746 125102 674752 125166
rect 674816 125164 674822 125166
rect 674816 125104 676320 125164
rect 674816 125102 674822 125104
rect 676047 124646 676113 124649
rect 676047 124644 676320 124646
rect 676047 124588 676052 124644
rect 676108 124588 676320 124644
rect 676047 124586 676320 124588
rect 676047 124583 676113 124586
rect 184431 124572 184497 124575
rect 184431 124570 190560 124572
rect 184431 124514 184436 124570
rect 184492 124514 190560 124570
rect 184431 124512 190560 124514
rect 184431 124509 184497 124512
rect 147375 124276 147441 124279
rect 143904 124274 147441 124276
rect 143904 124218 147380 124274
rect 147436 124218 147441 124274
rect 143904 124216 147441 124218
rect 147375 124213 147441 124216
rect 675951 124276 676017 124279
rect 675951 124274 676320 124276
rect 675951 124218 675956 124274
rect 676012 124218 676320 124274
rect 675951 124216 676320 124218
rect 675951 124213 676017 124216
rect 184335 123832 184401 123835
rect 647919 123832 647985 123835
rect 184335 123830 190560 123832
rect 184335 123774 184340 123830
rect 184396 123774 190560 123830
rect 184335 123772 190560 123774
rect 640194 123830 647985 123832
rect 640194 123774 647924 123830
rect 647980 123774 647985 123830
rect 640194 123772 647985 123774
rect 184335 123769 184401 123772
rect 640194 123358 640254 123772
rect 647919 123769 647985 123772
rect 676047 123684 676113 123687
rect 676047 123682 676320 123684
rect 676047 123626 676052 123682
rect 676108 123626 676320 123682
rect 676047 123624 676320 123626
rect 676047 123621 676113 123624
rect 184623 123092 184689 123095
rect 184623 123090 190560 123092
rect 184623 123034 184628 123090
rect 184684 123034 190560 123090
rect 184623 123032 190560 123034
rect 184623 123029 184689 123032
rect 143874 122500 143934 122988
rect 676290 122947 676350 123062
rect 676290 122942 676401 122947
rect 676290 122886 676340 122942
rect 676396 122886 676401 122942
rect 676290 122884 676401 122886
rect 676335 122881 676401 122884
rect 147471 122500 147537 122503
rect 143874 122498 147537 122500
rect 143874 122442 147476 122498
rect 147532 122442 147537 122498
rect 143874 122440 147537 122442
rect 147471 122437 147537 122440
rect 676143 122500 676209 122503
rect 676290 122500 676350 122692
rect 676143 122498 676350 122500
rect 676143 122442 676148 122498
rect 676204 122442 676350 122498
rect 676143 122440 676350 122442
rect 676143 122437 676209 122440
rect 184431 122204 184497 122207
rect 184431 122202 190560 122204
rect 184431 122146 184436 122202
rect 184492 122146 190560 122202
rect 184431 122144 190560 122146
rect 184431 122141 184497 122144
rect 647727 122056 647793 122059
rect 640194 122054 647793 122056
rect 640194 121998 647732 122054
rect 647788 121998 647793 122054
rect 640194 121996 647793 121998
rect 149295 121760 149361 121763
rect 143904 121758 149361 121760
rect 143904 121702 149300 121758
rect 149356 121702 149361 121758
rect 143904 121700 149361 121702
rect 149295 121697 149361 121700
rect 184527 121612 184593 121615
rect 184527 121610 190560 121612
rect 184527 121554 184532 121610
rect 184588 121554 190560 121610
rect 184527 121552 190560 121554
rect 184527 121549 184593 121552
rect 640194 121434 640254 121996
rect 647727 121993 647793 121996
rect 676290 121911 676350 122174
rect 676239 121906 676350 121911
rect 676239 121850 676244 121906
rect 676300 121850 676350 121906
rect 676239 121848 676350 121850
rect 676239 121845 676305 121848
rect 184335 120724 184401 120727
rect 184335 120722 190560 120724
rect 184335 120666 184340 120722
rect 184396 120666 190560 120722
rect 184335 120664 190560 120666
rect 184335 120661 184401 120664
rect 146991 120576 147057 120579
rect 143904 120574 147057 120576
rect 143904 120518 146996 120574
rect 147052 120518 147057 120574
rect 143904 120516 147057 120518
rect 146991 120513 147057 120516
rect 184527 120132 184593 120135
rect 184527 120130 190014 120132
rect 184527 120074 184532 120130
rect 184588 120074 190014 120130
rect 184527 120072 190014 120074
rect 184527 120069 184593 120072
rect 189954 120058 190014 120072
rect 189954 119998 190560 120058
rect 647919 119540 647985 119543
rect 640416 119538 647985 119540
rect 640416 119482 647924 119538
rect 647980 119482 647985 119538
rect 640416 119480 647985 119482
rect 647919 119477 647985 119480
rect 149199 119392 149265 119395
rect 143904 119390 149265 119392
rect 143904 119334 149204 119390
rect 149260 119334 149265 119390
rect 143904 119332 149265 119334
rect 149199 119329 149265 119332
rect 184623 119244 184689 119247
rect 184623 119242 190560 119244
rect 184623 119186 184628 119242
rect 184684 119186 190560 119242
rect 184623 119184 190560 119186
rect 184623 119181 184689 119184
rect 184431 118652 184497 118655
rect 184431 118650 190014 118652
rect 184431 118594 184436 118650
rect 184492 118594 190014 118650
rect 184431 118592 190014 118594
rect 184431 118589 184497 118592
rect 189954 118578 190014 118592
rect 189954 118518 190560 118578
rect 148911 118208 148977 118211
rect 143874 118206 148977 118208
rect 143874 118150 148916 118206
rect 148972 118150 148977 118206
rect 143874 118148 148977 118150
rect 143874 118104 143934 118148
rect 148911 118145 148977 118148
rect 184335 117764 184401 117767
rect 184335 117762 190560 117764
rect 184335 117706 184340 117762
rect 184396 117706 190560 117762
rect 184335 117704 190560 117706
rect 184335 117701 184401 117704
rect 646671 117616 646737 117619
rect 640416 117614 646737 117616
rect 640416 117558 646676 117614
rect 646732 117558 646737 117614
rect 640416 117556 646737 117558
rect 646671 117553 646737 117556
rect 184431 117024 184497 117027
rect 184431 117022 190014 117024
rect 184431 116966 184436 117022
rect 184492 116966 190014 117022
rect 184431 116964 190014 116966
rect 184431 116961 184497 116964
rect 189954 116950 190014 116964
rect 189954 116890 190560 116950
rect 149103 116876 149169 116879
rect 143904 116874 149169 116876
rect 143904 116818 149108 116874
rect 149164 116818 149169 116874
rect 143904 116816 149169 116818
rect 149103 116813 149169 116816
rect 184623 116284 184689 116287
rect 184623 116282 190560 116284
rect 184623 116226 184628 116282
rect 184684 116226 190560 116282
rect 184623 116224 190560 116226
rect 184623 116221 184689 116224
rect 149583 115692 149649 115695
rect 647919 115692 647985 115695
rect 143904 115690 149649 115692
rect 143904 115634 149588 115690
rect 149644 115634 149649 115690
rect 143904 115632 149649 115634
rect 640416 115690 647985 115692
rect 640416 115634 647924 115690
rect 647980 115634 647985 115690
rect 640416 115632 647985 115634
rect 149583 115629 149649 115632
rect 647919 115629 647985 115632
rect 184527 115396 184593 115399
rect 184527 115394 190560 115396
rect 184527 115338 184532 115394
rect 184588 115338 190560 115394
rect 184527 115336 190560 115338
rect 184527 115333 184593 115336
rect 184335 114804 184401 114807
rect 184335 114802 190560 114804
rect 184335 114746 184340 114802
rect 184396 114746 190560 114802
rect 184335 114744 190560 114746
rect 184335 114741 184401 114744
rect 149007 114508 149073 114511
rect 143904 114506 149073 114508
rect 143904 114450 149012 114506
rect 149068 114450 149073 114506
rect 143904 114448 149073 114450
rect 149007 114445 149073 114448
rect 674938 114298 674944 114362
rect 675008 114360 675014 114362
rect 675375 114360 675441 114363
rect 675008 114358 675441 114360
rect 675008 114302 675380 114358
rect 675436 114302 675441 114358
rect 675008 114300 675441 114302
rect 675008 114298 675014 114300
rect 675375 114297 675441 114300
rect 184431 113916 184497 113919
rect 184431 113914 190560 113916
rect 184431 113858 184436 113914
rect 184492 113858 190560 113914
rect 184431 113856 190560 113858
rect 184431 113853 184497 113856
rect 149487 113176 149553 113179
rect 143904 113174 149553 113176
rect 143904 113118 149492 113174
rect 149548 113118 149553 113174
rect 143904 113116 149553 113118
rect 149487 113113 149553 113116
rect 184527 113176 184593 113179
rect 640194 113176 640254 113738
rect 646575 113176 646641 113179
rect 184527 113174 190560 113176
rect 184527 113118 184532 113174
rect 184588 113118 190560 113174
rect 184527 113116 190560 113118
rect 640194 113174 646641 113176
rect 640194 113118 646580 113174
rect 646636 113118 646641 113174
rect 640194 113116 646641 113118
rect 184527 113113 184593 113116
rect 646575 113113 646641 113116
rect 184623 112436 184689 112439
rect 184623 112434 190560 112436
rect 184623 112378 184628 112434
rect 184684 112378 190560 112434
rect 184623 112376 190560 112378
rect 184623 112373 184689 112376
rect 675130 112226 675136 112290
rect 675200 112288 675206 112290
rect 675375 112288 675441 112291
rect 675200 112286 675441 112288
rect 675200 112230 675380 112286
rect 675436 112230 675441 112286
rect 675200 112228 675441 112230
rect 675200 112226 675206 112228
rect 675375 112225 675441 112228
rect 146895 111992 146961 111995
rect 143904 111990 146961 111992
rect 143904 111934 146900 111990
rect 146956 111934 146961 111990
rect 143904 111932 146961 111934
rect 146895 111929 146961 111932
rect 184431 111696 184497 111699
rect 184431 111694 190014 111696
rect 184431 111638 184436 111694
rect 184492 111638 190014 111694
rect 184431 111636 190014 111638
rect 184431 111633 184497 111636
rect 189954 111622 190014 111636
rect 189954 111562 190560 111622
rect 640386 111400 640446 111888
rect 647055 111400 647121 111403
rect 640386 111398 647121 111400
rect 640386 111342 647060 111398
rect 647116 111342 647121 111398
rect 640386 111340 647121 111342
rect 647055 111337 647121 111340
rect 148815 110956 148881 110959
rect 143904 110954 148881 110956
rect 143904 110898 148820 110954
rect 148876 110898 148881 110954
rect 143904 110896 148881 110898
rect 148815 110893 148881 110896
rect 184335 110956 184401 110959
rect 184335 110954 190560 110956
rect 184335 110898 184340 110954
rect 184396 110898 190560 110954
rect 184335 110896 190560 110898
rect 184335 110893 184401 110896
rect 184527 110216 184593 110219
rect 184527 110214 190014 110216
rect 184527 110158 184532 110214
rect 184588 110158 190014 110214
rect 184527 110156 190014 110158
rect 184527 110153 184593 110156
rect 189954 110142 190014 110156
rect 189954 110082 190560 110142
rect 143874 109476 143934 109668
rect 148335 109476 148401 109479
rect 143874 109474 148401 109476
rect 143874 109418 148340 109474
rect 148396 109418 148401 109474
rect 143874 109416 148401 109418
rect 640386 109476 640446 109890
rect 646671 109476 646737 109479
rect 640386 109474 646737 109476
rect 640386 109418 646676 109474
rect 646732 109418 646737 109474
rect 640386 109416 646737 109418
rect 148335 109413 148401 109416
rect 646671 109413 646737 109416
rect 148282 109266 148288 109330
rect 148352 109328 148358 109330
rect 148352 109268 190560 109328
rect 148352 109266 148358 109268
rect 184431 108736 184497 108739
rect 184431 108734 190014 108736
rect 184431 108678 184436 108734
rect 184492 108678 190014 108734
rect 184431 108676 190014 108678
rect 184431 108673 184497 108676
rect 189954 108662 190014 108676
rect 189954 108602 190560 108662
rect 148431 108440 148497 108443
rect 143904 108438 148497 108440
rect 143904 108382 148436 108438
rect 148492 108382 148497 108438
rect 143904 108380 148497 108382
rect 148431 108377 148497 108380
rect 674362 108082 674368 108146
rect 674432 108144 674438 108146
rect 675471 108144 675537 108147
rect 674432 108142 675537 108144
rect 674432 108086 675476 108142
rect 675532 108086 675537 108142
rect 674432 108084 675537 108086
rect 674432 108082 674438 108084
rect 675471 108081 675537 108084
rect 646767 107996 646833 107999
rect 640416 107994 646833 107996
rect 640416 107938 646772 107994
rect 646828 107938 646833 107994
rect 640416 107936 646833 107938
rect 646767 107933 646833 107936
rect 184335 107848 184401 107851
rect 184335 107846 190560 107848
rect 184335 107790 184340 107846
rect 184396 107790 190560 107846
rect 184335 107788 190560 107790
rect 184335 107785 184401 107788
rect 148623 107256 148689 107259
rect 143904 107254 148689 107256
rect 143904 107198 148628 107254
rect 148684 107198 148689 107254
rect 143904 107196 148689 107198
rect 148623 107193 148689 107196
rect 184527 107108 184593 107111
rect 184527 107106 190560 107108
rect 184527 107050 184532 107106
rect 184588 107050 190560 107106
rect 184527 107048 190560 107050
rect 184527 107045 184593 107048
rect 184431 106368 184497 106371
rect 669519 106368 669585 106371
rect 184431 106366 190560 106368
rect 184431 106310 184436 106366
rect 184492 106310 190560 106366
rect 184431 106308 190560 106310
rect 665346 106366 669585 106368
rect 665346 106310 669524 106366
rect 669580 106310 669585 106366
rect 665346 106308 669585 106310
rect 184431 106305 184497 106308
rect 665346 106082 665406 106308
rect 669519 106305 669585 106308
rect 674746 106306 674752 106370
rect 674816 106368 674822 106370
rect 675375 106368 675441 106371
rect 674816 106366 675441 106368
rect 674816 106310 675380 106366
rect 675436 106310 675441 106366
rect 674816 106308 675441 106310
rect 674816 106306 674822 106308
rect 675375 106305 675441 106308
rect 147951 106072 148017 106075
rect 645903 106072 645969 106075
rect 143904 106070 148017 106072
rect 143904 106014 147956 106070
rect 148012 106014 148017 106070
rect 143904 106012 148017 106014
rect 640416 106070 645969 106072
rect 640416 106014 645908 106070
rect 645964 106014 645969 106070
rect 640416 106012 645969 106014
rect 147951 106009 148017 106012
rect 645903 106009 645969 106012
rect 184335 105628 184401 105631
rect 184335 105626 190560 105628
rect 184335 105570 184340 105626
rect 184396 105570 190560 105626
rect 184335 105568 190560 105570
rect 184335 105565 184401 105568
rect 665346 105332 665406 105361
rect 668175 105332 668241 105335
rect 665346 105330 668241 105332
rect 665346 105274 668180 105330
rect 668236 105274 668241 105330
rect 665346 105272 668241 105274
rect 668175 105269 668241 105272
rect 665295 105184 665361 105187
rect 665295 105182 665406 105184
rect 665295 105126 665300 105182
rect 665356 105126 665406 105182
rect 665295 105121 665406 105126
rect 674554 105122 674560 105186
rect 674624 105184 674630 105186
rect 675375 105184 675441 105187
rect 674624 105182 675441 105184
rect 674624 105126 675380 105182
rect 675436 105126 675441 105182
rect 674624 105124 675441 105126
rect 674624 105122 674630 105124
rect 675375 105121 675441 105124
rect 665346 104996 665406 105121
rect 184527 104888 184593 104891
rect 184527 104886 190014 104888
rect 184527 104830 184532 104886
rect 184588 104830 190014 104886
rect 184527 104828 190014 104830
rect 184527 104825 184593 104828
rect 189954 104814 190014 104828
rect 189954 104754 190560 104814
rect 148047 104740 148113 104743
rect 143904 104738 148113 104740
rect 143904 104682 148052 104738
rect 148108 104682 148113 104738
rect 143904 104680 148113 104682
rect 148047 104677 148113 104680
rect 647919 104148 647985 104151
rect 640416 104146 647985 104148
rect 640416 104090 647924 104146
rect 647980 104090 647985 104146
rect 640416 104088 647985 104090
rect 647919 104085 647985 104088
rect 184623 104000 184689 104003
rect 184623 103998 190560 104000
rect 184623 103942 184628 103998
rect 184684 103942 190560 103998
rect 184623 103940 190560 103942
rect 184623 103937 184689 103940
rect 147663 103556 147729 103559
rect 143904 103554 147729 103556
rect 143904 103498 147668 103554
rect 147724 103498 147729 103554
rect 143904 103496 147729 103498
rect 147663 103493 147729 103496
rect 184335 103408 184401 103411
rect 184335 103406 190014 103408
rect 184335 103350 184340 103406
rect 184396 103350 190014 103406
rect 184335 103348 190014 103350
rect 184335 103345 184401 103348
rect 189954 103334 190014 103348
rect 189954 103274 190560 103334
rect 675663 103262 675729 103263
rect 675663 103258 675712 103262
rect 675776 103260 675782 103262
rect 675663 103202 675668 103258
rect 675663 103198 675712 103202
rect 675776 103200 675820 103260
rect 675776 103198 675782 103200
rect 675663 103197 675729 103198
rect 184527 102520 184593 102523
rect 184527 102518 190560 102520
rect 184527 102462 184532 102518
rect 184588 102462 190560 102518
rect 184527 102460 190560 102462
rect 184527 102457 184593 102460
rect 148527 102372 148593 102375
rect 143904 102370 148593 102372
rect 143904 102314 148532 102370
rect 148588 102314 148593 102370
rect 143904 102312 148593 102314
rect 148527 102309 148593 102312
rect 645135 102224 645201 102227
rect 640416 102222 645201 102224
rect 640416 102166 645140 102222
rect 645196 102166 645201 102222
rect 640416 102164 645201 102166
rect 645135 102161 645201 102164
rect 184431 101928 184497 101931
rect 184431 101926 190014 101928
rect 184431 101870 184436 101926
rect 184492 101870 190014 101926
rect 184431 101868 190014 101870
rect 184431 101865 184497 101868
rect 189954 101854 190014 101868
rect 189954 101794 190560 101854
rect 675375 101486 675441 101487
rect 675322 101484 675328 101486
rect 675284 101424 675328 101484
rect 675392 101482 675441 101486
rect 675436 101426 675441 101482
rect 675322 101422 675328 101424
rect 675392 101422 675441 101426
rect 675375 101421 675441 101422
rect 143874 100892 143934 101084
rect 184623 101040 184689 101043
rect 184623 101038 190560 101040
rect 184623 100982 184628 101038
rect 184684 100982 190560 101038
rect 184623 100980 190560 100982
rect 184623 100977 184689 100980
rect 149679 100892 149745 100895
rect 143874 100890 149745 100892
rect 143874 100834 149684 100890
rect 149740 100834 149745 100890
rect 143874 100832 149745 100834
rect 149679 100829 149745 100832
rect 184335 100300 184401 100303
rect 184335 100298 190014 100300
rect 184335 100242 184340 100298
rect 184396 100242 190014 100298
rect 184335 100240 190014 100242
rect 184335 100237 184401 100240
rect 189954 100226 190014 100240
rect 189954 100166 190560 100226
rect 148239 99856 148305 99859
rect 143904 99854 148305 99856
rect 143904 99798 148244 99854
rect 148300 99798 148305 99854
rect 143904 99796 148305 99798
rect 148239 99793 148305 99796
rect 640194 99708 640254 100270
rect 647919 99708 647985 99711
rect 640194 99706 647985 99708
rect 640194 99650 647924 99706
rect 647980 99650 647985 99706
rect 640194 99648 647985 99650
rect 647919 99645 647985 99648
rect 184431 99560 184497 99563
rect 184431 99558 190560 99560
rect 184431 99502 184436 99558
rect 184492 99502 190560 99558
rect 184431 99500 190560 99502
rect 184431 99497 184497 99500
rect 148143 98672 148209 98675
rect 143904 98670 148209 98672
rect 143904 98614 148148 98670
rect 148204 98614 148209 98670
rect 143904 98612 148209 98614
rect 148143 98609 148209 98612
rect 184527 98672 184593 98675
rect 184527 98670 190560 98672
rect 184527 98614 184532 98670
rect 184588 98614 190560 98670
rect 184527 98612 190560 98614
rect 184527 98609 184593 98612
rect 184623 98080 184689 98083
rect 640386 98080 640446 98420
rect 646959 98080 647025 98083
rect 184623 98078 190560 98080
rect 184623 98022 184628 98078
rect 184684 98022 190560 98078
rect 184623 98020 190560 98022
rect 640386 98078 647025 98080
rect 640386 98022 646964 98078
rect 647020 98022 647025 98078
rect 640386 98020 647025 98022
rect 184623 98017 184689 98020
rect 646959 98017 647025 98020
rect 148719 97488 148785 97491
rect 143904 97486 148785 97488
rect 143904 97430 148724 97486
rect 148780 97430 148785 97486
rect 143904 97428 148785 97430
rect 148719 97425 148785 97428
rect 184335 97192 184401 97195
rect 184335 97190 190560 97192
rect 184335 97134 184340 97190
rect 184396 97134 190560 97190
rect 184335 97132 190560 97134
rect 184335 97129 184401 97132
rect 184431 96452 184497 96455
rect 184431 96450 190560 96452
rect 184431 96394 184436 96450
rect 184492 96394 190560 96450
rect 184431 96392 190560 96394
rect 184431 96389 184497 96392
rect 143874 95712 143934 96200
rect 640386 96008 640446 96570
rect 645423 96008 645489 96011
rect 640386 96006 645489 96008
rect 640386 95950 645428 96006
rect 645484 95950 645489 96006
rect 640386 95948 645489 95950
rect 645423 95945 645489 95948
rect 149487 95712 149553 95715
rect 143874 95710 149553 95712
rect 143874 95654 149492 95710
rect 149548 95654 149553 95710
rect 143874 95652 149553 95654
rect 149487 95649 149553 95652
rect 184527 95712 184593 95715
rect 184527 95710 190560 95712
rect 184527 95654 184532 95710
rect 184588 95654 190560 95710
rect 184527 95652 190560 95654
rect 184527 95649 184593 95652
rect 147567 94972 147633 94975
rect 143904 94970 147633 94972
rect 143904 94914 147572 94970
rect 147628 94914 147633 94970
rect 143904 94912 147633 94914
rect 147567 94909 147633 94912
rect 184335 94972 184401 94975
rect 184335 94970 190014 94972
rect 184335 94914 184340 94970
rect 184396 94914 190014 94970
rect 184335 94912 190014 94914
rect 184335 94909 184401 94912
rect 189954 94898 190014 94912
rect 189954 94838 190560 94898
rect 184527 94232 184593 94235
rect 184527 94230 190560 94232
rect 184527 94174 184532 94230
rect 184588 94174 190560 94230
rect 184527 94172 190560 94174
rect 184527 94169 184593 94172
rect 640386 94084 640446 94646
rect 647727 94084 647793 94087
rect 640386 94082 647793 94084
rect 640386 94026 647732 94082
rect 647788 94026 647793 94082
rect 640386 94024 647793 94026
rect 647727 94021 647793 94024
rect 149199 93788 149265 93791
rect 143904 93786 149265 93788
rect 143904 93730 149204 93786
rect 149260 93730 149265 93786
rect 143904 93728 149265 93730
rect 149199 93725 149265 93728
rect 184431 93492 184497 93495
rect 184431 93490 190014 93492
rect 184431 93434 184436 93490
rect 184492 93434 190014 93490
rect 184431 93432 190014 93434
rect 184431 93429 184497 93432
rect 189954 93418 190014 93432
rect 189954 93358 190560 93418
rect 184335 92752 184401 92755
rect 647823 92752 647889 92755
rect 184335 92750 190560 92752
rect 184335 92694 184340 92750
rect 184396 92694 190560 92750
rect 184335 92692 190560 92694
rect 640416 92750 647889 92752
rect 640416 92694 647828 92750
rect 647884 92694 647889 92750
rect 640416 92692 647889 92694
rect 184335 92689 184401 92692
rect 647823 92689 647889 92692
rect 148911 92604 148977 92607
rect 143904 92602 148977 92604
rect 143904 92546 148916 92602
rect 148972 92546 148977 92602
rect 143904 92544 148977 92546
rect 148911 92541 148977 92544
rect 189954 91878 190560 91938
rect 184335 91864 184401 91867
rect 189954 91864 190014 91878
rect 184335 91862 190014 91864
rect 184335 91806 184340 91862
rect 184396 91806 190014 91862
rect 184335 91804 190014 91806
rect 184335 91801 184401 91804
rect 149007 91420 149073 91423
rect 143904 91418 149073 91420
rect 143904 91362 149012 91418
rect 149068 91362 149073 91418
rect 143904 91360 149073 91362
rect 149007 91357 149073 91360
rect 184431 91124 184497 91127
rect 184431 91122 190560 91124
rect 184431 91066 184436 91122
rect 184492 91066 190560 91122
rect 184431 91064 190560 91066
rect 184431 91061 184497 91064
rect 659343 90828 659409 90831
rect 640416 90826 659409 90828
rect 640416 90770 659348 90826
rect 659404 90770 659409 90826
rect 640416 90768 659409 90770
rect 659343 90765 659409 90768
rect 184527 90384 184593 90387
rect 184527 90382 190560 90384
rect 184527 90326 184532 90382
rect 184588 90326 190560 90382
rect 184527 90324 190560 90326
rect 184527 90321 184593 90324
rect 149103 90236 149169 90239
rect 143904 90234 149169 90236
rect 143904 90178 149108 90234
rect 149164 90178 149169 90234
rect 143904 90176 149169 90178
rect 149103 90173 149169 90176
rect 184623 89644 184689 89647
rect 184623 89642 190560 89644
rect 184623 89586 184628 89642
rect 184684 89586 190560 89642
rect 184623 89584 190560 89586
rect 184623 89581 184689 89584
rect 149295 89052 149361 89055
rect 143904 89050 149361 89052
rect 143904 88994 149300 89050
rect 149356 88994 149361 89050
rect 143904 88992 149361 88994
rect 149295 88989 149361 88992
rect 184335 88904 184401 88907
rect 645903 88904 645969 88907
rect 184335 88902 190560 88904
rect 184335 88846 184340 88902
rect 184396 88846 190560 88902
rect 184335 88844 190560 88846
rect 640416 88902 645969 88904
rect 640416 88846 645908 88902
rect 645964 88846 645969 88902
rect 640416 88844 645969 88846
rect 184335 88841 184401 88844
rect 645903 88841 645969 88844
rect 184527 88164 184593 88167
rect 184527 88162 190014 88164
rect 184527 88106 184532 88162
rect 184588 88106 190014 88162
rect 184527 88104 190014 88106
rect 184527 88101 184593 88104
rect 189954 88090 190014 88104
rect 189954 88030 190560 88090
rect 143874 87276 143934 87764
rect 149391 87276 149457 87279
rect 143874 87274 149457 87276
rect 143874 87218 149396 87274
rect 149452 87218 149457 87274
rect 143874 87216 149457 87218
rect 149391 87213 149457 87216
rect 184431 87276 184497 87279
rect 184431 87274 190560 87276
rect 184431 87218 184436 87274
rect 184492 87218 190560 87274
rect 184431 87216 190560 87218
rect 184431 87213 184497 87216
rect 647919 87128 647985 87131
rect 640386 87126 647985 87128
rect 640386 87070 647924 87126
rect 647980 87070 647985 87126
rect 640386 87068 647985 87070
rect 640386 86950 640446 87068
rect 647919 87065 647985 87068
rect 653679 86980 653745 86983
rect 653679 86978 656736 86980
rect 653679 86922 653684 86978
rect 653740 86922 656736 86978
rect 653679 86920 656736 86922
rect 653679 86917 653745 86920
rect 184623 86684 184689 86687
rect 184623 86682 190014 86684
rect 184623 86626 184628 86682
rect 184684 86626 190014 86682
rect 184623 86624 190014 86626
rect 184623 86621 184689 86624
rect 189954 86610 190014 86624
rect 189954 86550 190560 86610
rect 148815 86536 148881 86539
rect 143904 86534 148881 86536
rect 143904 86478 148820 86534
rect 148876 86478 148881 86534
rect 143904 86476 148881 86478
rect 148815 86473 148881 86476
rect 663279 86388 663345 86391
rect 663234 86386 663345 86388
rect 663234 86330 663284 86386
rect 663340 86330 663345 86386
rect 663234 86325 663345 86330
rect 650895 86240 650961 86243
rect 650895 86238 656736 86240
rect 650895 86182 650900 86238
rect 650956 86182 656736 86238
rect 663234 86210 663294 86325
rect 650895 86180 656736 86182
rect 650895 86177 650961 86180
rect 184335 85796 184401 85799
rect 184335 85794 190560 85796
rect 184335 85738 184340 85794
rect 184396 85738 190560 85794
rect 184335 85736 190560 85738
rect 184335 85733 184401 85736
rect 148335 85352 148401 85355
rect 143904 85350 148401 85352
rect 143904 85294 148340 85350
rect 148396 85294 148401 85350
rect 143904 85292 148401 85294
rect 148335 85289 148401 85292
rect 652335 85352 652401 85355
rect 652335 85350 656736 85352
rect 652335 85294 652340 85350
rect 652396 85294 656736 85350
rect 652335 85292 656736 85294
rect 652335 85289 652401 85292
rect 184431 85204 184497 85207
rect 184431 85202 190014 85204
rect 184431 85146 184436 85202
rect 184492 85146 190014 85202
rect 184431 85144 190014 85146
rect 184431 85141 184497 85144
rect 189954 85130 190014 85144
rect 189954 85070 190560 85130
rect 640194 84464 640254 85026
rect 663234 84763 663294 85322
rect 663234 84758 663345 84763
rect 663234 84702 663284 84758
rect 663340 84702 663345 84758
rect 663234 84700 663345 84702
rect 663279 84697 663345 84700
rect 645903 84464 645969 84467
rect 640194 84462 645969 84464
rect 640194 84406 645908 84462
rect 645964 84406 645969 84462
rect 640194 84404 645969 84406
rect 645903 84401 645969 84404
rect 184527 84316 184593 84319
rect 651759 84316 651825 84319
rect 184527 84314 190560 84316
rect 184527 84258 184532 84314
rect 184588 84258 190560 84314
rect 184527 84256 190560 84258
rect 651759 84314 656736 84316
rect 651759 84258 651764 84314
rect 651820 84258 656736 84314
rect 651759 84256 656736 84258
rect 184527 84253 184593 84256
rect 651759 84253 651825 84256
rect 148527 84168 148593 84171
rect 143904 84166 148593 84168
rect 143904 84110 148532 84166
rect 148588 84110 148593 84166
rect 143904 84108 148593 84110
rect 148527 84105 148593 84108
rect 663426 84023 663486 84582
rect 663426 84018 663537 84023
rect 663426 83962 663476 84018
rect 663532 83962 663537 84018
rect 663426 83960 663537 83962
rect 663471 83957 663537 83960
rect 189954 83442 190560 83502
rect 184335 83428 184401 83431
rect 189954 83428 190014 83442
rect 184335 83426 190014 83428
rect 184335 83370 184340 83426
rect 184396 83370 190014 83426
rect 184335 83368 190014 83370
rect 652239 83428 652305 83431
rect 652239 83426 656736 83428
rect 652239 83370 652244 83426
rect 652300 83370 656736 83426
rect 652239 83368 656736 83370
rect 184335 83365 184401 83368
rect 652239 83365 652305 83368
rect 143874 82392 143934 82880
rect 184527 82836 184593 82839
rect 184527 82834 190560 82836
rect 184527 82778 184532 82834
rect 184588 82778 190560 82834
rect 184527 82776 190560 82778
rect 184527 82773 184593 82776
rect 640386 82688 640446 83176
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 647919 82688 647985 82691
rect 640386 82686 647985 82688
rect 640386 82630 647924 82686
rect 647980 82630 647985 82686
rect 640386 82628 647985 82630
rect 647919 82625 647985 82628
rect 652431 82688 652497 82691
rect 652431 82686 656736 82688
rect 652431 82630 652436 82686
rect 652492 82630 656736 82686
rect 652431 82628 656736 82630
rect 652431 82625 652497 82628
rect 149583 82392 149649 82395
rect 143874 82390 149649 82392
rect 143874 82334 149588 82390
rect 149644 82334 149649 82390
rect 143874 82332 149649 82334
rect 149583 82329 149649 82332
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 184431 81948 184497 81951
rect 184431 81946 190560 81948
rect 184431 81890 184436 81946
rect 184492 81890 190560 81946
rect 184431 81888 190560 81890
rect 184431 81885 184497 81888
rect 148431 81652 148497 81655
rect 143904 81650 148497 81652
rect 143904 81594 148436 81650
rect 148492 81594 148497 81650
rect 143904 81592 148497 81594
rect 148431 81589 148497 81592
rect 662415 81652 662481 81655
rect 663042 81652 663102 81770
rect 662415 81650 663102 81652
rect 662415 81594 662420 81650
rect 662476 81594 663102 81650
rect 662415 81592 663102 81594
rect 662415 81589 662481 81592
rect 184623 81356 184689 81359
rect 184623 81354 190560 81356
rect 184623 81298 184628 81354
rect 184684 81298 190560 81354
rect 184623 81296 190560 81298
rect 184623 81293 184689 81296
rect 640386 81060 640446 81326
rect 647919 81060 647985 81063
rect 640386 81058 647985 81060
rect 640386 81002 647924 81058
rect 647980 81002 647985 81058
rect 640386 81000 647985 81002
rect 647919 80997 647985 81000
rect 148719 80468 148785 80471
rect 143904 80466 148785 80468
rect 143904 80410 148724 80466
rect 148780 80410 148785 80466
rect 143904 80408 148785 80410
rect 148719 80405 148785 80408
rect 184335 80468 184401 80471
rect 184335 80466 190560 80468
rect 184335 80410 184340 80466
rect 184396 80410 190560 80466
rect 184335 80408 190560 80410
rect 184335 80405 184401 80408
rect 184431 79876 184497 79879
rect 184431 79874 190014 79876
rect 184431 79818 184436 79874
rect 184492 79818 190014 79874
rect 184431 79816 190014 79818
rect 184431 79813 184497 79816
rect 189954 79802 190014 79816
rect 189954 79742 190560 79802
rect 645519 79432 645585 79435
rect 640416 79430 645585 79432
rect 640416 79374 645524 79430
rect 645580 79374 645585 79430
rect 640416 79372 645585 79374
rect 645519 79369 645585 79372
rect 149679 79284 149745 79287
rect 143904 79282 149745 79284
rect 143904 79226 149684 79282
rect 149740 79226 149745 79282
rect 143904 79224 149745 79226
rect 149679 79221 149745 79224
rect 184623 78988 184689 78991
rect 184623 78986 190560 78988
rect 184623 78930 184628 78986
rect 184684 78930 190560 78986
rect 184623 78928 190560 78930
rect 184623 78925 184689 78928
rect 184527 78248 184593 78251
rect 184527 78246 190014 78248
rect 184527 78190 184532 78246
rect 184588 78190 190014 78246
rect 184527 78188 190014 78190
rect 184527 78185 184593 78188
rect 189954 78174 190014 78188
rect 189954 78114 190560 78174
rect 148623 77952 148689 77955
rect 143904 77950 148689 77952
rect 143904 77894 148628 77950
rect 148684 77894 148689 77950
rect 143904 77892 148689 77894
rect 148623 77889 148689 77892
rect 184431 77508 184497 77511
rect 647919 77508 647985 77511
rect 184431 77506 190560 77508
rect 184431 77450 184436 77506
rect 184492 77450 190560 77506
rect 184431 77448 190560 77450
rect 640416 77506 647985 77508
rect 640416 77450 647924 77506
rect 647980 77450 647985 77506
rect 640416 77448 647985 77450
rect 184431 77445 184497 77448
rect 647919 77445 647985 77448
rect 149103 76768 149169 76771
rect 143904 76766 149169 76768
rect 143904 76710 149108 76766
rect 149164 76710 149169 76766
rect 143904 76708 149169 76710
rect 149103 76705 149169 76708
rect 184527 76768 184593 76771
rect 184527 76766 190014 76768
rect 184527 76710 184532 76766
rect 184588 76710 190014 76766
rect 184527 76708 190014 76710
rect 184527 76705 184593 76708
rect 189954 76694 190014 76708
rect 189954 76634 190560 76694
rect 184335 76028 184401 76031
rect 184335 76026 190560 76028
rect 184335 75970 184340 76026
rect 184396 75970 190560 76026
rect 184335 75968 190560 75970
rect 184335 75965 184401 75968
rect 149391 75584 149457 75587
rect 645999 75584 646065 75587
rect 143904 75582 149457 75584
rect 143904 75526 149396 75582
rect 149452 75526 149457 75582
rect 143904 75524 149457 75526
rect 640416 75582 646065 75584
rect 640416 75526 646004 75582
rect 646060 75526 646065 75582
rect 640416 75524 646065 75526
rect 149391 75521 149457 75524
rect 645999 75521 646065 75524
rect 184623 75140 184689 75143
rect 184623 75138 190560 75140
rect 184623 75082 184628 75138
rect 184684 75082 190560 75138
rect 184623 75080 190560 75082
rect 184623 75077 184689 75080
rect 184335 74400 184401 74403
rect 184335 74398 190560 74400
rect 184335 74342 184340 74398
rect 184396 74342 190560 74398
rect 184335 74340 190560 74342
rect 184335 74337 184401 74340
rect 143874 73808 143934 74296
rect 149583 73808 149649 73811
rect 143874 73806 149649 73808
rect 143874 73750 149588 73806
rect 149644 73750 149649 73806
rect 143874 73748 149649 73750
rect 149583 73745 149649 73748
rect 184431 73660 184497 73663
rect 647919 73660 647985 73663
rect 184431 73658 190560 73660
rect 184431 73602 184436 73658
rect 184492 73602 190560 73658
rect 184431 73600 190560 73602
rect 640416 73658 647985 73660
rect 640416 73602 647924 73658
rect 647980 73602 647985 73658
rect 640416 73600 647985 73602
rect 184431 73597 184497 73600
rect 647919 73597 647985 73600
rect 149007 73068 149073 73071
rect 143904 73066 149073 73068
rect 143904 73010 149012 73066
rect 149068 73010 149073 73066
rect 143904 73008 149073 73010
rect 149007 73005 149073 73008
rect 184527 72920 184593 72923
rect 184527 72918 190560 72920
rect 184527 72862 184532 72918
rect 184588 72862 190560 72918
rect 184527 72860 190560 72862
rect 184527 72857 184593 72860
rect 184623 72180 184689 72183
rect 184623 72178 190560 72180
rect 184623 72122 184628 72178
rect 184684 72122 190560 72178
rect 184623 72120 190560 72122
rect 184623 72117 184689 72120
rect 149199 72032 149265 72035
rect 143904 72030 149265 72032
rect 143904 71974 149204 72030
rect 149260 71974 149265 72030
rect 143904 71972 149265 71974
rect 149199 71969 149265 71972
rect 647151 71884 647217 71887
rect 640386 71882 647217 71884
rect 640386 71826 647156 71882
rect 647212 71826 647217 71882
rect 640386 71824 647217 71826
rect 640386 71706 640446 71824
rect 647151 71821 647217 71824
rect 184335 71440 184401 71443
rect 184335 71438 190014 71440
rect 184335 71382 184340 71438
rect 184396 71382 190014 71438
rect 184335 71380 190014 71382
rect 184335 71377 184401 71380
rect 189954 71366 190014 71380
rect 189954 71306 190560 71366
rect 149391 70848 149457 70851
rect 143904 70846 149457 70848
rect 143904 70790 149396 70846
rect 149452 70790 149457 70846
rect 143904 70788 149457 70790
rect 149391 70785 149457 70788
rect 184431 70552 184497 70555
rect 184431 70550 190560 70552
rect 184431 70494 184436 70550
rect 184492 70494 190560 70550
rect 184431 70492 190560 70494
rect 184431 70489 184497 70492
rect 184527 69960 184593 69963
rect 184527 69958 190014 69960
rect 184527 69902 184532 69958
rect 184588 69902 190014 69958
rect 184527 69900 190014 69902
rect 184527 69897 184593 69900
rect 189954 69886 190014 69900
rect 189954 69826 190560 69886
rect 640386 69664 640446 69856
rect 647919 69664 647985 69667
rect 640386 69662 647985 69664
rect 640386 69606 647924 69662
rect 647980 69606 647985 69662
rect 640386 69604 647985 69606
rect 647919 69601 647985 69604
rect 149295 69516 149361 69519
rect 143904 69514 149361 69516
rect 143904 69458 149300 69514
rect 149356 69458 149361 69514
rect 143904 69456 149361 69458
rect 149295 69453 149361 69456
rect 184335 69072 184401 69075
rect 184335 69070 190560 69072
rect 184335 69014 184340 69070
rect 184396 69014 190560 69070
rect 184335 69012 190560 69014
rect 184335 69009 184401 69012
rect 646863 68628 646929 68631
rect 640194 68626 646929 68628
rect 640194 68570 646868 68626
rect 646924 68570 646929 68626
rect 640194 68568 646929 68570
rect 184335 68480 184401 68483
rect 184335 68478 190014 68480
rect 184335 68422 184340 68478
rect 184396 68422 190014 68478
rect 184335 68420 190014 68422
rect 184335 68417 184401 68420
rect 189954 68406 190014 68420
rect 189954 68346 190560 68406
rect 149583 68332 149649 68335
rect 143904 68330 149649 68332
rect 143904 68274 149588 68330
rect 149644 68274 149649 68330
rect 143904 68272 149649 68274
rect 149583 68269 149649 68272
rect 640194 68006 640254 68568
rect 646863 68565 646929 68568
rect 184527 67592 184593 67595
rect 184527 67590 190560 67592
rect 184527 67534 184532 67590
rect 184588 67534 190560 67590
rect 184527 67532 190560 67534
rect 184527 67529 184593 67532
rect 149487 67148 149553 67151
rect 143904 67146 149553 67148
rect 143904 67090 149492 67146
rect 149548 67090 149553 67146
rect 143904 67088 149553 67090
rect 149487 67085 149553 67088
rect 184431 66852 184497 66855
rect 184431 66850 190560 66852
rect 184431 66794 184436 66850
rect 184492 66794 190560 66850
rect 184431 66792 190560 66794
rect 184431 66789 184497 66792
rect 645999 66260 646065 66263
rect 640194 66258 646065 66260
rect 640194 66202 646004 66258
rect 646060 66202 646065 66258
rect 640194 66200 646065 66202
rect 184335 66112 184401 66115
rect 184335 66110 190560 66112
rect 184335 66054 184340 66110
rect 184396 66054 190560 66110
rect 640194 66082 640254 66200
rect 645999 66197 646065 66200
rect 184335 66052 190560 66054
rect 184335 66049 184401 66052
rect 143874 65372 143934 65860
rect 149679 65372 149745 65375
rect 143874 65370 149745 65372
rect 143874 65314 149684 65370
rect 149740 65314 149745 65370
rect 143874 65312 149745 65314
rect 149679 65309 149745 65312
rect 184527 65224 184593 65227
rect 184527 65222 190560 65224
rect 184527 65166 184532 65222
rect 184588 65166 190560 65222
rect 184527 65164 190560 65166
rect 184527 65161 184593 65164
rect 149391 64632 149457 64635
rect 143904 64630 149457 64632
rect 143904 64574 149396 64630
rect 149452 64574 149457 64630
rect 143904 64572 149457 64574
rect 149391 64569 149457 64572
rect 184623 64632 184689 64635
rect 184623 64630 190014 64632
rect 184623 64574 184628 64630
rect 184684 64574 190014 64630
rect 184623 64572 190014 64574
rect 184623 64569 184689 64572
rect 189954 64558 190014 64572
rect 189954 64498 190560 64558
rect 647919 64188 647985 64191
rect 640416 64186 647985 64188
rect 640416 64130 647924 64186
rect 647980 64130 647985 64186
rect 640416 64128 647985 64130
rect 647919 64125 647985 64128
rect 184431 63744 184497 63747
rect 184431 63742 190560 63744
rect 184431 63686 184436 63742
rect 184492 63686 190560 63742
rect 184431 63684 190560 63686
rect 184431 63681 184497 63684
rect 149295 63448 149361 63451
rect 143904 63446 149361 63448
rect 143904 63390 149300 63446
rect 149356 63390 149361 63446
rect 143904 63388 149361 63390
rect 149295 63385 149361 63388
rect 184335 63152 184401 63155
rect 184335 63150 190014 63152
rect 184335 63094 184340 63150
rect 184396 63094 190014 63150
rect 184335 63092 190014 63094
rect 184335 63089 184401 63092
rect 189954 63078 190014 63092
rect 189954 63018 190560 63078
rect 149391 62264 149457 62267
rect 143904 62262 149457 62264
rect 143904 62206 149396 62262
rect 149452 62206 149457 62262
rect 143904 62204 149457 62206
rect 149391 62201 149457 62204
rect 184431 62264 184497 62267
rect 647919 62264 647985 62267
rect 184431 62262 190560 62264
rect 184431 62206 184436 62262
rect 184492 62206 190560 62262
rect 184431 62204 190560 62206
rect 640416 62262 647985 62264
rect 640416 62206 647924 62262
rect 647980 62206 647985 62262
rect 640416 62204 647985 62206
rect 184431 62201 184497 62204
rect 647919 62201 647985 62204
rect 184623 61524 184689 61527
rect 184623 61522 190014 61524
rect 184623 61466 184628 61522
rect 184684 61466 190014 61522
rect 184623 61464 190014 61466
rect 184623 61461 184689 61464
rect 189954 61450 190014 61464
rect 189954 61390 190560 61450
rect 143874 60636 143934 60976
rect 184527 60784 184593 60787
rect 184527 60782 190560 60784
rect 184527 60726 184532 60782
rect 184588 60726 190560 60782
rect 184527 60724 190560 60726
rect 184527 60721 184593 60724
rect 149487 60636 149553 60639
rect 143874 60634 149553 60636
rect 143874 60578 149492 60634
rect 149548 60578 149553 60634
rect 143874 60576 149553 60578
rect 149487 60573 149553 60576
rect 647055 60340 647121 60343
rect 640416 60338 647121 60340
rect 640416 60282 647060 60338
rect 647116 60282 647121 60338
rect 640416 60280 647121 60282
rect 647055 60277 647121 60280
rect 184335 60044 184401 60047
rect 184335 60042 190014 60044
rect 184335 59986 184340 60042
rect 184396 59986 190014 60042
rect 184335 59984 190014 59986
rect 184335 59981 184401 59984
rect 189954 59970 190014 59984
rect 189954 59910 190560 59970
rect 149391 59748 149457 59751
rect 143904 59746 149457 59748
rect 143904 59690 149396 59746
rect 149452 59690 149457 59746
rect 143904 59688 149457 59690
rect 149391 59685 149457 59688
rect 184431 59304 184497 59307
rect 184431 59302 190560 59304
rect 184431 59246 184436 59302
rect 184492 59246 190560 59302
rect 184431 59244 190560 59246
rect 184431 59241 184497 59244
rect 645999 59008 646065 59011
rect 640386 59006 646065 59008
rect 640386 58950 646004 59006
rect 646060 58950 646065 59006
rect 640386 58948 646065 58950
rect 149391 58564 149457 58567
rect 143904 58562 149457 58564
rect 143904 58506 149396 58562
rect 149452 58506 149457 58562
rect 143904 58504 149457 58506
rect 149391 58501 149457 58504
rect 184527 58416 184593 58419
rect 184527 58414 190560 58416
rect 184527 58358 184532 58414
rect 184588 58358 190560 58414
rect 640386 58386 640446 58948
rect 645999 58945 646065 58948
rect 184527 58356 190560 58358
rect 184527 58353 184593 58356
rect 184335 57676 184401 57679
rect 184335 57674 190560 57676
rect 184335 57618 184340 57674
rect 184396 57618 190560 57674
rect 184335 57616 190560 57618
rect 184335 57613 184401 57616
rect 149487 57380 149553 57383
rect 143904 57378 149553 57380
rect 143904 57322 149492 57378
rect 149548 57322 149553 57378
rect 143904 57320 149553 57322
rect 149487 57317 149553 57320
rect 646767 57084 646833 57087
rect 640386 57082 646833 57084
rect 640386 57026 646772 57082
rect 646828 57026 646833 57082
rect 640386 57024 646833 57026
rect 184335 56936 184401 56939
rect 184335 56934 190560 56936
rect 184335 56878 184340 56934
rect 184396 56878 190560 56934
rect 184335 56876 190560 56878
rect 184335 56873 184401 56876
rect 640386 56536 640446 57024
rect 646767 57021 646833 57024
rect 149391 56196 149457 56199
rect 143874 56194 149457 56196
rect 143874 56138 149396 56194
rect 149452 56138 149457 56194
rect 143874 56136 149457 56138
rect 143874 56092 143934 56136
rect 149391 56133 149457 56136
rect 184335 56196 184401 56199
rect 184335 56194 190560 56196
rect 184335 56138 184340 56194
rect 184396 56138 190560 56194
rect 184335 56136 190560 56138
rect 184335 56133 184401 56136
rect 184431 55456 184497 55459
rect 184431 55454 190560 55456
rect 184431 55398 184436 55454
rect 184492 55398 190560 55454
rect 184431 55396 190560 55398
rect 184431 55393 184497 55396
rect 149679 54864 149745 54867
rect 143904 54862 149745 54864
rect 143904 54806 149684 54862
rect 149740 54806 149745 54862
rect 143904 54804 149745 54806
rect 149679 54801 149745 54804
rect 184335 54716 184401 54719
rect 646479 54716 646545 54719
rect 184335 54714 190014 54716
rect 184335 54658 184340 54714
rect 184396 54658 190014 54714
rect 184335 54656 190014 54658
rect 184335 54653 184401 54656
rect 189954 54642 190014 54656
rect 640386 54714 646545 54716
rect 640386 54658 646484 54714
rect 646540 54658 646545 54714
rect 640386 54656 646545 54658
rect 189954 54582 190560 54642
rect 640386 54612 640446 54656
rect 646479 54653 646545 54656
rect 184335 53976 184401 53979
rect 184335 53974 190560 53976
rect 184335 53918 184340 53974
rect 184396 53918 190560 53974
rect 184335 53916 190560 53918
rect 184335 53913 184401 53916
rect 149391 53828 149457 53831
rect 143904 53826 149457 53828
rect 143904 53770 149396 53826
rect 149452 53770 149457 53826
rect 143904 53768 149457 53770
rect 149391 53765 149457 53768
rect 419727 47612 419793 47615
rect 492975 47612 493041 47615
rect 419727 47610 493041 47612
rect 419727 47554 419732 47610
rect 419788 47554 492980 47610
rect 493036 47554 493041 47610
rect 419727 47552 493041 47554
rect 419727 47549 419793 47552
rect 492975 47549 493041 47552
rect 406767 47464 406833 47467
rect 357830 47462 406833 47464
rect 357830 47406 406772 47462
rect 406828 47406 406833 47462
rect 357830 47404 406833 47406
rect 357830 42139 357890 47404
rect 406767 47401 406833 47404
rect 474447 47464 474513 47467
rect 562479 47464 562545 47467
rect 474447 47462 562545 47464
rect 474447 47406 474452 47462
rect 474508 47406 562484 47462
rect 562540 47406 562545 47462
rect 474447 47404 562545 47406
rect 474447 47401 474513 47404
rect 562479 47401 562545 47404
rect 357711 42136 357890 42139
rect 357668 42134 357890 42136
rect 357668 42078 357716 42134
rect 357772 42078 357890 42134
rect 357668 42076 357890 42078
rect 357711 42074 357890 42076
rect 357711 42073 357777 42074
rect 415503 41988 415569 41991
rect 434895 41988 434961 41991
rect 415503 41986 434961 41988
rect 415503 41930 415508 41986
rect 415564 41930 434900 41986
rect 434956 41930 434961 41986
rect 415503 41928 434961 41930
rect 415503 41925 415569 41928
rect 434895 41925 434961 41928
rect 187599 41840 187665 41843
rect 194319 41840 194385 41843
rect 302895 41840 302961 41843
rect 307215 41840 307281 41843
rect 416847 41840 416913 41843
rect 470319 41840 470385 41843
rect 518703 41842 518769 41843
rect 187599 41838 190170 41840
rect 187599 41782 187604 41838
rect 187660 41782 190170 41838
rect 187599 41780 190170 41782
rect 187599 41777 187665 41780
rect 190110 40406 190170 41780
rect 194319 41838 195014 41840
rect 194319 41782 194324 41838
rect 194380 41782 195014 41838
rect 194319 41780 195014 41782
rect 194319 41777 194385 41780
rect 194954 40568 195014 41780
rect 302895 41838 305114 41840
rect 302895 41782 302900 41838
rect 302956 41782 305114 41838
rect 302895 41780 305114 41782
rect 302895 41777 302961 41780
rect 305054 40804 305114 41780
rect 307215 41838 308090 41840
rect 307215 41782 307220 41838
rect 307276 41782 308090 41838
rect 307215 41780 308090 41782
rect 307215 41777 307281 41780
rect 308026 40956 308090 41780
rect 416847 41838 417627 41840
rect 416847 41782 416852 41838
rect 416908 41782 417627 41838
rect 416847 41780 417627 41782
rect 416847 41777 416913 41780
rect 337455 40956 337521 40959
rect 308026 40954 337521 40956
rect 308026 40898 337460 40954
rect 337516 40898 337521 40954
rect 308026 40896 337521 40898
rect 337455 40893 337521 40896
rect 331215 40804 331281 40807
rect 305054 40802 331281 40804
rect 305054 40746 331220 40802
rect 331276 40746 331281 40802
rect 305054 40744 331281 40746
rect 331215 40741 331281 40744
rect 417567 40656 417627 41780
rect 470319 41838 478110 41840
rect 470319 41782 470324 41838
rect 470380 41782 478110 41838
rect 470319 41780 478110 41782
rect 470319 41777 470385 41780
rect 420687 40656 420753 40659
rect 417567 40654 420753 40656
rect 417567 40598 420692 40654
rect 420748 40598 420753 40654
rect 417567 40596 420753 40598
rect 478050 40656 478110 41780
rect 518662 41838 518769 41842
rect 520335 41840 520401 41843
rect 518662 41782 518708 41838
rect 518764 41782 518769 41838
rect 518662 41777 518769 41782
rect 519077 41838 520401 41840
rect 519077 41782 520340 41838
rect 520396 41782 520401 41838
rect 519077 41780 520401 41782
rect 493935 40804 494001 40807
rect 518662 40804 518726 41777
rect 518842 41178 518848 41242
rect 518912 41240 518918 41242
rect 519077 41240 519137 41780
rect 520335 41777 520401 41780
rect 518912 41180 519137 41240
rect 518912 41178 518918 41180
rect 493935 40802 518726 40804
rect 493935 40746 493940 40802
rect 493996 40746 518726 40802
rect 493935 40744 518726 40746
rect 493935 40741 494001 40744
rect 545199 40656 545265 40659
rect 478050 40654 545265 40656
rect 478050 40598 545204 40654
rect 545260 40598 545265 40654
rect 478050 40596 545265 40598
rect 420687 40593 420753 40596
rect 545199 40593 545265 40596
rect 194954 40508 240629 40568
rect 584556 40510 584620 40516
rect 568545 40508 568551 40510
rect 216399 40406 216465 40409
rect 190110 40404 216465 40406
rect 190110 40348 216404 40404
rect 216460 40348 216465 40404
rect 190110 40346 216465 40348
rect 216399 40343 216465 40346
rect 240569 40254 240629 40508
rect 257342 40448 568551 40508
rect 257342 40254 257402 40448
rect 568545 40446 568551 40448
rect 568615 40446 568621 40510
rect 633615 40508 633681 40511
rect 584620 40506 633681 40508
rect 584620 40450 633620 40506
rect 633676 40450 633681 40506
rect 584620 40448 633681 40450
rect 584556 40440 584620 40446
rect 633615 40445 633681 40448
rect 240567 40248 240631 40254
rect 142287 40212 142353 40215
rect 142287 40210 142398 40212
rect 142287 40154 142292 40210
rect 142348 40154 142398 40210
rect 240567 40178 240631 40184
rect 257340 40248 257404 40254
rect 257340 40178 257404 40184
rect 506799 40212 506865 40215
rect 507130 40212 507136 40214
rect 506799 40210 507136 40212
rect 142287 40149 142398 40154
rect 506799 40154 506804 40210
rect 506860 40154 507136 40210
rect 506799 40152 507136 40154
rect 506799 40149 506865 40152
rect 507130 40150 507136 40152
rect 507200 40150 507206 40214
rect 142338 40064 142398 40149
rect 141753 40004 142398 40064
rect 141753 39886 141813 40004
<< via3 >>
rect 42112 968762 42176 968766
rect 42112 968706 42164 968762
rect 42164 968706 42176 968762
rect 42112 968702 42176 968706
rect 41728 967134 41792 967138
rect 41728 967078 41780 967134
rect 41780 967078 41792 967134
rect 41728 967074 41792 967078
rect 674368 966186 674432 966250
rect 674176 965742 674240 965806
rect 40576 965002 40640 965066
rect 674560 965002 674624 965066
rect 40768 963966 40832 964030
rect 40960 963374 41024 963438
rect 674752 963374 674816 963438
rect 41152 962782 41216 962846
rect 674944 962634 675008 962698
rect 41536 962190 41600 962254
rect 675712 962250 675776 962254
rect 675712 962194 675764 962250
rect 675764 962194 675776 962250
rect 675712 962190 675776 962194
rect 41344 959526 41408 959590
rect 40384 959082 40448 959146
rect 675136 959082 675200 959146
rect 676864 958342 676928 958406
rect 41920 957810 41984 957814
rect 41920 957754 41932 957810
rect 41932 957754 41984 957810
rect 41920 957750 41984 957754
rect 675328 957662 675392 957666
rect 675328 957606 675380 957662
rect 675380 957606 675392 957662
rect 675328 957602 675392 957606
rect 42304 957514 42368 957518
rect 42304 957458 42316 957514
rect 42316 957458 42368 957514
rect 42304 957454 42368 957458
rect 42496 956270 42560 956334
rect 675520 956034 675584 956038
rect 675520 955978 675572 956034
rect 675572 955978 675584 956034
rect 675520 955974 675584 955978
rect 677056 955974 677120 956038
rect 673984 953902 674048 953966
rect 677056 953310 677120 953374
rect 675904 951978 675968 952042
rect 42496 940434 42560 940498
rect 41728 939842 41792 939906
rect 41920 938880 41984 938944
rect 41536 938658 41600 938722
rect 42112 937770 42176 937834
rect 42304 936882 42368 936946
rect 674560 936734 674624 936798
rect 40384 936586 40448 936650
rect 673984 936586 674048 936650
rect 40576 935698 40640 935762
rect 40960 935698 41024 935762
rect 674368 935698 674432 935762
rect 674752 935254 674816 935318
rect 41344 935106 41408 935170
rect 675136 934662 675200 934726
rect 40768 934218 40832 934282
rect 41152 934218 41216 934282
rect 675904 934218 675968 934282
rect 674176 933774 674240 933838
rect 674944 933182 675008 933246
rect 675712 932664 675776 932728
rect 675520 932294 675584 932358
rect 675328 931702 675392 931766
rect 677056 931554 677120 931618
rect 676864 930962 676928 931026
rect 677248 930518 677312 930582
rect 673984 876350 674048 876414
rect 674176 876202 674240 876266
rect 674368 873982 674432 874046
rect 674560 869838 674624 869902
rect 675712 864718 675776 864722
rect 675712 864662 675764 864718
rect 675764 864662 675776 864718
rect 675712 864658 675776 864662
rect 674944 862882 675008 862946
rect 40768 816262 40832 816326
rect 41152 815226 41216 815290
rect 42112 814930 42176 814994
rect 41536 802054 41600 802118
rect 41344 801758 41408 801822
rect 41920 800546 41984 800610
rect 41728 800338 41792 800342
rect 41728 800282 41780 800338
rect 41780 800282 41792 800338
rect 41728 800278 41792 800282
rect 42304 800278 42368 800342
rect 42304 797466 42368 797530
rect 41728 796342 41792 796346
rect 41728 796286 41780 796342
rect 41780 796286 41792 796342
rect 41728 796282 41792 796286
rect 41920 794270 41984 794274
rect 41920 794214 41932 794270
rect 41932 794214 41984 794270
rect 41920 794210 41984 794214
rect 41344 790510 41408 790574
rect 41536 789178 41600 789242
rect 675328 787906 675392 787910
rect 675328 787850 675380 787906
rect 675380 787850 675392 787906
rect 675328 787846 675392 787850
rect 675136 786662 675200 786726
rect 675520 784798 675584 784802
rect 675520 784742 675532 784798
rect 675532 784742 675584 784798
rect 675520 784738 675584 784742
rect 676288 780594 676352 780658
rect 676864 779114 676928 779178
rect 677056 777486 677120 777550
rect 677056 777338 677120 777402
rect 675904 775414 675968 775478
rect 677056 774822 677120 774886
rect 674752 773638 674816 773702
rect 40768 773046 40832 773110
rect 40960 773046 41024 773110
rect 40576 772010 40640 772074
rect 41152 772010 41216 772074
rect 674176 758394 674240 758458
rect 40384 758186 40448 758250
rect 40960 758038 41024 758102
rect 675712 757802 675776 757866
rect 673984 757210 674048 757274
rect 42880 757122 42944 757126
rect 42880 757066 42932 757122
rect 42932 757066 42944 757122
rect 42880 757062 42944 757066
rect 674368 757062 674432 757126
rect 42496 756470 42560 756534
rect 674560 756322 674624 756386
rect 674944 755730 675008 755794
rect 677056 754102 677120 754166
rect 677440 753658 677504 753722
rect 42496 750994 42560 751058
rect 42880 749810 42944 749874
rect 40384 748626 40448 748690
rect 40960 748478 41024 748542
rect 674368 743150 674432 743214
rect 676096 742114 676160 742178
rect 674560 741670 674624 741734
rect 674944 740338 675008 740402
rect 675712 735514 675776 735518
rect 675712 735458 675724 735514
rect 675724 735458 675776 735514
rect 675712 735454 675776 735458
rect 677056 734418 677120 734482
rect 40768 729830 40832 729894
rect 40960 729830 41024 729894
rect 40576 728942 40640 729006
rect 40384 728794 40448 728858
rect 41728 722578 41792 722642
rect 40768 716954 40832 717018
rect 40384 716510 40448 716574
rect 43072 713994 43136 714058
rect 41920 713906 41984 713910
rect 41920 713850 41972 713906
rect 41972 713850 41984 713906
rect 41920 713846 41984 713850
rect 42880 713846 42944 713910
rect 675136 713402 675200 713466
rect 675904 712810 675968 712874
rect 675328 712218 675392 712282
rect 675520 712070 675584 712134
rect 41920 711626 41984 711690
rect 676288 711626 676352 711690
rect 674752 710738 674816 710802
rect 42880 709762 42944 709766
rect 42880 709706 42932 709762
rect 42932 709706 42944 709762
rect 42880 709702 42944 709706
rect 677248 709110 677312 709174
rect 676864 708518 676928 708582
rect 43072 707246 43136 707250
rect 43072 707190 43124 707246
rect 43124 707190 43136 707246
rect 43072 707186 43136 707190
rect 41728 706002 41792 706066
rect 40768 703634 40832 703698
rect 40384 703338 40448 703402
rect 675328 697922 675392 697926
rect 675328 697866 675380 697922
rect 675380 697866 675392 697922
rect 675328 697862 675392 697866
rect 676288 697270 676352 697334
rect 675520 696886 675584 696890
rect 675520 696830 675572 696886
rect 675572 696830 675584 696886
rect 675520 696826 675584 696830
rect 675136 694754 675200 694818
rect 676480 694162 676544 694226
rect 673984 690462 674048 690526
rect 676864 687354 676928 687418
rect 40768 686614 40832 686678
rect 40960 686614 41024 686678
rect 41152 685726 41216 685790
rect 40576 685578 40640 685642
rect 40576 672554 40640 672618
rect 40384 672406 40448 672470
rect 41728 670690 41792 670694
rect 41728 670634 41780 670690
rect 41780 670634 41792 670690
rect 41728 670630 41792 670634
rect 42496 670630 42560 670694
rect 42304 670038 42368 670102
rect 674560 668114 674624 668178
rect 674368 667078 674432 667142
rect 42304 666634 42368 666698
rect 674944 666634 675008 666698
rect 675712 666116 675776 666180
rect 42496 665154 42560 665218
rect 676096 665006 676160 665070
rect 41728 663438 41792 663442
rect 41728 663382 41780 663438
rect 41780 663382 41792 663438
rect 41728 663378 41792 663382
rect 677056 663378 677120 663442
rect 40576 660862 40640 660926
rect 40384 660270 40448 660334
rect 674944 652574 675008 652638
rect 674560 651538 674624 651602
rect 675712 649674 675776 649678
rect 675712 649618 675724 649674
rect 675724 649618 675776 649674
rect 675712 649614 675776 649618
rect 674176 645322 674240 645386
rect 40768 643398 40832 643462
rect 41152 642362 41216 642426
rect 675904 640290 675968 640354
rect 674752 638514 674816 638578
rect 41728 635776 41792 635840
rect 40384 629042 40448 629106
rect 42496 628006 42560 628070
rect 40576 627858 40640 627922
rect 41536 627918 41600 627922
rect 41536 627862 41548 627918
rect 41548 627862 41600 627918
rect 41536 627858 41600 627862
rect 42304 627710 42368 627774
rect 42880 627414 42944 627478
rect 675520 623122 675584 623186
rect 42496 622086 42560 622150
rect 675328 622086 675392 622150
rect 675136 621642 675200 621706
rect 42304 621494 42368 621558
rect 673984 621050 674048 621114
rect 41728 620962 41792 620966
rect 41728 620906 41780 620962
rect 41780 620906 41792 620962
rect 41728 620902 41792 620906
rect 676288 620310 676352 620374
rect 42880 620222 42944 620226
rect 42880 620166 42932 620222
rect 42932 620166 42944 620222
rect 42880 620162 42944 620166
rect 676480 619866 676544 619930
rect 41728 619126 41792 619190
rect 40576 618830 40640 618894
rect 676864 618830 676928 618894
rect 40384 616462 40448 616526
rect 41536 616018 41600 616082
rect 673984 607730 674048 607794
rect 41536 607582 41600 607646
rect 675136 606398 675200 606462
rect 674368 604770 674432 604834
rect 40768 600626 40832 600690
rect 41728 600478 41792 600542
rect 675328 600182 675392 600246
rect 41536 599738 41600 599802
rect 40576 599294 40640 599358
rect 676096 595298 676160 595362
rect 675520 593434 675584 593438
rect 675520 593378 675532 593434
rect 675532 593378 675584 593434
rect 675520 593374 675584 593378
rect 40384 585522 40448 585586
rect 40960 585374 41024 585438
rect 43072 584494 43136 584558
rect 42880 584198 42944 584262
rect 42880 578782 42944 578786
rect 42880 578726 42892 578782
rect 42892 578726 42944 578782
rect 42880 578722 42944 578726
rect 674560 577982 674624 578046
rect 43072 577538 43136 577602
rect 675904 577390 675968 577454
rect 674944 577242 675008 577306
rect 675712 576502 675776 576566
rect 674176 575910 674240 575974
rect 674752 575318 674816 575382
rect 40960 574430 41024 574494
rect 40384 573986 40448 574050
rect 674560 562590 674624 562654
rect 674944 561702 675008 561766
rect 674752 561406 674816 561470
rect 41728 558890 41792 558954
rect 676864 557558 676928 557622
rect 40384 557410 40448 557474
rect 40768 556670 40832 556734
rect 41728 556300 41792 556364
rect 40768 556078 40832 556142
rect 40576 555930 40640 555994
rect 40960 541574 41024 541638
rect 42496 541574 42560 541638
rect 41152 541426 41216 541490
rect 41728 541338 41792 541342
rect 41728 541282 41740 541338
rect 41740 541282 41792 541338
rect 41728 541278 41792 541282
rect 41920 541042 41984 541046
rect 41920 540986 41972 541042
rect 41972 540986 41984 541042
rect 41920 540982 41984 540986
rect 42304 540982 42368 541046
rect 42304 535654 42368 535718
rect 42496 535062 42560 535126
rect 675136 532990 675200 533054
rect 676096 532694 676160 532758
rect 673984 531806 674048 531870
rect 674368 531510 674432 531574
rect 40960 531362 41024 531426
rect 675328 530918 675392 530982
rect 41920 530682 41984 530686
rect 41920 530626 41972 530682
rect 41972 530626 41984 530682
rect 41920 530622 41984 530626
rect 675520 530326 675584 530390
rect 41728 529646 41792 529650
rect 41728 529590 41780 529646
rect 41780 529590 41792 529646
rect 41728 529586 41792 529590
rect 41152 526478 41216 526542
rect 674552 489182 674616 489246
rect 674360 487850 674424 487914
rect 674744 485926 674808 485990
rect 676864 483706 676928 483770
rect 40576 429834 40640 429898
rect 41728 429686 41792 429750
rect 40768 428502 40832 428566
rect 40768 427466 40832 427530
rect 41920 427170 41984 427234
rect 42304 426430 42368 426494
rect 40960 425986 41024 426050
rect 40384 425394 40448 425458
rect 41152 424506 41216 424570
rect 41344 423914 41408 423978
rect 41536 423470 41600 423534
rect 40576 421990 40640 422054
rect 41920 411246 41984 411250
rect 41920 411190 41972 411246
rect 41972 411190 41984 411246
rect 41920 411186 41984 411190
rect 40384 406006 40448 406070
rect 40576 403786 40640 403850
rect 41536 403046 41600 403110
rect 41344 402454 41408 402518
rect 40960 401862 41024 401926
rect 676672 400382 676736 400446
rect 674176 400234 674240 400298
rect 40768 399938 40832 400002
rect 41152 399494 41216 399558
rect 676480 399494 676544 399558
rect 674944 399198 675008 399262
rect 41920 398962 41984 398966
rect 41920 398906 41932 398962
rect 41932 398906 41984 398962
rect 41920 398902 41984 398906
rect 674368 398754 674432 398818
rect 675520 398162 675584 398226
rect 675904 397718 675968 397782
rect 675328 396830 675392 396894
rect 675136 396682 675200 396746
rect 676096 395942 676160 396006
rect 675712 395202 675776 395266
rect 676288 394610 676352 394674
rect 41128 390902 41192 390966
rect 41728 386470 41792 386534
rect 676480 385878 676544 385942
rect 675904 385582 675968 385646
rect 676672 384694 676736 384758
rect 41728 384398 41792 384462
rect 40768 384250 40832 384314
rect 41920 383954 41984 384018
rect 40960 383214 41024 383278
rect 674944 382918 675008 382982
rect 41344 382770 41408 382834
rect 675136 382770 675200 382834
rect 40384 382178 40448 382242
rect 675328 382178 675392 382242
rect 41152 381290 41216 381354
rect 675712 381202 675776 381206
rect 675712 381146 675764 381202
rect 675764 381146 675776 381202
rect 675712 381142 675776 381146
rect 41728 380994 41792 381058
rect 41536 380254 41600 380318
rect 674368 378774 674432 378838
rect 676288 377886 676352 377950
rect 676096 375666 676160 375730
rect 674176 373742 674240 373806
rect 675520 372026 675584 372030
rect 675520 371970 675572 372026
rect 675572 371970 675584 372026
rect 675520 371966 675584 371970
rect 41920 368178 41984 368182
rect 41920 368122 41972 368178
rect 41972 368122 41984 368178
rect 41920 368118 41984 368122
rect 40384 362790 40448 362854
rect 41536 359830 41600 359894
rect 41728 359446 41792 359450
rect 41728 359390 41780 359446
rect 41780 359390 41792 359446
rect 41728 359386 41792 359390
rect 41344 358646 41408 358710
rect 673984 358054 674048 358118
rect 674176 357018 674240 357082
rect 40768 356870 40832 356934
rect 41152 356426 41216 356490
rect 676096 356130 676160 356194
rect 40960 355538 41024 355602
rect 675904 355538 675968 355602
rect 674560 354946 674624 355010
rect 674944 353466 675008 353530
rect 674752 353022 674816 353086
rect 675520 351986 675584 352050
rect 675712 351468 675776 351532
rect 675136 351098 675200 351162
rect 40576 342662 40640 342726
rect 40768 341034 40832 341098
rect 41728 340812 41792 340876
rect 40576 340442 40640 340506
rect 41152 339554 41216 339618
rect 675904 339554 675968 339618
rect 40384 338962 40448 339026
rect 40960 338074 41024 338138
rect 41344 337482 41408 337546
rect 41536 337038 41600 337102
rect 675520 337098 675584 337102
rect 675520 337042 675532 337098
rect 675532 337042 675584 337098
rect 675520 337038 675584 337042
rect 675712 336506 675776 336510
rect 675712 336450 675764 336506
rect 675764 336450 675776 336506
rect 675712 336446 675776 336450
rect 674944 333486 675008 333550
rect 675136 330526 675200 330590
rect 674560 328306 674624 328370
rect 674752 326826 674816 326890
rect 41728 324962 41792 324966
rect 41728 324906 41780 324962
rect 41780 324906 41792 324962
rect 41728 324902 41792 324906
rect 40384 319722 40448 319786
rect 41536 316762 41600 316826
rect 41344 316022 41408 316086
rect 41152 315430 41216 315494
rect 40768 313654 40832 313718
rect 673984 313506 674048 313570
rect 40960 313210 41024 313274
rect 674368 312618 674432 312682
rect 674176 312470 674240 312534
rect 40576 312322 40640 312386
rect 673984 311730 674048 311794
rect 675904 311508 675968 311572
rect 674176 310990 674240 311054
rect 674560 309954 674624 310018
rect 675328 309066 675392 309130
rect 675136 308474 675200 308538
rect 674752 307734 674816 307798
rect 674944 306106 675008 306170
rect 675520 305514 675584 305578
rect 675712 304552 675776 304616
rect 40576 297818 40640 297882
rect 41728 297596 41792 297660
rect 40768 297226 40832 297290
rect 41152 296486 41216 296550
rect 41536 295746 41600 295810
rect 40960 294858 41024 294922
rect 40384 294266 40448 294330
rect 41344 293822 41408 293886
rect 675328 292846 675392 292850
rect 675328 292790 675380 292846
rect 675380 292790 675392 292846
rect 675328 292786 675392 292790
rect 675136 288494 675200 288558
rect 675712 287814 675776 287818
rect 675712 287758 675724 287814
rect 675724 287758 675776 287814
rect 675712 287754 675776 287758
rect 675520 287370 675584 287374
rect 675520 287314 675532 287370
rect 675532 287314 675584 287370
rect 675520 287310 675584 287314
rect 674944 285238 675008 285302
rect 674560 283610 674624 283674
rect 674752 281834 674816 281898
rect 41728 281746 41792 281750
rect 41728 281690 41780 281746
rect 41780 281690 41792 281746
rect 41728 281686 41792 281690
rect 42112 278578 42176 278642
rect 41536 276506 41600 276570
rect 41344 273546 41408 273610
rect 40384 272806 40448 272870
rect 41152 272362 41216 272426
rect 40576 270438 40640 270502
rect 40960 269994 41024 270058
rect 40768 269106 40832 269170
rect 674368 268514 674432 268578
rect 675520 267922 675584 267986
rect 673984 267478 674048 267542
rect 673984 267034 674048 267098
rect 674176 266442 674240 266506
rect 674176 265702 674240 265766
rect 675904 265554 675968 265618
rect 673984 264962 674048 265026
rect 674368 264962 674432 265026
rect 674560 264962 674624 265026
rect 675712 264074 675776 264138
rect 673984 263482 674048 263546
rect 674752 262742 674816 262806
rect 676288 261262 676352 261326
rect 674944 261114 675008 261178
rect 675136 260522 675200 260586
rect 676096 259782 676160 259846
rect 40576 254602 40640 254666
rect 41728 254454 41792 254518
rect 41920 253862 41984 253926
rect 40960 253270 41024 253334
rect 41536 252530 41600 252594
rect 40768 251642 40832 251706
rect 41152 251050 41216 251114
rect 41344 251050 41408 251114
rect 675904 249570 675968 249634
rect 675712 247558 675776 247562
rect 675712 247502 675724 247558
rect 675724 247502 675776 247558
rect 675712 247498 675776 247502
rect 676288 246610 676352 246674
rect 676096 245870 676160 245934
rect 148330 243354 148394 243418
rect 673984 243502 674048 243566
rect 675136 241874 675200 241938
rect 674944 240542 675008 240606
rect 41728 238382 41792 238386
rect 41728 238326 41780 238382
rect 41780 238326 41792 238382
rect 41728 238322 41792 238326
rect 674560 238174 674624 238238
rect 674752 236842 674816 236906
rect 41536 233290 41600 233354
rect 41152 230330 41216 230394
rect 41344 229738 41408 229802
rect 40960 228998 41024 229062
rect 40576 227370 40640 227434
rect 40768 226778 40832 226842
rect 41920 226246 41984 226250
rect 41920 226190 41972 226246
rect 41972 226190 41984 226246
rect 41920 226186 41984 226190
rect 675520 223374 675584 223438
rect 675904 222782 675968 222846
rect 674368 222634 674432 222698
rect 673984 221894 674048 221958
rect 674176 221302 674240 221366
rect 674176 220710 674240 220774
rect 675520 219970 675584 220034
rect 674752 219822 674816 219886
rect 674176 218934 674240 218998
rect 676288 218638 676352 218702
rect 675136 218342 675200 218406
rect 674560 217750 674624 217814
rect 676096 217010 676160 217074
rect 675712 216270 675776 216334
rect 674944 215826 675008 215890
rect 40576 211386 40640 211450
rect 40384 210942 40448 211006
rect 41728 210646 41792 210710
rect 41152 209906 41216 209970
rect 41536 209462 41600 209526
rect 40768 208426 40832 208490
rect 40960 207834 41024 207898
rect 41344 207834 41408 207898
rect 676096 205022 676160 205086
rect 675520 204342 675584 204346
rect 675520 204286 675532 204342
rect 675532 204286 675584 204342
rect 675520 204282 675584 204286
rect 676288 202654 676352 202718
rect 675712 201382 675776 201386
rect 675712 201326 675764 201382
rect 675764 201326 675776 201382
rect 675712 201322 675776 201326
rect 675136 198362 675200 198426
rect 674944 195254 675008 195318
rect 40384 195106 40448 195170
rect 674752 193478 674816 193542
rect 674560 191554 674624 191618
rect 41536 190074 41600 190138
rect 40960 187114 41024 187178
rect 41344 186670 41408 186734
rect 41152 185782 41216 185846
rect 40576 184006 40640 184070
rect 40768 183562 40832 183626
rect 41728 183030 41792 183034
rect 41728 182974 41780 183030
rect 41780 182974 41792 183030
rect 41728 182970 41792 182974
rect 675904 178382 675968 178446
rect 674368 177790 674432 177854
rect 673984 177198 674048 177262
rect 675520 176902 675584 176966
rect 674176 176310 674240 176374
rect 675520 175866 675584 175930
rect 674176 175718 674240 175782
rect 674752 174830 674816 174894
rect 674944 173350 675008 173414
rect 674560 172758 674624 172822
rect 148330 171722 148394 171786
rect 673984 170834 674048 170898
rect 675136 169946 675200 170010
rect 675328 169354 675392 169418
rect 675712 168762 675776 168826
rect 674944 153370 675008 153434
rect 148288 152778 148352 152842
rect 675328 152542 675392 152546
rect 675328 152486 675380 152542
rect 675380 152486 675392 152542
rect 675328 152482 675392 152486
rect 675136 151890 675200 151954
rect 675712 151358 675776 151362
rect 675712 151302 675724 151358
rect 675724 151302 675776 151358
rect 675712 151298 675776 151302
rect 673984 150262 674048 150326
rect 674752 148486 674816 148550
rect 674560 146562 674624 146626
rect 673368 133094 673432 133158
rect 674520 132058 674584 132122
rect 673176 131170 673240 131234
rect 674944 130134 675008 130198
rect 675712 129616 675776 129680
rect 675136 128654 675200 128718
rect 674368 128062 674432 128126
rect 675328 127618 675392 127682
rect 674560 125694 674624 125758
rect 674752 125102 674816 125166
rect 674944 114298 675008 114362
rect 675136 112226 675200 112290
rect 148288 109266 148352 109330
rect 674368 108082 674432 108146
rect 674752 106306 674816 106370
rect 674560 105122 674624 105186
rect 675712 103258 675776 103262
rect 675712 103202 675724 103258
rect 675724 103202 675776 103258
rect 675712 103198 675776 103202
rect 675328 101482 675392 101486
rect 675328 101426 675380 101482
rect 675380 101426 675392 101482
rect 675328 101422 675392 101426
rect 518848 41178 518912 41242
rect 568551 40446 568615 40510
rect 584556 40446 584620 40510
rect 240567 40184 240631 40248
rect 257340 40184 257404 40248
rect 507136 40150 507200 40214
<< metal4 >>
rect 42111 968766 42177 968767
rect 42111 968702 42112 968766
rect 42176 968702 42177 968766
rect 42111 968701 42177 968702
rect 41727 967138 41793 967139
rect 41727 967074 41728 967138
rect 41792 967074 41793 967138
rect 41727 967073 41793 967074
rect 40575 965066 40641 965067
rect 40575 965002 40576 965066
rect 40640 965002 40641 965066
rect 40575 965001 40641 965002
rect 40383 959146 40449 959147
rect 40383 959082 40384 959146
rect 40448 959082 40449 959146
rect 40383 959081 40449 959082
rect 40386 948837 40446 959081
rect 40578 949029 40638 965001
rect 40767 964030 40833 964031
rect 40767 963966 40768 964030
rect 40832 963966 40833 964030
rect 40767 963965 40833 963966
rect 40770 949221 40830 963965
rect 40959 963438 41025 963439
rect 40959 963374 40960 963438
rect 41024 963374 41025 963438
rect 40959 963373 41025 963374
rect 40962 949413 41022 963373
rect 41151 962846 41217 962847
rect 41151 962782 41152 962846
rect 41216 962782 41217 962846
rect 41151 962781 41217 962782
rect 41154 949605 41214 962781
rect 41535 962254 41601 962255
rect 41535 962190 41536 962254
rect 41600 962190 41601 962254
rect 41535 962189 41601 962190
rect 41343 959590 41409 959591
rect 41343 959526 41344 959590
rect 41408 959526 41409 959590
rect 41343 959525 41409 959526
rect 41346 949797 41406 959525
rect 41538 949989 41598 962189
rect 41730 950181 41790 967073
rect 41919 957814 41985 957815
rect 41919 957750 41920 957814
rect 41984 957750 41985 957814
rect 41919 957749 41985 957750
rect 41922 950373 41982 957749
rect 42114 950565 42174 968701
rect 674367 966250 674433 966251
rect 674367 966186 674368 966250
rect 674432 966186 674433 966250
rect 674367 966185 674433 966186
rect 674175 965806 674241 965807
rect 674175 965742 674176 965806
rect 674240 965742 674241 965806
rect 674175 965741 674241 965742
rect 42303 957518 42369 957519
rect 42303 957454 42304 957518
rect 42368 957454 42369 957518
rect 42303 957453 42369 957454
rect 42306 950757 42366 957453
rect 42495 956334 42561 956335
rect 42495 956270 42496 956334
rect 42560 956270 42561 956334
rect 42495 956269 42561 956270
rect 42498 950949 42558 956269
rect 673983 953966 674049 953967
rect 673983 953902 673984 953966
rect 674048 953902 674049 953966
rect 673983 953901 674049 953902
rect 673986 951188 674046 953901
rect 670580 951128 674046 951188
rect 42498 950889 45323 950949
rect 42306 950697 45131 950757
rect 42114 950505 44939 950565
rect 41922 950313 44747 950373
rect 41730 950121 44555 950181
rect 41538 949929 44363 949989
rect 41346 949737 44171 949797
rect 41154 949545 43979 949605
rect 40962 949353 43787 949413
rect 40770 949161 43595 949221
rect 40578 948969 43403 949029
rect 40386 948777 43211 948837
rect 43151 945534 43211 948777
rect 40386 945474 43211 945534
rect 40386 936651 40446 945474
rect 43343 945342 43403 948969
rect 40578 945282 43403 945342
rect 40383 936650 40449 936651
rect 40383 936586 40384 936650
rect 40448 936586 40449 936650
rect 40383 936585 40449 936586
rect 40578 935763 40638 945282
rect 43535 945150 43595 949161
rect 40770 945090 43595 945150
rect 40575 935762 40641 935763
rect 40575 935698 40576 935762
rect 40640 935698 40641 935762
rect 40575 935697 40641 935698
rect 40770 934283 40830 945090
rect 43727 944958 43787 949353
rect 40962 944898 43787 944958
rect 40962 935763 41022 944898
rect 43919 944766 43979 949545
rect 41154 944706 43979 944766
rect 40959 935762 41025 935763
rect 40959 935698 40960 935762
rect 41024 935698 41025 935762
rect 40959 935697 41025 935698
rect 41154 934283 41214 944706
rect 44111 944574 44171 949737
rect 41346 944514 44171 944574
rect 41346 935171 41406 944514
rect 44303 944382 44363 949929
rect 41538 944322 44363 944382
rect 41538 938723 41598 944322
rect 44495 944190 44555 950121
rect 41730 944130 44555 944190
rect 41730 939907 41790 944130
rect 44687 943998 44747 950313
rect 41922 943938 44747 943998
rect 41727 939906 41793 939907
rect 41727 939842 41728 939906
rect 41792 939842 41793 939906
rect 41727 939841 41793 939842
rect 41922 938945 41982 943938
rect 44879 943806 44939 950505
rect 42114 943746 44939 943806
rect 41919 938944 41985 938945
rect 41919 938880 41920 938944
rect 41984 938880 41985 938944
rect 41919 938879 41985 938880
rect 41535 938722 41601 938723
rect 41535 938658 41536 938722
rect 41600 938658 41601 938722
rect 41535 938657 41601 938658
rect 42114 937835 42174 943746
rect 45071 943614 45131 950697
rect 42306 943554 45131 943614
rect 42111 937834 42177 937835
rect 42111 937770 42112 937834
rect 42176 937770 42177 937834
rect 42111 937769 42177 937770
rect 42306 936947 42366 943554
rect 45263 943422 45323 950889
rect 42498 943362 45323 943422
rect 42498 940499 42558 943362
rect 42495 940498 42561 940499
rect 42495 940434 42496 940498
rect 42560 940434 42561 940498
rect 42495 940433 42561 940434
rect 670580 938452 670640 951128
rect 674178 950996 674238 965741
rect 670772 950936 674238 950996
rect 670772 938644 670832 950936
rect 674370 950804 674430 966185
rect 674559 965066 674625 965067
rect 674559 965002 674560 965066
rect 674624 965002 674625 965066
rect 674559 965001 674625 965002
rect 670964 950744 674430 950804
rect 670964 938836 671024 950744
rect 674562 950612 674622 965001
rect 674751 963438 674817 963439
rect 674751 963374 674752 963438
rect 674816 963374 674817 963438
rect 674751 963373 674817 963374
rect 671156 950552 674622 950612
rect 671156 939028 671216 950552
rect 674754 950420 674814 963373
rect 674943 962698 675009 962699
rect 674943 962634 674944 962698
rect 675008 962634 675009 962698
rect 674943 962633 675009 962634
rect 671348 950360 674814 950420
rect 671348 939220 671408 950360
rect 674946 950228 675006 962633
rect 675711 962254 675777 962255
rect 675711 962190 675712 962254
rect 675776 962190 675777 962254
rect 675711 962189 675777 962190
rect 675135 959146 675201 959147
rect 675135 959082 675136 959146
rect 675200 959082 675201 959146
rect 675135 959081 675201 959082
rect 671540 950168 675006 950228
rect 671540 939412 671600 950168
rect 675138 950036 675198 959081
rect 675327 957666 675393 957667
rect 675327 957602 675328 957666
rect 675392 957602 675393 957666
rect 675327 957601 675393 957602
rect 671732 949976 675198 950036
rect 671732 939604 671792 949976
rect 675330 949844 675390 957601
rect 675519 956038 675585 956039
rect 675519 955974 675520 956038
rect 675584 955974 675585 956038
rect 675519 955973 675585 955974
rect 671924 949784 675390 949844
rect 671924 939796 671984 949784
rect 675522 949652 675582 955973
rect 672116 949592 675582 949652
rect 672116 939988 672176 949592
rect 675714 949460 675774 962189
rect 676863 958406 676929 958407
rect 676863 958342 676864 958406
rect 676928 958342 676929 958406
rect 676863 958341 676929 958342
rect 675903 952042 675969 952043
rect 675903 951978 675904 952042
rect 675968 951978 675969 952042
rect 675903 951977 675969 951978
rect 672308 949400 675774 949460
rect 672308 940180 672368 949400
rect 675906 949268 675966 951977
rect 672500 949208 675966 949268
rect 672500 940372 672560 949208
rect 676866 948308 676926 958341
rect 677055 956038 677121 956039
rect 677055 955974 677056 956038
rect 677120 955974 677121 956038
rect 677055 955973 677121 955974
rect 677058 955407 677118 955973
rect 677058 955347 677310 955407
rect 677055 953374 677121 953375
rect 677055 953310 677056 953374
rect 677120 953310 677121 953374
rect 677055 953309 677121 953310
rect 673460 948248 676926 948308
rect 673460 941332 673520 948248
rect 677058 948116 677118 953309
rect 673652 948056 677118 948116
rect 673652 941524 673712 948056
rect 677250 947924 677310 955347
rect 673844 947864 677310 947924
rect 673844 941716 673904 947864
rect 673844 941656 677310 941716
rect 673652 941464 677118 941524
rect 673460 941272 676926 941332
rect 672500 940312 675966 940372
rect 672308 940120 675774 940180
rect 672116 939928 675582 939988
rect 671924 939736 675390 939796
rect 671732 939544 675198 939604
rect 671540 939352 675006 939412
rect 671348 939160 674814 939220
rect 671156 938968 674622 939028
rect 670964 938776 674430 938836
rect 670772 938584 674238 938644
rect 670580 938392 674046 938452
rect 42303 936946 42369 936947
rect 42303 936882 42304 936946
rect 42368 936882 42369 936946
rect 42303 936881 42369 936882
rect 673986 936651 674046 938392
rect 673983 936650 674049 936651
rect 673983 936586 673984 936650
rect 674048 936586 674049 936650
rect 673983 936585 674049 936586
rect 41343 935170 41409 935171
rect 41343 935106 41344 935170
rect 41408 935106 41409 935170
rect 41343 935105 41409 935106
rect 40767 934282 40833 934283
rect 40767 934218 40768 934282
rect 40832 934218 40833 934282
rect 40767 934217 40833 934218
rect 41151 934282 41217 934283
rect 41151 934218 41152 934282
rect 41216 934218 41217 934282
rect 41151 934217 41217 934218
rect 674178 933839 674238 938584
rect 674370 935763 674430 938776
rect 674562 936799 674622 938968
rect 674559 936798 674625 936799
rect 674559 936734 674560 936798
rect 674624 936734 674625 936798
rect 674559 936733 674625 936734
rect 674367 935762 674433 935763
rect 674367 935698 674368 935762
rect 674432 935698 674433 935762
rect 674367 935697 674433 935698
rect 674754 935319 674814 939160
rect 674751 935318 674817 935319
rect 674751 935254 674752 935318
rect 674816 935254 674817 935318
rect 674751 935253 674817 935254
rect 674175 933838 674241 933839
rect 674175 933774 674176 933838
rect 674240 933774 674241 933838
rect 674175 933773 674241 933774
rect 674946 933247 675006 939352
rect 675138 934727 675198 939544
rect 675135 934726 675201 934727
rect 675135 934662 675136 934726
rect 675200 934662 675201 934726
rect 675135 934661 675201 934662
rect 674943 933246 675009 933247
rect 674943 933182 674944 933246
rect 675008 933182 675009 933246
rect 674943 933181 675009 933182
rect 675330 931767 675390 939736
rect 675522 932359 675582 939928
rect 675714 932729 675774 940120
rect 675906 934283 675966 940312
rect 675903 934282 675969 934283
rect 675903 934218 675904 934282
rect 675968 934218 675969 934282
rect 675903 934217 675969 934218
rect 675711 932728 675777 932729
rect 675711 932664 675712 932728
rect 675776 932664 675777 932728
rect 675711 932663 675777 932664
rect 675519 932358 675585 932359
rect 675519 932294 675520 932358
rect 675584 932294 675585 932358
rect 675519 932293 675585 932294
rect 675327 931766 675393 931767
rect 675327 931702 675328 931766
rect 675392 931702 675393 931766
rect 675327 931701 675393 931702
rect 676866 931027 676926 941272
rect 677058 931619 677118 941464
rect 677055 931618 677121 931619
rect 677055 931554 677056 931618
rect 677120 931554 677121 931618
rect 677055 931553 677121 931554
rect 676863 931026 676929 931027
rect 676863 930962 676864 931026
rect 676928 930962 676929 931026
rect 676863 930961 676929 930962
rect 677250 930583 677310 941656
rect 677247 930582 677313 930583
rect 677247 930518 677248 930582
rect 677312 930518 677313 930582
rect 677247 930517 677313 930518
rect 673983 876414 674049 876415
rect 673983 876350 673984 876414
rect 674048 876350 674049 876414
rect 673983 876349 674049 876350
rect 40767 816326 40833 816327
rect 40767 816262 40768 816326
rect 40832 816262 40833 816326
rect 40767 816261 40833 816262
rect 40770 812190 40830 816261
rect 41151 815290 41217 815291
rect 41151 815226 41152 815290
rect 41216 815226 41217 815290
rect 41151 815225 41217 815226
rect 40770 812130 41022 812190
rect 40962 779088 41022 812130
rect 39932 779028 41022 779088
rect 39932 776137 39992 779028
rect 39932 776077 41022 776137
rect 40962 773111 41022 776077
rect 40767 773110 40833 773111
rect 40767 773046 40768 773110
rect 40832 773046 40833 773110
rect 40767 773045 40833 773046
rect 40959 773110 41025 773111
rect 40959 773046 40960 773110
rect 41024 773046 41025 773110
rect 40959 773045 41025 773046
rect 40575 772074 40641 772075
rect 40575 772010 40576 772074
rect 40640 772010 40641 772074
rect 40575 772009 40641 772010
rect 40383 758250 40449 758251
rect 40383 758186 40384 758250
rect 40448 758186 40449 758250
rect 40383 758185 40449 758186
rect 40386 748691 40446 758185
rect 40383 748690 40449 748691
rect 40383 748626 40384 748690
rect 40448 748626 40449 748690
rect 40383 748625 40449 748626
rect 40578 735908 40638 772009
rect 39974 735848 40638 735908
rect 40770 735854 40830 773045
rect 41154 772075 41214 815225
rect 42111 814994 42177 814995
rect 42111 814930 42112 814994
rect 42176 814930 42177 814994
rect 42111 814929 42177 814930
rect 41535 802118 41601 802119
rect 41535 802054 41536 802118
rect 41600 802054 41601 802118
rect 41535 802053 41601 802054
rect 41343 801822 41409 801823
rect 41343 801758 41344 801822
rect 41408 801758 41409 801822
rect 41343 801757 41409 801758
rect 41346 790575 41406 801757
rect 41343 790574 41409 790575
rect 41343 790510 41344 790574
rect 41408 790510 41409 790574
rect 41343 790509 41409 790510
rect 41538 789243 41598 802053
rect 41919 800610 41985 800611
rect 41919 800546 41920 800610
rect 41984 800546 41985 800610
rect 41919 800545 41985 800546
rect 41727 800342 41793 800343
rect 41727 800278 41728 800342
rect 41792 800278 41793 800342
rect 41727 800277 41793 800278
rect 41730 796347 41790 800277
rect 41727 796346 41793 796347
rect 41727 796282 41728 796346
rect 41792 796282 41793 796346
rect 41727 796281 41793 796282
rect 41922 794275 41982 800545
rect 41919 794274 41985 794275
rect 41919 794210 41920 794274
rect 41984 794210 41985 794274
rect 41919 794209 41985 794210
rect 41535 789242 41601 789243
rect 41535 789178 41536 789242
rect 41600 789178 41601 789242
rect 41535 789177 41601 789178
rect 42114 779238 42174 814929
rect 42303 800342 42369 800343
rect 42303 800278 42304 800342
rect 42368 800278 42369 800342
rect 42303 800277 42369 800278
rect 42306 797531 42366 800277
rect 42303 797530 42369 797531
rect 42303 797466 42304 797530
rect 42368 797466 42369 797530
rect 42303 797465 42369 797466
rect 42114 779178 42431 779238
rect 42371 776091 42431 779178
rect 42114 776031 42431 776091
rect 41151 772074 41217 772075
rect 41151 772010 41152 772074
rect 41216 772010 41217 772074
rect 41151 772009 41217 772010
rect 40959 758102 41025 758103
rect 40959 758038 40960 758102
rect 41024 758038 41025 758102
rect 40959 758037 41025 758038
rect 40962 748543 41022 758037
rect 40959 748542 41025 748543
rect 40959 748478 40960 748542
rect 41024 748478 41025 748542
rect 40959 748477 41025 748478
rect 42114 735876 42174 776031
rect 673986 772948 674046 876349
rect 674175 876266 674241 876267
rect 674175 876202 674176 876266
rect 674240 876202 674241 876266
rect 674175 876201 674241 876202
rect 670193 772888 674046 772948
rect 670193 760389 670253 772888
rect 674178 772756 674238 876201
rect 674367 874046 674433 874047
rect 674367 873982 674368 874046
rect 674432 873982 674433 874046
rect 674367 873981 674433 873982
rect 670385 772696 674238 772756
rect 670385 760581 670445 772696
rect 674370 772564 674430 873981
rect 674559 869902 674625 869903
rect 674559 869838 674560 869902
rect 674624 869838 674625 869902
rect 674559 869837 674625 869838
rect 670577 772504 674430 772564
rect 670577 760773 670637 772504
rect 674562 772372 674622 869837
rect 675711 864722 675777 864723
rect 675711 864658 675712 864722
rect 675776 864658 675777 864722
rect 675711 864657 675777 864658
rect 674943 862946 675009 862947
rect 674943 862882 674944 862946
rect 675008 862882 675009 862946
rect 674943 862881 675009 862882
rect 674751 773702 674817 773703
rect 674751 773638 674752 773702
rect 674816 773638 674817 773702
rect 674751 773637 674817 773638
rect 670769 772312 674622 772372
rect 670769 760965 670829 772312
rect 674754 772180 674814 773637
rect 670961 772120 674814 772180
rect 670961 761157 671021 772120
rect 674946 771988 675006 862881
rect 675327 787910 675393 787911
rect 675327 787846 675328 787910
rect 675392 787846 675393 787910
rect 675327 787845 675393 787846
rect 675135 786726 675201 786727
rect 675135 786662 675136 786726
rect 675200 786662 675201 786726
rect 675135 786661 675201 786662
rect 671153 771928 675006 771988
rect 671153 761349 671213 771928
rect 675138 771796 675198 786661
rect 671345 771736 675198 771796
rect 671345 761541 671405 771736
rect 675330 771604 675390 787845
rect 675519 784802 675585 784803
rect 675519 784738 675520 784802
rect 675584 784738 675585 784802
rect 675519 784737 675585 784738
rect 671537 771544 675390 771604
rect 671537 761733 671597 771544
rect 675522 771412 675582 784737
rect 671729 771352 675582 771412
rect 671729 761925 671789 771352
rect 675714 771220 675774 864657
rect 676287 780658 676353 780659
rect 676287 780594 676288 780658
rect 676352 780594 676353 780658
rect 676287 780593 676353 780594
rect 675903 775478 675969 775479
rect 675903 775414 675904 775478
rect 675968 775414 675969 775478
rect 675903 775413 675969 775414
rect 671921 771160 675774 771220
rect 671921 762117 671981 771160
rect 675906 771028 675966 775413
rect 676290 773116 676350 780593
rect 676863 779178 676929 779179
rect 676863 779114 676864 779178
rect 676928 779114 676929 779178
rect 676863 779113 676929 779114
rect 672113 770968 675966 771028
rect 676190 773056 676350 773116
rect 672113 762309 672173 770968
rect 676190 770744 676250 773056
rect 672497 770684 676250 770744
rect 672497 762693 672557 770684
rect 676866 770488 676926 779113
rect 677058 777551 677502 777585
rect 677055 777550 677502 777551
rect 677055 777486 677056 777550
rect 677120 777525 677502 777550
rect 677120 777486 677121 777525
rect 677055 777485 677121 777486
rect 677055 777402 677121 777403
rect 677055 777338 677056 777402
rect 677120 777338 677121 777402
rect 677055 777337 677121 777338
rect 677058 776919 677118 777337
rect 677058 776859 677310 776919
rect 677055 774886 677121 774887
rect 677055 774822 677056 774886
rect 677120 774822 677121 774886
rect 677055 774821 677121 774822
rect 673073 770428 676926 770488
rect 673073 763269 673133 770428
rect 677058 770296 677118 774821
rect 673265 770236 677118 770296
rect 673265 763461 673325 770236
rect 677250 770104 677310 776859
rect 673457 770044 677310 770104
rect 673457 763653 673517 770044
rect 677442 769912 677502 777525
rect 673649 769852 677502 769912
rect 673649 763845 673709 769852
rect 673649 763785 677502 763845
rect 673457 763593 677310 763653
rect 673265 763401 677118 763461
rect 673073 763209 676926 763269
rect 672497 762633 676350 762693
rect 672113 762249 675966 762309
rect 671921 762057 675774 762117
rect 671729 761865 675582 761925
rect 671537 761673 675390 761733
rect 671345 761481 675198 761541
rect 671153 761289 675006 761349
rect 670961 761097 674814 761157
rect 670769 760905 674622 760965
rect 670577 760713 674430 760773
rect 670385 760521 674238 760581
rect 670193 760329 674046 760389
rect 673986 757275 674046 760329
rect 674178 758459 674238 760521
rect 674175 758458 674241 758459
rect 674175 758394 674176 758458
rect 674240 758394 674241 758458
rect 674175 758393 674241 758394
rect 673983 757274 674049 757275
rect 673983 757210 673984 757274
rect 674048 757210 674049 757274
rect 673983 757209 674049 757210
rect 674370 757127 674430 760713
rect 42879 757126 42945 757127
rect 42879 757062 42880 757126
rect 42944 757062 42945 757126
rect 42879 757061 42945 757062
rect 674367 757126 674433 757127
rect 674367 757062 674368 757126
rect 674432 757062 674433 757126
rect 674367 757061 674433 757062
rect 42495 756534 42561 756535
rect 42495 756470 42496 756534
rect 42560 756470 42561 756534
rect 42495 756469 42561 756470
rect 42498 751059 42558 756469
rect 42495 751058 42561 751059
rect 42495 750994 42496 751058
rect 42560 750994 42561 751058
rect 42495 750993 42561 750994
rect 42882 749875 42942 757061
rect 674562 756387 674622 760905
rect 674559 756386 674625 756387
rect 674559 756322 674560 756386
rect 674624 756322 674625 756386
rect 674559 756321 674625 756322
rect 42879 749874 42945 749875
rect 42879 749810 42880 749874
rect 42944 749810 42945 749874
rect 42879 749809 42945 749810
rect 674367 743214 674433 743215
rect 674367 743150 674368 743214
rect 674432 743150 674433 743214
rect 674367 743149 674433 743150
rect 39974 732961 40034 735848
rect 40770 735794 41198 735854
rect 42114 735816 42522 735876
rect 41138 732973 41198 735794
rect 42462 732973 42522 735816
rect 40578 732961 40638 732973
rect 39974 732901 40638 732961
rect 40578 729007 40638 732901
rect 40770 732913 41198 732973
rect 42114 732913 42522 732973
rect 40770 729895 40830 732913
rect 40767 729894 40833 729895
rect 40767 729830 40768 729894
rect 40832 729830 40833 729894
rect 40767 729829 40833 729830
rect 40959 729894 41025 729895
rect 40959 729830 40960 729894
rect 41024 729830 41025 729894
rect 40959 729829 41025 729830
rect 40575 729006 40641 729007
rect 40575 728942 40576 729006
rect 40640 728942 40641 729006
rect 40575 728941 40641 728942
rect 40383 728858 40449 728859
rect 40383 728794 40384 728858
rect 40448 728794 40449 728858
rect 40383 728793 40449 728794
rect 40386 724305 40446 728793
rect 40386 724245 40638 724305
rect 40383 716574 40449 716575
rect 40383 716510 40384 716574
rect 40448 716510 40449 716574
rect 40383 716509 40449 716510
rect 40386 703403 40446 716509
rect 40383 703402 40449 703403
rect 40383 703338 40384 703402
rect 40448 703338 40449 703402
rect 40383 703337 40449 703338
rect 40578 693022 40638 724245
rect 40767 717018 40833 717019
rect 40767 716954 40768 717018
rect 40832 716954 40833 717018
rect 40767 716953 40833 716954
rect 40770 703699 40830 716953
rect 40767 703698 40833 703699
rect 40767 703634 40768 703698
rect 40832 703634 40833 703698
rect 40767 703633 40833 703634
rect 39888 692962 40638 693022
rect 40962 693043 41022 729829
rect 41727 722642 41793 722643
rect 41727 722578 41728 722642
rect 41792 722578 41793 722642
rect 41727 722577 41793 722578
rect 41730 706067 41790 722577
rect 41919 713910 41985 713911
rect 41919 713846 41920 713910
rect 41984 713846 41985 713910
rect 41919 713845 41985 713846
rect 41922 711691 41982 713845
rect 41919 711690 41985 711691
rect 41919 711626 41920 711690
rect 41984 711626 41985 711690
rect 41919 711625 41985 711626
rect 41727 706066 41793 706067
rect 41727 706002 41728 706066
rect 41792 706002 41793 706066
rect 41727 706001 41793 706002
rect 42114 693060 42174 732913
rect 674370 727960 674430 743149
rect 674559 741734 674625 741735
rect 674559 741670 674560 741734
rect 674624 741670 674625 741734
rect 674559 741669 674625 741670
rect 670894 727900 674430 727960
rect 670894 714305 670954 727900
rect 674562 727768 674622 741669
rect 671086 727708 674622 727768
rect 671086 714497 671146 727708
rect 674754 727576 674814 761097
rect 674946 755795 675006 761289
rect 674943 755794 675009 755795
rect 674943 755730 674944 755794
rect 675008 755730 675009 755794
rect 674943 755729 675009 755730
rect 674943 740402 675009 740403
rect 674943 740338 674944 740402
rect 675008 740338 675009 740402
rect 674943 740337 675009 740338
rect 671278 727516 674814 727576
rect 671278 714689 671338 727516
rect 674946 727384 675006 740337
rect 671470 727324 675006 727384
rect 671470 714881 671530 727324
rect 675138 727192 675198 761481
rect 671662 727132 675198 727192
rect 671662 715073 671722 727132
rect 675330 727000 675390 761673
rect 671854 726940 675390 727000
rect 671854 715265 671914 726940
rect 675522 726808 675582 761865
rect 675714 757867 675774 762057
rect 675711 757866 675777 757867
rect 675711 757802 675712 757866
rect 675776 757802 675777 757866
rect 675711 757801 675777 757802
rect 675711 735518 675777 735519
rect 675711 735454 675712 735518
rect 675776 735454 675777 735518
rect 675711 735453 675777 735454
rect 672046 726748 675582 726808
rect 672046 715457 672106 726748
rect 675714 726616 675774 735453
rect 672238 726556 675774 726616
rect 672238 715649 672298 726556
rect 675906 726424 675966 762249
rect 676095 742178 676161 742179
rect 676095 742114 676096 742178
rect 676160 742114 676161 742178
rect 676095 742113 676161 742114
rect 672430 726364 675966 726424
rect 672430 715841 672490 726364
rect 676098 726232 676158 742113
rect 672622 726172 676158 726232
rect 672622 716033 672682 726172
rect 676290 726040 676350 762633
rect 672814 725980 676350 726040
rect 672814 716225 672874 725980
rect 676866 725464 676926 763209
rect 677058 754167 677118 763401
rect 677055 754166 677121 754167
rect 677055 754102 677056 754166
rect 677120 754102 677121 754166
rect 677055 754101 677121 754102
rect 677055 734482 677121 734483
rect 677055 734418 677056 734482
rect 677120 734418 677121 734482
rect 677055 734417 677121 734418
rect 673390 725404 676926 725464
rect 673390 716801 673450 725404
rect 677058 725272 677118 734417
rect 673582 725212 677118 725272
rect 673582 716993 673642 725212
rect 677250 725080 677310 763593
rect 677442 753723 677502 763785
rect 677439 753722 677505 753723
rect 677439 753658 677440 753722
rect 677504 753658 677505 753722
rect 677439 753657 677505 753658
rect 673774 725020 677310 725080
rect 673774 717185 673834 725020
rect 673774 717125 677310 717185
rect 673582 716933 677118 716993
rect 673390 716741 676926 716801
rect 672814 716165 676350 716225
rect 672622 715973 676158 716033
rect 672430 715781 675966 715841
rect 672238 715589 675774 715649
rect 672046 715397 675582 715457
rect 671854 715205 675390 715265
rect 671662 715013 675198 715073
rect 671470 714821 675006 714881
rect 671278 714629 674814 714689
rect 671086 714437 674622 714497
rect 670894 714245 674430 714305
rect 43071 714058 43137 714059
rect 43071 713994 43072 714058
rect 43136 713994 43137 714058
rect 43071 713993 43137 713994
rect 42879 713910 42945 713911
rect 42879 713846 42880 713910
rect 42944 713846 42945 713910
rect 42879 713845 42945 713846
rect 42882 709767 42942 713845
rect 42879 709766 42945 709767
rect 42879 709702 42880 709766
rect 42944 709702 42945 709766
rect 42879 709701 42945 709702
rect 43074 707251 43134 713993
rect 43071 707250 43137 707251
rect 43071 707186 43072 707250
rect 43136 707186 43137 707250
rect 43071 707185 43137 707186
rect 40962 692983 41159 693043
rect 42114 693000 42445 693060
rect 39888 689831 39948 692962
rect 39888 689771 40638 689831
rect 41099 689801 41159 692983
rect 40578 685643 40638 689771
rect 40770 689741 41159 689801
rect 42114 689785 42174 689801
rect 42385 689785 42445 693000
rect 673983 690526 674049 690527
rect 673983 690462 673984 690526
rect 674048 690462 674049 690526
rect 673983 690461 674049 690462
rect 40770 686679 40830 689741
rect 42114 689725 42445 689785
rect 40767 686678 40833 686679
rect 40767 686614 40768 686678
rect 40832 686614 40833 686678
rect 40767 686613 40833 686614
rect 40959 686678 41025 686679
rect 40959 686614 40960 686678
rect 41024 686614 41025 686678
rect 40959 686613 41025 686614
rect 40575 685642 40641 685643
rect 40575 685578 40576 685642
rect 40640 685578 40641 685642
rect 40575 685577 40641 685578
rect 40575 672618 40641 672619
rect 40575 672554 40576 672618
rect 40640 672554 40641 672618
rect 40575 672553 40641 672554
rect 40383 672470 40449 672471
rect 40383 672406 40384 672470
rect 40448 672406 40449 672470
rect 40383 672405 40449 672406
rect 40386 660335 40446 672405
rect 40578 660927 40638 672553
rect 40575 660926 40641 660927
rect 40575 660862 40576 660926
rect 40640 660862 40641 660926
rect 40575 660861 40641 660862
rect 40383 660334 40449 660335
rect 40383 660270 40384 660334
rect 40448 660270 40449 660334
rect 40383 660269 40449 660270
rect 40962 659550 41022 686613
rect 41151 685790 41217 685791
rect 41151 685726 41152 685790
rect 41216 685726 41217 685790
rect 41151 685725 41217 685726
rect 40770 659490 41022 659550
rect 40770 649585 40830 659490
rect 39954 649525 40830 649585
rect 39954 646713 40014 649525
rect 39954 646653 40830 646713
rect 40770 643463 40830 646653
rect 40767 643462 40833 643463
rect 40767 643398 40768 643462
rect 40832 643398 40833 643462
rect 40767 643397 40833 643398
rect 41154 642427 41214 685725
rect 41727 670694 41793 670695
rect 41727 670630 41728 670694
rect 41792 670630 41793 670694
rect 41727 670629 41793 670630
rect 41730 663443 41790 670629
rect 41727 663442 41793 663443
rect 41727 663378 41728 663442
rect 41792 663378 41793 663442
rect 41727 663377 41793 663378
rect 42114 649613 42174 689725
rect 673986 683146 674046 690461
rect 669934 683086 674046 683146
rect 42495 670694 42561 670695
rect 42495 670630 42496 670694
rect 42560 670630 42561 670694
rect 42495 670629 42561 670630
rect 42303 670102 42369 670103
rect 42303 670038 42304 670102
rect 42368 670038 42369 670102
rect 42303 670037 42369 670038
rect 42306 666699 42366 670037
rect 42303 666698 42369 666699
rect 42303 666634 42304 666698
rect 42368 666634 42369 666698
rect 42303 666633 42369 666634
rect 42498 665219 42558 670629
rect 669934 669448 669994 683086
rect 674370 682762 674430 714245
rect 670318 682702 674430 682762
rect 670318 669832 670378 682702
rect 674562 682570 674622 714437
rect 674754 710803 674814 714629
rect 674751 710802 674817 710803
rect 674751 710738 674752 710802
rect 674816 710738 674817 710802
rect 674751 710737 674817 710738
rect 670510 682510 674622 682570
rect 670510 670024 670570 682510
rect 674946 682186 675006 714821
rect 675138 713467 675198 715013
rect 675135 713466 675201 713467
rect 675135 713402 675136 713466
rect 675200 713402 675201 713466
rect 675135 713401 675201 713402
rect 675330 712283 675390 715205
rect 675327 712282 675393 712283
rect 675327 712218 675328 712282
rect 675392 712218 675393 712282
rect 675327 712217 675393 712218
rect 675522 712135 675582 715397
rect 675519 712134 675585 712135
rect 675519 712070 675520 712134
rect 675584 712070 675585 712134
rect 675519 712069 675585 712070
rect 675327 697926 675393 697927
rect 675327 697862 675328 697926
rect 675392 697862 675393 697926
rect 675327 697861 675393 697862
rect 675135 694818 675201 694819
rect 675135 694754 675136 694818
rect 675200 694754 675201 694818
rect 675135 694753 675201 694754
rect 670894 682126 675006 682186
rect 670894 670408 670954 682126
rect 675138 681994 675198 694753
rect 671086 681934 675198 681994
rect 671086 670600 671146 681934
rect 675330 681802 675390 697861
rect 675519 696890 675585 696891
rect 675519 696826 675520 696890
rect 675584 696826 675585 696890
rect 675519 696825 675585 696826
rect 671278 681742 675390 681802
rect 671278 670792 671338 681742
rect 675522 681610 675582 696825
rect 671470 681550 675582 681610
rect 671470 670984 671530 681550
rect 675714 681418 675774 715589
rect 675906 712875 675966 715781
rect 675903 712874 675969 712875
rect 675903 712810 675904 712874
rect 675968 712810 675969 712874
rect 675903 712809 675969 712810
rect 671662 681358 675774 681418
rect 671662 671176 671722 681358
rect 676098 681034 676158 715973
rect 676290 711691 676350 716165
rect 676287 711690 676353 711691
rect 676287 711626 676288 711690
rect 676352 711626 676353 711690
rect 676287 711625 676353 711626
rect 676866 708583 676926 716741
rect 676863 708582 676929 708583
rect 676863 708518 676864 708582
rect 676928 708518 676929 708582
rect 676863 708517 676929 708518
rect 676287 697334 676353 697335
rect 676287 697270 676288 697334
rect 676352 697270 676353 697334
rect 676287 697269 676353 697270
rect 672046 680974 676158 681034
rect 672046 671560 672106 680974
rect 676290 680842 676350 697269
rect 676479 694226 676545 694227
rect 676479 694162 676480 694226
rect 676544 694162 676545 694226
rect 676479 694161 676545 694162
rect 672238 680782 676350 680842
rect 672238 671752 672298 680782
rect 676482 680650 676542 694161
rect 676863 687418 676929 687419
rect 676863 687354 676864 687418
rect 676928 687354 676929 687418
rect 676863 687353 676929 687354
rect 672430 680590 676542 680650
rect 672430 671944 672490 680590
rect 676866 680266 676926 687353
rect 672814 680206 676926 680266
rect 672814 672328 672874 680206
rect 677058 680074 677118 716933
rect 677250 709175 677310 717125
rect 677247 709174 677313 709175
rect 677247 709110 677248 709174
rect 677312 709110 677313 709174
rect 677247 709109 677313 709110
rect 673006 680014 677118 680074
rect 673006 672520 673066 680014
rect 673006 672460 677118 672520
rect 672814 672268 676926 672328
rect 672430 671884 676542 671944
rect 672238 671692 676350 671752
rect 672046 671500 676158 671560
rect 671662 671116 675774 671176
rect 671470 670924 675582 670984
rect 671278 670732 675390 670792
rect 671086 670540 675198 670600
rect 670894 670348 675006 670408
rect 670510 669964 674622 670024
rect 670318 669772 674430 669832
rect 669934 669388 674046 669448
rect 42495 665218 42561 665219
rect 42495 665154 42496 665218
rect 42560 665154 42561 665218
rect 42495 665153 42561 665154
rect 42114 649553 42522 649613
rect 42114 646628 42174 646634
rect 42462 646628 42522 649553
rect 42114 646568 42522 646628
rect 41151 642426 41217 642427
rect 41151 642362 41152 642426
rect 41216 642362 41217 642426
rect 41151 642361 41217 642362
rect 41727 635840 41793 635841
rect 41727 635776 41728 635840
rect 41792 635776 41793 635840
rect 41727 635775 41793 635776
rect 40383 629106 40449 629107
rect 40383 629042 40384 629106
rect 40448 629042 40449 629106
rect 40383 629041 40449 629042
rect 40386 616527 40446 629041
rect 40575 627922 40641 627923
rect 40575 627858 40576 627922
rect 40640 627858 40641 627922
rect 40575 627857 40641 627858
rect 41535 627922 41601 627923
rect 41535 627858 41536 627922
rect 41600 627858 41601 627922
rect 41535 627857 41601 627858
rect 40578 618895 40638 627857
rect 40575 618894 40641 618895
rect 40575 618830 40576 618894
rect 40640 618830 40641 618894
rect 40575 618829 40641 618830
rect 40383 616526 40449 616527
rect 40383 616462 40384 616526
rect 40448 616462 40449 616526
rect 40383 616461 40449 616462
rect 41538 616083 41598 627857
rect 41730 620967 41790 635775
rect 41727 620966 41793 620967
rect 41727 620902 41728 620966
rect 41792 620902 41793 620966
rect 41727 620901 41793 620902
rect 41727 619190 41793 619191
rect 41727 619126 41728 619190
rect 41792 619126 41793 619190
rect 41727 619125 41793 619126
rect 41535 616082 41601 616083
rect 41535 616018 41536 616082
rect 41600 616018 41601 616082
rect 41535 616017 41601 616018
rect 41535 607646 41601 607647
rect 41535 607582 41536 607646
rect 41600 607582 41601 607646
rect 41535 607581 41601 607582
rect 41538 606519 41598 607581
rect 41107 606459 41598 606519
rect 41107 603449 41167 606459
rect 41730 606347 41790 619125
rect 42114 606561 42174 646568
rect 673986 637800 674046 669388
rect 674370 667143 674430 669772
rect 674562 668179 674622 669964
rect 674559 668178 674625 668179
rect 674559 668114 674560 668178
rect 674624 668114 674625 668178
rect 674559 668113 674625 668114
rect 674367 667142 674433 667143
rect 674367 667078 674368 667142
rect 674432 667078 674433 667142
rect 674367 667077 674433 667078
rect 674946 666699 675006 670348
rect 674943 666698 675009 666699
rect 674943 666634 674944 666698
rect 675008 666634 675009 666698
rect 674943 666633 675009 666634
rect 674943 652638 675009 652639
rect 674943 652574 674944 652638
rect 675008 652574 675009 652638
rect 674943 652573 675009 652574
rect 674559 651602 674625 651603
rect 674559 651538 674560 651602
rect 674624 651538 674625 651602
rect 674559 651537 674625 651538
rect 674175 645386 674241 645387
rect 674175 645322 674176 645386
rect 674240 645322 674241 645386
rect 674175 645321 674241 645322
rect 670613 637740 674046 637800
rect 42495 628070 42561 628071
rect 42495 628006 42496 628070
rect 42560 628006 42561 628070
rect 42495 628005 42561 628006
rect 42303 627774 42369 627775
rect 42303 627710 42304 627774
rect 42368 627710 42369 627774
rect 42303 627709 42369 627710
rect 42306 621559 42366 627709
rect 42498 622151 42558 628005
rect 42879 627478 42945 627479
rect 42879 627414 42880 627478
rect 42944 627414 42945 627478
rect 42879 627413 42945 627414
rect 42495 622150 42561 622151
rect 42495 622086 42496 622150
rect 42560 622086 42561 622150
rect 42495 622085 42561 622086
rect 42303 621558 42369 621559
rect 42303 621494 42304 621558
rect 42368 621494 42369 621558
rect 42303 621493 42369 621494
rect 42882 620227 42942 627413
rect 670613 625612 670673 637740
rect 674178 637608 674238 645321
rect 670805 637548 674238 637608
rect 670805 625804 670865 637548
rect 674562 637224 674622 651537
rect 674751 638578 674817 638579
rect 674751 638514 674752 638578
rect 674816 638514 674817 638578
rect 674751 638513 674817 638514
rect 671189 637164 674622 637224
rect 671189 626188 671249 637164
rect 674754 637032 674814 638513
rect 671381 636972 674814 637032
rect 671381 626380 671441 636972
rect 674946 636840 675006 652573
rect 671573 636780 675006 636840
rect 671573 626572 671633 636780
rect 675138 636648 675198 670540
rect 671765 636588 675198 636648
rect 671765 626764 671825 636588
rect 675330 636456 675390 670732
rect 671957 636396 675390 636456
rect 671957 626956 672017 636396
rect 675522 636264 675582 670924
rect 675714 666181 675774 671116
rect 675711 666180 675777 666181
rect 675711 666116 675712 666180
rect 675776 666116 675777 666180
rect 675711 666115 675777 666116
rect 676098 665071 676158 671500
rect 676095 665070 676161 665071
rect 676095 665006 676096 665070
rect 676160 665006 676161 665070
rect 676095 665005 676161 665006
rect 675711 649678 675777 649679
rect 675711 649614 675712 649678
rect 675776 649614 675777 649678
rect 675711 649613 675777 649614
rect 672149 636204 675582 636264
rect 672149 627148 672209 636204
rect 675714 636072 675774 649613
rect 675903 640354 675969 640355
rect 675903 640290 675904 640354
rect 675968 640290 675969 640354
rect 675903 640289 675969 640290
rect 672341 636012 675774 636072
rect 672341 627340 672401 636012
rect 675906 635880 675966 640289
rect 672533 635820 675966 635880
rect 672533 627532 672593 635820
rect 676290 635496 676350 671692
rect 672917 635436 676350 635496
rect 672917 627916 672977 635436
rect 676482 635304 676542 671884
rect 673109 635244 676542 635304
rect 673109 628108 673169 635244
rect 676866 634920 676926 672268
rect 677058 663443 677118 672460
rect 677055 663442 677121 663443
rect 677055 663378 677056 663442
rect 677120 663378 677121 663442
rect 677055 663377 677121 663378
rect 673493 634860 676926 634920
rect 673493 628492 673553 634860
rect 673493 628432 676926 628492
rect 673109 628048 676542 628108
rect 672917 627856 676350 627916
rect 672533 627472 675966 627532
rect 672341 627280 675774 627340
rect 672149 627088 675582 627148
rect 671957 626896 675390 626956
rect 671765 626704 675198 626764
rect 671573 626512 675006 626572
rect 671381 626320 674814 626380
rect 671189 626128 674622 626188
rect 670805 625744 674238 625804
rect 670613 625552 674046 625612
rect 673986 621115 674046 625552
rect 673983 621114 674049 621115
rect 673983 621050 673984 621114
rect 674048 621050 674049 621114
rect 673983 621049 674049 621050
rect 42879 620226 42945 620227
rect 42879 620162 42880 620226
rect 42944 620162 42945 620226
rect 42879 620161 42945 620162
rect 673983 607794 674049 607795
rect 673983 607730 673984 607794
rect 674048 607730 674049 607794
rect 673983 607729 674049 607730
rect 42114 606501 42494 606561
rect 41247 606287 41790 606347
rect 41247 603636 41307 606287
rect 41247 603576 41790 603636
rect 41107 603389 41598 603449
rect 40767 600690 40833 600691
rect 40767 600626 40768 600690
rect 40832 600626 40833 600690
rect 40767 600625 40833 600626
rect 40575 599358 40641 599359
rect 40575 599294 40576 599358
rect 40640 599294 40641 599358
rect 40575 599293 40641 599294
rect 40383 585586 40449 585587
rect 40383 585522 40384 585586
rect 40448 585522 40449 585586
rect 40383 585521 40449 585522
rect 40386 574051 40446 585521
rect 40383 574050 40449 574051
rect 40383 573986 40384 574050
rect 40448 573986 40449 574050
rect 40383 573985 40449 573986
rect 40578 563732 40638 599293
rect 40770 563876 40830 600625
rect 41538 599803 41598 603389
rect 41730 600543 41790 603576
rect 42434 603468 42494 606501
rect 42114 603408 42494 603468
rect 41727 600542 41793 600543
rect 41727 600478 41728 600542
rect 41792 600478 41793 600542
rect 41727 600477 41793 600478
rect 41535 599802 41601 599803
rect 41535 599738 41536 599802
rect 41600 599738 41601 599802
rect 41535 599737 41601 599738
rect 40959 585438 41025 585439
rect 40959 585374 40960 585438
rect 41024 585374 41025 585438
rect 40959 585373 41025 585374
rect 40962 574495 41022 585373
rect 40959 574494 41025 574495
rect 40959 574430 40960 574494
rect 41024 574430 41025 574494
rect 40959 574429 41025 574430
rect 42114 563886 42174 603408
rect 673986 591326 674046 607729
rect 671315 591266 674046 591326
rect 43071 584558 43137 584559
rect 43071 584494 43072 584558
rect 43136 584494 43137 584558
rect 43071 584493 43137 584494
rect 42879 584262 42945 584263
rect 42879 584198 42880 584262
rect 42944 584198 42945 584262
rect 42879 584197 42945 584198
rect 42882 578787 42942 584197
rect 42879 578786 42945 578787
rect 42879 578722 42880 578786
rect 42944 578722 42945 578786
rect 42879 578721 42945 578722
rect 43074 577603 43134 584493
rect 671315 581376 671375 591266
rect 674178 591134 674238 625744
rect 674367 604834 674433 604835
rect 674367 604770 674368 604834
rect 674432 604770 674433 604834
rect 674367 604769 674433 604770
rect 671507 591074 674238 591134
rect 671507 581568 671567 591074
rect 674370 590942 674430 604769
rect 671699 590882 674430 590942
rect 671699 581760 671759 590882
rect 674562 590750 674622 626128
rect 671891 590690 674622 590750
rect 671891 581952 671951 590690
rect 674754 590558 674814 626320
rect 672083 590498 674814 590558
rect 672083 582144 672143 590498
rect 674946 590366 675006 626512
rect 675138 621707 675198 626704
rect 675330 622151 675390 626896
rect 675522 623187 675582 627088
rect 675519 623186 675585 623187
rect 675519 623122 675520 623186
rect 675584 623122 675585 623186
rect 675519 623121 675585 623122
rect 675327 622150 675393 622151
rect 675327 622086 675328 622150
rect 675392 622086 675393 622150
rect 675327 622085 675393 622086
rect 675135 621706 675201 621707
rect 675135 621642 675136 621706
rect 675200 621642 675201 621706
rect 675135 621641 675201 621642
rect 675135 606462 675201 606463
rect 675135 606398 675136 606462
rect 675200 606398 675201 606462
rect 675135 606397 675201 606398
rect 672275 590306 675006 590366
rect 672275 582336 672335 590306
rect 675138 590174 675198 606397
rect 675327 600246 675393 600247
rect 675327 600182 675328 600246
rect 675392 600182 675393 600246
rect 675327 600181 675393 600182
rect 672467 590114 675198 590174
rect 672467 582528 672527 590114
rect 675330 589982 675390 600181
rect 675519 593438 675585 593439
rect 675519 593374 675520 593438
rect 675584 593374 675585 593438
rect 675519 593373 675585 593374
rect 672659 589922 675390 589982
rect 672659 582720 672719 589922
rect 675522 589790 675582 593373
rect 672851 589730 675582 589790
rect 672851 582912 672911 589730
rect 675714 589598 675774 627280
rect 673043 589538 675774 589598
rect 673043 583104 673103 589538
rect 675906 589406 675966 627472
rect 676290 620375 676350 627856
rect 676287 620374 676353 620375
rect 676287 620310 676288 620374
rect 676352 620310 676353 620374
rect 676287 620309 676353 620310
rect 676482 619931 676542 628048
rect 676479 619930 676545 619931
rect 676479 619866 676480 619930
rect 676544 619866 676545 619930
rect 676479 619865 676545 619866
rect 676866 618895 676926 628432
rect 676863 618894 676929 618895
rect 676863 618830 676864 618894
rect 676928 618830 676929 618894
rect 676863 618829 676929 618830
rect 676095 595362 676161 595363
rect 676095 595298 676096 595362
rect 676160 595298 676161 595362
rect 676095 595297 676161 595298
rect 673235 589346 675966 589406
rect 673235 583296 673295 589346
rect 676098 589214 676158 595297
rect 673427 589154 676158 589214
rect 673427 583488 673487 589154
rect 673427 583428 676158 583488
rect 673235 583236 675966 583296
rect 673043 583044 675774 583104
rect 672851 582852 675582 582912
rect 672659 582660 675390 582720
rect 672467 582468 675198 582528
rect 672275 582276 675006 582336
rect 672083 582084 674814 582144
rect 671891 581892 674622 581952
rect 671699 581700 674430 581760
rect 671507 581508 674238 581568
rect 671315 581316 674046 581376
rect 43071 577602 43137 577603
rect 43071 577538 43072 577602
rect 43136 577538 43137 577602
rect 43071 577537 43137 577538
rect 40770 563816 41263 563876
rect 42114 563826 42630 563886
rect 40578 563672 41135 563732
rect 41075 560615 41135 563672
rect 40578 560555 41135 560615
rect 40383 557474 40449 557475
rect 40383 557410 40384 557474
rect 40448 557410 40449 557474
rect 40383 557409 40449 557410
rect 40386 550110 40446 557409
rect 40578 555995 40638 560555
rect 41203 560461 41263 563816
rect 40770 560401 41263 560461
rect 40770 556735 40830 560401
rect 42570 560327 42630 563826
rect 42114 560267 42630 560327
rect 41727 558954 41793 558955
rect 41727 558890 41728 558954
rect 41792 558890 41793 558954
rect 41727 558889 41793 558890
rect 40767 556734 40833 556735
rect 40767 556670 40768 556734
rect 40832 556670 40833 556734
rect 40767 556669 40833 556670
rect 41730 556365 41790 558889
rect 41727 556364 41793 556365
rect 41727 556300 41728 556364
rect 41792 556300 41793 556364
rect 41727 556299 41793 556300
rect 40767 556142 40833 556143
rect 40767 556078 40768 556142
rect 40832 556078 40833 556142
rect 40767 556077 40833 556078
rect 40575 555994 40641 555995
rect 40575 555930 40576 555994
rect 40640 555930 40641 555994
rect 40575 555929 40641 555930
rect 40386 550050 40638 550110
rect 40578 545453 40638 550050
rect 40770 545634 40830 556077
rect 40770 545574 41241 545634
rect 40578 545393 41090 545453
rect 41030 542284 41090 545393
rect 40578 542224 41090 542284
rect 40578 435736 40638 542224
rect 41181 542067 41241 545574
rect 42114 545613 42174 560267
rect 42114 545553 42467 545613
rect 42407 542127 42467 545553
rect 673986 545509 674046 581316
rect 674178 575975 674238 581508
rect 674175 575974 674241 575975
rect 674175 575910 674176 575974
rect 674240 575910 674241 575974
rect 674175 575909 674241 575910
rect 40770 542007 41241 542067
rect 42114 542067 42467 542127
rect 671910 545449 674046 545509
rect 40770 435893 40830 542007
rect 40959 541638 41025 541639
rect 40959 541574 40960 541638
rect 41024 541574 41025 541638
rect 40959 541573 41025 541574
rect 40962 531427 41022 541573
rect 41151 541490 41217 541491
rect 41151 541426 41152 541490
rect 41216 541426 41217 541490
rect 41151 541425 41217 541426
rect 40959 531426 41025 531427
rect 40959 531362 40960 531426
rect 41024 531362 41025 531426
rect 40959 531361 41025 531362
rect 41154 526543 41214 541425
rect 41727 541342 41793 541343
rect 41727 541278 41728 541342
rect 41792 541278 41793 541342
rect 41727 541277 41793 541278
rect 41730 529651 41790 541277
rect 41919 541046 41985 541047
rect 41919 540982 41920 541046
rect 41984 540982 41985 541046
rect 41919 540981 41985 540982
rect 41922 530687 41982 540981
rect 41919 530686 41985 530687
rect 41919 530622 41920 530686
rect 41984 530622 41985 530686
rect 41919 530621 41985 530622
rect 41727 529650 41793 529651
rect 41727 529586 41728 529650
rect 41792 529586 41793 529650
rect 41727 529585 41793 529586
rect 41151 526542 41217 526543
rect 41151 526478 41152 526542
rect 41216 526478 41217 526542
rect 41151 526477 41217 526478
rect 42114 435967 42174 542067
rect 42495 541638 42561 541639
rect 42495 541574 42496 541638
rect 42560 541574 42561 541638
rect 42495 541573 42561 541574
rect 42303 541046 42369 541047
rect 42303 540982 42304 541046
rect 42368 540982 42369 541046
rect 42303 540981 42369 540982
rect 42306 535719 42366 540981
rect 42303 535718 42369 535719
rect 42303 535654 42304 535718
rect 42368 535654 42369 535718
rect 42303 535653 42369 535654
rect 42498 535127 42558 541573
rect 671910 536326 671970 545449
rect 674370 545125 674430 581700
rect 674562 578047 674622 581892
rect 674559 578046 674625 578047
rect 674559 577982 674560 578046
rect 674624 577982 674625 578046
rect 674559 577981 674625 577982
rect 674754 575383 674814 582084
rect 674946 577307 675006 582276
rect 674943 577306 675009 577307
rect 674943 577242 674944 577306
rect 675008 577242 675009 577306
rect 674943 577241 675009 577242
rect 674751 575382 674817 575383
rect 674751 575318 674752 575382
rect 674816 575318 674817 575382
rect 674751 575317 674817 575318
rect 674559 562654 674625 562655
rect 674559 562590 674560 562654
rect 674624 562590 674625 562654
rect 674559 562589 674625 562590
rect 672294 545065 674430 545125
rect 672294 536710 672354 545065
rect 674562 544933 674622 562589
rect 674943 561766 675009 561767
rect 674943 561702 674944 561766
rect 675008 561702 675009 561766
rect 674943 561701 675009 561702
rect 674751 561470 674817 561471
rect 674751 561406 674752 561470
rect 674816 561406 674817 561470
rect 674751 561405 674817 561406
rect 672486 544873 674622 544933
rect 672486 536902 672546 544873
rect 674754 544741 674814 561405
rect 672678 544681 674814 544741
rect 672678 537094 672738 544681
rect 674946 544549 675006 561701
rect 672870 544489 675006 544549
rect 672870 537286 672930 544489
rect 675138 544357 675198 582468
rect 673062 544297 675198 544357
rect 673062 537478 673122 544297
rect 675330 544165 675390 582660
rect 673254 544105 675390 544165
rect 673254 537670 673314 544105
rect 675522 543973 675582 582852
rect 675714 576567 675774 583044
rect 675906 577455 675966 583236
rect 675903 577454 675969 577455
rect 675903 577390 675904 577454
rect 675968 577390 675969 577454
rect 675903 577389 675969 577390
rect 675711 576566 675777 576567
rect 675711 576502 675712 576566
rect 675776 576502 675777 576566
rect 675711 576501 675777 576502
rect 673446 543913 675582 543973
rect 673446 537862 673506 543913
rect 673446 537802 675582 537862
rect 673254 537610 675390 537670
rect 673062 537418 675198 537478
rect 672870 537226 675006 537286
rect 672678 537034 674814 537094
rect 672486 536842 674622 536902
rect 672294 536650 674430 536710
rect 671910 536266 674046 536326
rect 42495 535126 42561 535127
rect 42495 535062 42496 535126
rect 42560 535062 42561 535126
rect 42495 535061 42561 535062
rect 673986 531871 674046 536266
rect 673983 531870 674049 531871
rect 673983 531806 673984 531870
rect 674048 531806 674049 531870
rect 673983 531805 674049 531806
rect 674370 531575 674430 536650
rect 674367 531574 674433 531575
rect 674367 531510 674368 531574
rect 674432 531510 674433 531574
rect 674367 531509 674433 531510
rect 674562 501384 674622 536842
rect 674362 501324 674622 501384
rect 674362 487915 674422 501324
rect 674754 501225 674814 537034
rect 674554 501165 674814 501225
rect 674554 489247 674614 501165
rect 674946 501078 675006 537226
rect 675138 533055 675198 537418
rect 675135 533054 675201 533055
rect 675135 532990 675136 533054
rect 675200 532990 675201 533054
rect 675135 532989 675201 532990
rect 675330 530983 675390 537610
rect 675327 530982 675393 530983
rect 675327 530918 675328 530982
rect 675392 530918 675393 530982
rect 675327 530917 675393 530918
rect 675522 530391 675582 537802
rect 676098 532759 676158 583428
rect 676863 557622 676929 557623
rect 676863 557558 676864 557622
rect 676928 557558 676929 557622
rect 676863 557557 676929 557558
rect 676866 544149 676926 557557
rect 676269 544089 676926 544149
rect 676269 538249 676329 544089
rect 676269 538189 676926 538249
rect 676095 532758 676161 532759
rect 676095 532694 676096 532758
rect 676160 532694 676161 532758
rect 676095 532693 676161 532694
rect 675519 530390 675585 530391
rect 675519 530326 675520 530390
rect 675584 530326 675585 530390
rect 675519 530325 675585 530326
rect 674746 501018 675006 501078
rect 674551 489246 674617 489247
rect 674551 489182 674552 489246
rect 674616 489182 674617 489246
rect 674551 489181 674617 489182
rect 674359 487914 674425 487915
rect 674359 487850 674360 487914
rect 674424 487850 674425 487914
rect 674359 487849 674425 487850
rect 674746 485991 674806 501018
rect 676866 500557 676926 538189
rect 676137 500497 676926 500557
rect 676137 494483 676197 500497
rect 676137 494423 676926 494483
rect 674743 485990 674809 485991
rect 674743 485926 674744 485990
rect 674808 485926 674809 485990
rect 674743 485925 674809 485926
rect 676866 483771 676926 494423
rect 676863 483770 676929 483771
rect 676863 483706 676864 483770
rect 676928 483706 676929 483770
rect 676863 483705 676929 483706
rect 42114 435907 42516 435967
rect 40770 435833 41278 435893
rect 40578 435676 41137 435736
rect 41077 432326 41137 435676
rect 40578 432266 41137 432326
rect 40578 429899 40638 432266
rect 41218 432084 41278 435833
rect 40770 432024 41278 432084
rect 40575 429898 40641 429899
rect 40575 429834 40576 429898
rect 40640 429834 40641 429898
rect 40575 429833 40641 429834
rect 40770 428567 40830 432024
rect 42456 431836 42516 435907
rect 42114 431776 42516 431836
rect 41727 429750 41793 429751
rect 41727 429686 41728 429750
rect 41792 429686 41793 429750
rect 41727 429685 41793 429686
rect 40767 428566 40833 428567
rect 40767 428502 40768 428566
rect 40832 428502 40833 428566
rect 40767 428501 40833 428502
rect 40767 427530 40833 427531
rect 40767 427466 40768 427530
rect 40832 427466 40833 427530
rect 40767 427465 40833 427466
rect 40383 425458 40449 425459
rect 40383 425394 40384 425458
rect 40448 425394 40449 425458
rect 40383 425393 40449 425394
rect 40386 406071 40446 425393
rect 40575 422054 40641 422055
rect 40575 421990 40576 422054
rect 40640 421990 40641 422054
rect 40575 421989 40641 421990
rect 40383 406070 40449 406071
rect 40383 406006 40384 406070
rect 40448 406006 40449 406070
rect 40383 406005 40449 406006
rect 40578 403851 40638 421989
rect 40575 403850 40641 403851
rect 40575 403786 40576 403850
rect 40640 403786 40641 403850
rect 40575 403785 40641 403786
rect 40770 400003 40830 427465
rect 40959 426050 41025 426051
rect 40959 425986 40960 426050
rect 41024 425986 41025 426050
rect 40959 425985 41025 425986
rect 40962 401927 41022 425985
rect 41151 424570 41217 424571
rect 41151 424506 41152 424570
rect 41216 424506 41217 424570
rect 41151 424505 41217 424506
rect 40959 401926 41025 401927
rect 40959 401862 40960 401926
rect 41024 401862 41025 401926
rect 40959 401861 41025 401862
rect 40767 400002 40833 400003
rect 40767 399938 40768 400002
rect 40832 399938 40833 400002
rect 40767 399937 40833 399938
rect 41154 399559 41214 424505
rect 41343 423978 41409 423979
rect 41343 423914 41344 423978
rect 41408 423914 41409 423978
rect 41343 423913 41409 423914
rect 41346 402519 41406 423913
rect 41535 423534 41601 423535
rect 41535 423470 41536 423534
rect 41600 423470 41601 423534
rect 41535 423469 41601 423470
rect 41538 403111 41598 423469
rect 41535 403110 41601 403111
rect 41535 403046 41536 403110
rect 41600 403046 41601 403110
rect 41535 403045 41601 403046
rect 41343 402518 41409 402519
rect 41343 402454 41344 402518
rect 41408 402454 41409 402518
rect 41343 402453 41409 402454
rect 41151 399558 41217 399559
rect 41151 399494 41152 399558
rect 41216 399494 41217 399558
rect 41151 399493 41217 399494
rect 41730 392410 41790 429685
rect 42114 429150 42174 431776
rect 42114 429090 42558 429150
rect 41919 427234 41985 427235
rect 41919 427170 41920 427234
rect 41984 427170 41985 427234
rect 41919 427169 41985 427170
rect 41922 411251 41982 427169
rect 42303 426494 42369 426495
rect 42303 426430 42304 426494
rect 42368 426430 42369 426494
rect 42303 426429 42369 426430
rect 41919 411250 41985 411251
rect 41919 411186 41920 411250
rect 41984 411186 41985 411250
rect 41919 411185 41985 411186
rect 42306 409953 42366 426429
rect 41922 409893 42366 409953
rect 41922 398967 41982 409893
rect 42498 408990 42558 429090
rect 42114 408930 42558 408990
rect 41919 398966 41985 398967
rect 41919 398902 41920 398966
rect 41984 398902 41985 398966
rect 41919 398901 41985 398902
rect 42114 392602 42174 408930
rect 676671 400446 676737 400447
rect 676671 400382 676672 400446
rect 676736 400382 676737 400446
rect 676671 400381 676737 400382
rect 674175 400298 674241 400299
rect 674175 400234 674176 400298
rect 674240 400234 674241 400298
rect 674175 400233 674241 400234
rect 42114 392542 42426 392602
rect 41130 392350 41790 392410
rect 41130 390967 41190 392350
rect 41127 390966 41193 390967
rect 41127 390902 41128 390966
rect 41192 390902 41193 390966
rect 41127 390901 41193 390902
rect 42366 389109 42426 392542
rect 42114 389049 42426 389109
rect 41727 386534 41793 386535
rect 41727 386470 41728 386534
rect 41792 386470 41793 386534
rect 41727 386469 41793 386470
rect 41730 384645 41790 386469
rect 40578 384585 41790 384645
rect 40383 382242 40449 382243
rect 40383 382178 40384 382242
rect 40448 382178 40449 382242
rect 40383 382177 40449 382178
rect 40386 362855 40446 382177
rect 40383 362854 40449 362855
rect 40383 362790 40384 362854
rect 40448 362790 40449 362854
rect 40383 362789 40449 362790
rect 40578 349856 40638 384585
rect 41730 384463 41790 384585
rect 41727 384462 41793 384463
rect 41727 384398 41728 384462
rect 41792 384398 41793 384462
rect 41727 384397 41793 384398
rect 40767 384314 40833 384315
rect 40767 384250 40768 384314
rect 40832 384250 40833 384314
rect 40767 384249 40833 384250
rect 40770 356935 40830 384249
rect 41919 384018 41985 384019
rect 41919 383954 41920 384018
rect 41984 383954 41985 384018
rect 41919 383953 41985 383954
rect 40959 383278 41025 383279
rect 40959 383214 40960 383278
rect 41024 383214 41025 383278
rect 40959 383213 41025 383214
rect 40767 356934 40833 356935
rect 40767 356870 40768 356934
rect 40832 356870 40833 356934
rect 40767 356869 40833 356870
rect 40962 355603 41022 383213
rect 41343 382834 41409 382835
rect 41343 382770 41344 382834
rect 41408 382770 41409 382834
rect 41343 382769 41409 382770
rect 41151 381354 41217 381355
rect 41151 381290 41152 381354
rect 41216 381290 41217 381354
rect 41151 381289 41217 381290
rect 41154 356491 41214 381289
rect 41346 358711 41406 382769
rect 41727 381058 41793 381059
rect 41727 380994 41728 381058
rect 41792 380994 41793 381058
rect 41727 380993 41793 380994
rect 41535 380318 41601 380319
rect 41535 380254 41536 380318
rect 41600 380254 41601 380318
rect 41535 380253 41601 380254
rect 41538 359895 41598 380253
rect 41535 359894 41601 359895
rect 41535 359830 41536 359894
rect 41600 359830 41601 359894
rect 41535 359829 41601 359830
rect 41730 359451 41790 380993
rect 41922 368183 41982 383953
rect 41919 368182 41985 368183
rect 41919 368118 41920 368182
rect 41984 368118 41985 368182
rect 41919 368117 41985 368118
rect 41727 359450 41793 359451
rect 41727 359386 41728 359450
rect 41792 359386 41793 359450
rect 41727 359385 41793 359386
rect 41343 358710 41409 358711
rect 41343 358646 41344 358710
rect 41408 358646 41409 358710
rect 41343 358645 41409 358646
rect 41151 356490 41217 356491
rect 41151 356426 41152 356490
rect 41216 356426 41217 356490
rect 41151 356425 41217 356426
rect 40959 355602 41025 355603
rect 40959 355538 40960 355602
rect 41024 355538 41025 355602
rect 40959 355537 41025 355538
rect 40578 349796 41197 349856
rect 41137 346345 41197 349796
rect 42114 349841 42174 389049
rect 674178 373807 674238 400233
rect 676479 399558 676545 399559
rect 676479 399494 676480 399558
rect 676544 399494 676545 399558
rect 676479 399493 676545 399494
rect 674943 399262 675009 399263
rect 674943 399198 674944 399262
rect 675008 399198 675009 399262
rect 674943 399197 675009 399198
rect 674367 398818 674433 398819
rect 674367 398754 674368 398818
rect 674432 398754 674433 398818
rect 674367 398753 674433 398754
rect 674370 378839 674430 398753
rect 674946 382983 675006 399197
rect 675519 398226 675585 398227
rect 675519 398162 675520 398226
rect 675584 398162 675585 398226
rect 675519 398161 675585 398162
rect 675327 396894 675393 396895
rect 675327 396830 675328 396894
rect 675392 396830 675393 396894
rect 675327 396829 675393 396830
rect 675135 396746 675201 396747
rect 675135 396682 675136 396746
rect 675200 396682 675201 396746
rect 675135 396681 675201 396682
rect 674943 382982 675009 382983
rect 674943 382918 674944 382982
rect 675008 382918 675009 382982
rect 674943 382917 675009 382918
rect 675138 382835 675198 396681
rect 675135 382834 675201 382835
rect 675135 382770 675136 382834
rect 675200 382770 675201 382834
rect 675135 382769 675201 382770
rect 675330 382243 675390 396829
rect 675327 382242 675393 382243
rect 675327 382178 675328 382242
rect 675392 382178 675393 382242
rect 675327 382177 675393 382178
rect 674367 378838 674433 378839
rect 674367 378774 674368 378838
rect 674432 378774 674433 378838
rect 674367 378773 674433 378774
rect 674175 373806 674241 373807
rect 674175 373742 674176 373806
rect 674240 373742 674241 373806
rect 674175 373741 674241 373742
rect 675522 372031 675582 398161
rect 675903 397782 675969 397783
rect 675903 397718 675904 397782
rect 675968 397718 675969 397782
rect 675903 397717 675969 397718
rect 675711 395266 675777 395267
rect 675711 395202 675712 395266
rect 675776 395202 675777 395266
rect 675711 395201 675777 395202
rect 675714 381207 675774 395201
rect 675906 385647 675966 397717
rect 676095 396006 676161 396007
rect 676095 395942 676096 396006
rect 676160 395942 676161 396006
rect 676095 395941 676161 395942
rect 675903 385646 675969 385647
rect 675903 385582 675904 385646
rect 675968 385582 675969 385646
rect 675903 385581 675969 385582
rect 675711 381206 675777 381207
rect 675711 381142 675712 381206
rect 675776 381142 675777 381206
rect 675711 381141 675777 381142
rect 676098 375731 676158 395941
rect 676287 394674 676353 394675
rect 676287 394610 676288 394674
rect 676352 394610 676353 394674
rect 676287 394609 676353 394610
rect 676290 377951 676350 394609
rect 676482 385943 676542 399493
rect 676479 385942 676545 385943
rect 676479 385878 676480 385942
rect 676544 385878 676545 385942
rect 676479 385877 676545 385878
rect 676674 384759 676734 400381
rect 676671 384758 676737 384759
rect 676671 384694 676672 384758
rect 676736 384694 676737 384758
rect 676671 384693 676737 384694
rect 676287 377950 676353 377951
rect 676287 377886 676288 377950
rect 676352 377886 676353 377950
rect 676287 377885 676353 377886
rect 676095 375730 676161 375731
rect 676095 375666 676096 375730
rect 676160 375666 676161 375730
rect 676095 375665 676161 375666
rect 675519 372030 675585 372031
rect 675519 371966 675520 372030
rect 675584 371966 675585 372030
rect 675519 371965 675585 371966
rect 673983 358118 674049 358119
rect 673983 358054 673984 358118
rect 674048 358054 674049 358118
rect 673983 358053 674049 358054
rect 42114 349781 42549 349841
rect 42489 346415 42549 349781
rect 40578 346285 41197 346345
rect 42114 346355 42549 346415
rect 40578 342727 40638 346285
rect 40575 342726 40641 342727
rect 40575 342662 40576 342726
rect 40640 342662 40641 342726
rect 40575 342661 40641 342662
rect 40767 341098 40833 341099
rect 40767 341034 40768 341098
rect 40832 341034 40833 341098
rect 40767 341033 40833 341034
rect 40575 340506 40641 340507
rect 40575 340442 40576 340506
rect 40640 340442 40641 340506
rect 40575 340441 40641 340442
rect 40383 339026 40449 339027
rect 40383 338962 40384 339026
rect 40448 338962 40449 339026
rect 40383 338961 40449 338962
rect 40386 319787 40446 338961
rect 40383 319786 40449 319787
rect 40383 319722 40384 319786
rect 40448 319722 40449 319786
rect 40383 319721 40449 319722
rect 40578 312387 40638 340441
rect 40770 313719 40830 341033
rect 41727 340876 41793 340877
rect 41727 340812 41728 340876
rect 41792 340812 41793 340876
rect 41727 340811 41793 340812
rect 41151 339618 41217 339619
rect 41151 339554 41152 339618
rect 41216 339554 41217 339618
rect 41151 339553 41217 339554
rect 40959 338138 41025 338139
rect 40959 338074 40960 338138
rect 41024 338074 41025 338138
rect 40959 338073 41025 338074
rect 40767 313718 40833 313719
rect 40767 313654 40768 313718
rect 40832 313654 40833 313718
rect 40767 313653 40833 313654
rect 40962 313275 41022 338073
rect 41154 315495 41214 339553
rect 41343 337546 41409 337547
rect 41343 337482 41344 337546
rect 41408 337482 41409 337546
rect 41343 337481 41409 337482
rect 41346 316087 41406 337481
rect 41535 337102 41601 337103
rect 41535 337038 41536 337102
rect 41600 337038 41601 337102
rect 41535 337037 41601 337038
rect 41538 316827 41598 337037
rect 41730 324967 41790 340811
rect 41727 324966 41793 324967
rect 41727 324902 41728 324966
rect 41792 324902 41793 324966
rect 41727 324901 41793 324902
rect 41535 316826 41601 316827
rect 41535 316762 41536 316826
rect 41600 316762 41601 316826
rect 41535 316761 41601 316762
rect 41343 316086 41409 316087
rect 41343 316022 41344 316086
rect 41408 316022 41409 316086
rect 41343 316021 41409 316022
rect 41151 315494 41217 315495
rect 41151 315430 41152 315494
rect 41216 315430 41217 315494
rect 41151 315429 41217 315430
rect 40959 313274 41025 313275
rect 40959 313210 40960 313274
rect 41024 313210 41025 313274
rect 40959 313209 41025 313210
rect 40575 312386 40641 312387
rect 40575 312322 40576 312386
rect 40640 312322 40641 312386
rect 40575 312321 40641 312322
rect 42114 307171 42174 346355
rect 673986 313571 674046 358053
rect 674175 357082 674241 357083
rect 674175 357018 674176 357082
rect 674240 357018 674241 357082
rect 674175 357017 674241 357018
rect 673983 313570 674049 313571
rect 673983 313506 673984 313570
rect 674048 313506 674049 313570
rect 673983 313505 674049 313506
rect 674178 312535 674238 357017
rect 676095 356194 676161 356195
rect 676095 356130 676096 356194
rect 676160 356130 676161 356194
rect 676095 356129 676161 356130
rect 675903 355602 675969 355603
rect 675903 355538 675904 355602
rect 675968 355538 675969 355602
rect 675903 355537 675969 355538
rect 674559 355010 674625 355011
rect 674559 354946 674560 355010
rect 674624 354946 674625 355010
rect 674559 354945 674625 354946
rect 674562 328371 674622 354945
rect 674943 353530 675009 353531
rect 674943 353466 674944 353530
rect 675008 353466 675009 353530
rect 674943 353465 675009 353466
rect 674751 353086 674817 353087
rect 674751 353022 674752 353086
rect 674816 353022 674817 353086
rect 674751 353021 674817 353022
rect 674559 328370 674625 328371
rect 674559 328306 674560 328370
rect 674624 328306 674625 328370
rect 674559 328305 674625 328306
rect 674754 326891 674814 353021
rect 674946 333551 675006 353465
rect 675519 352050 675585 352051
rect 675519 351986 675520 352050
rect 675584 351986 675585 352050
rect 675519 351985 675585 351986
rect 675135 351162 675201 351163
rect 675135 351098 675136 351162
rect 675200 351098 675201 351162
rect 675135 351097 675201 351098
rect 674943 333550 675009 333551
rect 674943 333486 674944 333550
rect 675008 333486 675009 333550
rect 674943 333485 675009 333486
rect 675138 330591 675198 351097
rect 675522 337103 675582 351985
rect 675711 351532 675777 351533
rect 675711 351468 675712 351532
rect 675776 351468 675777 351532
rect 675711 351467 675777 351468
rect 675519 337102 675585 337103
rect 675519 337038 675520 337102
rect 675584 337038 675585 337102
rect 675519 337037 675585 337038
rect 675714 336511 675774 351467
rect 675906 339619 675966 355537
rect 675903 339618 675969 339619
rect 675903 339554 675904 339618
rect 675968 339554 675969 339618
rect 675903 339553 675969 339554
rect 676098 336990 676158 356129
rect 675906 336930 676158 336990
rect 675711 336510 675777 336511
rect 675711 336446 675712 336510
rect 675776 336446 675777 336510
rect 675711 336445 675777 336446
rect 675135 330590 675201 330591
rect 675135 330526 675136 330590
rect 675200 330526 675201 330590
rect 675135 330525 675201 330526
rect 674751 326890 674817 326891
rect 674751 326826 674752 326890
rect 674816 326826 674817 326890
rect 674751 326825 674817 326826
rect 674367 312682 674433 312683
rect 674367 312618 674368 312682
rect 674432 312618 674433 312682
rect 674367 312617 674433 312618
rect 674175 312534 674241 312535
rect 674175 312470 674176 312534
rect 674240 312470 674241 312534
rect 674175 312469 674241 312470
rect 673983 311794 674049 311795
rect 673983 311730 673984 311794
rect 674048 311730 674049 311794
rect 673983 311729 674049 311730
rect 42114 307111 42532 307171
rect 42472 303631 42532 307111
rect 42114 303571 42532 303631
rect 40575 297882 40641 297883
rect 40575 297818 40576 297882
rect 40640 297818 40641 297882
rect 40575 297817 40641 297818
rect 40383 294330 40449 294331
rect 40383 294266 40384 294330
rect 40448 294266 40449 294330
rect 40383 294265 40449 294266
rect 40386 272871 40446 294265
rect 40383 272870 40449 272871
rect 40383 272806 40384 272870
rect 40448 272806 40449 272870
rect 40383 272805 40449 272806
rect 40578 270503 40638 297817
rect 41727 297660 41793 297661
rect 41727 297596 41728 297660
rect 41792 297596 41793 297660
rect 41727 297595 41793 297596
rect 40767 297290 40833 297291
rect 40767 297226 40768 297290
rect 40832 297226 40833 297290
rect 40767 297225 40833 297226
rect 40575 270502 40641 270503
rect 40575 270438 40576 270502
rect 40640 270438 40641 270502
rect 40575 270437 40641 270438
rect 40770 269171 40830 297225
rect 41151 296550 41217 296551
rect 41151 296486 41152 296550
rect 41216 296486 41217 296550
rect 41151 296485 41217 296486
rect 40959 294922 41025 294923
rect 40959 294858 40960 294922
rect 41024 294858 41025 294922
rect 40959 294857 41025 294858
rect 40962 270059 41022 294857
rect 41154 272427 41214 296485
rect 41535 295810 41601 295811
rect 41535 295746 41536 295810
rect 41600 295746 41601 295810
rect 41535 295745 41601 295746
rect 41343 293886 41409 293887
rect 41343 293822 41344 293886
rect 41408 293822 41409 293886
rect 41343 293821 41409 293822
rect 41346 273611 41406 293821
rect 41538 276571 41598 295745
rect 41730 281751 41790 297595
rect 41727 281750 41793 281751
rect 41727 281686 41728 281750
rect 41792 281686 41793 281750
rect 41727 281685 41793 281686
rect 42114 278643 42174 303571
rect 42111 278642 42177 278643
rect 42111 278578 42112 278642
rect 42176 278578 42177 278642
rect 42111 278577 42177 278578
rect 41535 276570 41601 276571
rect 41535 276506 41536 276570
rect 41600 276506 41601 276570
rect 41535 276505 41601 276506
rect 41343 273610 41409 273611
rect 41343 273546 41344 273610
rect 41408 273546 41409 273610
rect 41343 273545 41409 273546
rect 41151 272426 41217 272427
rect 41151 272362 41152 272426
rect 41216 272362 41217 272426
rect 41151 272361 41217 272362
rect 40959 270058 41025 270059
rect 40959 269994 40960 270058
rect 41024 269994 41025 270058
rect 40959 269993 41025 269994
rect 40767 269170 40833 269171
rect 40767 269106 40768 269170
rect 40832 269106 40833 269170
rect 40767 269105 40833 269106
rect 673986 267543 674046 311729
rect 674175 311054 674241 311055
rect 674175 310990 674176 311054
rect 674240 310990 674241 311054
rect 674175 310989 674241 310990
rect 673983 267542 674049 267543
rect 673983 267478 673984 267542
rect 674048 267478 674049 267542
rect 673983 267477 674049 267478
rect 673983 267098 674049 267099
rect 673983 267034 673984 267098
rect 674048 267034 674049 267098
rect 673983 267033 674049 267034
rect 673986 265027 674046 267033
rect 674178 266507 674238 310989
rect 674370 268579 674430 312617
rect 675906 311573 675966 336930
rect 675903 311572 675969 311573
rect 675903 311508 675904 311572
rect 675968 311508 675969 311572
rect 675903 311507 675969 311508
rect 674559 310018 674625 310019
rect 674559 309954 674560 310018
rect 674624 309954 674625 310018
rect 674559 309953 674625 309954
rect 674562 283675 674622 309953
rect 675327 309130 675393 309131
rect 675327 309066 675328 309130
rect 675392 309066 675393 309130
rect 675327 309065 675393 309066
rect 675135 308538 675201 308539
rect 675135 308474 675136 308538
rect 675200 308474 675201 308538
rect 675135 308473 675201 308474
rect 674751 307798 674817 307799
rect 674751 307734 674752 307798
rect 674816 307734 674817 307798
rect 674751 307733 674817 307734
rect 674559 283674 674625 283675
rect 674559 283610 674560 283674
rect 674624 283610 674625 283674
rect 674559 283609 674625 283610
rect 674754 281899 674814 307733
rect 674943 306170 675009 306171
rect 674943 306106 674944 306170
rect 675008 306106 675009 306170
rect 674943 306105 675009 306106
rect 674946 285303 675006 306105
rect 675138 288559 675198 308473
rect 675330 292851 675390 309065
rect 675519 305578 675585 305579
rect 675519 305514 675520 305578
rect 675584 305514 675585 305578
rect 675519 305513 675585 305514
rect 675327 292850 675393 292851
rect 675327 292786 675328 292850
rect 675392 292786 675393 292850
rect 675327 292785 675393 292786
rect 675135 288558 675201 288559
rect 675135 288494 675136 288558
rect 675200 288494 675201 288558
rect 675135 288493 675201 288494
rect 675522 287375 675582 305513
rect 675711 304616 675777 304617
rect 675711 304552 675712 304616
rect 675776 304552 675777 304616
rect 675711 304551 675777 304552
rect 675714 287819 675774 304551
rect 675711 287818 675777 287819
rect 675711 287754 675712 287818
rect 675776 287754 675777 287818
rect 675711 287753 675777 287754
rect 675519 287374 675585 287375
rect 675519 287310 675520 287374
rect 675584 287310 675585 287374
rect 675519 287309 675585 287310
rect 674943 285302 675009 285303
rect 674943 285238 674944 285302
rect 675008 285238 675009 285302
rect 674943 285237 675009 285238
rect 674751 281898 674817 281899
rect 674751 281834 674752 281898
rect 674816 281834 674817 281898
rect 674751 281833 674817 281834
rect 674367 268578 674433 268579
rect 674367 268514 674368 268578
rect 674432 268514 674433 268578
rect 674367 268513 674433 268514
rect 675519 267986 675585 267987
rect 675519 267922 675520 267986
rect 675584 267922 675585 267986
rect 675519 267921 675585 267922
rect 674175 266506 674241 266507
rect 674175 266442 674176 266506
rect 674240 266442 674241 266506
rect 674175 266441 674241 266442
rect 674175 265766 674241 265767
rect 674175 265702 674176 265766
rect 674240 265702 674241 265766
rect 674175 265701 674241 265702
rect 673983 265026 674049 265027
rect 673983 264962 673984 265026
rect 674048 264962 674049 265026
rect 673983 264961 674049 264962
rect 673983 263546 674049 263547
rect 673983 263482 673984 263546
rect 674048 263482 674049 263546
rect 673983 263481 674049 263482
rect 40575 254666 40641 254667
rect 40575 254602 40576 254666
rect 40640 254602 40641 254666
rect 40575 254601 40641 254602
rect 40578 227435 40638 254601
rect 41727 254518 41793 254519
rect 41727 254454 41728 254518
rect 41792 254454 41793 254518
rect 41727 254453 41793 254454
rect 40959 253334 41025 253335
rect 40959 253270 40960 253334
rect 41024 253270 41025 253334
rect 40959 253269 41025 253270
rect 40767 251706 40833 251707
rect 40767 251642 40768 251706
rect 40832 251642 40833 251706
rect 40767 251641 40833 251642
rect 40575 227434 40641 227435
rect 40575 227370 40576 227434
rect 40640 227370 40641 227434
rect 40575 227369 40641 227370
rect 40770 226843 40830 251641
rect 40962 229063 41022 253269
rect 41535 252594 41601 252595
rect 41535 252530 41536 252594
rect 41600 252530 41601 252594
rect 41535 252529 41601 252530
rect 41151 251114 41217 251115
rect 41151 251050 41152 251114
rect 41216 251050 41217 251114
rect 41151 251049 41217 251050
rect 41343 251114 41409 251115
rect 41343 251050 41344 251114
rect 41408 251050 41409 251114
rect 41343 251049 41409 251050
rect 41154 230395 41214 251049
rect 41151 230394 41217 230395
rect 41151 230330 41152 230394
rect 41216 230330 41217 230394
rect 41151 230329 41217 230330
rect 41346 229803 41406 251049
rect 41538 233355 41598 252529
rect 41730 238387 41790 254453
rect 41919 253926 41985 253927
rect 41919 253862 41920 253926
rect 41984 253862 41985 253926
rect 41919 253861 41985 253862
rect 41727 238386 41793 238387
rect 41727 238322 41728 238386
rect 41792 238322 41793 238386
rect 41727 238321 41793 238322
rect 41535 233354 41601 233355
rect 41535 233290 41536 233354
rect 41600 233290 41601 233354
rect 41535 233289 41601 233290
rect 41343 229802 41409 229803
rect 41343 229738 41344 229802
rect 41408 229738 41409 229802
rect 41343 229737 41409 229738
rect 40959 229062 41025 229063
rect 40959 228998 40960 229062
rect 41024 228998 41025 229062
rect 40959 228997 41025 228998
rect 40767 226842 40833 226843
rect 40767 226778 40768 226842
rect 40832 226778 40833 226842
rect 40767 226777 40833 226778
rect 41922 226251 41982 253861
rect 673986 243567 674046 263481
rect 673983 243566 674049 243567
rect 673983 243502 673984 243566
rect 674048 243502 674049 243566
rect 673983 243501 674049 243502
rect 148329 243418 148395 243419
rect 148329 243354 148330 243418
rect 148394 243354 148395 243418
rect 148329 243353 148395 243354
rect 41919 226250 41985 226251
rect 41919 226186 41920 226250
rect 41984 226186 41985 226250
rect 41919 226185 41985 226186
rect 40575 211450 40641 211451
rect 40575 211386 40576 211450
rect 40640 211386 40641 211450
rect 40575 211385 40641 211386
rect 40383 211006 40449 211007
rect 40383 210942 40384 211006
rect 40448 210942 40449 211006
rect 40383 210941 40449 210942
rect 40386 195171 40446 210941
rect 40383 195170 40449 195171
rect 40383 195106 40384 195170
rect 40448 195106 40449 195170
rect 40383 195105 40449 195106
rect 40578 184071 40638 211385
rect 41727 210710 41793 210711
rect 41727 210646 41728 210710
rect 41792 210646 41793 210710
rect 41727 210645 41793 210646
rect 41151 209970 41217 209971
rect 41151 209906 41152 209970
rect 41216 209906 41217 209970
rect 41151 209905 41217 209906
rect 40767 208490 40833 208491
rect 40767 208426 40768 208490
rect 40832 208426 40833 208490
rect 40767 208425 40833 208426
rect 40575 184070 40641 184071
rect 40575 184006 40576 184070
rect 40640 184006 40641 184070
rect 40575 184005 40641 184006
rect 40770 183627 40830 208425
rect 40959 207898 41025 207899
rect 40959 207834 40960 207898
rect 41024 207834 41025 207898
rect 40959 207833 41025 207834
rect 40962 187179 41022 207833
rect 40959 187178 41025 187179
rect 40959 187114 40960 187178
rect 41024 187114 41025 187178
rect 40959 187113 41025 187114
rect 41154 185847 41214 209905
rect 41535 209526 41601 209527
rect 41535 209462 41536 209526
rect 41600 209462 41601 209526
rect 41535 209461 41601 209462
rect 41343 207898 41409 207899
rect 41343 207834 41344 207898
rect 41408 207834 41409 207898
rect 41343 207833 41409 207834
rect 41346 186735 41406 207833
rect 41538 190139 41598 209461
rect 41535 190138 41601 190139
rect 41535 190074 41536 190138
rect 41600 190074 41601 190138
rect 41535 190073 41601 190074
rect 41343 186734 41409 186735
rect 41343 186670 41344 186734
rect 41408 186670 41409 186734
rect 41343 186669 41409 186670
rect 41151 185846 41217 185847
rect 41151 185782 41152 185846
rect 41216 185782 41217 185846
rect 41151 185781 41217 185782
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 41730 183035 41790 210645
rect 41727 183034 41793 183035
rect 41727 182970 41728 183034
rect 41792 182970 41793 183034
rect 41727 182969 41793 182970
rect 148332 171787 148392 243353
rect 674178 232438 674238 265701
rect 674367 265026 674433 265027
rect 674367 264962 674368 265026
rect 674432 264962 674433 265026
rect 674367 264961 674433 264962
rect 674559 265026 674625 265027
rect 674559 264962 674560 265026
rect 674624 264962 674625 265026
rect 674559 264961 674625 264962
rect 674370 232696 674430 264961
rect 674562 238239 674622 264961
rect 674751 262806 674817 262807
rect 674751 262742 674752 262806
rect 674816 262742 674817 262806
rect 674751 262741 674817 262742
rect 674559 238238 674625 238239
rect 674559 238174 674560 238238
rect 674624 238174 674625 238238
rect 674559 238173 674625 238174
rect 674754 236907 674814 262741
rect 674943 261178 675009 261179
rect 674943 261114 674944 261178
rect 675008 261114 675009 261178
rect 674943 261113 675009 261114
rect 674946 240607 675006 261113
rect 675135 260586 675201 260587
rect 675135 260522 675136 260586
rect 675200 260522 675201 260586
rect 675135 260521 675201 260522
rect 675138 241939 675198 260521
rect 675135 241938 675201 241939
rect 675135 241874 675136 241938
rect 675200 241874 675201 241938
rect 675135 241873 675201 241874
rect 674943 240606 675009 240607
rect 674943 240542 674944 240606
rect 675008 240542 675009 240606
rect 674943 240541 675009 240542
rect 674751 236906 674817 236907
rect 674751 236842 674752 236906
rect 674816 236842 674817 236906
rect 674751 236841 674817 236842
rect 674370 232636 674873 232696
rect 674178 232378 674692 232438
rect 674632 224573 674692 232378
rect 674178 224513 674692 224573
rect 673983 221958 674049 221959
rect 673983 221894 673984 221958
rect 674048 221894 674049 221958
rect 673983 221893 674049 221894
rect 673986 186751 674046 221893
rect 674178 221367 674238 224513
rect 674813 224220 674873 232636
rect 675522 231587 675582 267921
rect 675903 265618 675969 265619
rect 675903 265554 675904 265618
rect 675968 265554 675969 265618
rect 675903 265553 675969 265554
rect 675711 264138 675777 264139
rect 675711 264074 675712 264138
rect 675776 264074 675777 264138
rect 675711 264073 675777 264074
rect 675714 247563 675774 264073
rect 675906 249635 675966 265553
rect 676287 261326 676353 261327
rect 676287 261262 676288 261326
rect 676352 261262 676353 261326
rect 676287 261261 676353 261262
rect 676095 259846 676161 259847
rect 676095 259782 676096 259846
rect 676160 259782 676161 259846
rect 676095 259781 676161 259782
rect 675903 249634 675969 249635
rect 675903 249570 675904 249634
rect 675968 249570 675969 249634
rect 675903 249569 675969 249570
rect 675711 247562 675777 247563
rect 675711 247498 675712 247562
rect 675776 247498 675777 247562
rect 675711 247497 675777 247498
rect 676098 245935 676158 259781
rect 676290 246675 676350 261261
rect 676287 246674 676353 246675
rect 676287 246610 676288 246674
rect 676352 246610 676353 246674
rect 676287 246609 676353 246610
rect 676095 245934 676161 245935
rect 676095 245870 676096 245934
rect 676160 245870 676161 245934
rect 676095 245869 676161 245870
rect 675522 231527 676101 231587
rect 676041 225728 676101 231527
rect 674370 224160 674873 224220
rect 675522 225668 676101 225728
rect 674370 222699 674430 224160
rect 675522 223439 675582 225668
rect 675519 223438 675585 223439
rect 675519 223374 675520 223438
rect 675584 223374 675585 223438
rect 675519 223373 675585 223374
rect 675903 222846 675969 222847
rect 675903 222782 675904 222846
rect 675968 222782 675969 222846
rect 675903 222781 675969 222782
rect 674367 222698 674433 222699
rect 674367 222634 674368 222698
rect 674432 222634 674433 222698
rect 674367 222633 674433 222634
rect 674175 221366 674241 221367
rect 674175 221302 674176 221366
rect 674240 221302 674241 221366
rect 674175 221301 674241 221302
rect 674175 220774 674241 220775
rect 674175 220710 674176 220774
rect 674240 220710 674241 220774
rect 674175 220709 674241 220710
rect 674178 218999 674238 220709
rect 675519 220034 675585 220035
rect 675519 219970 675520 220034
rect 675584 219970 675585 220034
rect 675519 219969 675585 219970
rect 674751 219886 674817 219887
rect 674751 219822 674752 219886
rect 674816 219822 674817 219886
rect 674751 219821 674817 219822
rect 674175 218998 674241 218999
rect 674175 218934 674176 218998
rect 674240 218934 674241 218998
rect 674175 218933 674241 218934
rect 673187 186691 674046 186751
rect 673187 180293 673247 186691
rect 674178 186548 674238 218933
rect 674559 217814 674625 217815
rect 674559 217750 674560 217814
rect 674624 217750 674625 217814
rect 674559 217749 674625 217750
rect 674562 191619 674622 217749
rect 674754 193543 674814 219821
rect 675135 218406 675201 218407
rect 675135 218342 675136 218406
rect 675200 218342 675201 218406
rect 675135 218341 675201 218342
rect 674943 215890 675009 215891
rect 674943 215826 674944 215890
rect 675008 215826 675009 215890
rect 674943 215825 675009 215826
rect 674946 195319 675006 215825
rect 675138 198427 675198 218341
rect 675522 204347 675582 219969
rect 675711 216334 675777 216335
rect 675711 216270 675712 216334
rect 675776 216270 675777 216334
rect 675711 216269 675777 216270
rect 675519 204346 675585 204347
rect 675519 204282 675520 204346
rect 675584 204282 675585 204346
rect 675519 204281 675585 204282
rect 675714 201387 675774 216269
rect 675711 201386 675777 201387
rect 675711 201322 675712 201386
rect 675776 201322 675777 201386
rect 675711 201321 675777 201322
rect 675135 198426 675201 198427
rect 675135 198362 675136 198426
rect 675200 198362 675201 198426
rect 675135 198361 675201 198362
rect 674943 195318 675009 195319
rect 674943 195254 674944 195318
rect 675008 195254 675009 195318
rect 674943 195253 675009 195254
rect 674751 193542 674817 193543
rect 674751 193478 674752 193542
rect 674816 193478 674817 193542
rect 674751 193477 674817 193478
rect 674559 191618 674625 191619
rect 674559 191554 674560 191618
rect 674624 191554 674625 191618
rect 674559 191553 674625 191554
rect 673356 186488 674238 186548
rect 673356 180531 673416 186488
rect 673356 180471 674238 180531
rect 673187 180233 674046 180293
rect 673986 177263 674046 180233
rect 673983 177262 674049 177263
rect 673983 177198 673984 177262
rect 674048 177198 674049 177262
rect 673983 177197 674049 177198
rect 674178 176375 674238 180471
rect 675906 178447 675966 222781
rect 676287 218702 676353 218703
rect 676287 218638 676288 218702
rect 676352 218638 676353 218702
rect 676287 218637 676353 218638
rect 676095 217074 676161 217075
rect 676095 217010 676096 217074
rect 676160 217010 676161 217074
rect 676095 217009 676161 217010
rect 676098 205087 676158 217009
rect 676095 205086 676161 205087
rect 676095 205022 676096 205086
rect 676160 205022 676161 205086
rect 676095 205021 676161 205022
rect 676290 202719 676350 218637
rect 676287 202718 676353 202719
rect 676287 202654 676288 202718
rect 676352 202654 676353 202718
rect 676287 202653 676353 202654
rect 675903 178446 675969 178447
rect 675903 178382 675904 178446
rect 675968 178382 675969 178446
rect 675903 178381 675969 178382
rect 674367 177854 674433 177855
rect 674367 177790 674368 177854
rect 674432 177790 674433 177854
rect 674367 177789 674433 177790
rect 674175 176374 674241 176375
rect 674175 176310 674176 176374
rect 674240 176310 674241 176374
rect 674175 176309 674241 176310
rect 674175 175782 674241 175783
rect 674175 175718 674176 175782
rect 674240 175718 674241 175782
rect 674175 175717 674241 175718
rect 148329 171786 148395 171787
rect 148329 171722 148330 171786
rect 148394 171722 148395 171786
rect 148329 171721 148395 171722
rect 673983 170898 674049 170899
rect 673983 170834 673984 170898
rect 674048 170834 674049 170898
rect 673983 170833 674049 170834
rect 148287 152842 148353 152843
rect 148287 152778 148288 152842
rect 148352 152778 148353 152842
rect 148287 152777 148353 152778
rect 148290 109331 148350 152777
rect 673986 150327 674046 170833
rect 673983 150326 674049 150327
rect 673983 150262 673984 150326
rect 674048 150262 674049 150326
rect 673983 150261 674049 150262
rect 674178 143082 674238 175717
rect 673178 143022 674238 143082
rect 673178 131235 673238 143022
rect 674370 142718 674430 177789
rect 675519 176966 675585 176967
rect 675519 176902 675520 176966
rect 675584 176902 675585 176966
rect 675519 176901 675585 176902
rect 675522 175931 675582 176901
rect 675519 175930 675585 175931
rect 675519 175866 675520 175930
rect 675584 175866 675585 175930
rect 675519 175865 675585 175866
rect 674751 174894 674817 174895
rect 674751 174830 674752 174894
rect 674816 174830 674817 174894
rect 674751 174829 674817 174830
rect 674559 172822 674625 172823
rect 674559 172758 674560 172822
rect 674624 172758 674625 172822
rect 674559 172757 674625 172758
rect 674562 146627 674622 172757
rect 674754 148551 674814 174829
rect 674943 173414 675009 173415
rect 674943 173350 674944 173414
rect 675008 173350 675009 173414
rect 674943 173349 675009 173350
rect 674946 153435 675006 173349
rect 675135 170010 675201 170011
rect 675135 169946 675136 170010
rect 675200 169946 675201 170010
rect 675135 169945 675201 169946
rect 674943 153434 675009 153435
rect 674943 153370 674944 153434
rect 675008 153370 675009 153434
rect 674943 153369 675009 153370
rect 675138 151955 675198 169945
rect 675327 169418 675393 169419
rect 675327 169354 675328 169418
rect 675392 169354 675393 169418
rect 675327 169353 675393 169354
rect 675330 152547 675390 169353
rect 675327 152546 675393 152547
rect 675327 152482 675328 152546
rect 675392 152482 675393 152546
rect 675327 152481 675393 152482
rect 675135 151954 675201 151955
rect 675135 151890 675136 151954
rect 675200 151890 675201 151954
rect 675135 151889 675201 151890
rect 674751 148550 674817 148551
rect 674751 148486 674752 148550
rect 674816 148486 674817 148550
rect 674751 148485 674817 148486
rect 674559 146626 674625 146627
rect 674559 146562 674560 146626
rect 674624 146562 674625 146626
rect 674559 146561 674625 146562
rect 673370 142658 674430 142718
rect 673370 133159 673430 142658
rect 675522 142115 675582 175865
rect 675711 168826 675777 168827
rect 675711 168762 675712 168826
rect 675776 168762 675777 168826
rect 675711 168761 675777 168762
rect 675714 151363 675774 168761
rect 675711 151362 675777 151363
rect 675711 151298 675712 151362
rect 675776 151298 675777 151362
rect 675711 151297 675777 151298
rect 674522 142055 675582 142115
rect 673367 133158 673433 133159
rect 673367 133094 673368 133158
rect 673432 133094 673433 133158
rect 673367 133093 673433 133094
rect 674522 132123 674582 142055
rect 674519 132122 674585 132123
rect 674519 132058 674520 132122
rect 674584 132058 674585 132122
rect 674519 132057 674585 132058
rect 673175 131234 673241 131235
rect 673175 131170 673176 131234
rect 673240 131170 673241 131234
rect 673175 131169 673241 131170
rect 674943 130198 675009 130199
rect 674943 130134 674944 130198
rect 675008 130134 675009 130198
rect 674943 130133 675009 130134
rect 674367 128126 674433 128127
rect 674367 128062 674368 128126
rect 674432 128062 674433 128126
rect 674367 128061 674433 128062
rect 148287 109330 148353 109331
rect 148287 109266 148288 109330
rect 148352 109266 148353 109330
rect 148287 109265 148353 109266
rect 674370 108147 674430 128061
rect 674559 125758 674625 125759
rect 674559 125694 674560 125758
rect 674624 125694 674625 125758
rect 674559 125693 674625 125694
rect 674367 108146 674433 108147
rect 674367 108082 674368 108146
rect 674432 108082 674433 108146
rect 674367 108081 674433 108082
rect 674562 105187 674622 125693
rect 674751 125166 674817 125167
rect 674751 125102 674752 125166
rect 674816 125102 674817 125166
rect 674751 125101 674817 125102
rect 674754 106371 674814 125101
rect 674946 114363 675006 130133
rect 675711 129680 675777 129681
rect 675711 129616 675712 129680
rect 675776 129616 675777 129680
rect 675711 129615 675777 129616
rect 675135 128718 675201 128719
rect 675135 128654 675136 128718
rect 675200 128654 675201 128718
rect 675135 128653 675201 128654
rect 674943 114362 675009 114363
rect 674943 114298 674944 114362
rect 675008 114298 675009 114362
rect 674943 114297 675009 114298
rect 675138 112291 675198 128653
rect 675327 127682 675393 127683
rect 675327 127618 675328 127682
rect 675392 127618 675393 127682
rect 675327 127617 675393 127618
rect 675135 112290 675201 112291
rect 675135 112226 675136 112290
rect 675200 112226 675201 112290
rect 675135 112225 675201 112226
rect 674751 106370 674817 106371
rect 674751 106306 674752 106370
rect 674816 106306 674817 106370
rect 674751 106305 674817 106306
rect 674559 105186 674625 105187
rect 674559 105122 674560 105186
rect 674624 105122 674625 105186
rect 674559 105121 674625 105122
rect 675330 101487 675390 127617
rect 675714 103263 675774 129615
rect 675711 103262 675777 103263
rect 675711 103198 675712 103262
rect 675776 103198 675777 103262
rect 675711 103197 675777 103198
rect 675327 101486 675393 101487
rect 675327 101422 675328 101486
rect 675392 101422 675393 101486
rect 675327 101421 675393 101422
rect 518847 41242 518913 41243
rect 518847 41178 518848 41242
rect 518912 41178 518913 41242
rect 518847 41177 518913 41178
rect 518850 40411 518910 41177
rect 568550 40510 568616 40511
rect 568550 40446 568551 40510
rect 568615 40508 568616 40510
rect 584555 40510 584621 40511
rect 584555 40508 584556 40510
rect 568615 40448 584556 40508
rect 568615 40446 568616 40448
rect 568550 40445 568616 40446
rect 584555 40446 584556 40448
rect 584620 40446 584621 40510
rect 584555 40445 584621 40446
rect 240566 40248 240632 40249
rect 240566 40184 240567 40248
rect 240631 40246 240632 40248
rect 257339 40248 257405 40249
rect 257339 40246 257340 40248
rect 240631 40186 257340 40246
rect 240631 40184 240632 40186
rect 240566 40183 240632 40184
rect 257339 40184 257340 40186
rect 257404 40184 257405 40248
rect 257339 40183 257405 40184
rect 507135 40150 507136 40175
rect 507200 40150 507201 40175
rect 507135 40149 507201 40150
<< via4 >>
rect 507050 40214 507286 40411
rect 507050 40175 507136 40214
rect 507136 40175 507200 40214
rect 507200 40175 507286 40214
rect 518762 40175 518998 40411
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 442854 19619 453734
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 182580 262883 187699 264182
rect 180738 260392 185857 261691
rect 180753 257779 185872 259078
rect 181613 255363 186732 256662
rect 414961 252857 419536 254186
rect 415323 250350 419898 251679
rect 415550 247873 420125 249202
rect 415867 245352 420442 246681
rect 184415 242851 188990 244180
rect 415565 240323 420140 241652
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 667620 66907 669733 74575
rect 671454 66982 673567 74650
rect 507008 40411 519040 40453
rect 507008 40175 507050 40411
rect 507286 40175 518762 40411
rect 518998 40175 519040 40411
rect 507008 40133 519040 40175
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use mgmt_core  soc ~/gits/caravel/maglef
timestamp 1624566096
transform 1 0 190434 0 1 53602
box 0 0 450000 168026
use storage  storage ~/gits/caravel/maglef
timestamp 1624446576
transform 1 0 52032 0 1 53156
box 1066 70 92000 191480
use gpio_control_block  gpio_control_bidir_1\[0\] ~/gits/caravel/maglef
timestamp 1624273664
transform -1 0 710203 0 1 121000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1624273664
transform -1 0 710203 0 1 166200
box -1620 -364 34000 13964
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level ~/gits/caravel/maglef
timestamp 1608587524
transform -1 0 145710 0 -1 50488
box 480 -400 3456 3800
use user_id_programming  user_id_value ~/gits/caravel/maglef
timestamp 1607107372
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use simple_por  por ~/gits/caravel/maglef
timestamp 1606790297
transform 1 0 654146 0 -1 112882
box 25 11 11344 8291
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1624273664
transform 1 0 7631 0 1 202600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1624273664
transform 1 0 7631 0 1 245800
box -1620 -364 34000 13964
use mgmt_protect  mgmt_buffers ~/gits/caravel/maglef
timestamp 1624984707
transform 1 0 192180 0 1 240036
box -2762 -2778 222734 26170
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1624273664
transform -1 0 710203 0 1 256400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1624273664
transform -1 0 710203 0 1 211200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[16\]
timestamp 1624273664
transform 1 0 7631 0 1 289000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1624273664
transform 1 0 7631 0 1 332200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1624273664
transform 1 0 7631 0 1 375400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1624273664
transform -1 0 710203 0 1 346400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1624273664
transform -1 0 710203 0 1 301400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1624273664
transform -1 0 710203 0 1 391600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1624273664
transform -1 0 710203 0 1 479800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1624273664
transform 1 0 7631 0 1 418600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1624273664
transform 1 0 7631 0 1 632600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1624273664
transform 1 0 7631 0 1 589400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1624273664
transform 1 0 7631 0 1 546200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1624273664
transform -1 0 710203 0 1 523800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1624273664
transform -1 0 710203 0 1 568800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1624273664
transform -1 0 710203 0 1 614000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1624273664
transform 1 0 7631 0 1 762200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1624273664
transform 1 0 7631 0 1 719000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1624273664
transform 1 0 7631 0 1 675800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1624273664
transform -1 0 710203 0 1 704200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[11\]
timestamp 1624273664
transform -1 0 710203 0 1 749200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1624273664
transform -1 0 710203 0 1 659000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1624273664
transform 1 0 7631 0 1 805400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1624273664
transform 0 1 97200 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1624273664
transform 1 0 7631 0 1 931224
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1624273664
transform 0 1 200000 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1624273664
transform 0 1 148600 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[16\]
timestamp 1624273664
transform 0 1 353400 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1624273664
transform 0 1 303000 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1624273664
transform 0 1 251400 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[14\]
timestamp 1624273664
transform 0 1 497800 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[15\]
timestamp 1624273664
transform 0 1 420800 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[13\]
timestamp 1624273664
transform 0 1 549200 -1 0 1030077
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[12\]
timestamp 1624273664
transform -1 0 710203 0 1 927600
box -1620 -364 34000 13964
use user_project_wrapper  mprj
timestamp 1624557694
transform 1 0 65308 0 1 278718
box -8576 -7506 592500 711442
use chip_io  padframe
timestamp 1624978002
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use caravel_power_routing  caravel_power_routing_0
timestamp 1625001417
transform 1 0 38561 0 1 38708
box -33118 599 673272 993231
<< labels >>
flabel metal5 s 187640 6598 200180 19088 0 FreeSans 16000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363580 19088 0 FreeSans 16000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308780 19088 0 FreeSans 16000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418380 19088 0 FreeSans 16000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473180 19088 0 FreeSans 16000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527980 19088 0 FreeSans 16000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113780 0 FreeSans 16000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696980 0 FreeSans 16000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741980 0 FreeSans 16000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786980 0 FreeSans 16000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876180 0 FreeSans 16000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965380 0 FreeSans 16000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628220 1018512 640760 1031002 0 FreeSans 16000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526420 1018512 538960 1031002 0 FreeSans 16000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475020 1018512 487560 1031002 0 FreeSans 16000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386020 1018512 398560 1031002 0 FreeSans 16000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284220 1018512 296760 1031002 0 FreeSans 16000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158980 0 FreeSans 16000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 232620 1018512 245160 1031002 0 FreeSans 16000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181220 1018512 193760 1031002 0 FreeSans 16000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 129820 1018512 142360 1031002 0 FreeSans 16000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78420 1018512 90960 1031002 0 FreeSans 16000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6598 956420 19088 968960 0 FreeSans 16000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786620 19088 799160 0 FreeSans 16000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743420 19088 755960 0 FreeSans 16000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700220 19088 712760 0 FreeSans 16000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657020 19088 669560 0 FreeSans 16000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613820 19088 626360 0 FreeSans 16000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203980 0 FreeSans 16000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570620 19088 583160 0 FreeSans 16000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527420 19088 539960 0 FreeSans 16000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399820 19088 412360 0 FreeSans 16000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356620 19088 369160 0 FreeSans 16000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313420 19088 325960 0 FreeSans 16000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270220 19088 282760 0 FreeSans 16000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227020 19088 239560 0 FreeSans 16000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183820 19088 196360 0 FreeSans 16000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249180 0 FreeSans 16000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294180 0 FreeSans 16000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339180 0 FreeSans 16000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384380 0 FreeSans 16000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561580 0 FreeSans 16000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606780 0 FreeSans 16000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651780 0 FreeSans 16000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 16000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 16000 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 16000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 16000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 16000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 16000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 16000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 16000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 16000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 16000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 16000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 16000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 16000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 16000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 16000 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 16000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 16000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 16000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 16000 0 0 0 vssio_2
port 62 nsew signal bidirectional
flabel metal2 s 579796 53602 579852 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[0]
port 63 nsew signal tristate
flabel metal2 s 597092 53602 597148 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[1]
port 64 nsew signal tristate
flabel metal2 s 614388 53602 614444 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[2]
port 65 nsew signal tristate
flabel metal2 s 631684 53602 631740 54402 0 FreeSans 16000 0 0 0 pwr_ctrl_out[3]
port 66 nsew signal tristate
flabel metal5 184920 263575 184920 263575 0 FreeSans 8000 0 0 0 vccd2_core
flabel metal5 182956 261182 182956 261182 0 FreeSans 8000 0 0 0 vssd2_core
flabel metal5 183201 258482 183201 258482 0 FreeSans 8000 0 0 0 vdda2_core
flabel metal5 183999 256028 183999 256028 0 FreeSans 8000 0 0 0 vssa2_core
flabel metal5 186454 243448 186454 243448 0 FreeSans 8000 0 0 0 vccd_core
flabel metal5 417916 240932 417916 240932 0 FreeSans 8000 0 0 0 vssd_core
flabel metal5 418100 245964 418100 245964 0 FreeSans 8000 0 0 0 vssa1_core
flabel metal5 417793 248603 417793 248603 0 FreeSans 8000 0 0 0 vdda1_core
flabel metal5 417486 250996 417486 250996 0 FreeSans 8000 0 0 0 vssd1_core
flabel metal5 417118 253512 417118 253512 0 FreeSans 8000 0 0 0 vccd1_core
flabel metal5 668612 70870 668612 70870 0 FreeSans 8000 90 0 0 vddio_core
flabel metal5 672443 71154 672443 71154 0 FreeSans 8000 90 0 0 vssio_core
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
