VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_io
  CLASS BLOCK ;
  FOREIGN chip_io ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 938.200 32.990 1000.900 95.440 ;
    END
  END clock
  PIN clock_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.635 208.565 936.915 210.965 ;
    END
  END clock_core
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.215 208.565 970.495 210.965 ;
    END
  END por
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1755.200 32.990 1817.900 95.440 ;
    END
  END flash_clk
  PIN flash_clk_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.835 208.565 1809.115 210.965 ;
    END
  END flash_clk_core
  PIN flash_clk_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.215 208.565 1787.495 210.965 ;
    END
  END flash_clk_ieb_core
  PIN flash_clk_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.475 208.565 1824.755 210.965 ;
    END
  END flash_clk_oeb_core
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1481.200 32.990 1543.900 95.440 ;
    END
  END flash_csb
  PIN flash_csb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.835 208.565 1535.115 210.965 ;
    END
  END flash_csb_core
  PIN flash_csb_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.215 208.565 1513.495 210.965 ;
    END
  END flash_csb_ieb_core
  PIN flash_csb_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.475 208.565 1550.755 210.965 ;
    END
  END flash_csb_oeb_core
  PIN flash_io0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2029.200 32.990 2091.900 95.440 ;
    END
  END flash_io0
  PIN flash_io0_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.635 208.565 2027.915 210.965 ;
    END
  END flash_io0_di_core
  PIN flash_io0_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.835 208.565 2083.115 210.965 ;
    END
  END flash_io0_do_core
  PIN flash_io0_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2046.150 220.900 2046.470 220.960 ;
        RECT 2061.330 220.900 2061.650 220.960 ;
        RECT 2076.970 220.900 2077.290 220.960 ;
        RECT 2046.150 220.760 2077.290 220.900 ;
        RECT 2046.150 220.700 2046.470 220.760 ;
        RECT 2061.330 220.700 2061.650 220.760 ;
        RECT 2076.970 220.700 2077.290 220.760 ;
      LAYER via ;
        RECT 2046.180 220.700 2046.440 220.960 ;
        RECT 2061.360 220.700 2061.620 220.960 ;
        RECT 2077.000 220.700 2077.260 220.960 ;
      LAYER met2 ;
        RECT 2046.180 220.670 2046.440 220.990 ;
        RECT 2061.360 220.670 2061.620 220.990 ;
        RECT 2077.000 220.670 2077.260 220.990 ;
        RECT 2046.240 210.965 2046.380 220.670 ;
        RECT 2061.420 210.965 2061.560 220.670 ;
        RECT 2077.060 210.965 2077.200 220.670 ;
        RECT 2046.035 209.100 2046.380 210.965 ;
        RECT 2061.215 209.100 2061.560 210.965 ;
        RECT 2076.855 209.100 2077.200 210.965 ;
        RECT 2046.035 208.565 2046.315 209.100 ;
        RECT 2061.215 208.565 2061.495 209.100 ;
        RECT 2076.855 208.565 2077.135 209.100 ;
    END
  END flash_io0_ieb_core
  PIN flash_io0_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2055.350 223.280 2055.670 223.340 ;
        RECT 2098.590 223.280 2098.910 223.340 ;
        RECT 2055.350 223.140 2098.910 223.280 ;
        RECT 2055.350 223.080 2055.670 223.140 ;
        RECT 2098.590 223.080 2098.910 223.140 ;
      LAYER via ;
        RECT 2055.380 223.080 2055.640 223.340 ;
        RECT 2098.620 223.080 2098.880 223.340 ;
      LAYER met2 ;
        RECT 2055.380 223.050 2055.640 223.370 ;
        RECT 2098.620 223.050 2098.880 223.370 ;
        RECT 2055.440 210.965 2055.580 223.050 ;
        RECT 2098.680 210.965 2098.820 223.050 ;
        RECT 2055.235 209.100 2055.580 210.965 ;
        RECT 2098.475 209.100 2098.820 210.965 ;
        RECT 2055.235 208.565 2055.515 209.100 ;
        RECT 2098.475 208.565 2098.755 209.100 ;
    END
  END flash_io0_oeb_core
  PIN flash_io1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2303.200 32.990 2365.900 95.440 ;
    END
  END flash_io1
  PIN flash_io1_di_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.635 208.565 2301.915 210.965 ;
    END
  END flash_io1_di_core
  PIN flash_io1_do_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.835 208.565 2357.115 210.965 ;
    END
  END flash_io1_do_core
  PIN flash_io1_ieb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2320.770 209.340 2321.090 209.400 ;
        RECT 2335.950 209.340 2336.270 209.400 ;
        RECT 2350.210 209.340 2350.530 209.400 ;
        RECT 2320.770 209.200 2350.530 209.340 ;
        RECT 2320.770 209.140 2321.090 209.200 ;
        RECT 2335.950 209.140 2336.270 209.200 ;
        RECT 2350.210 209.140 2350.530 209.200 ;
      LAYER via ;
        RECT 2320.800 209.140 2321.060 209.400 ;
        RECT 2335.980 209.140 2336.240 209.400 ;
        RECT 2350.240 209.140 2350.500 209.400 ;
      LAYER met2 ;
        RECT 2320.035 209.170 2320.315 210.965 ;
        RECT 2320.800 209.170 2321.060 209.430 ;
        RECT 2320.035 209.110 2321.060 209.170 ;
        RECT 2335.215 209.170 2335.495 210.965 ;
        RECT 2335.980 209.170 2336.240 209.430 ;
        RECT 2335.215 209.110 2336.240 209.170 ;
        RECT 2350.240 209.170 2350.500 209.430 ;
        RECT 2350.855 209.170 2351.135 210.965 ;
        RECT 2350.240 209.110 2351.135 209.170 ;
        RECT 2320.035 209.030 2321.000 209.110 ;
        RECT 2335.215 209.030 2336.180 209.110 ;
        RECT 2350.300 209.030 2351.135 209.110 ;
        RECT 2320.035 208.565 2320.315 209.030 ;
        RECT 2335.215 208.565 2335.495 209.030 ;
        RECT 2350.855 208.565 2351.135 209.030 ;
    END
  END flash_io1_ieb_core
  PIN flash_io1_oeb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2329.050 221.580 2329.370 221.640 ;
        RECT 2372.290 221.580 2372.610 221.640 ;
        RECT 2329.050 221.440 2372.610 221.580 ;
        RECT 2329.050 221.380 2329.370 221.440 ;
        RECT 2372.290 221.380 2372.610 221.440 ;
      LAYER via ;
        RECT 2329.080 221.380 2329.340 221.640 ;
        RECT 2372.320 221.380 2372.580 221.640 ;
      LAYER met2 ;
        RECT 2329.080 221.350 2329.340 221.670 ;
        RECT 2372.320 221.350 2372.580 221.670 ;
        RECT 2329.140 210.965 2329.280 221.350 ;
        RECT 2372.380 210.965 2372.520 221.350 ;
        RECT 2329.140 209.030 2329.515 210.965 ;
        RECT 2372.380 209.030 2372.755 210.965 ;
        RECT 2329.235 208.565 2329.515 209.030 ;
        RECT 2372.475 208.565 2372.755 209.030 ;
    END
  END flash_io1_oeb_core
  PIN gpio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2577.200 32.990 2639.900 95.440 ;
    END
  END gpio
  PIN gpio_in_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.635 208.565 2575.915 210.965 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.215 208.565 2609.495 210.965 ;
    END
  END gpio_inenb_core
  PIN gpio_mode0_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.235 208.565 2603.515 210.965 ;
    END
  END gpio_mode0_core
  PIN gpio_mode1_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2594.010 220.900 2594.330 220.960 ;
        RECT 2624.830 220.900 2625.150 220.960 ;
        RECT 2594.010 220.760 2625.150 220.900 ;
        RECT 2594.010 220.700 2594.330 220.760 ;
        RECT 2624.830 220.700 2625.150 220.760 ;
      LAYER via ;
        RECT 2594.040 220.700 2594.300 220.960 ;
        RECT 2624.860 220.700 2625.120 220.960 ;
      LAYER met2 ;
        RECT 2594.040 220.670 2594.300 220.990 ;
        RECT 2624.860 220.670 2625.120 220.990 ;
        RECT 2594.100 210.965 2594.240 220.670 ;
        RECT 2624.920 210.965 2625.060 220.670 ;
        RECT 2594.035 208.565 2594.315 210.965 ;
        RECT 2624.855 208.565 2625.135 210.965 ;
    END
  END gpio_mode1_core
  PIN gpio_out_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.835 208.565 2631.115 210.965 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.475 208.565 2646.755 210.965 ;
    END
  END gpio_outenb_core
  PIN vccd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 350.270 98.100 404.670 ;
    END
  END vccd_pad
  PIN vdda_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3121.110 34.055 3181.950 94.880 ;
    END
  END vdda_pad
  PIN vddio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 558.050 94.880 618.890 ;
    END
  END vddio_pad
  PIN vddio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4356.050 94.880 4416.890 ;
    END
  END vddio_pad2
  PIN vssa_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 401.110 34.055 461.950 94.880 ;
    END
  END vssa_pad
  PIN vssd_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1216.330 30.835 1270.730 98.100 ;
    END
  END vssd_pad
  PIN vssio_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2852.110 34.055 2912.950 94.880 ;
    END
  END vssio_pad
  PIN vssio_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1674.050 5093.120 1734.890 5153.945 ;
    END
  END vssio_pad2
  PIN mprj_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 506.200 3555.010 568.900 ;
    END
  END mprj_io[0]
  PIN mprj_io_analog_en[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 529.015 3379.435 529.295 ;
    END
  END mprj_io_analog_en[0]
  PIN mprj_io_analog_pol[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 535.455 3379.435 535.735 ;
    END
  END mprj_io_analog_pol[0]
  PIN mprj_io_analog_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 550.635 3379.435 550.915 ;
    END
  END mprj_io_analog_sel[0]
  PIN mprj_io_dm[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 532.235 3379.435 532.515 ;
    END
  END mprj_io_dm[0]
  PIN mprj_io_dm[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 523.035 3379.435 523.315 ;
    END
  END mprj_io_dm[1]
  PIN mprj_io_dm[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 553.855 3379.435 554.135 ;
    END
  END mprj_io_dm[2]
  PIN mprj_io_holdover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 557.075 3379.435 557.355 ;
    END
  END mprj_io_holdover[0]
  PIN mprj_io_ib_mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 572.255 3379.435 572.535 ;
    END
  END mprj_io_ib_mode_sel[0]
  PIN mprj_io_inp_dis[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 538.215 3379.435 538.495 ;
    END
  END mprj_io_inp_dis[0]
  PIN mprj_io_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 575.475 3379.435 575.755 ;
    END
  END mprj_io_oeb[0]
  PIN mprj_io_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 559.835 3379.435 560.115 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_slow_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 513.835 3379.435 514.115 ;
    END
  END mprj_io_slow_sel[0]
  PIN mprj_io_vtrip_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 569.035 3379.435 569.315 ;
    END
  END mprj_io_vtrip_sel[0]
  PIN mprj_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 504.635 3379.435 504.915 ;
    END
  END mprj_io_in[0]
  PIN mprj_analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3433.055 3379.435 3433.335 ;
    END
  END mprj_analog_io[3]
  PIN mprj_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3422.200 3555.010 3484.900 ;
    END
  END mprj_io[10]
  PIN mprj_io_analog_en[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3445.015 3379.435 3445.295 ;
    END
  END mprj_io_analog_en[10]
  PIN mprj_io_analog_pol[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3451.455 3379.435 3451.735 ;
    END
  END mprj_io_analog_pol[10]
  PIN mprj_io_analog_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3466.635 3379.435 3466.915 ;
    END
  END mprj_io_analog_sel[10]
  PIN mprj_io_dm[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3448.235 3379.435 3448.515 ;
    END
  END mprj_io_dm[30]
  PIN mprj_io_dm[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3439.035 3379.435 3439.315 ;
    END
  END mprj_io_dm[31]
  PIN mprj_io_dm[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3469.855 3379.435 3470.135 ;
    END
  END mprj_io_dm[32]
  PIN mprj_io_holdover[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3473.075 3379.435 3473.355 ;
    END
  END mprj_io_holdover[10]
  PIN mprj_io_ib_mode_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3488.255 3379.435 3488.535 ;
    END
  END mprj_io_ib_mode_sel[10]
  PIN mprj_io_inp_dis[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3454.215 3379.435 3454.495 ;
    END
  END mprj_io_inp_dis[10]
  PIN mprj_io_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3491.475 3379.435 3491.755 ;
    END
  END mprj_io_oeb[10]
  PIN mprj_io_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3475.835 3379.435 3476.115 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_slow_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3429.835 3379.435 3430.115 ;
    END
  END mprj_io_slow_sel[10]
  PIN mprj_io_vtrip_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3485.035 3379.435 3485.315 ;
    END
  END mprj_io_vtrip_sel[10]
  PIN mprj_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3420.635 3379.435 3420.915 ;
    END
  END mprj_io_in[10]
  PIN mprj_analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3658.055 3379.435 3658.335 ;
    END
  END mprj_analog_io[4]
  PIN mprj_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3647.200 3555.010 3709.900 ;
    END
  END mprj_io[11]
  PIN mprj_io_analog_en[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3670.015 3379.435 3670.295 ;
    END
  END mprj_io_analog_en[11]
  PIN mprj_io_analog_pol[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3676.455 3379.435 3676.735 ;
    END
  END mprj_io_analog_pol[11]
  PIN mprj_io_analog_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3691.635 3379.435 3691.915 ;
    END
  END mprj_io_analog_sel[11]
  PIN mprj_io_dm[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3673.235 3379.435 3673.515 ;
    END
  END mprj_io_dm[33]
  PIN mprj_io_dm[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3664.035 3379.435 3664.315 ;
    END
  END mprj_io_dm[34]
  PIN mprj_io_dm[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3694.855 3379.435 3695.135 ;
    END
  END mprj_io_dm[35]
  PIN mprj_io_holdover[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3698.075 3379.435 3698.355 ;
    END
  END mprj_io_holdover[11]
  PIN mprj_io_ib_mode_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3713.255 3379.435 3713.535 ;
    END
  END mprj_io_ib_mode_sel[11]
  PIN mprj_io_inp_dis[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3679.215 3379.435 3679.495 ;
    END
  END mprj_io_inp_dis[11]
  PIN mprj_io_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3716.475 3379.435 3716.755 ;
    END
  END mprj_io_oeb[11]
  PIN mprj_io_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3700.835 3379.435 3701.115 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_slow_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3654.835 3379.435 3655.115 ;
    END
  END mprj_io_slow_sel[11]
  PIN mprj_io_vtrip_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3710.035 3379.435 3710.315 ;
    END
  END mprj_io_vtrip_sel[11]
  PIN mprj_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3645.635 3379.435 3645.915 ;
    END
  END mprj_io_in[11]
  PIN mprj_analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3883.055 3379.435 3883.335 ;
    END
  END mprj_analog_io[5]
  PIN mprj_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3872.200 3555.010 3934.900 ;
    END
  END mprj_io[12]
  PIN mprj_io_analog_en[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3895.015 3379.435 3895.295 ;
    END
  END mprj_io_analog_en[12]
  PIN mprj_io_analog_pol[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3901.455 3379.435 3901.735 ;
    END
  END mprj_io_analog_pol[12]
  PIN mprj_io_analog_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3916.635 3379.435 3916.915 ;
    END
  END mprj_io_analog_sel[12]
  PIN mprj_io_dm[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3898.235 3379.435 3898.515 ;
    END
  END mprj_io_dm[36]
  PIN mprj_io_dm[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3889.035 3379.435 3889.315 ;
    END
  END mprj_io_dm[37]
  PIN mprj_io_dm[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3919.855 3379.435 3920.135 ;
    END
  END mprj_io_dm[38]
  PIN mprj_io_holdover[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3923.075 3379.435 3923.355 ;
    END
  END mprj_io_holdover[12]
  PIN mprj_io_ib_mode_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3938.255 3379.435 3938.535 ;
    END
  END mprj_io_ib_mode_sel[12]
  PIN mprj_io_inp_dis[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3904.215 3379.435 3904.495 ;
    END
  END mprj_io_inp_dis[12]
  PIN mprj_io_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3941.475 3379.435 3941.755 ;
    END
  END mprj_io_oeb[12]
  PIN mprj_io_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3925.835 3379.435 3926.115 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_slow_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3879.835 3379.435 3880.115 ;
    END
  END mprj_io_slow_sel[12]
  PIN mprj_io_vtrip_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3935.035 3379.435 3935.315 ;
    END
  END mprj_io_vtrip_sel[12]
  PIN mprj_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3870.635 3379.435 3870.915 ;
    END
  END mprj_io_in[12]
  PIN mprj_analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4329.055 3379.435 4329.335 ;
    END
  END mprj_analog_io[6]
  PIN mprj_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4318.200 3555.010 4380.900 ;
    END
  END mprj_io[13]
  PIN mprj_io_analog_en[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4341.015 3379.435 4341.295 ;
    END
  END mprj_io_analog_en[13]
  PIN mprj_io_analog_pol[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4347.455 3379.435 4347.735 ;
    END
  END mprj_io_analog_pol[13]
  PIN mprj_io_analog_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4362.635 3379.435 4362.915 ;
    END
  END mprj_io_analog_sel[13]
  PIN mprj_io_dm[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4344.235 3379.435 4344.515 ;
    END
  END mprj_io_dm[39]
  PIN mprj_io_dm[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4335.035 3379.435 4335.315 ;
    END
  END mprj_io_dm[40]
  PIN mprj_io_dm[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4365.855 3379.435 4366.135 ;
    END
  END mprj_io_dm[41]
  PIN mprj_io_holdover[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4369.075 3379.435 4369.355 ;
    END
  END mprj_io_holdover[13]
  PIN mprj_io_ib_mode_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4384.255 3379.435 4384.535 ;
    END
  END mprj_io_ib_mode_sel[13]
  PIN mprj_io_inp_dis[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4350.215 3379.435 4350.495 ;
    END
  END mprj_io_inp_dis[13]
  PIN mprj_io_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4387.475 3379.435 4387.755 ;
    END
  END mprj_io_oeb[13]
  PIN mprj_io_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4371.835 3379.435 4372.115 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_slow_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4325.835 3379.435 4326.115 ;
    END
  END mprj_io_slow_sel[13]
  PIN mprj_io_vtrip_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4381.035 3379.435 4381.315 ;
    END
  END mprj_io_vtrip_sel[13]
  PIN mprj_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4316.635 3379.435 4316.915 ;
    END
  END mprj_io_in[13]
  PIN mprj_analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4775.055 3379.435 4775.335 ;
    END
  END mprj_analog_io[7]
  PIN mprj_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 4764.200 3555.010 4826.900 ;
    END
  END mprj_io[14]
  PIN mprj_io_analog_en[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4787.015 3379.435 4787.295 ;
    END
  END mprj_io_analog_en[14]
  PIN mprj_io_analog_pol[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4793.455 3379.435 4793.735 ;
    END
  END mprj_io_analog_pol[14]
  PIN mprj_io_analog_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4808.635 3379.435 4808.915 ;
    END
  END mprj_io_analog_sel[14]
  PIN mprj_io_dm[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4790.235 3379.435 4790.515 ;
    END
  END mprj_io_dm[42]
  PIN mprj_io_dm[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4781.035 3379.435 4781.315 ;
    END
  END mprj_io_dm[43]
  PIN mprj_io_dm[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4811.855 3379.435 4812.135 ;
    END
  END mprj_io_dm[44]
  PIN mprj_io_holdover[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4815.075 3379.435 4815.355 ;
    END
  END mprj_io_holdover[14]
  PIN mprj_io_ib_mode_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4830.255 3379.435 4830.535 ;
    END
  END mprj_io_ib_mode_sel[14]
  PIN mprj_io_inp_dis[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4796.215 3379.435 4796.495 ;
    END
  END mprj_io_inp_dis[14]
  PIN mprj_io_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4833.475 3379.435 4833.755 ;
    END
  END mprj_io_oeb[14]
  PIN mprj_io_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4817.835 3379.435 4818.115 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_slow_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4771.835 3379.435 4772.115 ;
    END
  END mprj_io_slow_sel[14]
  PIN mprj_io_vtrip_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4827.035 3379.435 4827.315 ;
    END
  END mprj_io_vtrip_sel[14]
  PIN mprj_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 4762.635 3379.435 4762.915 ;
    END
  END mprj_io_in[14]
  PIN mprj_analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3192.665 4977.035 3192.945 4979.435 ;
    END
  END mprj_analog_io[8]
  PIN mprj_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3141.100 5092.560 3203.800 5155.010 ;
    END
  END mprj_io[15]
  PIN mprj_io_analog_en[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3180.705 4977.035 3180.985 4979.435 ;
    END
  END mprj_io_analog_en[15]
  PIN mprj_io_analog_pol[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3174.265 4977.035 3174.545 4979.435 ;
    END
  END mprj_io_analog_pol[15]
  PIN mprj_io_analog_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3159.085 4977.035 3159.365 4979.435 ;
    END
  END mprj_io_analog_sel[15]
  PIN mprj_io_dm[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3177.485 4977.035 3177.765 4979.435 ;
    END
  END mprj_io_dm[45]
  PIN mprj_io_dm[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3186.685 4977.035 3186.965 4979.435 ;
    END
  END mprj_io_dm[46]
  PIN mprj_io_dm[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3155.865 4977.035 3156.145 4979.435 ;
    END
  END mprj_io_dm[47]
  PIN mprj_io_holdover[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3152.645 4977.035 3152.925 4979.435 ;
    END
  END mprj_io_holdover[15]
  PIN mprj_io_ib_mode_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3137.465 4977.035 3137.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[15]
  PIN mprj_io_inp_dis[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3171.505 4977.035 3171.785 4979.435 ;
    END
  END mprj_io_inp_dis[15]
  PIN mprj_io_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3134.245 4977.035 3134.525 4979.435 ;
    END
  END mprj_io_oeb[15]
  PIN mprj_io_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3149.885 4977.035 3150.165 4979.435 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_slow_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3195.885 4977.035 3196.165 4979.435 ;
    END
  END mprj_io_slow_sel[15]
  PIN mprj_io_vtrip_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3140.685 4977.035 3140.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[15]
  PIN mprj_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3205.085 4977.035 3205.365 4979.435 ;
    END
  END mprj_io_in[15]
  PIN mprj_analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2683.665 4977.035 2683.945 4979.435 ;
    END
  END mprj_analog_io[9]
  PIN mprj_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2632.100 5092.560 2694.800 5155.010 ;
    END
  END mprj_io[16]
  PIN mprj_io_analog_en[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.705 4977.035 2671.985 4979.435 ;
    END
  END mprj_io_analog_en[16]
  PIN mprj_io_analog_pol[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.265 4977.035 2665.545 4979.435 ;
    END
  END mprj_io_analog_pol[16]
  PIN mprj_io_analog_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.085 4977.035 2650.365 4979.435 ;
    END
  END mprj_io_analog_sel[16]
  PIN mprj_io_dm[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.485 4977.035 2668.765 4979.435 ;
    END
  END mprj_io_dm[48]
  PIN mprj_io_dm[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2677.685 4977.035 2677.965 4979.435 ;
    END
  END mprj_io_dm[49]
  PIN mprj_io_dm[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.865 4977.035 2647.145 4979.435 ;
    END
  END mprj_io_dm[50]
  PIN mprj_io_holdover[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.645 4977.035 2643.925 4979.435 ;
    END
  END mprj_io_holdover[16]
  PIN mprj_io_ib_mode_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2628.465 4977.035 2628.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[16]
  PIN mprj_io_inp_dis[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.505 4977.035 2662.785 4979.435 ;
    END
  END mprj_io_inp_dis[16]
  PIN mprj_io_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.245 4977.035 2625.525 4979.435 ;
    END
  END mprj_io_oeb[16]
  PIN mprj_io_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2640.885 4977.035 2641.165 4979.435 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_slow_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2686.885 4977.035 2687.165 4979.435 ;
    END
  END mprj_io_slow_sel[16]
  PIN mprj_io_vtrip_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.685 4977.035 2631.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[16]
  PIN mprj_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.085 4977.035 2696.365 4979.435 ;
    END
  END mprj_io_in[16]
  PIN mprj_analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2426.665 4977.035 2426.945 4979.435 ;
    END
  END mprj_analog_io[10]
  PIN mprj_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2375.100 5092.560 2437.800 5155.010 ;
    END
  END mprj_io[17]
  PIN mprj_io_analog_en[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.705 4977.035 2414.985 4979.435 ;
    END
  END mprj_io_analog_en[17]
  PIN mprj_io_analog_pol[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.265 4977.035 2408.545 4979.435 ;
    END
  END mprj_io_analog_pol[17]
  PIN mprj_io_analog_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.085 4977.035 2393.365 4979.435 ;
    END
  END mprj_io_analog_sel[17]
  PIN mprj_io_dm[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.485 4977.035 2411.765 4979.435 ;
    END
  END mprj_io_dm[51]
  PIN mprj_io_dm[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.685 4977.035 2420.965 4979.435 ;
    END
  END mprj_io_dm[52]
  PIN mprj_io_dm[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.865 4977.035 2390.145 4979.435 ;
    END
  END mprj_io_dm[53]
  PIN mprj_io_holdover[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.645 4977.035 2386.925 4979.435 ;
    END
  END mprj_io_holdover[17]
  PIN mprj_io_ib_mode_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2371.465 4977.035 2371.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[17]
  PIN mprj_io_inp_dis[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.505 4977.035 2405.785 4979.435 ;
    END
  END mprj_io_inp_dis[17]
  PIN mprj_io_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.245 4977.035 2368.525 4979.435 ;
    END
  END mprj_io_oeb[17]
  PIN mprj_io_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2383.885 4977.035 2384.165 4979.435 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_slow_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.885 4977.035 2430.165 4979.435 ;
    END
  END mprj_io_slow_sel[17]
  PIN mprj_io_vtrip_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.685 4977.035 2374.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[17]
  PIN mprj_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.085 4977.035 2439.365 4979.435 ;
    END
  END mprj_io_in[17]
  PIN mprj_analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.665 4977.035 1981.945 4979.435 ;
    END
  END mprj_analog_io[11]
  PIN mprj_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1930.100 5092.560 1992.800 5155.010 ;
    END
  END mprj_io[18]
  PIN mprj_io_analog_en[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.705 4977.035 1969.985 4979.435 ;
    END
  END mprj_io_analog_en[18]
  PIN mprj_io_analog_pol[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.265 4977.035 1963.545 4979.435 ;
    END
  END mprj_io_analog_pol[18]
  PIN mprj_io_analog_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.085 4977.035 1948.365 4979.435 ;
    END
  END mprj_io_analog_sel[18]
  PIN mprj_io_dm[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.485 4977.035 1966.765 4979.435 ;
    END
  END mprj_io_dm[54]
  PIN mprj_io_dm[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.685 4977.035 1975.965 4979.435 ;
    END
  END mprj_io_dm[55]
  PIN mprj_io_dm[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.865 4977.035 1945.145 4979.435 ;
    END
  END mprj_io_dm[56]
  PIN mprj_io_holdover[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.645 4977.035 1941.925 4979.435 ;
    END
  END mprj_io_holdover[18]
  PIN mprj_io_ib_mode_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.465 4977.035 1926.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[18]
  PIN mprj_io_inp_dis[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1960.505 4977.035 1960.785 4979.435 ;
    END
  END mprj_io_inp_dis[18]
  PIN mprj_io_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.245 4977.035 1923.525 4979.435 ;
    END
  END mprj_io_oeb[18]
  PIN mprj_io_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.885 4977.035 1939.165 4979.435 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_slow_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.885 4977.035 1985.165 4979.435 ;
    END
  END mprj_io_slow_sel[18]
  PIN mprj_io_vtrip_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.685 4977.035 1929.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[18]
  PIN mprj_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.085 4977.035 1994.365 4979.435 ;
    END
  END mprj_io_in[18]
  PIN mprj_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 732.200 3555.010 794.900 ;
    END
  END mprj_io[1]
  PIN mprj_io_analog_en[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 755.015 3379.435 755.295 ;
    END
  END mprj_io_analog_en[1]
  PIN mprj_io_analog_pol[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 761.455 3379.435 761.735 ;
    END
  END mprj_io_analog_pol[1]
  PIN mprj_io_analog_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 776.635 3379.435 776.915 ;
    END
  END mprj_io_analog_sel[1]
  PIN mprj_io_dm[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 758.235 3379.435 758.515 ;
    END
  END mprj_io_dm[3]
  PIN mprj_io_dm[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 749.035 3379.435 749.315 ;
    END
  END mprj_io_dm[4]
  PIN mprj_io_dm[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 779.855 3379.435 780.135 ;
    END
  END mprj_io_dm[5]
  PIN mprj_io_holdover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 783.075 3379.435 783.355 ;
    END
  END mprj_io_holdover[1]
  PIN mprj_io_ib_mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 798.255 3379.435 798.535 ;
    END
  END mprj_io_ib_mode_sel[1]
  PIN mprj_io_inp_dis[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 764.215 3379.435 764.495 ;
    END
  END mprj_io_inp_dis[1]
  PIN mprj_io_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 801.475 3379.435 801.755 ;
    END
  END mprj_io_oeb[1]
  PIN mprj_io_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 785.835 3379.435 786.115 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_slow_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 739.835 3379.435 740.115 ;
    END
  END mprj_io_slow_sel[1]
  PIN mprj_io_vtrip_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 795.035 3379.435 795.315 ;
    END
  END mprj_io_vtrip_sel[1]
  PIN mprj_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 730.635 3379.435 730.915 ;
    END
  END mprj_io_in[1]
  PIN mprj_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 957.200 3555.010 1019.900 ;
    END
  END mprj_io[2]
  PIN mprj_io_analog_en[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 980.015 3379.435 980.295 ;
    END
  END mprj_io_analog_en[2]
  PIN mprj_io_analog_pol[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 986.455 3379.435 986.735 ;
    END
  END mprj_io_analog_pol[2]
  PIN mprj_io_analog_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1001.635 3379.435 1001.915 ;
    END
  END mprj_io_analog_sel[2]
  PIN mprj_io_dm[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 983.235 3379.435 983.515 ;
    END
  END mprj_io_dm[6]
  PIN mprj_io_dm[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 974.035 3379.435 974.315 ;
    END
  END mprj_io_dm[7]
  PIN mprj_io_dm[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1004.855 3379.435 1005.135 ;
    END
  END mprj_io_dm[8]
  PIN mprj_io_holdover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1008.075 3379.435 1008.355 ;
    END
  END mprj_io_holdover[2]
  PIN mprj_io_ib_mode_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1023.255 3379.435 1023.535 ;
    END
  END mprj_io_ib_mode_sel[2]
  PIN mprj_io_inp_dis[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 989.215 3379.435 989.495 ;
    END
  END mprj_io_inp_dis[2]
  PIN mprj_io_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1026.475 3379.435 1026.755 ;
    END
  END mprj_io_oeb[2]
  PIN mprj_io_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1010.835 3379.435 1011.115 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_slow_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 964.835 3379.435 965.115 ;
    END
  END mprj_io_slow_sel[2]
  PIN mprj_io_vtrip_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1020.035 3379.435 1020.315 ;
    END
  END mprj_io_vtrip_sel[2]
  PIN mprj_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 955.635 3379.435 955.915 ;
    END
  END mprj_io_in[2]
  PIN mprj_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1183.200 3555.010 1245.900 ;
    END
  END mprj_io[3]
  PIN mprj_io_analog_en[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1206.015 3379.435 1206.295 ;
    END
  END mprj_io_analog_en[3]
  PIN mprj_io_analog_pol[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1212.455 3379.435 1212.735 ;
    END
  END mprj_io_analog_pol[3]
  PIN mprj_io_analog_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1227.635 3379.435 1227.915 ;
    END
  END mprj_io_analog_sel[3]
  PIN mprj_io_dm[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1200.035 3379.435 1200.315 ;
    END
  END mprj_io_dm[10]
  PIN mprj_io_dm[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1230.855 3379.435 1231.135 ;
    END
  END mprj_io_dm[11]
  PIN mprj_io_dm[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1209.235 3379.435 1209.515 ;
    END
  END mprj_io_dm[9]
  PIN mprj_io_holdover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1234.075 3379.435 1234.355 ;
    END
  END mprj_io_holdover[3]
  PIN mprj_io_ib_mode_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1249.255 3379.435 1249.535 ;
    END
  END mprj_io_ib_mode_sel[3]
  PIN mprj_io_inp_dis[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1215.215 3379.435 1215.495 ;
    END
  END mprj_io_inp_dis[3]
  PIN mprj_io_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1252.475 3379.435 1252.755 ;
    END
  END mprj_io_oeb[3]
  PIN mprj_io_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1236.835 3379.435 1237.115 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_slow_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1190.835 3379.435 1191.115 ;
    END
  END mprj_io_slow_sel[3]
  PIN mprj_io_vtrip_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1246.035 3379.435 1246.315 ;
    END
  END mprj_io_vtrip_sel[3]
  PIN mprj_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1181.635 3379.435 1181.915 ;
    END
  END mprj_io_in[3]
  PIN mprj_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1408.200 3555.010 1470.900 ;
    END
  END mprj_io[4]
  PIN mprj_io_analog_en[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1431.015 3379.435 1431.295 ;
    END
  END mprj_io_analog_en[4]
  PIN mprj_io_analog_pol[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1437.455 3379.435 1437.735 ;
    END
  END mprj_io_analog_pol[4]
  PIN mprj_io_analog_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1452.635 3379.435 1452.915 ;
    END
  END mprj_io_analog_sel[4]
  PIN mprj_io_dm[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1434.235 3379.435 1434.515 ;
    END
  END mprj_io_dm[12]
  PIN mprj_io_dm[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1425.035 3379.435 1425.315 ;
    END
  END mprj_io_dm[13]
  PIN mprj_io_dm[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1455.855 3379.435 1456.135 ;
    END
  END mprj_io_dm[14]
  PIN mprj_io_holdover[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1459.075 3379.435 1459.355 ;
    END
  END mprj_io_holdover[4]
  PIN mprj_io_ib_mode_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1474.255 3379.435 1474.535 ;
    END
  END mprj_io_ib_mode_sel[4]
  PIN mprj_io_inp_dis[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1440.215 3379.435 1440.495 ;
    END
  END mprj_io_inp_dis[4]
  PIN mprj_io_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1477.475 3379.435 1477.755 ;
    END
  END mprj_io_oeb[4]
  PIN mprj_io_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1461.835 3379.435 1462.115 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_slow_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1415.835 3379.435 1416.115 ;
    END
  END mprj_io_slow_sel[4]
  PIN mprj_io_vtrip_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1471.035 3379.435 1471.315 ;
    END
  END mprj_io_vtrip_sel[4]
  PIN mprj_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1406.635 3379.435 1406.915 ;
    END
  END mprj_io_in[4]
  PIN mprj_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1633.200 3555.010 1695.900 ;
    END
  END mprj_io[5]
  PIN mprj_io_analog_en[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1656.015 3379.435 1656.295 ;
    END
  END mprj_io_analog_en[5]
  PIN mprj_io_analog_pol[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1662.455 3379.435 1662.735 ;
    END
  END mprj_io_analog_pol[5]
  PIN mprj_io_analog_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1677.635 3379.435 1677.915 ;
    END
  END mprj_io_analog_sel[5]
  PIN mprj_io_dm[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1659.235 3379.435 1659.515 ;
    END
  END mprj_io_dm[15]
  PIN mprj_io_dm[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1650.035 3379.435 1650.315 ;
    END
  END mprj_io_dm[16]
  PIN mprj_io_dm[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1680.855 3379.435 1681.135 ;
    END
  END mprj_io_dm[17]
  PIN mprj_io_holdover[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1684.075 3379.435 1684.355 ;
    END
  END mprj_io_holdover[5]
  PIN mprj_io_ib_mode_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1699.255 3379.435 1699.535 ;
    END
  END mprj_io_ib_mode_sel[5]
  PIN mprj_io_inp_dis[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1665.215 3379.435 1665.495 ;
    END
  END mprj_io_inp_dis[5]
  PIN mprj_io_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1702.475 3379.435 1702.755 ;
    END
  END mprj_io_oeb[5]
  PIN mprj_io_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1686.835 3379.435 1687.115 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_slow_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1640.835 3379.435 1641.115 ;
    END
  END mprj_io_slow_sel[5]
  PIN mprj_io_vtrip_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1696.035 3379.435 1696.315 ;
    END
  END mprj_io_vtrip_sel[5]
  PIN mprj_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1631.635 3379.435 1631.915 ;
    END
  END mprj_io_in[5]
  PIN mprj_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 1859.200 3555.010 1921.900 ;
    END
  END mprj_io[6]
  PIN mprj_io_analog_en[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1882.015 3379.435 1882.295 ;
    END
  END mprj_io_analog_en[6]
  PIN mprj_io_analog_pol[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1888.455 3379.435 1888.735 ;
    END
  END mprj_io_analog_pol[6]
  PIN mprj_io_analog_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1903.635 3379.435 1903.915 ;
    END
  END mprj_io_analog_sel[6]
  PIN mprj_io_dm[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1885.235 3379.435 1885.515 ;
    END
  END mprj_io_dm[18]
  PIN mprj_io_dm[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1876.035 3379.435 1876.315 ;
    END
  END mprj_io_dm[19]
  PIN mprj_io_dm[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1906.855 3379.435 1907.135 ;
    END
  END mprj_io_dm[20]
  PIN mprj_io_holdover[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1910.075 3379.435 1910.355 ;
    END
  END mprj_io_holdover[6]
  PIN mprj_io_ib_mode_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1925.255 3379.435 1925.535 ;
    END
  END mprj_io_ib_mode_sel[6]
  PIN mprj_io_inp_dis[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1891.215 3379.435 1891.495 ;
    END
  END mprj_io_inp_dis[6]
  PIN mprj_io_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1928.475 3379.435 1928.755 ;
    END
  END mprj_io_oeb[6]
  PIN mprj_io_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1912.835 3379.435 1913.115 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_slow_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1866.835 3379.435 1867.115 ;
    END
  END mprj_io_slow_sel[6]
  PIN mprj_io_vtrip_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1922.035 3379.435 1922.315 ;
    END
  END mprj_io_vtrip_sel[6]
  PIN mprj_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 1857.635 3379.435 1857.915 ;
    END
  END mprj_io_in[6]
  PIN mprj_analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2756.055 3379.435 2756.335 ;
    END
  END mprj_analog_io[0]
  PIN mprj_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2745.200 3555.010 2807.900 ;
    END
  END mprj_io[7]
  PIN mprj_io_analog_en[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2768.015 3379.435 2768.295 ;
    END
  END mprj_io_analog_en[7]
  PIN mprj_io_analog_pol[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2774.455 3379.435 2774.735 ;
    END
  END mprj_io_analog_pol[7]
  PIN mprj_io_analog_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2789.635 3379.435 2789.915 ;
    END
  END mprj_io_analog_sel[7]
  PIN mprj_io_dm[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2771.235 3379.435 2771.515 ;
    END
  END mprj_io_dm[21]
  PIN mprj_io_dm[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2762.035 3379.435 2762.315 ;
    END
  END mprj_io_dm[22]
  PIN mprj_io_dm[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2792.855 3379.435 2793.135 ;
    END
  END mprj_io_dm[23]
  PIN mprj_io_holdover[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2796.075 3379.435 2796.355 ;
    END
  END mprj_io_holdover[7]
  PIN mprj_io_ib_mode_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2811.255 3379.435 2811.535 ;
    END
  END mprj_io_ib_mode_sel[7]
  PIN mprj_io_inp_dis[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2777.215 3379.435 2777.495 ;
    END
  END mprj_io_inp_dis[7]
  PIN mprj_io_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2814.475 3379.435 2814.755 ;
    END
  END mprj_io_oeb[7]
  PIN mprj_io_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2798.835 3379.435 2799.115 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_slow_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2752.835 3379.435 2753.115 ;
    END
  END mprj_io_slow_sel[7]
  PIN mprj_io_vtrip_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2808.035 3379.435 2808.315 ;
    END
  END mprj_io_vtrip_sel[7]
  PIN mprj_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2743.635 3379.435 2743.915 ;
    END
  END mprj_io_in[7]
  PIN mprj_analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2982.055 3379.435 2982.335 ;
    END
  END mprj_analog_io[1]
  PIN mprj_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 2971.200 3555.010 3033.900 ;
    END
  END mprj_io[8]
  PIN mprj_io_analog_en[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2994.015 3379.435 2994.295 ;
    END
  END mprj_io_analog_en[8]
  PIN mprj_io_analog_pol[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3000.455 3379.435 3000.735 ;
    END
  END mprj_io_analog_pol[8]
  PIN mprj_io_analog_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3015.635 3379.435 3015.915 ;
    END
  END mprj_io_analog_sel[8]
  PIN mprj_io_dm[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2997.235 3379.435 2997.515 ;
    END
  END mprj_io_dm[24]
  PIN mprj_io_dm[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2988.035 3379.435 2988.315 ;
    END
  END mprj_io_dm[25]
  PIN mprj_io_dm[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3018.855 3379.435 3019.135 ;
    END
  END mprj_io_dm[26]
  PIN mprj_io_holdover[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3022.075 3379.435 3022.355 ;
    END
  END mprj_io_holdover[8]
  PIN mprj_io_ib_mode_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3037.255 3379.435 3037.535 ;
    END
  END mprj_io_ib_mode_sel[8]
  PIN mprj_io_inp_dis[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3003.215 3379.435 3003.495 ;
    END
  END mprj_io_inp_dis[8]
  PIN mprj_io_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3040.475 3379.435 3040.755 ;
    END
  END mprj_io_oeb[8]
  PIN mprj_io_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3024.835 3379.435 3025.115 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_slow_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2978.835 3379.435 2979.115 ;
    END
  END mprj_io_slow_sel[8]
  PIN mprj_io_vtrip_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3034.035 3379.435 3034.315 ;
    END
  END mprj_io_vtrip_sel[8]
  PIN mprj_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 2969.635 3379.435 2969.915 ;
    END
  END mprj_io_in[8]
  PIN mprj_analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3207.055 3379.435 3207.335 ;
    END
  END mprj_analog_io[2]
  PIN mprj_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3492.560 3196.200 3555.010 3258.900 ;
    END
  END mprj_io[9]
  PIN mprj_io_analog_en[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3219.015 3379.435 3219.295 ;
    END
  END mprj_io_analog_en[9]
  PIN mprj_io_analog_pol[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3225.455 3379.435 3225.735 ;
    END
  END mprj_io_analog_pol[9]
  PIN mprj_io_analog_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3240.635 3379.435 3240.915 ;
    END
  END mprj_io_analog_sel[9]
  PIN mprj_io_dm[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3222.235 3379.435 3222.515 ;
    END
  END mprj_io_dm[27]
  PIN mprj_io_dm[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3213.035 3379.435 3213.315 ;
    END
  END mprj_io_dm[28]
  PIN mprj_io_dm[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3243.855 3379.435 3244.135 ;
    END
  END mprj_io_dm[29]
  PIN mprj_io_holdover[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3247.075 3379.435 3247.355 ;
    END
  END mprj_io_holdover[9]
  PIN mprj_io_ib_mode_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3262.255 3379.435 3262.535 ;
    END
  END mprj_io_ib_mode_sel[9]
  PIN mprj_io_inp_dis[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3228.215 3379.435 3228.495 ;
    END
  END mprj_io_inp_dis[9]
  PIN mprj_io_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3265.475 3379.435 3265.755 ;
    END
  END mprj_io_oeb[9]
  PIN mprj_io_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3249.835 3379.435 3250.115 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_slow_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3203.835 3379.435 3204.115 ;
    END
  END mprj_io_slow_sel[9]
  PIN mprj_io_vtrip_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3259.035 3379.435 3259.315 ;
    END
  END mprj_io_vtrip_sel[9]
  PIN mprj_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3377.035 3194.635 3379.435 3194.915 ;
    END
  END mprj_io_in[9]
  PIN mprj_analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.665 4977.035 1472.945 4979.435 ;
    END
  END mprj_analog_io[12]
  PIN mprj_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1421.100 5092.560 1483.800 5155.010 ;
    END
  END mprj_io[19]
  PIN mprj_io_analog_en[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.705 4977.035 1460.985 4979.435 ;
    END
  END mprj_io_analog_en[19]
  PIN mprj_io_analog_pol[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.265 4977.035 1454.545 4979.435 ;
    END
  END mprj_io_analog_pol[19]
  PIN mprj_io_analog_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.085 4977.035 1439.365 4979.435 ;
    END
  END mprj_io_analog_sel[19]
  PIN mprj_io_dm[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.485 4977.035 1457.765 4979.435 ;
    END
  END mprj_io_dm[57]
  PIN mprj_io_dm[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.685 4977.035 1466.965 4979.435 ;
    END
  END mprj_io_dm[58]
  PIN mprj_io_dm[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.865 4977.035 1436.145 4979.435 ;
    END
  END mprj_io_dm[59]
  PIN mprj_io_holdover[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.645 4977.035 1432.925 4979.435 ;
    END
  END mprj_io_holdover[19]
  PIN mprj_io_ib_mode_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.465 4977.035 1417.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[19]
  PIN mprj_io_inp_dis[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.505 4977.035 1451.785 4979.435 ;
    END
  END mprj_io_inp_dis[19]
  PIN mprj_io_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.245 4977.035 1414.525 4979.435 ;
    END
  END mprj_io_oeb[19]
  PIN mprj_io_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.885 4977.035 1430.165 4979.435 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_slow_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.885 4977.035 1476.165 4979.435 ;
    END
  END mprj_io_slow_sel[19]
  PIN mprj_io_vtrip_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.685 4977.035 1420.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[19]
  PIN mprj_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.085 4977.035 1485.365 4979.435 ;
    END
  END mprj_io_in[19]
  PIN mprj_analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3120.665 210.965 3120.945 ;
    END
  END mprj_analog_io[22]
  PIN mprj_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3069.100 95.440 3131.800 ;
    END
  END mprj_io[29]
  PIN mprj_io_analog_en[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3108.705 210.965 3108.985 ;
    END
  END mprj_io_analog_en[29]
  PIN mprj_io_analog_pol[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3102.265 210.965 3102.545 ;
    END
  END mprj_io_analog_pol[29]
  PIN mprj_io_analog_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3087.085 210.965 3087.365 ;
    END
  END mprj_io_analog_sel[29]
  PIN mprj_io_dm[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3105.485 210.965 3105.765 ;
    END
  END mprj_io_dm[87]
  PIN mprj_io_dm[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3114.685 210.965 3114.965 ;
    END
  END mprj_io_dm[88]
  PIN mprj_io_dm[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3083.865 210.965 3084.145 ;
    END
  END mprj_io_dm[89]
  PIN mprj_io_holdover[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3080.645 210.965 3080.925 ;
    END
  END mprj_io_holdover[29]
  PIN mprj_io_ib_mode_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3065.465 210.965 3065.745 ;
    END
  END mprj_io_ib_mode_sel[29]
  PIN mprj_io_inp_dis[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3099.505 210.965 3099.785 ;
    END
  END mprj_io_inp_dis[29]
  PIN mprj_io_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3062.245 210.965 3062.525 ;
    END
  END mprj_io_oeb[29]
  PIN mprj_io_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3077.885 210.965 3078.165 ;
    END
  END mprj_io_out[29]
  PIN mprj_io_slow_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3123.885 210.965 3124.165 ;
    END
  END mprj_io_slow_sel[29]
  PIN mprj_io_vtrip_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3068.685 210.965 3068.965 ;
    END
  END mprj_io_vtrip_sel[29]
  PIN mprj_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3133.085 210.965 3133.365 ;
    END
  END mprj_io_in[29]
  PIN mprj_analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2904.665 210.965 2904.945 ;
    END
  END mprj_analog_io[23]
  PIN mprj_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2853.100 95.440 2915.800 ;
    END
  END mprj_io[30]
  PIN mprj_io_analog_en[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2892.705 210.965 2892.985 ;
    END
  END mprj_io_analog_en[30]
  PIN mprj_io_analog_pol[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2886.265 210.965 2886.545 ;
    END
  END mprj_io_analog_pol[30]
  PIN mprj_io_analog_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2871.085 210.965 2871.365 ;
    END
  END mprj_io_analog_sel[30]
  PIN mprj_io_dm[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2889.485 210.965 2889.765 ;
    END
  END mprj_io_dm[90]
  PIN mprj_io_dm[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2898.685 210.965 2898.965 ;
    END
  END mprj_io_dm[91]
  PIN mprj_io_dm[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2867.865 210.965 2868.145 ;
    END
  END mprj_io_dm[92]
  PIN mprj_io_holdover[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2864.645 210.965 2864.925 ;
    END
  END mprj_io_holdover[30]
  PIN mprj_io_ib_mode_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2849.465 210.965 2849.745 ;
    END
  END mprj_io_ib_mode_sel[30]
  PIN mprj_io_inp_dis[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2883.505 210.965 2883.785 ;
    END
  END mprj_io_inp_dis[30]
  PIN mprj_io_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2846.245 210.965 2846.525 ;
    END
  END mprj_io_oeb[30]
  PIN mprj_io_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2861.885 210.965 2862.165 ;
    END
  END mprj_io_out[30]
  PIN mprj_io_slow_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2907.885 210.965 2908.165 ;
    END
  END mprj_io_slow_sel[30]
  PIN mprj_io_vtrip_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2852.685 210.965 2852.965 ;
    END
  END mprj_io_vtrip_sel[30]
  PIN mprj_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2917.085 210.965 2917.365 ;
    END
  END mprj_io_in[30]
  PIN mprj_analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2688.665 210.965 2688.945 ;
    END
  END mprj_analog_io[24]
  PIN mprj_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 2637.100 95.440 2699.800 ;
    END
  END mprj_io[31]
  PIN mprj_io_analog_en[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2676.705 210.965 2676.985 ;
    END
  END mprj_io_analog_en[31]
  PIN mprj_io_analog_pol[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2670.265 210.965 2670.545 ;
    END
  END mprj_io_analog_pol[31]
  PIN mprj_io_analog_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2655.085 210.965 2655.365 ;
    END
  END mprj_io_analog_sel[31]
  PIN mprj_io_dm[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2673.485 210.965 2673.765 ;
    END
  END mprj_io_dm[93]
  PIN mprj_io_dm[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2682.685 210.965 2682.965 ;
    END
  END mprj_io_dm[94]
  PIN mprj_io_dm[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2651.865 210.965 2652.145 ;
    END
  END mprj_io_dm[95]
  PIN mprj_io_holdover[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2648.645 210.965 2648.925 ;
    END
  END mprj_io_holdover[31]
  PIN mprj_io_ib_mode_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2633.465 210.965 2633.745 ;
    END
  END mprj_io_ib_mode_sel[31]
  PIN mprj_io_inp_dis[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2667.505 210.965 2667.785 ;
    END
  END mprj_io_inp_dis[31]
  PIN mprj_io_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2630.245 210.965 2630.525 ;
    END
  END mprj_io_oeb[31]
  PIN mprj_io_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2645.885 210.965 2646.165 ;
    END
  END mprj_io_out[31]
  PIN mprj_io_slow_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2691.885 210.965 2692.165 ;
    END
  END mprj_io_slow_sel[31]
  PIN mprj_io_vtrip_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2636.685 210.965 2636.965 ;
    END
  END mprj_io_vtrip_sel[31]
  PIN mprj_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2701.085 210.965 2701.365 ;
    END
  END mprj_io_in[31]
  PIN mprj_analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2050.665 210.965 2050.945 ;
    END
  END mprj_analog_io[25]
  PIN mprj_io[32]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1999.100 95.440 2061.800 ;
    END
  END mprj_io[32]
  PIN mprj_io_analog_en[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2038.705 210.965 2038.985 ;
    END
  END mprj_io_analog_en[32]
  PIN mprj_io_analog_pol[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2032.265 210.965 2032.545 ;
    END
  END mprj_io_analog_pol[32]
  PIN mprj_io_analog_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2017.085 210.965 2017.365 ;
    END
  END mprj_io_analog_sel[32]
  PIN mprj_io_dm[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2035.485 210.965 2035.765 ;
    END
  END mprj_io_dm[96]
  PIN mprj_io_dm[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2044.685 210.965 2044.965 ;
    END
  END mprj_io_dm[97]
  PIN mprj_io_dm[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2013.865 210.965 2014.145 ;
    END
  END mprj_io_dm[98]
  PIN mprj_io_holdover[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2010.645 210.965 2010.925 ;
    END
  END mprj_io_holdover[32]
  PIN mprj_io_ib_mode_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1995.465 210.965 1995.745 ;
    END
  END mprj_io_ib_mode_sel[32]
  PIN mprj_io_inp_dis[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2029.505 210.965 2029.785 ;
    END
  END mprj_io_inp_dis[32]
  PIN mprj_io_oeb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1992.245 210.965 1992.525 ;
    END
  END mprj_io_oeb[32]
  PIN mprj_io_out[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2007.885 210.965 2008.165 ;
    END
  END mprj_io_out[32]
  PIN mprj_io_slow_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2053.885 210.965 2054.165 ;
    END
  END mprj_io_slow_sel[32]
  PIN mprj_io_vtrip_sel[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1998.685 210.965 1998.965 ;
    END
  END mprj_io_vtrip_sel[32]
  PIN mprj_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 2063.085 210.965 2063.365 ;
    END
  END mprj_io_in[32]
  PIN mprj_analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1834.665 210.965 1834.945 ;
    END
  END mprj_analog_io[26]
  PIN mprj_io[33]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1783.100 95.440 1845.800 ;
    END
  END mprj_io[33]
  PIN mprj_io_analog_en[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1822.705 210.965 1822.985 ;
    END
  END mprj_io_analog_en[33]
  PIN mprj_io_analog_pol[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1816.265 210.965 1816.545 ;
    END
  END mprj_io_analog_pol[33]
  PIN mprj_io_analog_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1801.085 210.965 1801.365 ;
    END
  END mprj_io_analog_sel[33]
  PIN mprj_io_dm[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1828.685 210.965 1828.965 ;
    END
  END mprj_io_dm[100]
  PIN mprj_io_dm[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1797.865 210.965 1798.145 ;
    END
  END mprj_io_dm[101]
  PIN mprj_io_dm[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1819.485 210.965 1819.765 ;
    END
  END mprj_io_dm[99]
  PIN mprj_io_holdover[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1794.645 210.965 1794.925 ;
    END
  END mprj_io_holdover[33]
  PIN mprj_io_ib_mode_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1779.465 210.965 1779.745 ;
    END
  END mprj_io_ib_mode_sel[33]
  PIN mprj_io_inp_dis[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1813.505 210.965 1813.785 ;
    END
  END mprj_io_inp_dis[33]
  PIN mprj_io_oeb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1776.245 210.965 1776.525 ;
    END
  END mprj_io_oeb[33]
  PIN mprj_io_out[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1791.885 210.965 1792.165 ;
    END
  END mprj_io_out[33]
  PIN mprj_io_slow_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1837.885 210.965 1838.165 ;
    END
  END mprj_io_slow_sel[33]
  PIN mprj_io_vtrip_sel[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1782.685 210.965 1782.965 ;
    END
  END mprj_io_vtrip_sel[33]
  PIN mprj_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1847.085 210.965 1847.365 ;
    END
  END mprj_io_in[33]
  PIN mprj_analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1618.665 210.965 1618.945 ;
    END
  END mprj_analog_io[27]
  PIN mprj_io[34]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1567.100 95.440 1629.800 ;
    END
  END mprj_io[34]
  PIN mprj_io_analog_en[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1606.705 210.965 1606.985 ;
    END
  END mprj_io_analog_en[34]
  PIN mprj_io_analog_pol[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1600.265 210.965 1600.545 ;
    END
  END mprj_io_analog_pol[34]
  PIN mprj_io_analog_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1585.085 210.965 1585.365 ;
    END
  END mprj_io_analog_sel[34]
  PIN mprj_io_dm[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1603.485 210.965 1603.765 ;
    END
  END mprj_io_dm[102]
  PIN mprj_io_dm[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1612.685 210.965 1612.965 ;
    END
  END mprj_io_dm[103]
  PIN mprj_io_dm[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1581.865 210.965 1582.145 ;
    END
  END mprj_io_dm[104]
  PIN mprj_io_holdover[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1578.645 210.965 1578.925 ;
    END
  END mprj_io_holdover[34]
  PIN mprj_io_ib_mode_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1563.465 210.965 1563.745 ;
    END
  END mprj_io_ib_mode_sel[34]
  PIN mprj_io_inp_dis[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1597.505 210.965 1597.785 ;
    END
  END mprj_io_inp_dis[34]
  PIN mprj_io_oeb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1560.245 210.965 1560.525 ;
    END
  END mprj_io_oeb[34]
  PIN mprj_io_out[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1575.885 210.965 1576.165 ;
    END
  END mprj_io_out[34]
  PIN mprj_io_slow_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1621.885 210.965 1622.165 ;
    END
  END mprj_io_slow_sel[34]
  PIN mprj_io_vtrip_sel[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1566.685 210.965 1566.965 ;
    END
  END mprj_io_vtrip_sel[34]
  PIN mprj_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1631.085 210.965 1631.365 ;
    END
  END mprj_io_in[34]
  PIN mprj_analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1402.665 210.965 1402.945 ;
    END
  END mprj_analog_io[28]
  PIN mprj_io[35]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1351.100 95.440 1413.800 ;
    END
  END mprj_io[35]
  PIN mprj_io_analog_en[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1390.705 210.965 1390.985 ;
    END
  END mprj_io_analog_en[35]
  PIN mprj_io_analog_pol[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1384.265 210.965 1384.545 ;
    END
  END mprj_io_analog_pol[35]
  PIN mprj_io_analog_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1369.085 210.965 1369.365 ;
    END
  END mprj_io_analog_sel[35]
  PIN mprj_io_dm[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1387.485 210.965 1387.765 ;
    END
  END mprj_io_dm[105]
  PIN mprj_io_dm[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1396.685 210.965 1396.965 ;
    END
  END mprj_io_dm[106]
  PIN mprj_io_dm[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1365.865 210.965 1366.145 ;
    END
  END mprj_io_dm[107]
  PIN mprj_io_holdover[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1362.645 210.965 1362.925 ;
    END
  END mprj_io_holdover[35]
  PIN mprj_io_ib_mode_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1347.465 210.965 1347.745 ;
    END
  END mprj_io_ib_mode_sel[35]
  PIN mprj_io_inp_dis[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1381.505 210.965 1381.785 ;
    END
  END mprj_io_inp_dis[35]
  PIN mprj_io_oeb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1344.245 210.965 1344.525 ;
    END
  END mprj_io_oeb[35]
  PIN mprj_io_out[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1359.885 210.965 1360.165 ;
    END
  END mprj_io_out[35]
  PIN mprj_io_slow_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1405.885 210.965 1406.165 ;
    END
  END mprj_io_slow_sel[35]
  PIN mprj_io_vtrip_sel[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1350.685 210.965 1350.965 ;
    END
  END mprj_io_vtrip_sel[35]
  PIN mprj_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1415.085 210.965 1415.365 ;
    END
  END mprj_io_in[35]
  PIN mprj_io[36]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 1135.100 95.440 1197.800 ;
    END
  END mprj_io[36]
  PIN mprj_io_analog_en[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1174.705 210.965 1174.985 ;
    END
  END mprj_io_analog_en[36]
  PIN mprj_io_analog_pol[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1168.265 210.965 1168.545 ;
    END
  END mprj_io_analog_pol[36]
  PIN mprj_io_analog_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1153.085 210.965 1153.365 ;
    END
  END mprj_io_analog_sel[36]
  PIN mprj_io_dm[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1171.485 210.965 1171.765 ;
    END
  END mprj_io_dm[108]
  PIN mprj_io_dm[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1180.685 210.965 1180.965 ;
    END
  END mprj_io_dm[109]
  PIN mprj_io_dm[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1149.865 210.965 1150.145 ;
    END
  END mprj_io_dm[110]
  PIN mprj_io_holdover[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1146.645 210.965 1146.925 ;
    END
  END mprj_io_holdover[36]
  PIN mprj_io_ib_mode_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1131.465 210.965 1131.745 ;
    END
  END mprj_io_ib_mode_sel[36]
  PIN mprj_io_inp_dis[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1165.505 210.965 1165.785 ;
    END
  END mprj_io_inp_dis[36]
  PIN mprj_io_oeb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1128.245 210.965 1128.525 ;
    END
  END mprj_io_oeb[36]
  PIN mprj_io_out[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1143.885 210.965 1144.165 ;
    END
  END mprj_io_out[36]
  PIN mprj_io_slow_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1189.885 210.965 1190.165 ;
    END
  END mprj_io_slow_sel[36]
  PIN mprj_io_vtrip_sel[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1134.685 210.965 1134.965 ;
    END
  END mprj_io_vtrip_sel[36]
  PIN mprj_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 1199.085 210.965 1199.365 ;
    END
  END mprj_io_in[36]
  PIN mprj_io[37]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 919.100 95.440 981.800 ;
    END
  END mprj_io[37]
  PIN mprj_io_analog_en[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 958.705 210.965 958.985 ;
    END
  END mprj_io_analog_en[37]
  PIN mprj_io_analog_pol[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 952.265 210.965 952.545 ;
    END
  END mprj_io_analog_pol[37]
  PIN mprj_io_analog_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 937.085 210.965 937.365 ;
    END
  END mprj_io_analog_sel[37]
  PIN mprj_io_dm[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 955.485 210.965 955.765 ;
    END
  END mprj_io_dm[111]
  PIN mprj_io_dm[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 964.685 210.965 964.965 ;
    END
  END mprj_io_dm[112]
  PIN mprj_io_dm[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 933.865 210.965 934.145 ;
    END
  END mprj_io_dm[113]
  PIN mprj_io_holdover[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 930.645 210.965 930.925 ;
    END
  END mprj_io_holdover[37]
  PIN mprj_io_ib_mode_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 915.465 210.965 915.745 ;
    END
  END mprj_io_ib_mode_sel[37]
  PIN mprj_io_inp_dis[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 949.505 210.965 949.785 ;
    END
  END mprj_io_inp_dis[37]
  PIN mprj_io_oeb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 912.245 210.965 912.525 ;
    END
  END mprj_io_oeb[37]
  PIN mprj_io_out[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 927.885 210.965 928.165 ;
    END
  END mprj_io_out[37]
  PIN mprj_io_slow_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 973.885 210.965 974.165 ;
    END
  END mprj_io_slow_sel[37]
  PIN mprj_io_vtrip_sel[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 918.685 210.965 918.965 ;
    END
  END mprj_io_vtrip_sel[37]
  PIN mprj_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 983.085 210.965 983.365 ;
    END
  END mprj_io_in[37]
  PIN mprj_analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.665 4977.035 1214.945 4979.435 ;
    END
  END mprj_analog_io[13]
  PIN mprj_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1163.100 5092.560 1225.800 5155.010 ;
    END
  END mprj_io[20]
  PIN mprj_io_analog_en[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.705 4977.035 1202.985 4979.435 ;
    END
  END mprj_io_analog_en[20]
  PIN mprj_io_analog_pol[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.265 4977.035 1196.545 4979.435 ;
    END
  END mprj_io_analog_pol[20]
  PIN mprj_io_analog_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.085 4977.035 1181.365 4979.435 ;
    END
  END mprj_io_analog_sel[20]
  PIN mprj_io_dm[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.485 4977.035 1199.765 4979.435 ;
    END
  END mprj_io_dm[60]
  PIN mprj_io_dm[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.685 4977.035 1208.965 4979.435 ;
    END
  END mprj_io_dm[61]
  PIN mprj_io_dm[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.865 4977.035 1178.145 4979.435 ;
    END
  END mprj_io_dm[62]
  PIN mprj_io_holdover[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.645 4977.035 1174.925 4979.435 ;
    END
  END mprj_io_holdover[20]
  PIN mprj_io_ib_mode_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.465 4977.035 1159.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[20]
  PIN mprj_io_inp_dis[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.505 4977.035 1193.785 4979.435 ;
    END
  END mprj_io_inp_dis[20]
  PIN mprj_io_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.245 4977.035 1156.525 4979.435 ;
    END
  END mprj_io_oeb[20]
  PIN mprj_io_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.885 4977.035 1172.165 4979.435 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_slow_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.885 4977.035 1218.165 4979.435 ;
    END
  END mprj_io_slow_sel[20]
  PIN mprj_io_vtrip_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.685 4977.035 1162.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[20]
  PIN mprj_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.085 4977.035 1227.365 4979.435 ;
    END
  END mprj_io_in[20]
  PIN mprj_analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.665 4977.035 957.945 4979.435 ;
    END
  END mprj_analog_io[14]
  PIN mprj_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 906.100 5092.560 968.800 5155.010 ;
    END
  END mprj_io[21]
  PIN mprj_io_analog_en[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.705 4977.035 945.985 4979.435 ;
    END
  END mprj_io_analog_en[21]
  PIN mprj_io_analog_pol[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.265 4977.035 939.545 4979.435 ;
    END
  END mprj_io_analog_pol[21]
  PIN mprj_io_analog_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.085 4977.035 924.365 4979.435 ;
    END
  END mprj_io_analog_sel[21]
  PIN mprj_io_dm[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.485 4977.035 942.765 4979.435 ;
    END
  END mprj_io_dm[63]
  PIN mprj_io_dm[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.685 4977.035 951.965 4979.435 ;
    END
  END mprj_io_dm[64]
  PIN mprj_io_dm[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.865 4977.035 921.145 4979.435 ;
    END
  END mprj_io_dm[65]
  PIN mprj_io_holdover[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.645 4977.035 917.925 4979.435 ;
    END
  END mprj_io_holdover[21]
  PIN mprj_io_ib_mode_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.465 4977.035 902.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[21]
  PIN mprj_io_inp_dis[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.505 4977.035 936.785 4979.435 ;
    END
  END mprj_io_inp_dis[21]
  PIN mprj_io_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.245 4977.035 899.525 4979.435 ;
    END
  END mprj_io_oeb[21]
  PIN mprj_io_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.885 4977.035 915.165 4979.435 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_slow_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.885 4977.035 961.165 4979.435 ;
    END
  END mprj_io_slow_sel[21]
  PIN mprj_io_vtrip_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.685 4977.035 905.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[21]
  PIN mprj_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.085 4977.035 970.365 4979.435 ;
    END
  END mprj_io_in[21]
  PIN mprj_analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.665 4977.035 700.945 4979.435 ;
    END
  END mprj_analog_io[15]
  PIN mprj_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 649.100 5092.560 711.800 5155.010 ;
    END
  END mprj_io[22]
  PIN mprj_io_analog_en[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.705 4977.035 688.985 4979.435 ;
    END
  END mprj_io_analog_en[22]
  PIN mprj_io_analog_pol[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.265 4977.035 682.545 4979.435 ;
    END
  END mprj_io_analog_pol[22]
  PIN mprj_io_analog_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.085 4977.035 667.365 4979.435 ;
    END
  END mprj_io_analog_sel[22]
  PIN mprj_io_dm[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.485 4977.035 685.765 4979.435 ;
    END
  END mprj_io_dm[66]
  PIN mprj_io_dm[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.685 4977.035 694.965 4979.435 ;
    END
  END mprj_io_dm[67]
  PIN mprj_io_dm[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.865 4977.035 664.145 4979.435 ;
    END
  END mprj_io_dm[68]
  PIN mprj_io_holdover[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.645 4977.035 660.925 4979.435 ;
    END
  END mprj_io_holdover[22]
  PIN mprj_io_ib_mode_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.465 4977.035 645.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[22]
  PIN mprj_io_inp_dis[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.505 4977.035 679.785 4979.435 ;
    END
  END mprj_io_inp_dis[22]
  PIN mprj_io_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.245 4977.035 642.525 4979.435 ;
    END
  END mprj_io_oeb[22]
  PIN mprj_io_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.885 4977.035 658.165 4979.435 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_slow_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.885 4977.035 704.165 4979.435 ;
    END
  END mprj_io_slow_sel[22]
  PIN mprj_io_vtrip_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.685 4977.035 648.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[22]
  PIN mprj_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.085 4977.035 713.365 4979.435 ;
    END
  END mprj_io_in[22]
  PIN mprj_analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.665 4977.035 443.945 4979.435 ;
    END
  END mprj_analog_io[16]
  PIN mprj_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 392.100 5092.560 454.800 5155.010 ;
    END
  END mprj_io[23]
  PIN mprj_io_analog_en[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.705 4977.035 431.985 4979.435 ;
    END
  END mprj_io_analog_en[23]
  PIN mprj_io_analog_pol[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.265 4977.035 425.545 4979.435 ;
    END
  END mprj_io_analog_pol[23]
  PIN mprj_io_analog_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.085 4977.035 410.365 4979.435 ;
    END
  END mprj_io_analog_sel[23]
  PIN mprj_io_dm[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.485 4977.035 428.765 4979.435 ;
    END
  END mprj_io_dm[69]
  PIN mprj_io_dm[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.685 4977.035 437.965 4979.435 ;
    END
  END mprj_io_dm[70]
  PIN mprj_io_dm[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.865 4977.035 407.145 4979.435 ;
    END
  END mprj_io_dm[71]
  PIN mprj_io_holdover[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.645 4977.035 403.925 4979.435 ;
    END
  END mprj_io_holdover[23]
  PIN mprj_io_ib_mode_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.465 4977.035 388.745 4979.435 ;
    END
  END mprj_io_ib_mode_sel[23]
  PIN mprj_io_inp_dis[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.505 4977.035 422.785 4979.435 ;
    END
  END mprj_io_inp_dis[23]
  PIN mprj_io_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.245 4977.035 385.525 4979.435 ;
    END
  END mprj_io_oeb[23]
  PIN mprj_io_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.885 4977.035 401.165 4979.435 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_slow_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.885 4977.035 447.165 4979.435 ;
    END
  END mprj_io_slow_sel[23]
  PIN mprj_io_vtrip_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.685 4977.035 391.965 4979.435 ;
    END
  END mprj_io_vtrip_sel[23]
  PIN mprj_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.085 4977.035 456.365 4979.435 ;
    END
  END mprj_io_in[23]
  PIN mprj_analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4833.665 210.965 4833.945 ;
    END
  END mprj_analog_io[17]
  PIN mprj_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 4782.100 95.440 4844.800 ;
    END
  END mprj_io[24]
  PIN mprj_io_analog_en[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4821.705 210.965 4821.985 ;
    END
  END mprj_io_analog_en[24]
  PIN mprj_io_analog_pol[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4815.265 210.965 4815.545 ;
    END
  END mprj_io_analog_pol[24]
  PIN mprj_io_analog_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4800.085 210.965 4800.365 ;
    END
  END mprj_io_analog_sel[24]
  PIN mprj_io_dm[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4818.485 210.965 4818.765 ;
    END
  END mprj_io_dm[72]
  PIN mprj_io_dm[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4827.685 210.965 4827.965 ;
    END
  END mprj_io_dm[73]
  PIN mprj_io_dm[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4796.865 210.965 4797.145 ;
    END
  END mprj_io_dm[74]
  PIN mprj_io_holdover[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4793.645 210.965 4793.925 ;
    END
  END mprj_io_holdover[24]
  PIN mprj_io_ib_mode_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4778.465 210.965 4778.745 ;
    END
  END mprj_io_ib_mode_sel[24]
  PIN mprj_io_inp_dis[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4812.505 210.965 4812.785 ;
    END
  END mprj_io_inp_dis[24]
  PIN mprj_io_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4775.245 210.965 4775.525 ;
    END
  END mprj_io_oeb[24]
  PIN mprj_io_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4790.885 210.965 4791.165 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_slow_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4836.885 210.965 4837.165 ;
    END
  END mprj_io_slow_sel[24]
  PIN mprj_io_vtrip_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4781.685 210.965 4781.965 ;
    END
  END mprj_io_vtrip_sel[24]
  PIN mprj_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 4846.085 210.965 4846.365 ;
    END
  END mprj_io_in[24]
  PIN mprj_analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3984.665 210.965 3984.945 ;
    END
  END mprj_analog_io[18]
  PIN mprj_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3933.100 95.440 3995.800 ;
    END
  END mprj_io[25]
  PIN mprj_io_analog_en[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3972.705 210.965 3972.985 ;
    END
  END mprj_io_analog_en[25]
  PIN mprj_io_analog_pol[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3966.265 210.965 3966.545 ;
    END
  END mprj_io_analog_pol[25]
  PIN mprj_io_analog_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3951.085 210.965 3951.365 ;
    END
  END mprj_io_analog_sel[25]
  PIN mprj_io_dm[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3969.485 210.965 3969.765 ;
    END
  END mprj_io_dm[75]
  PIN mprj_io_dm[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3978.685 210.965 3978.965 ;
    END
  END mprj_io_dm[76]
  PIN mprj_io_dm[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3947.865 210.965 3948.145 ;
    END
  END mprj_io_dm[77]
  PIN mprj_io_holdover[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3944.645 210.965 3944.925 ;
    END
  END mprj_io_holdover[25]
  PIN mprj_io_ib_mode_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3929.465 210.965 3929.745 ;
    END
  END mprj_io_ib_mode_sel[25]
  PIN mprj_io_inp_dis[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3963.505 210.965 3963.785 ;
    END
  END mprj_io_inp_dis[25]
  PIN mprj_io_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3926.245 210.965 3926.525 ;
    END
  END mprj_io_oeb[25]
  PIN mprj_io_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3941.885 210.965 3942.165 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_slow_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3987.885 210.965 3988.165 ;
    END
  END mprj_io_slow_sel[25]
  PIN mprj_io_vtrip_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3932.685 210.965 3932.965 ;
    END
  END mprj_io_vtrip_sel[25]
  PIN mprj_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3997.085 210.965 3997.365 ;
    END
  END mprj_io_in[25]
  PIN mprj_analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3768.665 210.965 3768.945 ;
    END
  END mprj_analog_io[19]
  PIN mprj_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3717.100 95.440 3779.800 ;
    END
  END mprj_io[26]
  PIN mprj_io_analog_en[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3756.705 210.965 3756.985 ;
    END
  END mprj_io_analog_en[26]
  PIN mprj_io_analog_pol[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3750.265 210.965 3750.545 ;
    END
  END mprj_io_analog_pol[26]
  PIN mprj_io_analog_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3735.085 210.965 3735.365 ;
    END
  END mprj_io_analog_sel[26]
  PIN mprj_io_dm[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3753.485 210.965 3753.765 ;
    END
  END mprj_io_dm[78]
  PIN mprj_io_dm[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3762.685 210.965 3762.965 ;
    END
  END mprj_io_dm[79]
  PIN mprj_io_dm[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3731.865 210.965 3732.145 ;
    END
  END mprj_io_dm[80]
  PIN mprj_io_holdover[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3728.645 210.965 3728.925 ;
    END
  END mprj_io_holdover[26]
  PIN mprj_io_ib_mode_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3713.465 210.965 3713.745 ;
    END
  END mprj_io_ib_mode_sel[26]
  PIN mprj_io_inp_dis[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3747.505 210.965 3747.785 ;
    END
  END mprj_io_inp_dis[26]
  PIN mprj_io_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3710.245 210.965 3710.525 ;
    END
  END mprj_io_oeb[26]
  PIN mprj_io_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3725.885 210.965 3726.165 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_slow_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3771.885 210.965 3772.165 ;
    END
  END mprj_io_slow_sel[26]
  PIN mprj_io_vtrip_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3716.685 210.965 3716.965 ;
    END
  END mprj_io_vtrip_sel[26]
  PIN mprj_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3781.085 210.965 3781.365 ;
    END
  END mprj_io_in[26]
  PIN mprj_analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3552.665 210.965 3552.945 ;
    END
  END mprj_analog_io[20]
  PIN mprj_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3501.100 95.440 3563.800 ;
    END
  END mprj_io[27]
  PIN mprj_io_analog_en[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3540.705 210.965 3540.985 ;
    END
  END mprj_io_analog_en[27]
  PIN mprj_io_analog_pol[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3534.265 210.965 3534.545 ;
    END
  END mprj_io_analog_pol[27]
  PIN mprj_io_analog_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3519.085 210.965 3519.365 ;
    END
  END mprj_io_analog_sel[27]
  PIN mprj_io_dm[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3537.485 210.965 3537.765 ;
    END
  END mprj_io_dm[81]
  PIN mprj_io_dm[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3546.685 210.965 3546.965 ;
    END
  END mprj_io_dm[82]
  PIN mprj_io_dm[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3515.865 210.965 3516.145 ;
    END
  END mprj_io_dm[83]
  PIN mprj_io_holdover[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3512.645 210.965 3512.925 ;
    END
  END mprj_io_holdover[27]
  PIN mprj_io_ib_mode_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3497.465 210.965 3497.745 ;
    END
  END mprj_io_ib_mode_sel[27]
  PIN mprj_io_inp_dis[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3531.505 210.965 3531.785 ;
    END
  END mprj_io_inp_dis[27]
  PIN mprj_io_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3494.245 210.965 3494.525 ;
    END
  END mprj_io_oeb[27]
  PIN mprj_io_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3509.885 210.965 3510.165 ;
    END
  END mprj_io_out[27]
  PIN mprj_io_slow_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3555.885 210.965 3556.165 ;
    END
  END mprj_io_slow_sel[27]
  PIN mprj_io_vtrip_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3500.685 210.965 3500.965 ;
    END
  END mprj_io_vtrip_sel[27]
  PIN mprj_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3565.085 210.965 3565.365 ;
    END
  END mprj_io_in[27]
  PIN mprj_analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3336.665 210.965 3336.945 ;
    END
  END mprj_analog_io[21]
  PIN mprj_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.990 3285.100 95.440 3347.800 ;
    END
  END mprj_io[28]
  PIN mprj_io_analog_en[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3324.705 210.965 3324.985 ;
    END
  END mprj_io_analog_en[28]
  PIN mprj_io_analog_pol[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3318.265 210.965 3318.545 ;
    END
  END mprj_io_analog_pol[28]
  PIN mprj_io_analog_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3303.085 210.965 3303.365 ;
    END
  END mprj_io_analog_sel[28]
  PIN mprj_io_dm[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3321.485 210.965 3321.765 ;
    END
  END mprj_io_dm[84]
  PIN mprj_io_dm[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3330.685 210.965 3330.965 ;
    END
  END mprj_io_dm[85]
  PIN mprj_io_dm[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3299.865 210.965 3300.145 ;
    END
  END mprj_io_dm[86]
  PIN mprj_io_holdover[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3296.645 210.965 3296.925 ;
    END
  END mprj_io_holdover[28]
  PIN mprj_io_ib_mode_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3281.465 210.965 3281.745 ;
    END
  END mprj_io_ib_mode_sel[28]
  PIN mprj_io_inp_dis[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3315.505 210.965 3315.785 ;
    END
  END mprj_io_inp_dis[28]
  PIN mprj_io_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3278.245 210.965 3278.525 ;
    END
  END mprj_io_oeb[28]
  PIN mprj_io_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3293.885 210.965 3294.165 ;
    END
  END mprj_io_out[28]
  PIN mprj_io_slow_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3339.885 210.965 3340.165 ;
    END
  END mprj_io_slow_sel[28]
  PIN mprj_io_vtrip_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3284.685 210.965 3284.965 ;
    END
  END mprj_io_vtrip_sel[28]
  PIN mprj_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.565 3349.085 210.965 3349.365 ;
    END
  END mprj_io_in[28]
  PIN porb_h
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1423.310 4976.480 1423.630 4976.540 ;
        RECT 1444.930 4976.480 1445.250 4976.540 ;
        RECT 1423.310 4976.340 1445.250 4976.480 ;
        RECT 1423.310 4976.280 1423.630 4976.340 ;
        RECT 1444.930 4976.280 1445.250 4976.340 ;
        RECT 651.430 4976.140 651.750 4976.200 ;
        RECT 673.050 4976.140 673.370 4976.200 ;
        RECT 651.430 4976.000 673.370 4976.140 ;
        RECT 651.430 4975.940 651.750 4976.000 ;
        RECT 673.050 4975.940 673.370 4976.000 ;
        RECT 2634.490 4976.140 2634.810 4976.200 ;
        RECT 2656.110 4976.140 2656.430 4976.200 ;
        RECT 2634.490 4976.000 2656.430 4976.140 ;
        RECT 2634.490 4975.940 2634.810 4976.000 ;
        RECT 2656.110 4975.940 2656.430 4976.000 ;
        RECT 394.290 4967.980 394.610 4968.040 ;
        RECT 415.910 4967.980 416.230 4968.040 ;
        RECT 394.290 4967.840 416.230 4967.980 ;
        RECT 394.290 4967.780 394.610 4967.840 ;
        RECT 415.910 4967.780 416.230 4967.840 ;
        RECT 1443.090 4967.300 1443.410 4967.360 ;
        RECT 1444.930 4967.300 1445.250 4967.360 ;
        RECT 1932.530 4967.300 1932.850 4967.360 ;
        RECT 1953.230 4967.300 1953.550 4967.360 ;
        RECT 1443.090 4967.160 1953.550 4967.300 ;
        RECT 1443.090 4967.100 1443.410 4967.160 ;
        RECT 1444.930 4967.100 1445.250 4967.160 ;
        RECT 1932.530 4967.100 1932.850 4967.160 ;
        RECT 1953.230 4967.100 1953.550 4967.160 ;
        RECT 415.910 4966.960 416.230 4967.020 ;
        RECT 651.430 4966.960 651.750 4967.020 ;
        RECT 908.570 4966.960 908.890 4967.020 ;
        RECT 930.190 4966.960 930.510 4967.020 ;
        RECT 1165.250 4966.960 1165.570 4967.020 ;
        RECT 1186.870 4966.960 1187.190 4967.020 ;
        RECT 415.910 4966.820 1187.190 4966.960 ;
        RECT 415.910 4966.760 416.230 4966.820 ;
        RECT 651.430 4966.760 651.750 4966.820 ;
        RECT 908.570 4966.760 908.890 4966.820 ;
        RECT 930.190 4966.760 930.510 4966.820 ;
        RECT 1165.250 4966.760 1165.570 4966.820 ;
        RECT 1186.870 4966.760 1187.190 4966.820 ;
        RECT 1954.610 4966.960 1954.930 4967.020 ;
        RECT 2377.350 4966.960 2377.670 4967.020 ;
        RECT 2398.970 4966.960 2399.290 4967.020 ;
        RECT 2634.490 4966.960 2634.810 4967.020 ;
        RECT 3143.250 4966.960 3143.570 4967.020 ;
        RECT 3164.870 4966.960 3165.190 4967.020 ;
        RECT 1954.610 4966.820 3165.190 4966.960 ;
        RECT 1954.610 4966.760 1954.930 4966.820 ;
        RECT 2377.350 4966.760 2377.670 4966.820 ;
        RECT 2398.970 4966.760 2399.290 4966.820 ;
        RECT 2634.490 4966.760 2634.810 4966.820 ;
        RECT 3143.250 4966.760 3143.570 4966.820 ;
        RECT 3164.870 4966.760 3165.190 4966.820 ;
        RECT 1186.960 4966.620 1187.100 4966.760 ;
        RECT 1443.090 4966.620 1443.410 4966.680 ;
        RECT 1186.960 4966.480 1443.410 4966.620 ;
        RECT 1443.090 4966.420 1443.410 4966.480 ;
        RECT 218.110 4965.600 218.430 4965.660 ;
        RECT 394.290 4965.600 394.610 4965.660 ;
        RECT 218.110 4965.460 394.610 4965.600 ;
        RECT 218.110 4965.400 218.430 4965.460 ;
        RECT 394.290 4965.400 394.610 4965.460 ;
        RECT 3164.870 4964.920 3165.190 4964.980 ;
        RECT 3371.870 4964.920 3372.190 4964.980 ;
        RECT 3164.870 4964.780 3372.190 4964.920 ;
        RECT 3164.870 4964.720 3165.190 4964.780 ;
        RECT 3371.870 4964.720 3372.190 4964.780 ;
        RECT 3371.870 4837.080 3372.190 4837.140 ;
        RECT 3376.010 4837.080 3376.330 4837.140 ;
        RECT 3371.870 4836.940 3376.330 4837.080 ;
        RECT 3371.870 4836.880 3372.190 4836.940 ;
        RECT 3376.010 4836.880 3376.330 4836.940 ;
        RECT 3376.010 4826.540 3376.330 4826.600 ;
        RECT 3376.930 4826.540 3377.250 4826.600 ;
        RECT 3376.010 4826.400 3377.250 4826.540 ;
        RECT 3376.010 4826.340 3376.330 4826.400 ;
        RECT 3376.930 4826.340 3377.250 4826.400 ;
        RECT 208.910 4806.820 209.230 4806.880 ;
        RECT 211.670 4806.820 211.990 4806.880 ;
        RECT 218.110 4806.820 218.430 4806.880 ;
        RECT 208.910 4806.680 218.430 4806.820 ;
        RECT 208.910 4806.620 209.230 4806.680 ;
        RECT 211.670 4806.620 211.990 4806.680 ;
        RECT 218.110 4806.620 218.430 4806.680 ;
        RECT 3375.090 4379.100 3375.410 4379.160 ;
        RECT 3376.930 4379.100 3377.250 4379.160 ;
        RECT 3375.090 4378.960 3377.250 4379.100 ;
        RECT 3375.090 4378.900 3375.410 4378.960 ;
        RECT 3376.930 4378.900 3377.250 4378.960 ;
        RECT 208.910 3959.880 209.230 3959.940 ;
        RECT 212.590 3959.880 212.910 3959.940 ;
        RECT 208.910 3959.740 212.910 3959.880 ;
        RECT 208.910 3959.680 209.230 3959.740 ;
        RECT 212.590 3959.680 212.910 3959.740 ;
        RECT 208.910 3933.360 209.230 3933.420 ;
        RECT 211.670 3933.360 211.990 3933.420 ;
        RECT 208.910 3933.220 211.990 3933.360 ;
        RECT 208.910 3933.160 209.230 3933.220 ;
        RECT 211.670 3933.160 211.990 3933.220 ;
        RECT 3376.010 3933.020 3376.330 3933.080 ;
        RECT 3376.930 3933.020 3377.250 3933.080 ;
        RECT 3376.010 3932.880 3377.250 3933.020 ;
        RECT 3376.010 3932.820 3376.330 3932.880 ;
        RECT 3376.930 3932.820 3377.250 3932.880 ;
        RECT 3376.010 3913.640 3376.330 3913.700 ;
        RECT 3376.930 3913.640 3377.250 3913.700 ;
        RECT 3376.010 3913.500 3377.250 3913.640 ;
        RECT 3376.010 3913.440 3376.330 3913.500 ;
        RECT 3376.930 3913.440 3377.250 3913.500 ;
        RECT 208.910 3738.540 209.230 3738.600 ;
        RECT 211.670 3738.540 211.990 3738.600 ;
        RECT 208.910 3738.400 211.990 3738.540 ;
        RECT 208.910 3738.340 209.230 3738.400 ;
        RECT 211.670 3738.340 211.990 3738.400 ;
        RECT 208.910 3719.160 209.230 3719.220 ;
        RECT 211.670 3719.160 211.990 3719.220 ;
        RECT 208.910 3719.020 211.990 3719.160 ;
        RECT 208.910 3718.960 209.230 3719.020 ;
        RECT 211.670 3718.960 211.990 3719.020 ;
        RECT 3375.550 3705.220 3375.870 3705.280 ;
        RECT 3377.850 3705.220 3378.170 3705.280 ;
        RECT 3375.550 3705.080 3378.170 3705.220 ;
        RECT 3375.550 3705.020 3375.870 3705.080 ;
        RECT 3377.850 3705.020 3378.170 3705.080 ;
        RECT 3375.550 3685.160 3375.870 3685.220 ;
        RECT 3376.930 3685.160 3377.250 3685.220 ;
        RECT 3375.550 3685.020 3377.250 3685.160 ;
        RECT 3375.550 3684.960 3375.870 3685.020 ;
        RECT 3376.930 3684.960 3377.250 3685.020 ;
        RECT 211.670 3528.900 211.990 3529.160 ;
        RECT 211.760 3527.800 211.900 3528.900 ;
        RECT 208.910 3527.740 209.230 3527.800 ;
        RECT 211.670 3527.740 211.990 3527.800 ;
        RECT 208.910 3527.600 211.990 3527.740 ;
        RECT 208.910 3527.540 209.230 3527.600 ;
        RECT 211.670 3527.540 211.990 3527.600 ;
        RECT 3375.090 3479.800 3375.410 3479.860 ;
        RECT 3376.930 3479.800 3377.250 3479.860 ;
        RECT 3375.090 3479.660 3377.250 3479.800 ;
        RECT 3375.090 3479.600 3375.410 3479.660 ;
        RECT 3376.930 3479.600 3377.250 3479.660 ;
        RECT 3375.090 3460.420 3375.410 3460.480 ;
        RECT 3376.930 3460.420 3377.250 3460.480 ;
        RECT 3375.090 3460.280 3377.250 3460.420 ;
        RECT 3375.090 3460.220 3375.410 3460.280 ;
        RECT 3376.930 3460.220 3377.250 3460.280 ;
        RECT 3375.550 3370.800 3375.870 3371.060 ;
        RECT 3375.640 3370.040 3375.780 3370.800 ;
        RECT 3375.550 3369.780 3375.870 3370.040 ;
        RECT 3375.550 3257.100 3375.870 3257.160 ;
        RECT 3376.930 3257.100 3377.250 3257.160 ;
        RECT 3375.550 3256.960 3377.250 3257.100 ;
        RECT 3375.550 3256.900 3375.870 3256.960 ;
        RECT 3376.930 3256.900 3377.250 3256.960 ;
        RECT 3375.550 3237.380 3375.870 3237.440 ;
        RECT 3376.930 3237.380 3377.250 3237.440 ;
        RECT 3375.550 3237.240 3377.250 3237.380 ;
        RECT 3375.550 3237.180 3375.870 3237.240 ;
        RECT 3376.930 3237.180 3377.250 3237.240 ;
        RECT 208.910 3069.420 209.230 3069.480 ;
        RECT 211.670 3069.420 211.990 3069.480 ;
        RECT 208.910 3069.280 211.990 3069.420 ;
        RECT 208.910 3069.220 209.230 3069.280 ;
        RECT 211.670 3069.220 211.990 3069.280 ;
        RECT 3375.550 3028.960 3375.870 3029.020 ;
        RECT 3377.850 3028.960 3378.170 3029.020 ;
        RECT 3375.550 3028.820 3378.170 3028.960 ;
        RECT 3375.550 3028.760 3375.870 3028.820 ;
        RECT 3377.850 3028.760 3378.170 3028.820 ;
        RECT 3375.550 3009.240 3375.870 3009.300 ;
        RECT 3376.930 3009.240 3377.250 3009.300 ;
        RECT 3375.550 3009.100 3377.250 3009.240 ;
        RECT 3375.550 3009.040 3375.870 3009.100 ;
        RECT 3376.930 3009.040 3377.250 3009.100 ;
        RECT 3375.550 2807.620 3375.870 2807.680 ;
        RECT 3376.930 2807.620 3377.250 2807.680 ;
        RECT 3375.550 2807.480 3377.250 2807.620 ;
        RECT 3375.550 2807.420 3375.870 2807.480 ;
        RECT 3376.930 2807.420 3377.250 2807.480 ;
        RECT 3375.550 2785.860 3375.870 2785.920 ;
        RECT 3376.930 2785.860 3377.250 2785.920 ;
        RECT 3375.550 2785.720 3377.250 2785.860 ;
        RECT 3375.550 2785.660 3375.870 2785.720 ;
        RECT 3376.930 2785.660 3377.250 2785.720 ;
        RECT 3375.550 1694.120 3375.870 1694.180 ;
        RECT 3376.930 1694.120 3377.250 1694.180 ;
        RECT 3375.550 1693.980 3377.250 1694.120 ;
        RECT 3375.550 1693.920 3375.870 1693.980 ;
        RECT 3376.930 1693.920 3377.250 1693.980 ;
        RECT 3375.090 1671.340 3375.410 1671.400 ;
        RECT 3376.930 1671.340 3377.250 1671.400 ;
        RECT 3375.090 1671.200 3377.250 1671.340 ;
        RECT 3375.090 1671.140 3375.410 1671.200 ;
        RECT 3376.930 1671.140 3377.250 1671.200 ;
        RECT 208.910 1593.820 209.230 1593.880 ;
        RECT 211.670 1593.820 211.990 1593.880 ;
        RECT 208.910 1593.680 211.990 1593.820 ;
        RECT 208.910 1593.620 209.230 1593.680 ;
        RECT 211.670 1593.620 211.990 1593.680 ;
        RECT 208.910 1567.640 209.230 1567.700 ;
        RECT 211.670 1567.640 211.990 1567.700 ;
        RECT 208.910 1567.500 211.990 1567.640 ;
        RECT 208.910 1567.440 209.230 1567.500 ;
        RECT 211.670 1567.440 211.990 1567.500 ;
        RECT 3375.090 1470.740 3375.410 1470.800 ;
        RECT 3376.930 1470.740 3377.250 1470.800 ;
        RECT 3375.090 1470.600 3377.250 1470.740 ;
        RECT 3375.090 1470.540 3375.410 1470.600 ;
        RECT 3376.930 1470.540 3377.250 1470.600 ;
        RECT 208.910 1372.820 209.230 1372.880 ;
        RECT 211.670 1372.820 211.990 1372.880 ;
        RECT 208.910 1372.680 211.990 1372.820 ;
        RECT 208.910 1372.620 209.230 1372.680 ;
        RECT 211.670 1372.620 211.990 1372.680 ;
        RECT 208.910 1353.100 209.230 1353.160 ;
        RECT 211.670 1353.100 211.990 1353.160 ;
        RECT 208.910 1352.960 211.990 1353.100 ;
        RECT 208.910 1352.900 209.230 1352.960 ;
        RECT 211.670 1352.900 211.990 1352.960 ;
        RECT 3375.550 1243.960 3375.870 1244.020 ;
        RECT 3376.930 1243.960 3377.250 1244.020 ;
        RECT 3375.550 1243.820 3377.250 1243.960 ;
        RECT 3375.550 1243.760 3375.870 1243.820 ;
        RECT 3376.930 1243.760 3377.250 1243.820 ;
        RECT 208.910 1162.020 209.230 1162.080 ;
        RECT 211.670 1162.020 211.990 1162.080 ;
        RECT 208.910 1161.880 211.990 1162.020 ;
        RECT 208.910 1161.820 209.230 1161.880 ;
        RECT 211.670 1161.820 211.990 1161.880 ;
        RECT 208.910 1135.500 209.230 1135.560 ;
        RECT 211.670 1135.500 211.990 1135.560 ;
        RECT 208.910 1135.360 211.990 1135.500 ;
        RECT 208.910 1135.300 209.230 1135.360 ;
        RECT 211.670 1135.300 211.990 1135.360 ;
        RECT 3375.550 1017.520 3375.870 1017.580 ;
        RECT 3376.470 1017.520 3376.790 1017.580 ;
        RECT 3375.550 1017.380 3376.790 1017.520 ;
        RECT 3375.550 1017.320 3375.870 1017.380 ;
        RECT 3376.470 1017.320 3376.790 1017.380 ;
        RECT 208.910 940.680 209.230 940.740 ;
        RECT 211.670 940.680 211.990 940.740 ;
        RECT 208.910 940.540 211.990 940.680 ;
        RECT 208.910 940.480 209.230 940.540 ;
        RECT 211.670 940.480 211.990 940.540 ;
        RECT 208.910 920.960 209.230 921.020 ;
        RECT 211.670 920.960 211.990 921.020 ;
        RECT 208.910 920.820 211.990 920.960 ;
        RECT 208.910 920.760 209.230 920.820 ;
        RECT 211.670 920.760 211.990 920.820 ;
        RECT 3375.090 565.660 3375.410 565.720 ;
        RECT 3376.930 565.660 3377.250 565.720 ;
        RECT 3375.090 565.520 3377.250 565.660 ;
        RECT 3375.090 565.460 3375.410 565.520 ;
        RECT 3376.930 565.460 3377.250 565.520 ;
        RECT 3375.090 544.240 3375.410 544.300 ;
        RECT 3376.930 544.240 3377.250 544.300 ;
        RECT 3375.090 544.100 3377.250 544.240 ;
        RECT 3375.090 544.040 3375.410 544.100 ;
        RECT 3376.930 544.040 3377.250 544.100 ;
        RECT 2637.250 224.980 2637.570 225.040 ;
        RECT 3375.090 224.980 3375.410 225.040 ;
        RECT 2637.250 224.840 3375.410 224.980 ;
        RECT 2637.250 224.780 2637.570 224.840 ;
        RECT 3375.090 224.780 3375.410 224.840 ;
        RECT 2067.770 221.920 2068.090 221.980 ;
        RECT 2089.390 221.920 2089.710 221.980 ;
        RECT 2341.470 221.920 2341.790 221.980 ;
        RECT 2363.090 221.920 2363.410 221.980 ;
        RECT 2615.630 221.920 2615.950 221.980 ;
        RECT 2637.250 221.920 2637.570 221.980 ;
        RECT 2067.770 221.780 2637.570 221.920 ;
        RECT 2067.770 221.720 2068.090 221.780 ;
        RECT 2089.390 221.720 2089.710 221.780 ;
        RECT 2341.470 221.720 2341.790 221.780 ;
        RECT 2363.090 221.720 2363.410 221.780 ;
        RECT 2615.630 221.720 2615.950 221.780 ;
        RECT 2637.250 221.720 2637.570 221.780 ;
        RECT 998.270 221.580 998.590 221.640 ;
        RECT 1519.450 221.580 1519.770 221.640 ;
        RECT 1541.070 221.580 1541.390 221.640 ;
        RECT 1793.610 221.580 1793.930 221.640 ;
        RECT 1815.230 221.580 1815.550 221.640 ;
        RECT 2067.860 221.580 2068.000 221.720 ;
        RECT 998.270 221.440 2068.000 221.580 ;
        RECT 998.270 221.380 998.590 221.440 ;
        RECT 1519.450 221.380 1519.770 221.440 ;
        RECT 1541.070 221.380 1541.390 221.440 ;
        RECT 1793.610 221.380 1793.930 221.440 ;
        RECT 1815.230 221.380 1815.550 221.440 ;
        RECT 211.670 210.360 211.990 210.420 ;
        RECT 725.490 210.360 725.810 210.420 ;
        RECT 211.670 210.220 725.810 210.360 ;
        RECT 211.670 210.160 211.990 210.220 ;
        RECT 725.490 210.160 725.810 210.220 ;
        RECT 930.650 209.340 930.970 209.400 ;
        RECT 976.190 209.340 976.510 209.400 ;
        RECT 997.810 209.340 998.130 209.400 ;
        RECT 930.650 209.200 998.130 209.340 ;
        RECT 930.650 209.140 930.970 209.200 ;
        RECT 976.190 209.140 976.510 209.200 ;
        RECT 997.810 209.140 998.130 209.200 ;
        RECT 725.490 207.300 725.810 207.360 ;
        RECT 930.650 207.300 930.970 207.360 ;
        RECT 725.490 207.160 930.970 207.300 ;
        RECT 725.490 207.100 725.810 207.160 ;
        RECT 930.650 207.100 930.970 207.160 ;
      LAYER via ;
        RECT 1423.340 4976.280 1423.600 4976.540 ;
        RECT 1444.960 4976.280 1445.220 4976.540 ;
        RECT 651.460 4975.940 651.720 4976.200 ;
        RECT 673.080 4975.940 673.340 4976.200 ;
        RECT 2634.520 4975.940 2634.780 4976.200 ;
        RECT 2656.140 4975.940 2656.400 4976.200 ;
        RECT 394.320 4967.780 394.580 4968.040 ;
        RECT 415.940 4967.780 416.200 4968.040 ;
        RECT 1443.120 4967.100 1443.380 4967.360 ;
        RECT 1444.960 4967.100 1445.220 4967.360 ;
        RECT 1932.560 4967.100 1932.820 4967.360 ;
        RECT 1953.260 4967.100 1953.520 4967.360 ;
        RECT 415.940 4966.760 416.200 4967.020 ;
        RECT 651.460 4966.760 651.720 4967.020 ;
        RECT 908.600 4966.760 908.860 4967.020 ;
        RECT 930.220 4966.760 930.480 4967.020 ;
        RECT 1165.280 4966.760 1165.540 4967.020 ;
        RECT 1186.900 4966.760 1187.160 4967.020 ;
        RECT 1954.640 4966.760 1954.900 4967.020 ;
        RECT 2377.380 4966.760 2377.640 4967.020 ;
        RECT 2399.000 4966.760 2399.260 4967.020 ;
        RECT 2634.520 4966.760 2634.780 4967.020 ;
        RECT 3143.280 4966.760 3143.540 4967.020 ;
        RECT 3164.900 4966.760 3165.160 4967.020 ;
        RECT 1443.120 4966.420 1443.380 4966.680 ;
        RECT 218.140 4965.400 218.400 4965.660 ;
        RECT 394.320 4965.400 394.580 4965.660 ;
        RECT 3164.900 4964.720 3165.160 4964.980 ;
        RECT 3371.900 4964.720 3372.160 4964.980 ;
        RECT 3371.900 4836.880 3372.160 4837.140 ;
        RECT 3376.040 4836.880 3376.300 4837.140 ;
        RECT 3376.040 4826.340 3376.300 4826.600 ;
        RECT 3376.960 4826.340 3377.220 4826.600 ;
        RECT 208.940 4806.620 209.200 4806.880 ;
        RECT 211.700 4806.620 211.960 4806.880 ;
        RECT 218.140 4806.620 218.400 4806.880 ;
        RECT 3375.120 4378.900 3375.380 4379.160 ;
        RECT 3376.960 4378.900 3377.220 4379.160 ;
        RECT 208.940 3959.680 209.200 3959.940 ;
        RECT 212.620 3959.680 212.880 3959.940 ;
        RECT 208.940 3933.160 209.200 3933.420 ;
        RECT 211.700 3933.160 211.960 3933.420 ;
        RECT 3376.040 3932.820 3376.300 3933.080 ;
        RECT 3376.960 3932.820 3377.220 3933.080 ;
        RECT 3376.040 3913.440 3376.300 3913.700 ;
        RECT 3376.960 3913.440 3377.220 3913.700 ;
        RECT 208.940 3738.340 209.200 3738.600 ;
        RECT 211.700 3738.340 211.960 3738.600 ;
        RECT 208.940 3718.960 209.200 3719.220 ;
        RECT 211.700 3718.960 211.960 3719.220 ;
        RECT 3375.580 3705.020 3375.840 3705.280 ;
        RECT 3377.880 3705.020 3378.140 3705.280 ;
        RECT 3375.580 3684.960 3375.840 3685.220 ;
        RECT 3376.960 3684.960 3377.220 3685.220 ;
        RECT 211.700 3528.900 211.960 3529.160 ;
        RECT 208.940 3527.540 209.200 3527.800 ;
        RECT 211.700 3527.540 211.960 3527.800 ;
        RECT 3375.120 3479.600 3375.380 3479.860 ;
        RECT 3376.960 3479.600 3377.220 3479.860 ;
        RECT 3375.120 3460.220 3375.380 3460.480 ;
        RECT 3376.960 3460.220 3377.220 3460.480 ;
        RECT 3375.580 3370.800 3375.840 3371.060 ;
        RECT 3375.580 3369.780 3375.840 3370.040 ;
        RECT 3375.580 3256.900 3375.840 3257.160 ;
        RECT 3376.960 3256.900 3377.220 3257.160 ;
        RECT 3375.580 3237.180 3375.840 3237.440 ;
        RECT 3376.960 3237.180 3377.220 3237.440 ;
        RECT 208.940 3069.220 209.200 3069.480 ;
        RECT 211.700 3069.220 211.960 3069.480 ;
        RECT 3375.580 3028.760 3375.840 3029.020 ;
        RECT 3377.880 3028.760 3378.140 3029.020 ;
        RECT 3375.580 3009.040 3375.840 3009.300 ;
        RECT 3376.960 3009.040 3377.220 3009.300 ;
        RECT 3375.580 2807.420 3375.840 2807.680 ;
        RECT 3376.960 2807.420 3377.220 2807.680 ;
        RECT 3375.580 2785.660 3375.840 2785.920 ;
        RECT 3376.960 2785.660 3377.220 2785.920 ;
        RECT 3375.580 1693.920 3375.840 1694.180 ;
        RECT 3376.960 1693.920 3377.220 1694.180 ;
        RECT 3375.120 1671.140 3375.380 1671.400 ;
        RECT 3376.960 1671.140 3377.220 1671.400 ;
        RECT 208.940 1593.620 209.200 1593.880 ;
        RECT 211.700 1593.620 211.960 1593.880 ;
        RECT 208.940 1567.440 209.200 1567.700 ;
        RECT 211.700 1567.440 211.960 1567.700 ;
        RECT 3375.120 1470.540 3375.380 1470.800 ;
        RECT 3376.960 1470.540 3377.220 1470.800 ;
        RECT 208.940 1372.620 209.200 1372.880 ;
        RECT 211.700 1372.620 211.960 1372.880 ;
        RECT 208.940 1352.900 209.200 1353.160 ;
        RECT 211.700 1352.900 211.960 1353.160 ;
        RECT 3375.580 1243.760 3375.840 1244.020 ;
        RECT 3376.960 1243.760 3377.220 1244.020 ;
        RECT 208.940 1161.820 209.200 1162.080 ;
        RECT 211.700 1161.820 211.960 1162.080 ;
        RECT 208.940 1135.300 209.200 1135.560 ;
        RECT 211.700 1135.300 211.960 1135.560 ;
        RECT 3375.580 1017.320 3375.840 1017.580 ;
        RECT 3376.500 1017.320 3376.760 1017.580 ;
        RECT 208.940 940.480 209.200 940.740 ;
        RECT 211.700 940.480 211.960 940.740 ;
        RECT 208.940 920.760 209.200 921.020 ;
        RECT 211.700 920.760 211.960 921.020 ;
        RECT 3375.120 565.460 3375.380 565.720 ;
        RECT 3376.960 565.460 3377.220 565.720 ;
        RECT 3375.120 544.040 3375.380 544.300 ;
        RECT 3376.960 544.040 3377.220 544.300 ;
        RECT 2637.280 224.780 2637.540 225.040 ;
        RECT 3375.120 224.780 3375.380 225.040 ;
        RECT 2067.800 221.720 2068.060 221.980 ;
        RECT 2089.420 221.720 2089.680 221.980 ;
        RECT 2341.500 221.720 2341.760 221.980 ;
        RECT 2363.120 221.720 2363.380 221.980 ;
        RECT 2615.660 221.720 2615.920 221.980 ;
        RECT 2637.280 221.720 2637.540 221.980 ;
        RECT 998.300 221.380 998.560 221.640 ;
        RECT 1519.480 221.380 1519.740 221.640 ;
        RECT 1541.100 221.380 1541.360 221.640 ;
        RECT 1793.640 221.380 1793.900 221.640 ;
        RECT 1815.260 221.380 1815.520 221.640 ;
        RECT 211.700 210.160 211.960 210.420 ;
        RECT 725.520 210.160 725.780 210.420 ;
        RECT 930.680 209.140 930.940 209.400 ;
        RECT 976.220 209.140 976.480 209.400 ;
        RECT 997.840 209.140 998.100 209.400 ;
        RECT 725.520 207.100 725.780 207.360 ;
        RECT 930.680 207.100 930.940 207.360 ;
      LAYER met2 ;
        RECT 394.445 4977.260 394.725 4979.435 ;
        RECT 416.065 4977.260 416.345 4979.435 ;
        RECT 394.380 4977.035 394.725 4977.260 ;
        RECT 416.000 4977.035 416.345 4977.260 ;
        RECT 651.445 4977.035 651.725 4979.435 ;
        RECT 673.065 4977.035 673.345 4979.435 ;
        RECT 908.445 4977.330 908.725 4979.435 ;
        RECT 930.065 4977.330 930.345 4979.435 ;
        RECT 1165.445 4977.330 1165.725 4979.435 ;
        RECT 1187.065 4977.330 1187.345 4979.435 ;
        RECT 908.445 4977.035 908.800 4977.330 ;
        RECT 930.065 4977.035 930.420 4977.330 ;
        RECT 394.380 4968.070 394.520 4977.035 ;
        RECT 416.000 4968.070 416.140 4977.035 ;
        RECT 651.520 4976.230 651.660 4977.035 ;
        RECT 673.140 4976.230 673.280 4977.035 ;
        RECT 651.460 4975.910 651.720 4976.230 ;
        RECT 673.080 4975.910 673.340 4976.230 ;
        RECT 394.320 4967.750 394.580 4968.070 ;
        RECT 415.940 4967.750 416.200 4968.070 ;
        RECT 394.380 4965.690 394.520 4967.750 ;
        RECT 416.000 4967.050 416.140 4967.750 ;
        RECT 651.520 4967.050 651.660 4975.910 ;
        RECT 908.660 4967.050 908.800 4977.035 ;
        RECT 930.280 4967.050 930.420 4977.035 ;
        RECT 1165.340 4977.035 1165.725 4977.330 ;
        RECT 1186.960 4977.035 1187.345 4977.330 ;
        RECT 1423.445 4977.260 1423.725 4979.435 ;
        RECT 1445.065 4977.260 1445.345 4979.435 ;
        RECT 1423.400 4977.035 1423.725 4977.260 ;
        RECT 1445.020 4977.035 1445.345 4977.260 ;
        RECT 1932.445 4977.260 1932.725 4979.435 ;
        RECT 1954.065 4977.330 1954.345 4979.435 ;
        RECT 1932.445 4977.035 1932.760 4977.260 ;
        RECT 1165.340 4967.050 1165.480 4977.035 ;
        RECT 1186.960 4967.050 1187.100 4977.035 ;
        RECT 1423.400 4976.570 1423.540 4977.035 ;
        RECT 1445.020 4976.570 1445.160 4977.035 ;
        RECT 1423.340 4976.250 1423.600 4976.570 ;
        RECT 1444.960 4976.250 1445.220 4976.570 ;
        RECT 1445.020 4967.390 1445.160 4976.250 ;
        RECT 1932.620 4967.390 1932.760 4977.035 ;
        RECT 1953.320 4977.190 1954.345 4977.330 ;
        RECT 2377.445 4977.260 2377.725 4979.435 ;
        RECT 2399.065 4977.260 2399.345 4979.435 ;
        RECT 1953.320 4967.390 1953.460 4977.190 ;
        RECT 1954.065 4977.035 1954.345 4977.190 ;
        RECT 2377.440 4977.035 2377.725 4977.260 ;
        RECT 2399.060 4977.035 2399.345 4977.260 ;
        RECT 2634.445 4977.035 2634.725 4979.435 ;
        RECT 2656.065 4977.035 2656.345 4979.435 ;
        RECT 3143.445 4977.330 3143.725 4979.435 ;
        RECT 3165.065 4977.330 3165.345 4979.435 ;
        RECT 3143.340 4977.035 3143.725 4977.330 ;
        RECT 3164.960 4977.035 3165.345 4977.330 ;
        RECT 1443.120 4967.070 1443.380 4967.390 ;
        RECT 1444.960 4967.070 1445.220 4967.390 ;
        RECT 1932.560 4967.070 1932.820 4967.390 ;
        RECT 1953.260 4967.130 1953.520 4967.390 ;
        RECT 1953.260 4967.070 1954.840 4967.130 ;
        RECT 415.940 4966.730 416.200 4967.050 ;
        RECT 651.460 4966.730 651.720 4967.050 ;
        RECT 908.600 4966.730 908.860 4967.050 ;
        RECT 930.220 4966.730 930.480 4967.050 ;
        RECT 1165.280 4966.730 1165.540 4967.050 ;
        RECT 1186.900 4966.730 1187.160 4967.050 ;
        RECT 1443.180 4966.710 1443.320 4967.070 ;
        RECT 1953.320 4967.050 1954.840 4967.070 ;
        RECT 2377.440 4967.050 2377.580 4977.035 ;
        RECT 2399.060 4967.050 2399.200 4977.035 ;
        RECT 2634.580 4976.230 2634.720 4977.035 ;
        RECT 2656.200 4976.230 2656.340 4977.035 ;
        RECT 2634.520 4975.910 2634.780 4976.230 ;
        RECT 2656.140 4975.910 2656.400 4976.230 ;
        RECT 2634.580 4967.050 2634.720 4975.910 ;
        RECT 3143.340 4967.050 3143.480 4977.035 ;
        RECT 3164.960 4967.050 3165.100 4977.035 ;
        RECT 1953.320 4966.990 1954.900 4967.050 ;
        RECT 1954.640 4966.730 1954.900 4966.990 ;
        RECT 2377.380 4966.730 2377.640 4967.050 ;
        RECT 2399.000 4966.730 2399.260 4967.050 ;
        RECT 2634.520 4966.730 2634.780 4967.050 ;
        RECT 3143.280 4966.730 3143.540 4967.050 ;
        RECT 3164.900 4966.730 3165.160 4967.050 ;
        RECT 1443.120 4966.390 1443.380 4966.710 ;
        RECT 218.140 4965.370 218.400 4965.690 ;
        RECT 394.320 4965.370 394.580 4965.690 ;
        RECT 218.200 4806.910 218.340 4965.370 ;
        RECT 3164.960 4965.010 3165.100 4966.730 ;
        RECT 3164.900 4964.690 3165.160 4965.010 ;
        RECT 3371.900 4964.690 3372.160 4965.010 ;
        RECT 3371.960 4837.170 3372.100 4964.690 ;
        RECT 3371.900 4836.850 3372.160 4837.170 ;
        RECT 3376.040 4836.850 3376.300 4837.170 ;
        RECT 3376.100 4826.630 3376.240 4836.850 ;
        RECT 3376.040 4826.370 3376.300 4826.630 ;
        RECT 3375.180 4826.310 3376.300 4826.370 ;
        RECT 3376.960 4826.310 3377.220 4826.630 ;
        RECT 3375.180 4826.230 3376.240 4826.310 ;
        RECT 3375.180 4816.270 3375.320 4826.230 ;
        RECT 3377.020 4824.555 3377.160 4826.310 ;
        RECT 3377.020 4824.415 3379.435 4824.555 ;
        RECT 3377.035 4824.275 3379.435 4824.415 ;
        RECT 3375.180 4816.130 3375.780 4816.270 ;
        RECT 208.940 4806.590 209.200 4806.910 ;
        RECT 211.700 4806.590 211.960 4806.910 ;
        RECT 218.140 4806.590 218.400 4806.910 ;
        RECT 209.000 4806.345 209.140 4806.590 ;
        RECT 208.565 4806.065 210.965 4806.345 ;
        RECT 211.760 4786.930 211.900 4806.590 ;
        RECT 3375.640 4800.530 3375.780 4816.130 ;
        RECT 3377.035 4802.795 3379.435 4802.935 ;
        RECT 3377.020 4802.655 3379.435 4802.795 ;
        RECT 3377.020 4800.530 3377.160 4802.655 ;
        RECT 3375.640 4800.390 3377.160 4800.530 ;
        RECT 209.000 4786.790 212.820 4786.930 ;
        RECT 209.000 4784.725 209.140 4786.790 ;
        RECT 208.565 4784.445 210.965 4784.725 ;
        RECT 212.680 3959.970 212.820 4786.790 ;
        RECT 3375.640 4767.970 3375.780 4800.390 ;
        RECT 3375.180 4767.830 3375.780 4767.970 ;
        RECT 3375.180 4379.190 3375.320 4767.830 ;
        RECT 3375.120 4378.870 3375.380 4379.190 ;
        RECT 3376.960 4378.870 3377.220 4379.190 ;
        RECT 3377.020 4378.555 3377.160 4378.870 ;
        RECT 3377.020 4378.275 3379.435 4378.555 ;
        RECT 3377.020 4376.210 3377.160 4378.275 ;
        RECT 3376.560 4376.070 3377.160 4376.210 ;
        RECT 3376.560 4356.490 3376.700 4376.070 ;
        RECT 3377.035 4356.795 3379.435 4356.935 ;
        RECT 3377.020 4356.655 3379.435 4356.795 ;
        RECT 3377.020 4356.490 3377.160 4356.655 ;
        RECT 3376.100 4356.350 3377.160 4356.490 ;
        RECT 208.940 3959.650 209.200 3959.970 ;
        RECT 212.620 3959.650 212.880 3959.970 ;
        RECT 209.000 3957.345 209.140 3959.650 ;
        RECT 208.565 3957.065 210.965 3957.345 ;
        RECT 212.680 3946.870 212.820 3959.650 ;
        RECT 211.760 3946.730 212.820 3946.870 ;
        RECT 208.565 3935.445 210.965 3935.725 ;
        RECT 208.610 3935.430 209.140 3935.445 ;
        RECT 209.000 3933.450 209.140 3935.430 ;
        RECT 211.760 3933.450 211.900 3946.730 ;
        RECT 208.940 3933.130 209.200 3933.450 ;
        RECT 211.700 3933.130 211.960 3933.450 ;
        RECT 208.565 3741.065 210.965 3741.345 ;
        RECT 209.000 3738.630 209.140 3741.065 ;
        RECT 211.760 3738.630 211.900 3933.130 ;
        RECT 3376.100 3933.110 3376.240 4356.350 ;
        RECT 3376.040 3932.790 3376.300 3933.110 ;
        RECT 3376.960 3932.790 3377.220 3933.110 ;
        RECT 3376.100 3913.730 3376.240 3932.790 ;
        RECT 3377.020 3932.555 3377.160 3932.790 ;
        RECT 3377.020 3932.415 3379.435 3932.555 ;
        RECT 3377.035 3932.275 3379.435 3932.415 ;
        RECT 3376.040 3913.410 3376.300 3913.730 ;
        RECT 3376.960 3913.410 3377.220 3913.730 ;
        RECT 3376.100 3913.130 3376.240 3913.410 ;
        RECT 3375.640 3912.990 3376.240 3913.130 ;
        RECT 208.940 3738.310 209.200 3738.630 ;
        RECT 211.700 3738.310 211.960 3738.630 ;
        RECT 208.565 3719.445 210.965 3719.725 ;
        RECT 209.000 3719.250 209.140 3719.445 ;
        RECT 211.760 3719.250 211.900 3738.310 ;
        RECT 208.940 3718.930 209.200 3719.250 ;
        RECT 211.700 3718.930 211.960 3719.250 ;
        RECT 211.760 3529.190 211.900 3718.930 ;
        RECT 3375.640 3705.310 3375.780 3912.990 ;
        RECT 3377.020 3910.935 3377.160 3913.410 ;
        RECT 3377.020 3910.795 3379.435 3910.935 ;
        RECT 3377.035 3910.655 3379.435 3910.795 ;
        RECT 3377.035 3707.415 3379.435 3707.555 ;
        RECT 3377.020 3707.275 3379.435 3707.415 ;
        RECT 3377.020 3705.370 3377.160 3707.275 ;
        RECT 3377.020 3705.310 3378.080 3705.370 ;
        RECT 3375.580 3704.990 3375.840 3705.310 ;
        RECT 3377.020 3705.230 3378.140 3705.310 ;
        RECT 3377.880 3704.990 3378.140 3705.230 ;
        RECT 3375.640 3685.250 3375.780 3704.990 ;
        RECT 3377.035 3685.795 3379.435 3685.935 ;
        RECT 3377.020 3685.655 3379.435 3685.795 ;
        RECT 3377.020 3685.250 3377.160 3685.655 ;
        RECT 3375.580 3684.930 3375.840 3685.250 ;
        RECT 3376.960 3684.930 3377.220 3685.250 ;
        RECT 211.700 3528.870 211.960 3529.190 ;
        RECT 208.940 3527.510 209.200 3527.830 ;
        RECT 211.700 3527.510 211.960 3527.830 ;
        RECT 209.000 3525.345 209.140 3527.510 ;
        RECT 208.565 3525.065 210.965 3525.345 ;
        RECT 211.760 3512.170 211.900 3527.510 ;
        RECT 211.300 3512.030 211.900 3512.170 ;
        RECT 208.610 3503.725 209.140 3503.770 ;
        RECT 208.565 3503.445 210.965 3503.725 ;
        RECT 209.000 3503.090 209.140 3503.445 ;
        RECT 211.300 3503.090 211.440 3512.030 ;
        RECT 209.000 3502.950 211.900 3503.090 ;
        RECT 208.565 3309.065 210.965 3309.345 ;
        RECT 209.460 3308.610 209.600 3309.065 ;
        RECT 211.760 3308.610 211.900 3502.950 ;
        RECT 3375.640 3479.970 3375.780 3684.930 ;
        RECT 3377.035 3482.415 3379.435 3482.555 ;
        RECT 3375.180 3479.890 3375.780 3479.970 ;
        RECT 3377.020 3482.275 3379.435 3482.415 ;
        RECT 3377.020 3479.890 3377.160 3482.275 ;
        RECT 3375.120 3479.830 3375.780 3479.890 ;
        RECT 3375.120 3479.570 3375.380 3479.830 ;
        RECT 3376.960 3479.570 3377.220 3479.890 ;
        RECT 3375.180 3460.510 3375.320 3479.570 ;
        RECT 3377.035 3460.860 3379.435 3460.935 ;
        RECT 3377.020 3460.655 3379.435 3460.860 ;
        RECT 3377.020 3460.510 3377.160 3460.655 ;
        RECT 3375.120 3460.190 3375.380 3460.510 ;
        RECT 3376.960 3460.190 3377.220 3460.510 ;
        RECT 3375.180 3415.570 3375.320 3460.190 ;
        RECT 3375.180 3415.430 3375.780 3415.570 ;
        RECT 3375.640 3371.090 3375.780 3415.430 ;
        RECT 3375.580 3370.770 3375.840 3371.090 ;
        RECT 3375.580 3369.750 3375.840 3370.070 ;
        RECT 209.460 3308.470 211.900 3308.610 ;
        RECT 208.565 3287.445 210.965 3287.725 ;
        RECT 208.610 3287.390 209.140 3287.445 ;
        RECT 209.000 3286.850 209.140 3287.390 ;
        RECT 211.300 3286.850 211.440 3308.470 ;
        RECT 209.000 3286.710 211.440 3286.850 ;
        RECT 211.300 3270.670 211.440 3286.710 ;
        RECT 211.300 3270.530 211.900 3270.670 ;
        RECT 211.760 3095.770 211.900 3270.530 ;
        RECT 3375.640 3257.190 3375.780 3369.750 ;
        RECT 3375.580 3256.870 3375.840 3257.190 ;
        RECT 3376.960 3256.870 3377.220 3257.190 ;
        RECT 3375.640 3237.470 3375.780 3256.870 ;
        RECT 3377.020 3256.555 3377.160 3256.870 ;
        RECT 3377.020 3256.415 3379.435 3256.555 ;
        RECT 3377.035 3256.275 3379.435 3256.415 ;
        RECT 3375.580 3237.150 3375.840 3237.470 ;
        RECT 3376.960 3237.150 3377.220 3237.470 ;
        RECT 209.000 3095.630 211.900 3095.770 ;
        RECT 209.000 3093.345 209.140 3095.630 ;
        RECT 208.565 3093.065 210.965 3093.345 ;
        RECT 208.565 3071.445 210.965 3071.725 ;
        RECT 209.000 3069.510 209.140 3071.445 ;
        RECT 211.760 3069.510 211.900 3095.630 ;
        RECT 208.940 3069.190 209.200 3069.510 ;
        RECT 211.700 3069.190 211.960 3069.510 ;
        RECT 211.760 2880.495 211.900 3069.190 ;
        RECT 3375.640 3029.050 3375.780 3237.150 ;
        RECT 3377.020 3234.935 3377.160 3237.150 ;
        RECT 3377.020 3234.795 3379.435 3234.935 ;
        RECT 3377.035 3234.655 3379.435 3234.795 ;
        RECT 3377.035 3031.415 3379.435 3031.555 ;
        RECT 3377.020 3031.275 3379.435 3031.415 ;
        RECT 3377.020 3029.170 3377.160 3031.275 ;
        RECT 3377.020 3029.050 3378.080 3029.170 ;
        RECT 3375.580 3028.730 3375.840 3029.050 ;
        RECT 3377.020 3029.030 3378.140 3029.050 ;
        RECT 3377.880 3028.730 3378.140 3029.030 ;
        RECT 3375.640 3009.330 3375.780 3028.730 ;
        RECT 3377.035 3009.795 3379.435 3009.935 ;
        RECT 3377.020 3009.655 3379.435 3009.795 ;
        RECT 3377.020 3009.330 3377.160 3009.655 ;
        RECT 3375.580 3009.010 3375.840 3009.330 ;
        RECT 3376.960 3009.010 3377.220 3009.330 ;
        RECT 211.300 2880.355 211.900 2880.495 ;
        RECT 208.565 2877.065 210.965 2877.345 ;
        RECT 209.460 2876.810 209.600 2877.065 ;
        RECT 211.300 2876.810 211.440 2880.355 ;
        RECT 209.460 2876.670 211.440 2876.810 ;
        RECT 208.610 2855.725 209.600 2855.730 ;
        RECT 208.565 2855.445 210.965 2855.725 ;
        RECT 209.460 2855.050 209.600 2855.445 ;
        RECT 211.300 2855.050 211.440 2876.670 ;
        RECT 209.460 2854.910 211.440 2855.050 ;
        RECT 211.300 2787.670 211.440 2854.910 ;
        RECT 3375.640 2807.710 3375.780 3009.010 ;
        RECT 3375.580 2807.390 3375.840 2807.710 ;
        RECT 3376.960 2807.390 3377.220 2807.710 ;
        RECT 211.300 2787.530 211.900 2787.670 ;
        RECT 211.760 2663.970 211.900 2787.530 ;
        RECT 3375.640 2785.950 3375.780 2807.390 ;
        RECT 3377.020 2805.555 3377.160 2807.390 ;
        RECT 3377.020 2805.340 3379.435 2805.555 ;
        RECT 3377.035 2805.275 3379.435 2805.340 ;
        RECT 3375.580 2785.630 3375.840 2785.950 ;
        RECT 3376.960 2785.630 3377.220 2785.950 ;
        RECT 3377.020 2783.935 3377.160 2785.630 ;
        RECT 3377.020 2783.795 3379.435 2783.935 ;
        RECT 3377.035 2783.655 3379.435 2783.795 ;
        RECT 209.000 2663.830 211.900 2663.970 ;
        RECT 209.000 2661.345 209.140 2663.830 ;
        RECT 208.565 2661.065 210.965 2661.345 ;
        RECT 208.565 2639.445 210.965 2639.725 ;
        RECT 209.460 2637.450 209.600 2639.445 ;
        RECT 211.300 2637.450 211.440 2663.830 ;
        RECT 209.460 2637.310 211.440 2637.450 ;
        RECT 211.300 2024.090 211.440 2637.310 ;
        RECT 209.460 2023.950 211.440 2024.090 ;
        RECT 209.460 2023.410 209.600 2023.950 ;
        RECT 208.610 2023.345 209.600 2023.410 ;
        RECT 208.565 2023.065 210.965 2023.345 ;
        RECT 208.565 2001.445 210.965 2001.725 ;
        RECT 209.000 2000.970 209.140 2001.445 ;
        RECT 211.300 2000.970 211.440 2023.950 ;
        RECT 209.000 2000.830 211.440 2000.970 ;
        RECT 211.300 1811.930 211.440 2000.830 ;
        RECT 3376.100 1919.910 3377.160 1920.050 ;
        RECT 3376.100 1897.865 3376.240 1919.910 ;
        RECT 3377.020 1919.555 3377.160 1919.910 ;
        RECT 3377.020 1919.300 3379.435 1919.555 ;
        RECT 3377.035 1919.275 3379.435 1919.300 ;
        RECT 3377.035 1897.865 3379.435 1897.935 ;
        RECT 3376.100 1897.725 3379.435 1897.865 ;
        RECT 3376.100 1869.970 3376.240 1897.725 ;
        RECT 3377.035 1897.655 3379.435 1897.725 ;
        RECT 3375.640 1869.830 3376.240 1869.970 ;
        RECT 211.300 1811.790 211.900 1811.930 ;
        RECT 211.760 1807.850 211.900 1811.790 ;
        RECT 209.460 1807.710 211.900 1807.850 ;
        RECT 209.460 1807.345 209.600 1807.710 ;
        RECT 208.565 1807.065 210.965 1807.345 ;
        RECT 208.610 1807.030 209.600 1807.065 ;
        RECT 208.565 1785.655 210.965 1785.725 ;
        RECT 211.300 1785.655 211.440 1807.710 ;
        RECT 208.565 1785.515 211.900 1785.655 ;
        RECT 208.565 1785.445 210.965 1785.515 ;
        RECT 211.760 1593.910 211.900 1785.515 ;
        RECT 3375.640 1694.210 3375.780 1869.830 ;
        RECT 3375.580 1693.890 3375.840 1694.210 ;
        RECT 3376.960 1693.890 3377.220 1694.210 ;
        RECT 3377.020 1693.555 3377.160 1693.890 ;
        RECT 3377.020 1693.275 3379.435 1693.555 ;
        RECT 3377.020 1690.890 3377.160 1693.275 ;
        RECT 3376.560 1690.750 3377.160 1690.890 ;
        RECT 3376.560 1671.850 3376.700 1690.750 ;
        RECT 3377.035 1671.850 3379.435 1671.935 ;
        RECT 3376.560 1671.710 3379.435 1671.850 ;
        RECT 3377.020 1671.655 3379.435 1671.710 ;
        RECT 3377.020 1671.430 3377.160 1671.655 ;
        RECT 3375.120 1671.110 3375.380 1671.430 ;
        RECT 3376.960 1671.110 3377.220 1671.430 ;
        RECT 208.940 1593.590 209.200 1593.910 ;
        RECT 211.700 1593.590 211.960 1593.910 ;
        RECT 209.000 1591.345 209.140 1593.590 ;
        RECT 208.565 1591.065 210.965 1591.345 ;
        RECT 208.565 1569.445 210.965 1569.725 ;
        RECT 209.000 1567.730 209.140 1569.445 ;
        RECT 211.760 1567.730 211.900 1593.590 ;
        RECT 208.940 1567.410 209.200 1567.730 ;
        RECT 211.700 1567.410 211.960 1567.730 ;
        RECT 208.610 1375.345 209.140 1375.370 ;
        RECT 208.565 1375.065 210.965 1375.345 ;
        RECT 209.000 1372.910 209.140 1375.065 ;
        RECT 211.760 1372.910 211.900 1567.410 ;
        RECT 3375.180 1470.830 3375.320 1671.110 ;
        RECT 3375.120 1470.510 3375.380 1470.830 ;
        RECT 3376.960 1470.510 3377.220 1470.830 ;
        RECT 3377.020 1468.555 3377.160 1470.510 ;
        RECT 3377.020 1468.530 3379.435 1468.555 ;
        RECT 3376.560 1468.390 3379.435 1468.530 ;
        RECT 3376.560 1446.770 3376.700 1468.390 ;
        RECT 3377.035 1468.275 3379.435 1468.390 ;
        RECT 3377.035 1446.770 3379.435 1446.935 ;
        RECT 3376.560 1446.655 3379.435 1446.770 ;
        RECT 3376.560 1446.630 3377.160 1446.655 ;
        RECT 3377.020 1444.050 3377.160 1446.630 ;
        RECT 3375.640 1443.910 3377.160 1444.050 ;
        RECT 208.940 1372.590 209.200 1372.910 ;
        RECT 211.700 1372.590 211.960 1372.910 ;
        RECT 208.565 1353.445 210.965 1353.725 ;
        RECT 209.000 1353.190 209.140 1353.445 ;
        RECT 211.760 1353.190 211.900 1372.590 ;
        RECT 208.940 1352.870 209.200 1353.190 ;
        RECT 211.700 1352.870 211.960 1353.190 ;
        RECT 211.760 1162.110 211.900 1352.870 ;
        RECT 3375.640 1244.050 3375.780 1443.910 ;
        RECT 3375.580 1243.730 3375.840 1244.050 ;
        RECT 3376.960 1243.730 3377.220 1244.050 ;
        RECT 3375.640 1242.070 3375.780 1243.730 ;
        RECT 3377.020 1243.555 3377.160 1243.730 ;
        RECT 3377.020 1243.380 3379.435 1243.555 ;
        RECT 3377.035 1243.275 3379.435 1243.380 ;
        RECT 3375.640 1241.930 3376.700 1242.070 ;
        RECT 3376.560 1221.865 3376.700 1241.930 ;
        RECT 3377.035 1221.865 3379.435 1221.935 ;
        RECT 3376.560 1221.725 3379.435 1221.865 ;
        RECT 3376.560 1218.970 3376.700 1221.725 ;
        RECT 3377.035 1221.655 3379.435 1221.725 ;
        RECT 3375.640 1218.830 3376.700 1218.970 ;
        RECT 208.940 1161.790 209.200 1162.110 ;
        RECT 211.700 1161.790 211.960 1162.110 ;
        RECT 209.000 1159.345 209.140 1161.790 ;
        RECT 208.565 1159.065 210.965 1159.345 ;
        RECT 208.565 1137.445 210.965 1137.725 ;
        RECT 209.000 1135.590 209.140 1137.445 ;
        RECT 211.760 1135.590 211.900 1161.790 ;
        RECT 208.940 1135.270 209.200 1135.590 ;
        RECT 211.700 1135.270 211.960 1135.590 ;
        RECT 208.565 943.065 210.965 943.345 ;
        RECT 209.000 940.770 209.140 943.065 ;
        RECT 211.760 940.770 211.900 1135.270 ;
        RECT 3375.640 1017.610 3375.780 1218.830 ;
        RECT 3376.560 1017.610 3376.700 1017.900 ;
        RECT 3375.580 1017.290 3375.840 1017.610 ;
        RECT 3376.500 1017.485 3376.760 1017.610 ;
        RECT 3377.035 1017.485 3379.435 1017.555 ;
        RECT 3376.500 1017.345 3379.435 1017.485 ;
        RECT 3376.500 1017.290 3376.760 1017.345 ;
        RECT 3376.560 995.930 3376.700 1017.290 ;
        RECT 3377.035 1017.275 3379.435 1017.345 ;
        RECT 3377.035 995.930 3379.435 995.935 ;
        RECT 3375.640 995.790 3379.435 995.930 ;
        RECT 208.940 940.450 209.200 940.770 ;
        RECT 211.700 940.450 211.960 940.770 ;
        RECT 208.565 921.445 210.965 921.725 ;
        RECT 209.000 921.050 209.140 921.445 ;
        RECT 211.760 921.050 211.900 940.450 ;
        RECT 208.940 920.730 209.200 921.050 ;
        RECT 211.700 920.730 211.960 921.050 ;
        RECT 211.760 210.450 211.900 920.730 ;
        RECT 3375.640 793.290 3375.780 995.790 ;
        RECT 3377.035 995.655 3379.435 995.790 ;
        RECT 3375.640 793.150 3376.700 793.290 ;
        RECT 3376.560 791.930 3376.700 793.150 ;
        RECT 3377.035 792.540 3379.435 792.555 ;
        RECT 3377.020 792.275 3379.435 792.540 ;
        RECT 3377.020 791.930 3377.160 792.275 ;
        RECT 3376.560 791.790 3377.160 791.930 ;
        RECT 3376.560 770.850 3376.700 791.790 ;
        RECT 3377.035 770.850 3379.435 770.935 ;
        RECT 3375.640 770.710 3379.435 770.850 ;
        RECT 3375.640 710.770 3375.780 770.710 ;
        RECT 3377.035 770.655 3379.435 770.710 ;
        RECT 3375.180 710.630 3375.780 710.770 ;
        RECT 3375.180 565.750 3375.320 710.630 ;
        RECT 3377.035 566.415 3379.435 566.555 ;
        RECT 3377.020 566.275 3379.435 566.415 ;
        RECT 3377.020 565.750 3377.160 566.275 ;
        RECT 3375.120 565.430 3375.380 565.750 ;
        RECT 3376.960 565.430 3377.220 565.750 ;
        RECT 3375.180 544.330 3375.320 565.430 ;
        RECT 3377.035 544.795 3379.435 544.935 ;
        RECT 3377.020 544.655 3379.435 544.795 ;
        RECT 3377.020 544.330 3377.160 544.655 ;
        RECT 3375.120 544.010 3375.380 544.330 ;
        RECT 3376.960 544.010 3377.220 544.330 ;
        RECT 3375.180 225.070 3375.320 544.010 ;
        RECT 2637.280 224.750 2637.540 225.070 ;
        RECT 3375.120 224.750 3375.380 225.070 ;
        RECT 2637.340 222.010 2637.480 224.750 ;
        RECT 2067.800 221.690 2068.060 222.010 ;
        RECT 2089.420 221.690 2089.680 222.010 ;
        RECT 2341.500 221.690 2341.760 222.010 ;
        RECT 2363.120 221.690 2363.380 222.010 ;
        RECT 2615.660 221.690 2615.920 222.010 ;
        RECT 2637.280 221.690 2637.540 222.010 ;
        RECT 998.300 221.350 998.560 221.670 ;
        RECT 1519.480 221.350 1519.740 221.670 ;
        RECT 1541.100 221.350 1541.360 221.670 ;
        RECT 1793.640 221.350 1793.900 221.670 ;
        RECT 1815.260 221.350 1815.520 221.670 ;
        RECT 998.360 210.965 998.500 221.350 ;
        RECT 1519.540 210.965 1519.680 221.350 ;
        RECT 1541.160 210.965 1541.300 221.350 ;
        RECT 1793.700 210.965 1793.840 221.350 ;
        RECT 1815.320 210.965 1815.460 221.350 ;
        RECT 2067.860 210.965 2068.000 221.690 ;
        RECT 2089.480 210.965 2089.620 221.690 ;
        RECT 211.700 210.130 211.960 210.450 ;
        RECT 725.520 210.130 725.780 210.450 ;
        RECT 725.580 207.390 725.720 210.130 ;
        RECT 930.680 209.110 930.940 209.430 ;
        RECT 976.220 209.170 976.480 209.430 ;
        RECT 976.655 209.170 976.935 210.965 ;
        RECT 976.220 209.110 976.935 209.170 ;
        RECT 997.840 209.170 998.100 209.430 ;
        RECT 998.275 209.170 998.555 210.965 ;
        RECT 997.840 209.110 998.555 209.170 ;
        RECT 930.740 207.390 930.880 209.110 ;
        RECT 976.280 209.030 976.935 209.110 ;
        RECT 997.900 209.030 998.555 209.110 ;
        RECT 1519.540 209.030 1519.935 210.965 ;
        RECT 1541.160 209.030 1541.555 210.965 ;
        RECT 976.655 208.565 976.935 209.030 ;
        RECT 998.275 208.565 998.555 209.030 ;
        RECT 1519.655 208.565 1519.935 209.030 ;
        RECT 1541.275 208.565 1541.555 209.030 ;
        RECT 1793.655 208.565 1793.935 210.965 ;
        RECT 1815.275 208.565 1815.555 210.965 ;
        RECT 2067.655 209.100 2068.000 210.965 ;
        RECT 2089.275 209.100 2089.620 210.965 ;
        RECT 2341.560 210.965 2341.700 221.690 ;
        RECT 2363.180 210.965 2363.320 221.690 ;
        RECT 2615.720 210.965 2615.860 221.690 ;
        RECT 2637.340 210.965 2637.480 221.690 ;
        RECT 2067.655 208.565 2067.935 209.100 ;
        RECT 2089.275 208.565 2089.555 209.100 ;
        RECT 2341.560 209.030 2341.935 210.965 ;
        RECT 2363.180 209.030 2363.555 210.965 ;
        RECT 2341.655 208.565 2341.935 209.030 ;
        RECT 2363.275 208.565 2363.555 209.030 ;
        RECT 2615.655 208.565 2615.935 210.965 ;
        RECT 2637.275 208.565 2637.555 210.965 ;
        RECT 725.520 207.070 725.780 207.390 ;
        RECT 930.680 207.070 930.940 207.390 ;
        RECT 725.580 201.010 725.720 207.070 ;
        RECT 725.515 200.870 725.720 201.010 ;
        RECT 725.515 200.000 725.655 200.870 ;
        RECT 725.455 198.530 725.715 200.000 ;
    END
  END porb_h
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 683.565 35.715 720.750 91.545 ;
    END
  END resetb
  PIN resetb_core_h
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 708.335 190.155 709.065 200.000 ;
        RECT 708.335 189.855 709.365 190.155 ;
        RECT 708.335 189.555 709.100 189.855 ;
        RECT 709.365 189.555 709.830 189.855 ;
        RECT 708.335 189.090 709.830 189.555 ;
        RECT 709.100 185.230 709.830 189.090 ;
    END
  END resetb_core_h
  PIN vdda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 468.035 181.615 663.965 185.065 ;
    END
  END vdda
  PIN vssa
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 143.265 964.910 143.595 ;
    END
  END vssa
  PIN vssd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 467.730 158.370 664.270 158.415 ;
        RECT 467.730 153.810 664.345 158.370 ;
        RECT 467.730 153.765 664.270 153.810 ;
    END
  END vssd
  PIN vccd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 4548.330 3557.165 4602.730 ;
    END
  END vccd1_pad
  PIN vdda1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 4099.110 3553.945 4159.950 ;
    END
  END vdda1_pad
  PIN vdda1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2526.110 3553.945 2586.950 ;
    END
  END vdda1_pad2
  PIN vssa1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2885.050 5093.120 2945.890 5153.945 ;
    END
  END vssa1_pad
  PIN vssa1_pad2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3493.120 2085.110 3553.945 2145.950 ;
    END
  END vssa1_pad2
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3396.885 2151.730 3401.535 2300.270 ;
    END
  END vccd1
  PIN vdda1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3402.935 2152.035 3406.385 2299.965 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3444.405 2151.730 3444.735 2771.910 ;
    END
  END vssa1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 3390.000 2349.500 3429.600 2373.500 ;
    END
  END vssd1
  PIN vssd1_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3489.900 2309.330 3557.165 2363.730 ;
    END
  END vssd1_pad
  PIN vccd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 4570.270 98.100 4624.670 ;
    END
  END vccd2_pad
  PIN vdda2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 2422.050 94.880 2482.890 ;
    END
  END vdda2_pad
  PIN vssa2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 34.055 4145.050 94.880 4205.890 ;
    END
  END vssa2_pad
  PIN vccd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 192.515 2277.730 197.965 2416.270 ;
    END
  END vccd
  PIN vccd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 186.465 2277.730 191.115 2416.270 ;
    END
  END vccd2
  PIN vdda2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 181.615 2278.035 185.065 2415.965 ;
    END
  END vdda2
  PIN vddio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 164.665 2277.730 168.115 2416.270 ;
    END
  END vddio
  PIN vssa2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.265 2035.090 143.595 2628.610 ;
    END
  END vssa2
  PIN vssd2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.400 2204.500 198.000 2228.500 ;
    END
  END vssd2
  PIN vssd2_pad
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 30.835 2214.270 98.100 2268.670 ;
    END
  END vssd2_pad
  PIN vssio
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.035 2279.000 24.215 2280.465 ;
        RECT 0.000 2277.730 24.215 2279.000 ;
    END
  END vssio
  OBS
      LAYER nwell ;
        RECT 380.585 5161.545 461.435 5166.975 ;
        RECT 380.585 5158.475 388.515 5161.545 ;
        RECT 447.970 5158.475 461.435 5161.545 ;
        RECT 380.585 5158.230 461.435 5158.475 ;
        RECT 637.585 5161.545 718.435 5166.975 ;
        RECT 637.585 5158.475 645.515 5161.545 ;
        RECT 704.970 5158.475 718.435 5161.545 ;
        RECT 637.585 5158.230 718.435 5158.475 ;
        RECT 894.585 5161.545 975.435 5166.975 ;
        RECT 894.585 5158.475 902.515 5161.545 ;
        RECT 961.970 5158.475 975.435 5161.545 ;
        RECT 894.585 5158.230 975.435 5158.475 ;
        RECT 1151.585 5161.545 1232.435 5166.975 ;
        RECT 1151.585 5158.475 1159.515 5161.545 ;
        RECT 1218.970 5158.475 1232.435 5161.545 ;
        RECT 1151.585 5158.230 1232.435 5158.475 ;
        RECT 1409.585 5161.545 1490.435 5166.975 ;
        RECT 1409.585 5158.475 1417.515 5161.545 ;
        RECT 1476.970 5158.475 1490.435 5161.545 ;
        RECT 1409.585 5158.230 1490.435 5158.475 ;
        RECT 1918.585 5161.545 1999.435 5166.975 ;
        RECT 1918.585 5158.475 1926.515 5161.545 ;
        RECT 1985.970 5158.475 1999.435 5161.545 ;
        RECT 1918.585 5158.230 1999.435 5158.475 ;
        RECT 2363.585 5161.545 2444.435 5166.975 ;
        RECT 2363.585 5158.475 2371.515 5161.545 ;
        RECT 2430.970 5158.475 2444.435 5161.545 ;
        RECT 2363.585 5158.230 2444.435 5158.475 ;
        RECT 2620.585 5161.545 2701.435 5166.975 ;
        RECT 2620.585 5158.475 2628.515 5161.545 ;
        RECT 2687.970 5158.475 2701.435 5161.545 ;
        RECT 2620.585 5158.230 2701.435 5158.475 ;
        RECT 3129.585 5161.545 3210.435 5166.975 ;
        RECT 3129.585 5158.475 3137.515 5161.545 ;
        RECT 3196.970 5158.475 3210.435 5161.545 ;
        RECT 3129.585 5158.230 3210.435 5158.475 ;
        RECT 380.585 5156.515 461.440 5158.230 ;
        RECT 380.585 5134.690 387.385 5156.515 ;
        RECT 459.630 5134.690 461.440 5156.515 ;
        RECT 380.585 5132.880 461.440 5134.690 ;
        RECT 637.585 5156.515 718.440 5158.230 ;
        RECT 637.585 5134.690 644.385 5156.515 ;
        RECT 716.630 5134.690 718.440 5156.515 ;
        RECT 637.585 5132.880 718.440 5134.690 ;
        RECT 894.585 5156.515 975.440 5158.230 ;
        RECT 894.585 5134.690 901.385 5156.515 ;
        RECT 973.630 5134.690 975.440 5156.515 ;
        RECT 894.585 5132.880 975.440 5134.690 ;
        RECT 1151.585 5156.515 1232.440 5158.230 ;
        RECT 1151.585 5134.690 1158.385 5156.515 ;
        RECT 1230.630 5134.690 1232.440 5156.515 ;
        RECT 1151.585 5132.880 1232.440 5134.690 ;
        RECT 1409.585 5156.515 1490.440 5158.230 ;
        RECT 1409.585 5134.690 1416.385 5156.515 ;
        RECT 1488.630 5134.690 1490.440 5156.515 ;
        RECT 1409.585 5132.880 1490.440 5134.690 ;
        RECT 1918.585 5156.515 1999.440 5158.230 ;
        RECT 1918.585 5134.690 1925.385 5156.515 ;
        RECT 1997.630 5134.690 1999.440 5156.515 ;
        RECT 1918.585 5132.880 1999.440 5134.690 ;
        RECT 2363.585 5156.515 2444.440 5158.230 ;
        RECT 2363.585 5134.690 2370.385 5156.515 ;
        RECT 2442.630 5134.690 2444.440 5156.515 ;
        RECT 2363.585 5132.880 2444.440 5134.690 ;
        RECT 2620.585 5156.515 2701.440 5158.230 ;
        RECT 2620.585 5134.690 2627.385 5156.515 ;
        RECT 2699.630 5134.690 2701.440 5156.515 ;
        RECT 2620.585 5132.880 2701.440 5134.690 ;
        RECT 3129.585 5156.515 3210.440 5158.230 ;
        RECT 3129.585 5134.690 3136.385 5156.515 ;
        RECT 3208.630 5134.690 3210.440 5156.515 ;
        RECT 3129.585 5132.880 3210.440 5134.690 ;
      LAYER pwell ;
        RECT 380.710 5128.685 461.290 5132.565 ;
        RECT 637.710 5128.685 718.290 5132.565 ;
        RECT 894.710 5128.685 975.290 5132.565 ;
        RECT 1151.710 5128.685 1232.290 5132.565 ;
        RECT 1409.710 5128.685 1490.290 5132.565 ;
        RECT 1918.710 5128.685 1999.290 5132.565 ;
        RECT 2363.710 5128.685 2444.290 5132.565 ;
        RECT 2620.710 5128.685 2701.290 5132.565 ;
        RECT 3129.710 5128.685 3210.290 5132.565 ;
      LAYER nwell ;
        RECT 427.040 5128.380 461.440 5128.385 ;
        RECT 684.040 5128.380 718.440 5128.385 ;
        RECT 941.040 5128.380 975.440 5128.385 ;
        RECT 1198.040 5128.380 1232.440 5128.385 ;
        RECT 1456.040 5128.380 1490.440 5128.385 ;
        RECT 1965.040 5128.380 1999.440 5128.385 ;
        RECT 2410.040 5128.380 2444.440 5128.385 ;
        RECT 2667.040 5128.380 2701.440 5128.385 ;
        RECT 3176.040 5128.380 3210.440 5128.385 ;
        RECT 380.585 5118.665 461.440 5128.380 ;
        RECT 637.585 5118.665 718.440 5128.380 ;
        RECT 894.585 5118.665 975.440 5128.380 ;
        RECT 1151.585 5118.665 1232.440 5128.380 ;
        RECT 1409.585 5118.665 1490.440 5128.380 ;
        RECT 1918.585 5118.665 1999.440 5128.380 ;
        RECT 2363.585 5118.665 2444.440 5128.380 ;
        RECT 2620.585 5118.665 2701.440 5128.380 ;
        RECT 3129.585 5118.665 3210.440 5128.380 ;
      LAYER pwell ;
        RECT 380.785 5117.315 421.245 5118.355 ;
        RECT 447.910 5117.315 461.290 5118.355 ;
        RECT 380.785 5113.135 461.290 5117.315 ;
        RECT 380.785 5091.550 386.735 5113.135 ;
        RECT 458.865 5091.550 461.290 5113.135 ;
        RECT 380.785 5089.965 461.290 5091.550 ;
        RECT 380.785 5084.255 386.215 5089.965 ;
        RECT 420.385 5088.820 461.290 5089.965 ;
        RECT 433.880 5087.520 461.290 5088.820 ;
        RECT 457.770 5085.985 461.290 5087.520 ;
        RECT 420.385 5084.255 461.290 5085.985 ;
        RECT 380.785 5083.975 461.290 5084.255 ;
        RECT 637.785 5117.315 678.245 5118.355 ;
        RECT 704.910 5117.315 718.290 5118.355 ;
        RECT 637.785 5113.135 718.290 5117.315 ;
        RECT 637.785 5091.550 643.735 5113.135 ;
        RECT 715.865 5091.550 718.290 5113.135 ;
        RECT 637.785 5089.965 718.290 5091.550 ;
        RECT 637.785 5084.255 643.215 5089.965 ;
        RECT 677.385 5088.820 718.290 5089.965 ;
        RECT 690.880 5087.520 718.290 5088.820 ;
        RECT 714.770 5085.985 718.290 5087.520 ;
        RECT 677.385 5084.255 718.290 5085.985 ;
        RECT 637.785 5083.975 718.290 5084.255 ;
        RECT 894.785 5117.315 935.245 5118.355 ;
        RECT 961.910 5117.315 975.290 5118.355 ;
        RECT 894.785 5113.135 975.290 5117.315 ;
        RECT 894.785 5091.550 900.735 5113.135 ;
        RECT 972.865 5091.550 975.290 5113.135 ;
        RECT 894.785 5089.965 975.290 5091.550 ;
        RECT 894.785 5084.255 900.215 5089.965 ;
        RECT 934.385 5088.820 975.290 5089.965 ;
        RECT 947.880 5087.520 975.290 5088.820 ;
        RECT 971.770 5085.985 975.290 5087.520 ;
        RECT 934.385 5084.255 975.290 5085.985 ;
        RECT 894.785 5083.975 975.290 5084.255 ;
        RECT 1151.785 5117.315 1192.245 5118.355 ;
        RECT 1218.910 5117.315 1232.290 5118.355 ;
        RECT 1151.785 5113.135 1232.290 5117.315 ;
        RECT 1151.785 5091.550 1157.735 5113.135 ;
        RECT 1229.865 5091.550 1232.290 5113.135 ;
        RECT 1151.785 5089.965 1232.290 5091.550 ;
        RECT 1151.785 5084.255 1157.215 5089.965 ;
        RECT 1191.385 5088.820 1232.290 5089.965 ;
        RECT 1204.880 5087.520 1232.290 5088.820 ;
        RECT 1228.770 5085.985 1232.290 5087.520 ;
        RECT 1191.385 5084.255 1232.290 5085.985 ;
        RECT 1151.785 5083.975 1232.290 5084.255 ;
        RECT 1409.785 5117.315 1450.245 5118.355 ;
        RECT 1476.910 5117.315 1490.290 5118.355 ;
        RECT 1409.785 5113.135 1490.290 5117.315 ;
        RECT 1409.785 5091.550 1415.735 5113.135 ;
        RECT 1487.865 5091.550 1490.290 5113.135 ;
        RECT 1409.785 5089.965 1490.290 5091.550 ;
        RECT 1409.785 5084.255 1415.215 5089.965 ;
        RECT 1449.385 5088.820 1490.290 5089.965 ;
        RECT 1462.880 5087.520 1490.290 5088.820 ;
        RECT 1486.770 5085.985 1490.290 5087.520 ;
        RECT 1449.385 5084.255 1490.290 5085.985 ;
        RECT 1409.785 5083.975 1490.290 5084.255 ;
        RECT 1918.785 5117.315 1959.245 5118.355 ;
        RECT 1985.910 5117.315 1999.290 5118.355 ;
        RECT 1918.785 5113.135 1999.290 5117.315 ;
        RECT 1918.785 5091.550 1924.735 5113.135 ;
        RECT 1996.865 5091.550 1999.290 5113.135 ;
        RECT 1918.785 5089.965 1999.290 5091.550 ;
        RECT 1918.785 5084.255 1924.215 5089.965 ;
        RECT 1958.385 5088.820 1999.290 5089.965 ;
        RECT 1971.880 5087.520 1999.290 5088.820 ;
        RECT 1995.770 5085.985 1999.290 5087.520 ;
        RECT 1958.385 5084.255 1999.290 5085.985 ;
        RECT 1918.785 5083.975 1999.290 5084.255 ;
        RECT 2363.785 5117.315 2404.245 5118.355 ;
        RECT 2430.910 5117.315 2444.290 5118.355 ;
        RECT 2363.785 5113.135 2444.290 5117.315 ;
        RECT 2363.785 5091.550 2369.735 5113.135 ;
        RECT 2441.865 5091.550 2444.290 5113.135 ;
        RECT 2363.785 5089.965 2444.290 5091.550 ;
        RECT 2363.785 5084.255 2369.215 5089.965 ;
        RECT 2403.385 5088.820 2444.290 5089.965 ;
        RECT 2416.880 5087.520 2444.290 5088.820 ;
        RECT 2440.770 5085.985 2444.290 5087.520 ;
        RECT 2403.385 5084.255 2444.290 5085.985 ;
        RECT 2363.785 5083.975 2444.290 5084.255 ;
        RECT 2620.785 5117.315 2661.245 5118.355 ;
        RECT 2687.910 5117.315 2701.290 5118.355 ;
        RECT 2620.785 5113.135 2701.290 5117.315 ;
        RECT 2620.785 5091.550 2626.735 5113.135 ;
        RECT 2698.865 5091.550 2701.290 5113.135 ;
        RECT 2620.785 5089.965 2701.290 5091.550 ;
        RECT 2620.785 5084.255 2626.215 5089.965 ;
        RECT 2660.385 5088.820 2701.290 5089.965 ;
        RECT 2673.880 5087.520 2701.290 5088.820 ;
        RECT 2697.770 5085.985 2701.290 5087.520 ;
        RECT 2660.385 5084.255 2701.290 5085.985 ;
        RECT 2620.785 5083.975 2701.290 5084.255 ;
        RECT 3129.785 5117.315 3170.245 5118.355 ;
        RECT 3196.910 5117.315 3210.290 5118.355 ;
        RECT 3129.785 5113.135 3210.290 5117.315 ;
        RECT 3129.785 5091.550 3135.735 5113.135 ;
        RECT 3207.865 5091.550 3210.290 5113.135 ;
        RECT 3129.785 5089.965 3210.290 5091.550 ;
        RECT 3129.785 5084.255 3135.215 5089.965 ;
        RECT 3169.385 5088.820 3210.290 5089.965 ;
        RECT 3182.880 5087.520 3210.290 5088.820 ;
        RECT 3206.770 5085.985 3210.290 5087.520 ;
        RECT 3169.385 5084.255 3210.290 5085.985 ;
        RECT 3129.785 5083.975 3210.290 5084.255 ;
        RECT 380.785 5083.260 426.840 5083.975 ;
        RECT 637.785 5083.260 683.840 5083.975 ;
        RECT 894.785 5083.260 940.840 5083.975 ;
        RECT 1151.785 5083.260 1197.840 5083.975 ;
        RECT 1409.785 5083.260 1455.840 5083.975 ;
        RECT 1918.785 5083.260 1964.840 5083.975 ;
        RECT 2363.785 5083.260 2409.840 5083.975 ;
        RECT 2620.785 5083.260 2666.840 5083.975 ;
        RECT 3129.785 5083.260 3175.840 5083.975 ;
        RECT 380.785 5082.955 427.590 5083.260 ;
        RECT 380.785 5080.935 390.300 5082.955 ;
      LAYER nwell ;
        RECT 427.940 5082.245 461.670 5083.165 ;
        RECT 443.650 5081.735 461.670 5082.245 ;
        RECT 380.585 5079.820 383.795 5080.400 ;
        RECT 380.585 5076.485 386.975 5079.820 ;
        RECT 380.880 5076.280 386.975 5076.485 ;
        RECT 380.880 5075.740 389.420 5076.280 ;
        RECT 380.880 5074.660 389.495 5075.740 ;
        RECT 380.880 5073.580 385.530 5074.660 ;
        RECT 460.240 5072.345 461.670 5081.735 ;
      LAYER pwell ;
        RECT 637.785 5082.955 684.590 5083.260 ;
        RECT 637.785 5080.935 647.300 5082.955 ;
      LAYER nwell ;
        RECT 684.940 5082.245 718.670 5083.165 ;
        RECT 700.650 5081.735 718.670 5082.245 ;
        RECT 637.585 5079.820 640.795 5080.400 ;
        RECT 637.585 5076.485 643.975 5079.820 ;
        RECT 637.880 5076.280 643.975 5076.485 ;
        RECT 637.880 5075.740 646.420 5076.280 ;
        RECT 637.880 5074.660 646.495 5075.740 ;
        RECT 637.880 5073.580 642.530 5074.660 ;
        RECT 717.240 5072.345 718.670 5081.735 ;
      LAYER pwell ;
        RECT 894.785 5082.955 941.590 5083.260 ;
        RECT 894.785 5080.935 904.300 5082.955 ;
      LAYER nwell ;
        RECT 941.940 5082.245 975.670 5083.165 ;
        RECT 957.650 5081.735 975.670 5082.245 ;
        RECT 894.585 5079.820 897.795 5080.400 ;
        RECT 894.585 5076.485 900.975 5079.820 ;
        RECT 894.880 5076.280 900.975 5076.485 ;
        RECT 894.880 5075.740 903.420 5076.280 ;
        RECT 894.880 5074.660 903.495 5075.740 ;
        RECT 894.880 5073.580 899.530 5074.660 ;
        RECT 974.240 5072.345 975.670 5081.735 ;
      LAYER pwell ;
        RECT 1151.785 5082.955 1198.590 5083.260 ;
        RECT 1151.785 5080.935 1161.300 5082.955 ;
      LAYER nwell ;
        RECT 1198.940 5082.245 1232.670 5083.165 ;
        RECT 1214.650 5081.735 1232.670 5082.245 ;
        RECT 1151.585 5079.820 1154.795 5080.400 ;
        RECT 1151.585 5076.485 1157.975 5079.820 ;
        RECT 1151.880 5076.280 1157.975 5076.485 ;
        RECT 1151.880 5075.740 1160.420 5076.280 ;
        RECT 1151.880 5074.660 1160.495 5075.740 ;
        RECT 1151.880 5073.580 1156.530 5074.660 ;
        RECT 1231.240 5072.345 1232.670 5081.735 ;
      LAYER pwell ;
        RECT 1409.785 5082.955 1456.590 5083.260 ;
        RECT 1409.785 5080.935 1419.300 5082.955 ;
      LAYER nwell ;
        RECT 1456.940 5082.245 1490.670 5083.165 ;
        RECT 1472.650 5081.735 1490.670 5082.245 ;
        RECT 1409.585 5079.820 1412.795 5080.400 ;
        RECT 1409.585 5076.485 1415.975 5079.820 ;
        RECT 1409.880 5076.280 1415.975 5076.485 ;
        RECT 1409.880 5075.740 1418.420 5076.280 ;
        RECT 1409.880 5074.660 1418.495 5075.740 ;
        RECT 1409.880 5073.580 1414.530 5074.660 ;
        RECT 1489.240 5072.345 1490.670 5081.735 ;
      LAYER pwell ;
        RECT 1918.785 5082.955 1965.590 5083.260 ;
        RECT 1918.785 5080.935 1928.300 5082.955 ;
      LAYER nwell ;
        RECT 1965.940 5082.245 1999.670 5083.165 ;
        RECT 1981.650 5081.735 1999.670 5082.245 ;
        RECT 1918.585 5079.820 1921.795 5080.400 ;
        RECT 1918.585 5076.485 1924.975 5079.820 ;
        RECT 1918.880 5076.280 1924.975 5076.485 ;
        RECT 1918.880 5075.740 1927.420 5076.280 ;
        RECT 1918.880 5074.660 1927.495 5075.740 ;
        RECT 1918.880 5073.580 1923.530 5074.660 ;
        RECT 1998.240 5072.345 1999.670 5081.735 ;
      LAYER pwell ;
        RECT 2363.785 5082.955 2410.590 5083.260 ;
        RECT 2363.785 5080.935 2373.300 5082.955 ;
      LAYER nwell ;
        RECT 2410.940 5082.245 2444.670 5083.165 ;
        RECT 2426.650 5081.735 2444.670 5082.245 ;
        RECT 2363.585 5079.820 2366.795 5080.400 ;
        RECT 2363.585 5076.485 2369.975 5079.820 ;
        RECT 2363.880 5076.280 2369.975 5076.485 ;
        RECT 2363.880 5075.740 2372.420 5076.280 ;
        RECT 2363.880 5074.660 2372.495 5075.740 ;
        RECT 2363.880 5073.580 2368.530 5074.660 ;
        RECT 2443.240 5072.345 2444.670 5081.735 ;
      LAYER pwell ;
        RECT 2620.785 5082.955 2667.590 5083.260 ;
        RECT 2620.785 5080.935 2630.300 5082.955 ;
      LAYER nwell ;
        RECT 2667.940 5082.245 2701.670 5083.165 ;
        RECT 2683.650 5081.735 2701.670 5082.245 ;
        RECT 2620.585 5079.820 2623.795 5080.400 ;
        RECT 2620.585 5076.485 2626.975 5079.820 ;
        RECT 2620.880 5076.280 2626.975 5076.485 ;
        RECT 2620.880 5075.740 2629.420 5076.280 ;
        RECT 2620.880 5074.660 2629.495 5075.740 ;
        RECT 2620.880 5073.580 2625.530 5074.660 ;
        RECT 2700.240 5072.345 2701.670 5081.735 ;
      LAYER pwell ;
        RECT 3129.785 5082.955 3176.590 5083.260 ;
        RECT 3129.785 5080.935 3139.300 5082.955 ;
      LAYER nwell ;
        RECT 3176.940 5082.245 3210.670 5083.165 ;
        RECT 3192.650 5081.735 3210.670 5082.245 ;
        RECT 3129.585 5079.820 3132.795 5080.400 ;
        RECT 3129.585 5076.485 3135.975 5079.820 ;
        RECT 3129.880 5076.280 3135.975 5076.485 ;
        RECT 3129.880 5075.740 3138.420 5076.280 ;
        RECT 3129.880 5074.660 3138.495 5075.740 ;
        RECT 3129.880 5073.580 3134.530 5074.660 ;
        RECT 3209.240 5072.345 3210.670 5081.735 ;
        RECT 427.940 5071.165 461.670 5072.345 ;
        RECT 684.940 5071.165 718.670 5072.345 ;
        RECT 941.940 5071.165 975.670 5072.345 ;
        RECT 1198.940 5071.165 1232.670 5072.345 ;
        RECT 1456.940 5071.165 1490.670 5072.345 ;
        RECT 1965.940 5071.165 1999.670 5072.345 ;
        RECT 2410.940 5071.165 2444.670 5072.345 ;
        RECT 2667.940 5071.165 2701.670 5072.345 ;
        RECT 3176.940 5071.165 3210.670 5072.345 ;
        RECT 380.285 5067.805 405.815 5069.235 ;
        RECT 380.285 5050.340 381.715 5067.805 ;
        RECT 460.240 5061.775 461.670 5071.165 ;
        RECT 443.650 5061.265 461.670 5061.775 ;
        RECT 427.940 5060.595 461.670 5061.265 ;
        RECT 460.125 5054.045 461.670 5060.595 ;
        RECT 451.335 5053.195 461.670 5054.045 ;
        RECT 380.285 5049.020 384.810 5050.340 ;
        RECT 380.285 5048.770 394.535 5049.020 ;
        RECT 380.285 5048.180 391.460 5048.770 ;
        RECT 380.285 5046.020 381.715 5048.180 ;
        RECT 380.285 5044.590 404.515 5046.020 ;
        RECT 460.125 5040.050 461.670 5053.195 ;
        RECT 637.285 5067.805 662.815 5069.235 ;
        RECT 637.285 5050.340 638.715 5067.805 ;
        RECT 717.240 5061.775 718.670 5071.165 ;
        RECT 700.650 5061.265 718.670 5061.775 ;
        RECT 684.940 5060.595 718.670 5061.265 ;
        RECT 717.125 5054.045 718.670 5060.595 ;
        RECT 708.335 5053.195 718.670 5054.045 ;
        RECT 637.285 5049.020 641.810 5050.340 ;
        RECT 637.285 5048.770 651.535 5049.020 ;
        RECT 637.285 5048.180 648.460 5048.770 ;
        RECT 637.285 5046.020 638.715 5048.180 ;
        RECT 637.285 5044.590 661.515 5046.020 ;
        RECT 717.125 5040.050 718.670 5053.195 ;
        RECT 894.285 5067.805 919.815 5069.235 ;
        RECT 894.285 5050.340 895.715 5067.805 ;
        RECT 974.240 5061.775 975.670 5071.165 ;
        RECT 957.650 5061.265 975.670 5061.775 ;
        RECT 941.940 5060.595 975.670 5061.265 ;
        RECT 974.125 5054.045 975.670 5060.595 ;
        RECT 965.335 5053.195 975.670 5054.045 ;
        RECT 894.285 5049.020 898.810 5050.340 ;
        RECT 894.285 5048.770 908.535 5049.020 ;
        RECT 894.285 5048.180 905.460 5048.770 ;
        RECT 894.285 5046.020 895.715 5048.180 ;
        RECT 894.285 5044.590 918.515 5046.020 ;
        RECT 974.125 5040.050 975.670 5053.195 ;
        RECT 1151.285 5067.805 1176.815 5069.235 ;
        RECT 1151.285 5050.340 1152.715 5067.805 ;
        RECT 1231.240 5061.775 1232.670 5071.165 ;
        RECT 1214.650 5061.265 1232.670 5061.775 ;
        RECT 1198.940 5060.595 1232.670 5061.265 ;
        RECT 1231.125 5054.045 1232.670 5060.595 ;
        RECT 1222.335 5053.195 1232.670 5054.045 ;
        RECT 1151.285 5049.020 1155.810 5050.340 ;
        RECT 1151.285 5048.770 1165.535 5049.020 ;
        RECT 1151.285 5048.180 1162.460 5048.770 ;
        RECT 1151.285 5046.020 1152.715 5048.180 ;
        RECT 1151.285 5044.590 1175.515 5046.020 ;
        RECT 1231.125 5040.050 1232.670 5053.195 ;
        RECT 1409.285 5067.805 1434.815 5069.235 ;
        RECT 1409.285 5050.340 1410.715 5067.805 ;
        RECT 1489.240 5061.775 1490.670 5071.165 ;
        RECT 1472.650 5061.265 1490.670 5061.775 ;
        RECT 1456.940 5060.595 1490.670 5061.265 ;
        RECT 1489.125 5054.045 1490.670 5060.595 ;
        RECT 1480.335 5053.195 1490.670 5054.045 ;
        RECT 1409.285 5049.020 1413.810 5050.340 ;
        RECT 1409.285 5048.770 1423.535 5049.020 ;
        RECT 1409.285 5048.180 1420.460 5048.770 ;
        RECT 1409.285 5046.020 1410.715 5048.180 ;
        RECT 1409.285 5044.590 1433.515 5046.020 ;
        RECT 1489.125 5040.050 1490.670 5053.195 ;
        RECT 1918.285 5067.805 1943.815 5069.235 ;
        RECT 1918.285 5050.340 1919.715 5067.805 ;
        RECT 1998.240 5061.775 1999.670 5071.165 ;
        RECT 1981.650 5061.265 1999.670 5061.775 ;
        RECT 1965.940 5060.595 1999.670 5061.265 ;
        RECT 1998.125 5054.045 1999.670 5060.595 ;
        RECT 1989.335 5053.195 1999.670 5054.045 ;
        RECT 1918.285 5049.020 1922.810 5050.340 ;
        RECT 1918.285 5048.770 1932.535 5049.020 ;
        RECT 1918.285 5048.180 1929.460 5048.770 ;
        RECT 1918.285 5046.020 1919.715 5048.180 ;
        RECT 1918.285 5044.590 1942.515 5046.020 ;
        RECT 1998.125 5040.050 1999.670 5053.195 ;
        RECT 2363.285 5067.805 2388.815 5069.235 ;
        RECT 2363.285 5050.340 2364.715 5067.805 ;
        RECT 2443.240 5061.775 2444.670 5071.165 ;
        RECT 2426.650 5061.265 2444.670 5061.775 ;
        RECT 2410.940 5060.595 2444.670 5061.265 ;
        RECT 2443.125 5054.045 2444.670 5060.595 ;
        RECT 2434.335 5053.195 2444.670 5054.045 ;
        RECT 2363.285 5049.020 2367.810 5050.340 ;
        RECT 2363.285 5048.770 2377.535 5049.020 ;
        RECT 2363.285 5048.180 2374.460 5048.770 ;
        RECT 2363.285 5046.020 2364.715 5048.180 ;
        RECT 2363.285 5044.590 2387.515 5046.020 ;
        RECT 2443.125 5040.050 2444.670 5053.195 ;
        RECT 2620.285 5067.805 2645.815 5069.235 ;
        RECT 2620.285 5050.340 2621.715 5067.805 ;
        RECT 2700.240 5061.775 2701.670 5071.165 ;
        RECT 2683.650 5061.265 2701.670 5061.775 ;
        RECT 2667.940 5060.595 2701.670 5061.265 ;
        RECT 2700.125 5054.045 2701.670 5060.595 ;
        RECT 2691.335 5053.195 2701.670 5054.045 ;
        RECT 2620.285 5049.020 2624.810 5050.340 ;
        RECT 2620.285 5048.770 2634.535 5049.020 ;
        RECT 2620.285 5048.180 2631.460 5048.770 ;
        RECT 2620.285 5046.020 2621.715 5048.180 ;
        RECT 2620.285 5044.590 2644.515 5046.020 ;
        RECT 2700.125 5040.050 2701.670 5053.195 ;
        RECT 3129.285 5067.805 3154.815 5069.235 ;
        RECT 3129.285 5050.340 3130.715 5067.805 ;
        RECT 3209.240 5061.775 3210.670 5071.165 ;
        RECT 3192.650 5061.265 3210.670 5061.775 ;
        RECT 3176.940 5060.595 3210.670 5061.265 ;
        RECT 3209.125 5054.045 3210.670 5060.595 ;
        RECT 3200.335 5053.195 3210.670 5054.045 ;
        RECT 3129.285 5049.020 3133.810 5050.340 ;
        RECT 3129.285 5048.770 3143.535 5049.020 ;
        RECT 3129.285 5048.180 3140.460 5048.770 ;
        RECT 3129.285 5046.020 3130.715 5048.180 ;
        RECT 3129.285 5044.590 3153.515 5046.020 ;
        RECT 3209.125 5040.050 3210.670 5053.195 ;
        RECT 451.335 5038.620 461.670 5040.050 ;
        RECT 708.335 5038.620 718.670 5040.050 ;
        RECT 965.335 5038.620 975.670 5040.050 ;
        RECT 1222.335 5038.620 1232.670 5040.050 ;
        RECT 1480.335 5038.620 1490.670 5040.050 ;
        RECT 1989.335 5038.620 1999.670 5040.050 ;
        RECT 2434.335 5038.620 2444.670 5040.050 ;
        RECT 2691.335 5038.620 2701.670 5040.050 ;
        RECT 3200.335 5038.620 3210.670 5040.050 ;
        RECT 429.915 5022.265 461.450 5024.055 ;
        RECT 686.915 5022.265 718.450 5024.055 ;
        RECT 943.915 5022.265 975.450 5024.055 ;
        RECT 1200.915 5022.265 1232.450 5024.055 ;
        RECT 1458.915 5022.265 1490.450 5024.055 ;
        RECT 1967.915 5022.265 1999.450 5024.055 ;
        RECT 2412.915 5022.265 2444.450 5024.055 ;
        RECT 2669.915 5022.265 2701.450 5024.055 ;
        RECT 3178.915 5022.265 3210.450 5024.055 ;
        RECT 439.275 5020.410 461.450 5022.265 ;
        RECT 696.275 5020.410 718.450 5022.265 ;
        RECT 953.275 5020.410 975.450 5022.265 ;
        RECT 1210.275 5020.410 1232.450 5022.265 ;
        RECT 1468.275 5020.410 1490.450 5022.265 ;
        RECT 1977.275 5020.410 1999.450 5022.265 ;
        RECT 2422.275 5020.410 2444.450 5022.265 ;
        RECT 2679.275 5020.410 2701.450 5022.265 ;
        RECT 3188.275 5020.410 3210.450 5022.265 ;
        RECT 445.830 5017.785 461.450 5020.410 ;
        RECT 702.830 5017.785 718.450 5020.410 ;
        RECT 959.830 5017.785 975.450 5020.410 ;
        RECT 1216.830 5017.785 1232.450 5020.410 ;
        RECT 1474.830 5017.785 1490.450 5020.410 ;
        RECT 1983.830 5017.785 1999.450 5020.410 ;
        RECT 2428.830 5017.785 2444.450 5020.410 ;
        RECT 2685.830 5017.785 2701.450 5020.410 ;
        RECT 3194.830 5017.785 3210.450 5020.410 ;
        RECT 445.830 5011.080 461.450 5013.345 ;
        RECT 702.830 5011.080 718.450 5013.345 ;
        RECT 959.830 5011.080 975.450 5013.345 ;
        RECT 1216.830 5011.080 1232.450 5013.345 ;
        RECT 1474.830 5011.080 1490.450 5013.345 ;
        RECT 1983.830 5011.080 1999.450 5013.345 ;
        RECT 2428.830 5011.080 2444.450 5013.345 ;
        RECT 2685.830 5011.080 2701.450 5013.345 ;
        RECT 3194.830 5011.080 3210.450 5013.345 ;
        RECT 385.580 5007.155 461.450 5011.080 ;
        RECT 642.580 5007.155 718.450 5011.080 ;
        RECT 899.580 5007.155 975.450 5011.080 ;
        RECT 1156.580 5007.155 1232.450 5011.080 ;
        RECT 1414.580 5007.155 1490.450 5011.080 ;
        RECT 1923.580 5007.155 1999.450 5011.080 ;
        RECT 2368.580 5007.155 2444.450 5011.080 ;
        RECT 2625.580 5007.155 2701.450 5011.080 ;
        RECT 3134.580 5007.155 3210.450 5011.080 ;
        RECT 380.585 4993.665 384.110 4997.325 ;
        RECT 637.585 4993.665 641.110 4997.325 ;
        RECT 894.585 4993.665 898.110 4997.325 ;
        RECT 1151.585 4993.665 1155.110 4997.325 ;
        RECT 1409.585 4993.665 1413.110 4997.325 ;
        RECT 1918.585 4993.665 1922.110 4997.325 ;
        RECT 2363.585 4993.665 2367.110 4997.325 ;
        RECT 2620.585 4993.665 2624.110 4997.325 ;
        RECT 3129.585 4993.665 3133.110 4997.325 ;
        RECT 1678.860 4988.685 1737.965 4990.205 ;
        RECT 2889.860 4988.685 2948.965 4990.205 ;
        RECT 29.770 4851.435 55.120 4851.440 ;
        RECT 21.025 4849.630 55.120 4851.435 ;
        RECT 21.025 4837.970 31.485 4849.630 ;
        RECT 21.025 4778.515 26.455 4837.970 ;
        RECT 29.525 4778.515 31.485 4837.970 ;
        RECT 21.025 4777.385 31.485 4778.515 ;
        RECT 53.310 4777.385 55.120 4849.630 ;
        RECT 21.025 4770.585 55.120 4777.385 ;
      LAYER pwell ;
        RECT 55.435 4770.710 59.315 4851.290 ;
      LAYER nwell ;
        RECT 59.615 4817.040 69.335 4851.440 ;
      LAYER pwell ;
        RECT 69.645 4848.865 104.025 4851.290 ;
        RECT 69.645 4837.910 74.865 4848.865 ;
      LAYER nwell ;
        RECT 59.620 4770.585 69.335 4817.040 ;
      LAYER pwell ;
        RECT 70.685 4811.245 74.865 4837.910 ;
        RECT 69.645 4776.735 74.865 4811.245 ;
        RECT 96.450 4847.770 104.025 4848.865 ;
        RECT 96.450 4823.880 100.480 4847.770 ;
        RECT 96.450 4810.385 99.180 4823.880 ;
        RECT 102.015 4816.840 104.025 4847.770 ;
      LAYER nwell ;
        RECT 104.835 4850.240 149.380 4851.670 ;
        RECT 104.835 4833.650 106.265 4850.240 ;
        RECT 104.835 4817.940 105.755 4833.650 ;
        RECT 115.655 4817.940 116.835 4850.240 ;
        RECT 126.225 4850.125 149.380 4850.240 ;
        RECT 126.225 4833.650 127.405 4850.125 ;
        RECT 133.955 4841.335 134.805 4850.125 ;
        RECT 147.950 4841.335 149.380 4850.125 ;
        RECT 126.735 4817.940 127.405 4833.650 ;
        RECT 163.945 4835.830 170.215 4851.450 ;
        RECT 174.655 4835.830 180.845 4851.450 ;
        RECT 163.945 4829.275 167.590 4835.830 ;
        RECT 163.945 4819.915 165.735 4829.275 ;
      LAYER pwell ;
        RECT 104.740 4816.840 105.045 4817.590 ;
        RECT 102.015 4810.385 105.045 4816.840 ;
        RECT 96.450 4776.735 98.035 4810.385 ;
        RECT 69.645 4776.215 98.035 4776.735 ;
        RECT 103.745 4780.300 105.045 4810.385 ;
        RECT 103.745 4776.215 107.065 4780.300 ;
      LAYER nwell ;
        RECT 112.260 4779.420 113.340 4779.495 ;
        RECT 111.720 4776.975 113.340 4779.420 ;
      LAYER pwell ;
        RECT 69.645 4770.785 107.065 4776.215 ;
      LAYER nwell ;
        RECT 108.180 4775.530 113.340 4776.975 ;
        RECT 108.180 4773.795 114.420 4775.530 ;
        RECT 107.600 4770.880 114.420 4773.795 ;
        RECT 118.765 4771.715 120.195 4795.815 ;
        RECT 138.980 4781.460 139.230 4784.535 ;
        RECT 138.980 4774.810 139.820 4781.460 ;
        RECT 137.660 4771.715 139.820 4774.810 ;
        RECT 141.980 4771.715 143.410 4794.515 ;
        RECT 176.920 4775.580 180.845 4835.830 ;
        RECT 3393.665 4834.890 3397.325 4838.415 ;
        RECT 3444.590 4837.285 3469.235 4838.715 ;
        RECT 3476.485 4838.120 3480.400 4838.415 ;
        RECT 107.600 4770.585 111.515 4770.880 ;
        RECT 118.765 4770.285 143.410 4771.715 ;
        RECT 190.675 4770.585 194.335 4774.110 ;
        RECT 3407.155 4773.170 3411.080 4833.420 ;
        RECT 3444.590 4814.485 3446.020 4837.285 ;
        RECT 3448.180 4834.190 3450.340 4837.285 ;
        RECT 3448.180 4827.540 3449.020 4834.190 ;
        RECT 3448.770 4824.465 3449.020 4827.540 ;
        RECT 3467.805 4813.185 3469.235 4837.285 ;
        RECT 3473.580 4835.205 3480.400 4838.120 ;
        RECT 3473.580 4833.470 3479.820 4835.205 ;
        RECT 3474.660 4832.025 3479.820 4833.470 ;
      LAYER pwell ;
        RECT 3480.935 4832.785 3518.355 4838.215 ;
      LAYER nwell ;
        RECT 3474.660 4829.580 3476.280 4832.025 ;
        RECT 3474.660 4829.505 3475.740 4829.580 ;
      LAYER pwell ;
        RECT 3480.935 4828.700 3484.255 4832.785 ;
        RECT 3482.955 4798.615 3484.255 4828.700 ;
        RECT 3489.965 4832.265 3518.355 4832.785 ;
        RECT 3489.965 4798.615 3491.550 4832.265 ;
        RECT 3482.955 4792.160 3485.985 4798.615 ;
        RECT 3482.955 4791.410 3483.260 4792.160 ;
      LAYER nwell ;
        RECT 3422.265 4779.725 3424.055 4789.085 ;
        RECT 3420.410 4773.170 3424.055 4779.725 ;
        RECT 3407.155 4757.550 3413.345 4773.170 ;
        RECT 3417.785 4757.550 3424.055 4773.170 ;
        RECT 3460.595 4775.350 3461.265 4791.060 ;
        RECT 3438.620 4758.875 3440.050 4767.665 ;
        RECT 3453.195 4758.875 3454.045 4767.665 ;
        RECT 3460.595 4758.875 3461.775 4775.350 ;
        RECT 3438.620 4758.760 3461.775 4758.875 ;
        RECT 3471.165 4758.760 3472.345 4791.060 ;
        RECT 3482.245 4775.350 3483.165 4791.060 ;
        RECT 3481.735 4758.760 3483.165 4775.350 ;
        RECT 3438.620 4757.330 3483.165 4758.760 ;
      LAYER pwell ;
        RECT 3483.975 4761.230 3485.985 4792.160 ;
        RECT 3488.820 4785.120 3491.550 4798.615 ;
        RECT 3487.520 4761.230 3491.550 4785.120 ;
        RECT 3483.975 4760.135 3491.550 4761.230 ;
        RECT 3513.135 4797.755 3518.355 4832.265 ;
        RECT 3513.135 4771.090 3517.315 4797.755 ;
      LAYER nwell ;
        RECT 3518.665 4791.960 3528.380 4838.415 ;
      LAYER pwell ;
        RECT 3513.135 4760.135 3518.355 4771.090 ;
        RECT 3483.975 4757.710 3518.355 4760.135 ;
      LAYER nwell ;
        RECT 3518.665 4757.560 3528.385 4791.960 ;
      LAYER pwell ;
        RECT 3528.685 4757.710 3532.565 4838.290 ;
      LAYER nwell ;
        RECT 3532.880 4831.615 3566.975 4838.415 ;
        RECT 3532.880 4759.370 3534.690 4831.615 ;
        RECT 3556.515 4830.485 3566.975 4831.615 ;
        RECT 3556.515 4771.030 3558.475 4830.485 ;
        RECT 3561.545 4771.030 3566.975 4830.485 ;
        RECT 3556.515 4759.370 3566.975 4771.030 ;
        RECT 3532.880 4757.565 3566.975 4759.370 ;
        RECT 3532.880 4757.560 3558.230 4757.565 ;
        RECT 197.795 4360.860 199.315 4419.965 ;
        RECT 3393.665 4388.890 3397.325 4392.415 ;
        RECT 3444.590 4391.285 3469.235 4392.715 ;
        RECT 3476.485 4392.120 3480.400 4392.415 ;
      LAYER pwell ;
        RECT 176.210 4352.495 199.065 4360.285 ;
      LAYER nwell ;
        RECT 3407.155 4327.170 3411.080 4387.420 ;
        RECT 3444.590 4368.485 3446.020 4391.285 ;
        RECT 3448.180 4388.190 3450.340 4391.285 ;
        RECT 3448.180 4381.540 3449.020 4388.190 ;
        RECT 3448.770 4378.465 3449.020 4381.540 ;
        RECT 3467.805 4367.185 3469.235 4391.285 ;
        RECT 3473.580 4389.205 3480.400 4392.120 ;
        RECT 3473.580 4387.470 3479.820 4389.205 ;
        RECT 3474.660 4386.025 3479.820 4387.470 ;
      LAYER pwell ;
        RECT 3480.935 4386.785 3518.355 4392.215 ;
      LAYER nwell ;
        RECT 3474.660 4383.580 3476.280 4386.025 ;
        RECT 3474.660 4383.505 3475.740 4383.580 ;
      LAYER pwell ;
        RECT 3480.935 4382.700 3484.255 4386.785 ;
        RECT 3482.955 4352.615 3484.255 4382.700 ;
        RECT 3489.965 4386.265 3518.355 4386.785 ;
        RECT 3489.965 4352.615 3491.550 4386.265 ;
        RECT 3482.955 4346.160 3485.985 4352.615 ;
        RECT 3482.955 4345.410 3483.260 4346.160 ;
      LAYER nwell ;
        RECT 3422.265 4333.725 3424.055 4343.085 ;
        RECT 3420.410 4327.170 3424.055 4333.725 ;
        RECT 3407.155 4311.550 3413.345 4327.170 ;
        RECT 3417.785 4311.550 3424.055 4327.170 ;
        RECT 3460.595 4329.350 3461.265 4345.060 ;
        RECT 3438.620 4312.875 3440.050 4321.665 ;
        RECT 3453.195 4312.875 3454.045 4321.665 ;
        RECT 3460.595 4312.875 3461.775 4329.350 ;
        RECT 3438.620 4312.760 3461.775 4312.875 ;
        RECT 3471.165 4312.760 3472.345 4345.060 ;
        RECT 3482.245 4329.350 3483.165 4345.060 ;
        RECT 3481.735 4312.760 3483.165 4329.350 ;
        RECT 3438.620 4311.330 3483.165 4312.760 ;
      LAYER pwell ;
        RECT 3483.975 4315.230 3485.985 4346.160 ;
        RECT 3488.820 4339.120 3491.550 4352.615 ;
        RECT 3487.520 4315.230 3491.550 4339.120 ;
        RECT 3483.975 4314.135 3491.550 4315.230 ;
        RECT 3513.135 4351.755 3518.355 4386.265 ;
        RECT 3513.135 4325.090 3517.315 4351.755 ;
      LAYER nwell ;
        RECT 3518.665 4345.960 3528.380 4392.415 ;
      LAYER pwell ;
        RECT 3513.135 4314.135 3518.355 4325.090 ;
        RECT 3483.975 4311.710 3518.355 4314.135 ;
      LAYER nwell ;
        RECT 3518.665 4311.560 3528.385 4345.960 ;
      LAYER pwell ;
        RECT 3528.685 4311.710 3532.565 4392.290 ;
      LAYER nwell ;
        RECT 3532.880 4385.615 3566.975 4392.415 ;
        RECT 3532.880 4313.370 3534.690 4385.615 ;
        RECT 3556.515 4384.485 3566.975 4385.615 ;
        RECT 3556.515 4325.030 3558.475 4384.485 ;
        RECT 3561.545 4325.030 3566.975 4384.485 ;
        RECT 3556.515 4313.370 3566.975 4325.030 ;
        RECT 3532.880 4311.565 3566.975 4313.370 ;
        RECT 3532.880 4311.560 3558.230 4311.565 ;
        RECT 197.795 4149.860 199.315 4208.965 ;
      LAYER pwell ;
        RECT 3388.935 4155.715 3411.790 4163.505 ;
      LAYER nwell ;
        RECT 3388.685 4096.035 3390.205 4155.140 ;
        RECT 29.770 4002.435 55.120 4002.440 ;
        RECT 21.025 4000.630 55.120 4002.435 ;
        RECT 21.025 3988.970 31.485 4000.630 ;
        RECT 21.025 3929.515 26.455 3988.970 ;
        RECT 29.525 3929.515 31.485 3988.970 ;
        RECT 21.025 3928.385 31.485 3929.515 ;
        RECT 53.310 3928.385 55.120 4000.630 ;
        RECT 21.025 3921.585 55.120 3928.385 ;
      LAYER pwell ;
        RECT 55.435 3921.710 59.315 4002.290 ;
      LAYER nwell ;
        RECT 59.615 3968.040 69.335 4002.440 ;
      LAYER pwell ;
        RECT 69.645 3999.865 104.025 4002.290 ;
        RECT 69.645 3988.910 74.865 3999.865 ;
      LAYER nwell ;
        RECT 59.620 3921.585 69.335 3968.040 ;
      LAYER pwell ;
        RECT 70.685 3962.245 74.865 3988.910 ;
        RECT 69.645 3927.735 74.865 3962.245 ;
        RECT 96.450 3998.770 104.025 3999.865 ;
        RECT 96.450 3974.880 100.480 3998.770 ;
        RECT 96.450 3961.385 99.180 3974.880 ;
        RECT 102.015 3967.840 104.025 3998.770 ;
      LAYER nwell ;
        RECT 104.835 4001.240 149.380 4002.670 ;
        RECT 104.835 3984.650 106.265 4001.240 ;
        RECT 104.835 3968.940 105.755 3984.650 ;
        RECT 115.655 3968.940 116.835 4001.240 ;
        RECT 126.225 4001.125 149.380 4001.240 ;
        RECT 126.225 3984.650 127.405 4001.125 ;
        RECT 133.955 3992.335 134.805 4001.125 ;
        RECT 147.950 3992.335 149.380 4001.125 ;
        RECT 126.735 3968.940 127.405 3984.650 ;
        RECT 163.945 3986.830 170.215 4002.450 ;
        RECT 174.655 3986.830 180.845 4002.450 ;
        RECT 163.945 3980.275 167.590 3986.830 ;
        RECT 163.945 3970.915 165.735 3980.275 ;
      LAYER pwell ;
        RECT 104.740 3967.840 105.045 3968.590 ;
        RECT 102.015 3961.385 105.045 3967.840 ;
        RECT 96.450 3927.735 98.035 3961.385 ;
        RECT 69.645 3927.215 98.035 3927.735 ;
        RECT 103.745 3931.300 105.045 3961.385 ;
        RECT 103.745 3927.215 107.065 3931.300 ;
      LAYER nwell ;
        RECT 112.260 3930.420 113.340 3930.495 ;
        RECT 111.720 3927.975 113.340 3930.420 ;
      LAYER pwell ;
        RECT 69.645 3921.785 107.065 3927.215 ;
      LAYER nwell ;
        RECT 108.180 3926.530 113.340 3927.975 ;
        RECT 108.180 3924.795 114.420 3926.530 ;
        RECT 107.600 3921.880 114.420 3924.795 ;
        RECT 118.765 3922.715 120.195 3946.815 ;
        RECT 138.980 3932.460 139.230 3935.535 ;
        RECT 138.980 3925.810 139.820 3932.460 ;
        RECT 137.660 3922.715 139.820 3925.810 ;
        RECT 141.980 3922.715 143.410 3945.515 ;
        RECT 176.920 3926.580 180.845 3986.830 ;
        RECT 3393.665 3942.890 3397.325 3946.415 ;
        RECT 3444.590 3945.285 3469.235 3946.715 ;
        RECT 3476.485 3946.120 3480.400 3946.415 ;
        RECT 107.600 3921.585 111.515 3921.880 ;
        RECT 118.765 3921.285 143.410 3922.715 ;
        RECT 190.675 3921.585 194.335 3925.110 ;
        RECT 3407.155 3881.170 3411.080 3941.420 ;
        RECT 3444.590 3922.485 3446.020 3945.285 ;
        RECT 3448.180 3942.190 3450.340 3945.285 ;
        RECT 3448.180 3935.540 3449.020 3942.190 ;
        RECT 3448.770 3932.465 3449.020 3935.540 ;
        RECT 3467.805 3921.185 3469.235 3945.285 ;
        RECT 3473.580 3943.205 3480.400 3946.120 ;
        RECT 3473.580 3941.470 3479.820 3943.205 ;
        RECT 3474.660 3940.025 3479.820 3941.470 ;
      LAYER pwell ;
        RECT 3480.935 3940.785 3518.355 3946.215 ;
      LAYER nwell ;
        RECT 3474.660 3937.580 3476.280 3940.025 ;
        RECT 3474.660 3937.505 3475.740 3937.580 ;
      LAYER pwell ;
        RECT 3480.935 3936.700 3484.255 3940.785 ;
        RECT 3482.955 3906.615 3484.255 3936.700 ;
        RECT 3489.965 3940.265 3518.355 3940.785 ;
        RECT 3489.965 3906.615 3491.550 3940.265 ;
        RECT 3482.955 3900.160 3485.985 3906.615 ;
        RECT 3482.955 3899.410 3483.260 3900.160 ;
      LAYER nwell ;
        RECT 3422.265 3887.725 3424.055 3897.085 ;
        RECT 3420.410 3881.170 3424.055 3887.725 ;
        RECT 3407.155 3865.550 3413.345 3881.170 ;
        RECT 3417.785 3865.550 3424.055 3881.170 ;
        RECT 3460.595 3883.350 3461.265 3899.060 ;
        RECT 3438.620 3866.875 3440.050 3875.665 ;
        RECT 3453.195 3866.875 3454.045 3875.665 ;
        RECT 3460.595 3866.875 3461.775 3883.350 ;
        RECT 3438.620 3866.760 3461.775 3866.875 ;
        RECT 3471.165 3866.760 3472.345 3899.060 ;
        RECT 3482.245 3883.350 3483.165 3899.060 ;
        RECT 3481.735 3866.760 3483.165 3883.350 ;
        RECT 3438.620 3865.330 3483.165 3866.760 ;
      LAYER pwell ;
        RECT 3483.975 3869.230 3485.985 3900.160 ;
        RECT 3488.820 3893.120 3491.550 3906.615 ;
        RECT 3487.520 3869.230 3491.550 3893.120 ;
        RECT 3483.975 3868.135 3491.550 3869.230 ;
        RECT 3513.135 3905.755 3518.355 3940.265 ;
        RECT 3513.135 3879.090 3517.315 3905.755 ;
      LAYER nwell ;
        RECT 3518.665 3899.960 3528.380 3946.415 ;
      LAYER pwell ;
        RECT 3513.135 3868.135 3518.355 3879.090 ;
        RECT 3483.975 3865.710 3518.355 3868.135 ;
      LAYER nwell ;
        RECT 3518.665 3865.560 3528.385 3899.960 ;
      LAYER pwell ;
        RECT 3528.685 3865.710 3532.565 3946.290 ;
      LAYER nwell ;
        RECT 3532.880 3939.615 3566.975 3946.415 ;
        RECT 3532.880 3867.370 3534.690 3939.615 ;
        RECT 3556.515 3938.485 3566.975 3939.615 ;
        RECT 3556.515 3879.030 3558.475 3938.485 ;
        RECT 3561.545 3879.030 3566.975 3938.485 ;
        RECT 3556.515 3867.370 3566.975 3879.030 ;
        RECT 3532.880 3865.565 3566.975 3867.370 ;
        RECT 3532.880 3865.560 3558.230 3865.565 ;
        RECT 29.770 3786.435 55.120 3786.440 ;
        RECT 21.025 3784.630 55.120 3786.435 ;
        RECT 21.025 3772.970 31.485 3784.630 ;
        RECT 21.025 3713.515 26.455 3772.970 ;
        RECT 29.525 3713.515 31.485 3772.970 ;
        RECT 21.025 3712.385 31.485 3713.515 ;
        RECT 53.310 3712.385 55.120 3784.630 ;
        RECT 21.025 3705.585 55.120 3712.385 ;
      LAYER pwell ;
        RECT 55.435 3705.710 59.315 3786.290 ;
      LAYER nwell ;
        RECT 59.615 3752.040 69.335 3786.440 ;
      LAYER pwell ;
        RECT 69.645 3783.865 104.025 3786.290 ;
        RECT 69.645 3772.910 74.865 3783.865 ;
      LAYER nwell ;
        RECT 59.620 3705.585 69.335 3752.040 ;
      LAYER pwell ;
        RECT 70.685 3746.245 74.865 3772.910 ;
        RECT 69.645 3711.735 74.865 3746.245 ;
        RECT 96.450 3782.770 104.025 3783.865 ;
        RECT 96.450 3758.880 100.480 3782.770 ;
        RECT 96.450 3745.385 99.180 3758.880 ;
        RECT 102.015 3751.840 104.025 3782.770 ;
      LAYER nwell ;
        RECT 104.835 3785.240 149.380 3786.670 ;
        RECT 104.835 3768.650 106.265 3785.240 ;
        RECT 104.835 3752.940 105.755 3768.650 ;
        RECT 115.655 3752.940 116.835 3785.240 ;
        RECT 126.225 3785.125 149.380 3785.240 ;
        RECT 126.225 3768.650 127.405 3785.125 ;
        RECT 133.955 3776.335 134.805 3785.125 ;
        RECT 147.950 3776.335 149.380 3785.125 ;
        RECT 126.735 3752.940 127.405 3768.650 ;
        RECT 163.945 3770.830 170.215 3786.450 ;
        RECT 174.655 3770.830 180.845 3786.450 ;
        RECT 163.945 3764.275 167.590 3770.830 ;
        RECT 163.945 3754.915 165.735 3764.275 ;
      LAYER pwell ;
        RECT 104.740 3751.840 105.045 3752.590 ;
        RECT 102.015 3745.385 105.045 3751.840 ;
        RECT 96.450 3711.735 98.035 3745.385 ;
        RECT 69.645 3711.215 98.035 3711.735 ;
        RECT 103.745 3715.300 105.045 3745.385 ;
        RECT 103.745 3711.215 107.065 3715.300 ;
      LAYER nwell ;
        RECT 112.260 3714.420 113.340 3714.495 ;
        RECT 111.720 3711.975 113.340 3714.420 ;
      LAYER pwell ;
        RECT 69.645 3705.785 107.065 3711.215 ;
      LAYER nwell ;
        RECT 108.180 3710.530 113.340 3711.975 ;
        RECT 108.180 3708.795 114.420 3710.530 ;
        RECT 107.600 3705.880 114.420 3708.795 ;
        RECT 118.765 3706.715 120.195 3730.815 ;
        RECT 138.980 3716.460 139.230 3719.535 ;
        RECT 138.980 3709.810 139.820 3716.460 ;
        RECT 137.660 3706.715 139.820 3709.810 ;
        RECT 141.980 3706.715 143.410 3729.515 ;
        RECT 176.920 3710.580 180.845 3770.830 ;
        RECT 3393.665 3717.890 3397.325 3721.415 ;
        RECT 3444.590 3720.285 3469.235 3721.715 ;
        RECT 3476.485 3721.120 3480.400 3721.415 ;
        RECT 107.600 3705.585 111.515 3705.880 ;
        RECT 118.765 3705.285 143.410 3706.715 ;
        RECT 190.675 3705.585 194.335 3709.110 ;
        RECT 3407.155 3656.170 3411.080 3716.420 ;
        RECT 3444.590 3697.485 3446.020 3720.285 ;
        RECT 3448.180 3717.190 3450.340 3720.285 ;
        RECT 3448.180 3710.540 3449.020 3717.190 ;
        RECT 3448.770 3707.465 3449.020 3710.540 ;
        RECT 3467.805 3696.185 3469.235 3720.285 ;
        RECT 3473.580 3718.205 3480.400 3721.120 ;
        RECT 3473.580 3716.470 3479.820 3718.205 ;
        RECT 3474.660 3715.025 3479.820 3716.470 ;
      LAYER pwell ;
        RECT 3480.935 3715.785 3518.355 3721.215 ;
      LAYER nwell ;
        RECT 3474.660 3712.580 3476.280 3715.025 ;
        RECT 3474.660 3712.505 3475.740 3712.580 ;
      LAYER pwell ;
        RECT 3480.935 3711.700 3484.255 3715.785 ;
        RECT 3482.955 3681.615 3484.255 3711.700 ;
        RECT 3489.965 3715.265 3518.355 3715.785 ;
        RECT 3489.965 3681.615 3491.550 3715.265 ;
        RECT 3482.955 3675.160 3485.985 3681.615 ;
        RECT 3482.955 3674.410 3483.260 3675.160 ;
      LAYER nwell ;
        RECT 3422.265 3662.725 3424.055 3672.085 ;
        RECT 3420.410 3656.170 3424.055 3662.725 ;
        RECT 3407.155 3640.550 3413.345 3656.170 ;
        RECT 3417.785 3640.550 3424.055 3656.170 ;
        RECT 3460.595 3658.350 3461.265 3674.060 ;
        RECT 3438.620 3641.875 3440.050 3650.665 ;
        RECT 3453.195 3641.875 3454.045 3650.665 ;
        RECT 3460.595 3641.875 3461.775 3658.350 ;
        RECT 3438.620 3641.760 3461.775 3641.875 ;
        RECT 3471.165 3641.760 3472.345 3674.060 ;
        RECT 3482.245 3658.350 3483.165 3674.060 ;
        RECT 3481.735 3641.760 3483.165 3658.350 ;
        RECT 3438.620 3640.330 3483.165 3641.760 ;
      LAYER pwell ;
        RECT 3483.975 3644.230 3485.985 3675.160 ;
        RECT 3488.820 3668.120 3491.550 3681.615 ;
        RECT 3487.520 3644.230 3491.550 3668.120 ;
        RECT 3483.975 3643.135 3491.550 3644.230 ;
        RECT 3513.135 3680.755 3518.355 3715.265 ;
        RECT 3513.135 3654.090 3517.315 3680.755 ;
      LAYER nwell ;
        RECT 3518.665 3674.960 3528.380 3721.415 ;
      LAYER pwell ;
        RECT 3513.135 3643.135 3518.355 3654.090 ;
        RECT 3483.975 3640.710 3518.355 3643.135 ;
      LAYER nwell ;
        RECT 3518.665 3640.560 3528.385 3674.960 ;
      LAYER pwell ;
        RECT 3528.685 3640.710 3532.565 3721.290 ;
      LAYER nwell ;
        RECT 3532.880 3714.615 3566.975 3721.415 ;
        RECT 3532.880 3642.370 3534.690 3714.615 ;
        RECT 3556.515 3713.485 3566.975 3714.615 ;
        RECT 3556.515 3654.030 3558.475 3713.485 ;
        RECT 3561.545 3654.030 3566.975 3713.485 ;
        RECT 3556.515 3642.370 3566.975 3654.030 ;
        RECT 3532.880 3640.565 3566.975 3642.370 ;
        RECT 3532.880 3640.560 3558.230 3640.565 ;
        RECT 29.770 3570.435 55.120 3570.440 ;
        RECT 21.025 3568.630 55.120 3570.435 ;
        RECT 21.025 3556.970 31.485 3568.630 ;
        RECT 21.025 3497.515 26.455 3556.970 ;
        RECT 29.525 3497.515 31.485 3556.970 ;
        RECT 21.025 3496.385 31.485 3497.515 ;
        RECT 53.310 3496.385 55.120 3568.630 ;
        RECT 21.025 3489.585 55.120 3496.385 ;
      LAYER pwell ;
        RECT 55.435 3489.710 59.315 3570.290 ;
      LAYER nwell ;
        RECT 59.615 3536.040 69.335 3570.440 ;
      LAYER pwell ;
        RECT 69.645 3567.865 104.025 3570.290 ;
        RECT 69.645 3556.910 74.865 3567.865 ;
      LAYER nwell ;
        RECT 59.620 3489.585 69.335 3536.040 ;
      LAYER pwell ;
        RECT 70.685 3530.245 74.865 3556.910 ;
        RECT 69.645 3495.735 74.865 3530.245 ;
        RECT 96.450 3566.770 104.025 3567.865 ;
        RECT 96.450 3542.880 100.480 3566.770 ;
        RECT 96.450 3529.385 99.180 3542.880 ;
        RECT 102.015 3535.840 104.025 3566.770 ;
      LAYER nwell ;
        RECT 104.835 3569.240 149.380 3570.670 ;
        RECT 104.835 3552.650 106.265 3569.240 ;
        RECT 104.835 3536.940 105.755 3552.650 ;
        RECT 115.655 3536.940 116.835 3569.240 ;
        RECT 126.225 3569.125 149.380 3569.240 ;
        RECT 126.225 3552.650 127.405 3569.125 ;
        RECT 133.955 3560.335 134.805 3569.125 ;
        RECT 147.950 3560.335 149.380 3569.125 ;
        RECT 126.735 3536.940 127.405 3552.650 ;
        RECT 163.945 3554.830 170.215 3570.450 ;
        RECT 174.655 3554.830 180.845 3570.450 ;
        RECT 163.945 3548.275 167.590 3554.830 ;
        RECT 163.945 3538.915 165.735 3548.275 ;
      LAYER pwell ;
        RECT 104.740 3535.840 105.045 3536.590 ;
        RECT 102.015 3529.385 105.045 3535.840 ;
        RECT 96.450 3495.735 98.035 3529.385 ;
        RECT 69.645 3495.215 98.035 3495.735 ;
        RECT 103.745 3499.300 105.045 3529.385 ;
        RECT 103.745 3495.215 107.065 3499.300 ;
      LAYER nwell ;
        RECT 112.260 3498.420 113.340 3498.495 ;
        RECT 111.720 3495.975 113.340 3498.420 ;
      LAYER pwell ;
        RECT 69.645 3489.785 107.065 3495.215 ;
      LAYER nwell ;
        RECT 108.180 3494.530 113.340 3495.975 ;
        RECT 108.180 3492.795 114.420 3494.530 ;
        RECT 107.600 3489.880 114.420 3492.795 ;
        RECT 118.765 3490.715 120.195 3514.815 ;
        RECT 138.980 3500.460 139.230 3503.535 ;
        RECT 138.980 3493.810 139.820 3500.460 ;
        RECT 137.660 3490.715 139.820 3493.810 ;
        RECT 141.980 3490.715 143.410 3513.515 ;
        RECT 176.920 3494.580 180.845 3554.830 ;
        RECT 107.600 3489.585 111.515 3489.880 ;
        RECT 118.765 3489.285 143.410 3490.715 ;
        RECT 190.675 3489.585 194.335 3493.110 ;
        RECT 3393.665 3492.890 3397.325 3496.415 ;
        RECT 3444.590 3495.285 3469.235 3496.715 ;
        RECT 3476.485 3496.120 3480.400 3496.415 ;
        RECT 3407.155 3431.170 3411.080 3491.420 ;
        RECT 3444.590 3472.485 3446.020 3495.285 ;
        RECT 3448.180 3492.190 3450.340 3495.285 ;
        RECT 3448.180 3485.540 3449.020 3492.190 ;
        RECT 3448.770 3482.465 3449.020 3485.540 ;
        RECT 3467.805 3471.185 3469.235 3495.285 ;
        RECT 3473.580 3493.205 3480.400 3496.120 ;
        RECT 3473.580 3491.470 3479.820 3493.205 ;
        RECT 3474.660 3490.025 3479.820 3491.470 ;
      LAYER pwell ;
        RECT 3480.935 3490.785 3518.355 3496.215 ;
      LAYER nwell ;
        RECT 3474.660 3487.580 3476.280 3490.025 ;
        RECT 3474.660 3487.505 3475.740 3487.580 ;
      LAYER pwell ;
        RECT 3480.935 3486.700 3484.255 3490.785 ;
        RECT 3482.955 3456.615 3484.255 3486.700 ;
        RECT 3489.965 3490.265 3518.355 3490.785 ;
        RECT 3489.965 3456.615 3491.550 3490.265 ;
        RECT 3482.955 3450.160 3485.985 3456.615 ;
        RECT 3482.955 3449.410 3483.260 3450.160 ;
      LAYER nwell ;
        RECT 3422.265 3437.725 3424.055 3447.085 ;
        RECT 3420.410 3431.170 3424.055 3437.725 ;
        RECT 3407.155 3415.550 3413.345 3431.170 ;
        RECT 3417.785 3415.550 3424.055 3431.170 ;
        RECT 3460.595 3433.350 3461.265 3449.060 ;
        RECT 3438.620 3416.875 3440.050 3425.665 ;
        RECT 3453.195 3416.875 3454.045 3425.665 ;
        RECT 3460.595 3416.875 3461.775 3433.350 ;
        RECT 3438.620 3416.760 3461.775 3416.875 ;
        RECT 3471.165 3416.760 3472.345 3449.060 ;
        RECT 3482.245 3433.350 3483.165 3449.060 ;
        RECT 3481.735 3416.760 3483.165 3433.350 ;
        RECT 3438.620 3415.330 3483.165 3416.760 ;
      LAYER pwell ;
        RECT 3483.975 3419.230 3485.985 3450.160 ;
        RECT 3488.820 3443.120 3491.550 3456.615 ;
        RECT 3487.520 3419.230 3491.550 3443.120 ;
        RECT 3483.975 3418.135 3491.550 3419.230 ;
        RECT 3513.135 3455.755 3518.355 3490.265 ;
        RECT 3513.135 3429.090 3517.315 3455.755 ;
      LAYER nwell ;
        RECT 3518.665 3449.960 3528.380 3496.415 ;
      LAYER pwell ;
        RECT 3513.135 3418.135 3518.355 3429.090 ;
        RECT 3483.975 3415.710 3518.355 3418.135 ;
      LAYER nwell ;
        RECT 3518.665 3415.560 3528.385 3449.960 ;
      LAYER pwell ;
        RECT 3528.685 3415.710 3532.565 3496.290 ;
      LAYER nwell ;
        RECT 3532.880 3489.615 3566.975 3496.415 ;
        RECT 3532.880 3417.370 3534.690 3489.615 ;
        RECT 3556.515 3488.485 3566.975 3489.615 ;
        RECT 3556.515 3429.030 3558.475 3488.485 ;
        RECT 3561.545 3429.030 3566.975 3488.485 ;
        RECT 3556.515 3417.370 3566.975 3429.030 ;
        RECT 3532.880 3415.565 3566.975 3417.370 ;
        RECT 3532.880 3415.560 3558.230 3415.565 ;
        RECT 29.770 3354.435 55.120 3354.440 ;
        RECT 21.025 3352.630 55.120 3354.435 ;
        RECT 21.025 3340.970 31.485 3352.630 ;
        RECT 21.025 3281.515 26.455 3340.970 ;
        RECT 29.525 3281.515 31.485 3340.970 ;
        RECT 21.025 3280.385 31.485 3281.515 ;
        RECT 53.310 3280.385 55.120 3352.630 ;
        RECT 21.025 3273.585 55.120 3280.385 ;
      LAYER pwell ;
        RECT 55.435 3273.710 59.315 3354.290 ;
      LAYER nwell ;
        RECT 59.615 3320.040 69.335 3354.440 ;
      LAYER pwell ;
        RECT 69.645 3351.865 104.025 3354.290 ;
        RECT 69.645 3340.910 74.865 3351.865 ;
      LAYER nwell ;
        RECT 59.620 3273.585 69.335 3320.040 ;
      LAYER pwell ;
        RECT 70.685 3314.245 74.865 3340.910 ;
        RECT 69.645 3279.735 74.865 3314.245 ;
        RECT 96.450 3350.770 104.025 3351.865 ;
        RECT 96.450 3326.880 100.480 3350.770 ;
        RECT 96.450 3313.385 99.180 3326.880 ;
        RECT 102.015 3319.840 104.025 3350.770 ;
      LAYER nwell ;
        RECT 104.835 3353.240 149.380 3354.670 ;
        RECT 104.835 3336.650 106.265 3353.240 ;
        RECT 104.835 3320.940 105.755 3336.650 ;
        RECT 115.655 3320.940 116.835 3353.240 ;
        RECT 126.225 3353.125 149.380 3353.240 ;
        RECT 126.225 3336.650 127.405 3353.125 ;
        RECT 133.955 3344.335 134.805 3353.125 ;
        RECT 147.950 3344.335 149.380 3353.125 ;
        RECT 126.735 3320.940 127.405 3336.650 ;
        RECT 163.945 3338.830 170.215 3354.450 ;
        RECT 174.655 3338.830 180.845 3354.450 ;
        RECT 163.945 3332.275 167.590 3338.830 ;
        RECT 163.945 3322.915 165.735 3332.275 ;
      LAYER pwell ;
        RECT 104.740 3319.840 105.045 3320.590 ;
        RECT 102.015 3313.385 105.045 3319.840 ;
        RECT 96.450 3279.735 98.035 3313.385 ;
        RECT 69.645 3279.215 98.035 3279.735 ;
        RECT 103.745 3283.300 105.045 3313.385 ;
        RECT 103.745 3279.215 107.065 3283.300 ;
      LAYER nwell ;
        RECT 112.260 3282.420 113.340 3282.495 ;
        RECT 111.720 3279.975 113.340 3282.420 ;
      LAYER pwell ;
        RECT 69.645 3273.785 107.065 3279.215 ;
      LAYER nwell ;
        RECT 108.180 3278.530 113.340 3279.975 ;
        RECT 108.180 3276.795 114.420 3278.530 ;
        RECT 107.600 3273.880 114.420 3276.795 ;
        RECT 118.765 3274.715 120.195 3298.815 ;
        RECT 138.980 3284.460 139.230 3287.535 ;
        RECT 138.980 3277.810 139.820 3284.460 ;
        RECT 137.660 3274.715 139.820 3277.810 ;
        RECT 141.980 3274.715 143.410 3297.515 ;
        RECT 176.920 3278.580 180.845 3338.830 ;
        RECT 107.600 3273.585 111.515 3273.880 ;
        RECT 118.765 3273.285 143.410 3274.715 ;
        RECT 190.675 3273.585 194.335 3277.110 ;
        RECT 3393.665 3266.890 3397.325 3270.415 ;
        RECT 3444.590 3269.285 3469.235 3270.715 ;
        RECT 3476.485 3270.120 3480.400 3270.415 ;
        RECT 3407.155 3205.170 3411.080 3265.420 ;
        RECT 3444.590 3246.485 3446.020 3269.285 ;
        RECT 3448.180 3266.190 3450.340 3269.285 ;
        RECT 3448.180 3259.540 3449.020 3266.190 ;
        RECT 3448.770 3256.465 3449.020 3259.540 ;
        RECT 3467.805 3245.185 3469.235 3269.285 ;
        RECT 3473.580 3267.205 3480.400 3270.120 ;
        RECT 3473.580 3265.470 3479.820 3267.205 ;
        RECT 3474.660 3264.025 3479.820 3265.470 ;
      LAYER pwell ;
        RECT 3480.935 3264.785 3518.355 3270.215 ;
      LAYER nwell ;
        RECT 3474.660 3261.580 3476.280 3264.025 ;
        RECT 3474.660 3261.505 3475.740 3261.580 ;
      LAYER pwell ;
        RECT 3480.935 3260.700 3484.255 3264.785 ;
        RECT 3482.955 3230.615 3484.255 3260.700 ;
        RECT 3489.965 3264.265 3518.355 3264.785 ;
        RECT 3489.965 3230.615 3491.550 3264.265 ;
        RECT 3482.955 3224.160 3485.985 3230.615 ;
        RECT 3482.955 3223.410 3483.260 3224.160 ;
      LAYER nwell ;
        RECT 3422.265 3211.725 3424.055 3221.085 ;
        RECT 3420.410 3205.170 3424.055 3211.725 ;
        RECT 3407.155 3189.550 3413.345 3205.170 ;
        RECT 3417.785 3189.550 3424.055 3205.170 ;
        RECT 3460.595 3207.350 3461.265 3223.060 ;
        RECT 3438.620 3190.875 3440.050 3199.665 ;
        RECT 3453.195 3190.875 3454.045 3199.665 ;
        RECT 3460.595 3190.875 3461.775 3207.350 ;
        RECT 3438.620 3190.760 3461.775 3190.875 ;
        RECT 3471.165 3190.760 3472.345 3223.060 ;
        RECT 3482.245 3207.350 3483.165 3223.060 ;
        RECT 3481.735 3190.760 3483.165 3207.350 ;
        RECT 3438.620 3189.330 3483.165 3190.760 ;
      LAYER pwell ;
        RECT 3483.975 3193.230 3485.985 3224.160 ;
        RECT 3488.820 3217.120 3491.550 3230.615 ;
        RECT 3487.520 3193.230 3491.550 3217.120 ;
        RECT 3483.975 3192.135 3491.550 3193.230 ;
        RECT 3513.135 3229.755 3518.355 3264.265 ;
        RECT 3513.135 3203.090 3517.315 3229.755 ;
      LAYER nwell ;
        RECT 3518.665 3223.960 3528.380 3270.415 ;
      LAYER pwell ;
        RECT 3513.135 3192.135 3518.355 3203.090 ;
        RECT 3483.975 3189.710 3518.355 3192.135 ;
      LAYER nwell ;
        RECT 3518.665 3189.560 3528.385 3223.960 ;
      LAYER pwell ;
        RECT 3528.685 3189.710 3532.565 3270.290 ;
      LAYER nwell ;
        RECT 3532.880 3263.615 3566.975 3270.415 ;
        RECT 3532.880 3191.370 3534.690 3263.615 ;
        RECT 3556.515 3262.485 3566.975 3263.615 ;
        RECT 3556.515 3203.030 3558.475 3262.485 ;
        RECT 3561.545 3203.030 3566.975 3262.485 ;
        RECT 3556.515 3191.370 3566.975 3203.030 ;
        RECT 3532.880 3189.565 3566.975 3191.370 ;
        RECT 3532.880 3189.560 3558.230 3189.565 ;
        RECT 29.770 3138.435 55.120 3138.440 ;
        RECT 21.025 3136.630 55.120 3138.435 ;
        RECT 21.025 3124.970 31.485 3136.630 ;
        RECT 21.025 3065.515 26.455 3124.970 ;
        RECT 29.525 3065.515 31.485 3124.970 ;
        RECT 21.025 3064.385 31.485 3065.515 ;
        RECT 53.310 3064.385 55.120 3136.630 ;
        RECT 21.025 3057.585 55.120 3064.385 ;
      LAYER pwell ;
        RECT 55.435 3057.710 59.315 3138.290 ;
      LAYER nwell ;
        RECT 59.615 3104.040 69.335 3138.440 ;
      LAYER pwell ;
        RECT 69.645 3135.865 104.025 3138.290 ;
        RECT 69.645 3124.910 74.865 3135.865 ;
      LAYER nwell ;
        RECT 59.620 3057.585 69.335 3104.040 ;
      LAYER pwell ;
        RECT 70.685 3098.245 74.865 3124.910 ;
        RECT 69.645 3063.735 74.865 3098.245 ;
        RECT 96.450 3134.770 104.025 3135.865 ;
        RECT 96.450 3110.880 100.480 3134.770 ;
        RECT 96.450 3097.385 99.180 3110.880 ;
        RECT 102.015 3103.840 104.025 3134.770 ;
      LAYER nwell ;
        RECT 104.835 3137.240 149.380 3138.670 ;
        RECT 104.835 3120.650 106.265 3137.240 ;
        RECT 104.835 3104.940 105.755 3120.650 ;
        RECT 115.655 3104.940 116.835 3137.240 ;
        RECT 126.225 3137.125 149.380 3137.240 ;
        RECT 126.225 3120.650 127.405 3137.125 ;
        RECT 133.955 3128.335 134.805 3137.125 ;
        RECT 147.950 3128.335 149.380 3137.125 ;
        RECT 126.735 3104.940 127.405 3120.650 ;
        RECT 163.945 3122.830 170.215 3138.450 ;
        RECT 174.655 3122.830 180.845 3138.450 ;
        RECT 163.945 3116.275 167.590 3122.830 ;
        RECT 163.945 3106.915 165.735 3116.275 ;
      LAYER pwell ;
        RECT 104.740 3103.840 105.045 3104.590 ;
        RECT 102.015 3097.385 105.045 3103.840 ;
        RECT 96.450 3063.735 98.035 3097.385 ;
        RECT 69.645 3063.215 98.035 3063.735 ;
        RECT 103.745 3067.300 105.045 3097.385 ;
        RECT 103.745 3063.215 107.065 3067.300 ;
      LAYER nwell ;
        RECT 112.260 3066.420 113.340 3066.495 ;
        RECT 111.720 3063.975 113.340 3066.420 ;
      LAYER pwell ;
        RECT 69.645 3057.785 107.065 3063.215 ;
      LAYER nwell ;
        RECT 108.180 3062.530 113.340 3063.975 ;
        RECT 108.180 3060.795 114.420 3062.530 ;
        RECT 107.600 3057.880 114.420 3060.795 ;
        RECT 118.765 3058.715 120.195 3082.815 ;
        RECT 138.980 3068.460 139.230 3071.535 ;
        RECT 138.980 3061.810 139.820 3068.460 ;
        RECT 137.660 3058.715 139.820 3061.810 ;
        RECT 141.980 3058.715 143.410 3081.515 ;
        RECT 176.920 3062.580 180.845 3122.830 ;
        RECT 107.600 3057.585 111.515 3057.880 ;
        RECT 118.765 3057.285 143.410 3058.715 ;
        RECT 190.675 3057.585 194.335 3061.110 ;
        RECT 3393.665 3041.890 3397.325 3045.415 ;
        RECT 3444.590 3044.285 3469.235 3045.715 ;
        RECT 3476.485 3045.120 3480.400 3045.415 ;
        RECT 3407.155 2980.170 3411.080 3040.420 ;
        RECT 3444.590 3021.485 3446.020 3044.285 ;
        RECT 3448.180 3041.190 3450.340 3044.285 ;
        RECT 3448.180 3034.540 3449.020 3041.190 ;
        RECT 3448.770 3031.465 3449.020 3034.540 ;
        RECT 3467.805 3020.185 3469.235 3044.285 ;
        RECT 3473.580 3042.205 3480.400 3045.120 ;
        RECT 3473.580 3040.470 3479.820 3042.205 ;
        RECT 3474.660 3039.025 3479.820 3040.470 ;
      LAYER pwell ;
        RECT 3480.935 3039.785 3518.355 3045.215 ;
      LAYER nwell ;
        RECT 3474.660 3036.580 3476.280 3039.025 ;
        RECT 3474.660 3036.505 3475.740 3036.580 ;
      LAYER pwell ;
        RECT 3480.935 3035.700 3484.255 3039.785 ;
        RECT 3482.955 3005.615 3484.255 3035.700 ;
        RECT 3489.965 3039.265 3518.355 3039.785 ;
        RECT 3489.965 3005.615 3491.550 3039.265 ;
        RECT 3482.955 2999.160 3485.985 3005.615 ;
        RECT 3482.955 2998.410 3483.260 2999.160 ;
      LAYER nwell ;
        RECT 3422.265 2986.725 3424.055 2996.085 ;
        RECT 3420.410 2980.170 3424.055 2986.725 ;
        RECT 3407.155 2964.550 3413.345 2980.170 ;
        RECT 3417.785 2964.550 3424.055 2980.170 ;
        RECT 3460.595 2982.350 3461.265 2998.060 ;
        RECT 3438.620 2965.875 3440.050 2974.665 ;
        RECT 3453.195 2965.875 3454.045 2974.665 ;
        RECT 3460.595 2965.875 3461.775 2982.350 ;
        RECT 3438.620 2965.760 3461.775 2965.875 ;
        RECT 3471.165 2965.760 3472.345 2998.060 ;
        RECT 3482.245 2982.350 3483.165 2998.060 ;
        RECT 3481.735 2965.760 3483.165 2982.350 ;
        RECT 3438.620 2964.330 3483.165 2965.760 ;
      LAYER pwell ;
        RECT 3483.975 2968.230 3485.985 2999.160 ;
        RECT 3488.820 2992.120 3491.550 3005.615 ;
        RECT 3487.520 2968.230 3491.550 2992.120 ;
        RECT 3483.975 2967.135 3491.550 2968.230 ;
        RECT 3513.135 3004.755 3518.355 3039.265 ;
        RECT 3513.135 2978.090 3517.315 3004.755 ;
      LAYER nwell ;
        RECT 3518.665 2998.960 3528.380 3045.415 ;
      LAYER pwell ;
        RECT 3513.135 2967.135 3518.355 2978.090 ;
        RECT 3483.975 2964.710 3518.355 2967.135 ;
      LAYER nwell ;
        RECT 3518.665 2964.560 3528.385 2998.960 ;
      LAYER pwell ;
        RECT 3528.685 2964.710 3532.565 3045.290 ;
      LAYER nwell ;
        RECT 3532.880 3038.615 3566.975 3045.415 ;
        RECT 3532.880 2966.370 3534.690 3038.615 ;
        RECT 3556.515 3037.485 3566.975 3038.615 ;
        RECT 3556.515 2978.030 3558.475 3037.485 ;
        RECT 3561.545 2978.030 3566.975 3037.485 ;
        RECT 3556.515 2966.370 3566.975 2978.030 ;
        RECT 3532.880 2964.565 3566.975 2966.370 ;
        RECT 3532.880 2964.560 3558.230 2964.565 ;
        RECT 29.770 2922.435 55.120 2922.440 ;
        RECT 21.025 2920.630 55.120 2922.435 ;
        RECT 21.025 2908.970 31.485 2920.630 ;
        RECT 21.025 2849.515 26.455 2908.970 ;
        RECT 29.525 2849.515 31.485 2908.970 ;
        RECT 21.025 2848.385 31.485 2849.515 ;
        RECT 53.310 2848.385 55.120 2920.630 ;
        RECT 21.025 2841.585 55.120 2848.385 ;
      LAYER pwell ;
        RECT 55.435 2841.710 59.315 2922.290 ;
      LAYER nwell ;
        RECT 59.615 2888.040 69.335 2922.440 ;
      LAYER pwell ;
        RECT 69.645 2919.865 104.025 2922.290 ;
        RECT 69.645 2908.910 74.865 2919.865 ;
      LAYER nwell ;
        RECT 59.620 2841.585 69.335 2888.040 ;
      LAYER pwell ;
        RECT 70.685 2882.245 74.865 2908.910 ;
        RECT 69.645 2847.735 74.865 2882.245 ;
        RECT 96.450 2918.770 104.025 2919.865 ;
        RECT 96.450 2894.880 100.480 2918.770 ;
        RECT 96.450 2881.385 99.180 2894.880 ;
        RECT 102.015 2887.840 104.025 2918.770 ;
      LAYER nwell ;
        RECT 104.835 2921.240 149.380 2922.670 ;
        RECT 104.835 2904.650 106.265 2921.240 ;
        RECT 104.835 2888.940 105.755 2904.650 ;
        RECT 115.655 2888.940 116.835 2921.240 ;
        RECT 126.225 2921.125 149.380 2921.240 ;
        RECT 126.225 2904.650 127.405 2921.125 ;
        RECT 133.955 2912.335 134.805 2921.125 ;
        RECT 147.950 2912.335 149.380 2921.125 ;
        RECT 126.735 2888.940 127.405 2904.650 ;
        RECT 163.945 2906.830 170.215 2922.450 ;
        RECT 174.655 2906.830 180.845 2922.450 ;
        RECT 163.945 2900.275 167.590 2906.830 ;
        RECT 163.945 2890.915 165.735 2900.275 ;
      LAYER pwell ;
        RECT 104.740 2887.840 105.045 2888.590 ;
        RECT 102.015 2881.385 105.045 2887.840 ;
        RECT 96.450 2847.735 98.035 2881.385 ;
        RECT 69.645 2847.215 98.035 2847.735 ;
        RECT 103.745 2851.300 105.045 2881.385 ;
        RECT 103.745 2847.215 107.065 2851.300 ;
      LAYER nwell ;
        RECT 112.260 2850.420 113.340 2850.495 ;
        RECT 111.720 2847.975 113.340 2850.420 ;
      LAYER pwell ;
        RECT 69.645 2841.785 107.065 2847.215 ;
      LAYER nwell ;
        RECT 108.180 2846.530 113.340 2847.975 ;
        RECT 108.180 2844.795 114.420 2846.530 ;
        RECT 107.600 2841.880 114.420 2844.795 ;
        RECT 118.765 2842.715 120.195 2866.815 ;
        RECT 138.980 2852.460 139.230 2855.535 ;
        RECT 138.980 2845.810 139.820 2852.460 ;
        RECT 137.660 2842.715 139.820 2845.810 ;
        RECT 141.980 2842.715 143.410 2865.515 ;
        RECT 176.920 2846.580 180.845 2906.830 ;
        RECT 107.600 2841.585 111.515 2841.880 ;
        RECT 118.765 2841.285 143.410 2842.715 ;
        RECT 190.675 2841.585 194.335 2845.110 ;
        RECT 3393.665 2815.890 3397.325 2819.415 ;
        RECT 3444.590 2818.285 3469.235 2819.715 ;
        RECT 3476.485 2819.120 3480.400 2819.415 ;
        RECT 3407.155 2754.170 3411.080 2814.420 ;
        RECT 3444.590 2795.485 3446.020 2818.285 ;
        RECT 3448.180 2815.190 3450.340 2818.285 ;
        RECT 3448.180 2808.540 3449.020 2815.190 ;
        RECT 3448.770 2805.465 3449.020 2808.540 ;
        RECT 3467.805 2794.185 3469.235 2818.285 ;
        RECT 3473.580 2816.205 3480.400 2819.120 ;
        RECT 3473.580 2814.470 3479.820 2816.205 ;
        RECT 3474.660 2813.025 3479.820 2814.470 ;
      LAYER pwell ;
        RECT 3480.935 2813.785 3518.355 2819.215 ;
      LAYER nwell ;
        RECT 3474.660 2810.580 3476.280 2813.025 ;
        RECT 3474.660 2810.505 3475.740 2810.580 ;
      LAYER pwell ;
        RECT 3480.935 2809.700 3484.255 2813.785 ;
        RECT 3482.955 2779.615 3484.255 2809.700 ;
        RECT 3489.965 2813.265 3518.355 2813.785 ;
        RECT 3489.965 2779.615 3491.550 2813.265 ;
        RECT 3482.955 2773.160 3485.985 2779.615 ;
        RECT 3482.955 2772.410 3483.260 2773.160 ;
      LAYER nwell ;
        RECT 3422.265 2760.725 3424.055 2770.085 ;
        RECT 3420.410 2754.170 3424.055 2760.725 ;
        RECT 3407.155 2738.550 3413.345 2754.170 ;
        RECT 3417.785 2738.550 3424.055 2754.170 ;
        RECT 3460.595 2756.350 3461.265 2772.060 ;
        RECT 3438.620 2739.875 3440.050 2748.665 ;
        RECT 3453.195 2739.875 3454.045 2748.665 ;
        RECT 3460.595 2739.875 3461.775 2756.350 ;
        RECT 3438.620 2739.760 3461.775 2739.875 ;
        RECT 3471.165 2739.760 3472.345 2772.060 ;
        RECT 3482.245 2756.350 3483.165 2772.060 ;
        RECT 3481.735 2739.760 3483.165 2756.350 ;
        RECT 3438.620 2738.330 3483.165 2739.760 ;
      LAYER pwell ;
        RECT 3483.975 2742.230 3485.985 2773.160 ;
        RECT 3488.820 2766.120 3491.550 2779.615 ;
        RECT 3487.520 2742.230 3491.550 2766.120 ;
        RECT 3483.975 2741.135 3491.550 2742.230 ;
        RECT 3513.135 2778.755 3518.355 2813.265 ;
        RECT 3513.135 2752.090 3517.315 2778.755 ;
      LAYER nwell ;
        RECT 3518.665 2772.960 3528.380 2819.415 ;
      LAYER pwell ;
        RECT 3513.135 2741.135 3518.355 2752.090 ;
        RECT 3483.975 2738.710 3518.355 2741.135 ;
      LAYER nwell ;
        RECT 3518.665 2738.560 3528.385 2772.960 ;
      LAYER pwell ;
        RECT 3528.685 2738.710 3532.565 2819.290 ;
      LAYER nwell ;
        RECT 3532.880 2812.615 3566.975 2819.415 ;
        RECT 3532.880 2740.370 3534.690 2812.615 ;
        RECT 3556.515 2811.485 3566.975 2812.615 ;
        RECT 3556.515 2752.030 3558.475 2811.485 ;
        RECT 3561.545 2752.030 3566.975 2811.485 ;
        RECT 3556.515 2740.370 3566.975 2752.030 ;
        RECT 3532.880 2738.565 3566.975 2740.370 ;
        RECT 3532.880 2738.560 3558.230 2738.565 ;
        RECT 29.770 2706.435 55.120 2706.440 ;
        RECT 21.025 2704.630 55.120 2706.435 ;
        RECT 21.025 2692.970 31.485 2704.630 ;
        RECT 21.025 2633.515 26.455 2692.970 ;
        RECT 29.525 2633.515 31.485 2692.970 ;
        RECT 21.025 2632.385 31.485 2633.515 ;
        RECT 53.310 2632.385 55.120 2704.630 ;
        RECT 21.025 2625.585 55.120 2632.385 ;
      LAYER pwell ;
        RECT 55.435 2625.710 59.315 2706.290 ;
      LAYER nwell ;
        RECT 59.615 2672.040 69.335 2706.440 ;
      LAYER pwell ;
        RECT 69.645 2703.865 104.025 2706.290 ;
        RECT 69.645 2692.910 74.865 2703.865 ;
      LAYER nwell ;
        RECT 59.620 2625.585 69.335 2672.040 ;
      LAYER pwell ;
        RECT 70.685 2666.245 74.865 2692.910 ;
        RECT 69.645 2631.735 74.865 2666.245 ;
        RECT 96.450 2702.770 104.025 2703.865 ;
        RECT 96.450 2678.880 100.480 2702.770 ;
        RECT 96.450 2665.385 99.180 2678.880 ;
        RECT 102.015 2671.840 104.025 2702.770 ;
      LAYER nwell ;
        RECT 104.835 2705.240 149.380 2706.670 ;
        RECT 104.835 2688.650 106.265 2705.240 ;
        RECT 104.835 2672.940 105.755 2688.650 ;
        RECT 115.655 2672.940 116.835 2705.240 ;
        RECT 126.225 2705.125 149.380 2705.240 ;
        RECT 126.225 2688.650 127.405 2705.125 ;
        RECT 133.955 2696.335 134.805 2705.125 ;
        RECT 147.950 2696.335 149.380 2705.125 ;
        RECT 126.735 2672.940 127.405 2688.650 ;
        RECT 163.945 2690.830 170.215 2706.450 ;
        RECT 174.655 2690.830 180.845 2706.450 ;
        RECT 163.945 2684.275 167.590 2690.830 ;
        RECT 163.945 2674.915 165.735 2684.275 ;
      LAYER pwell ;
        RECT 104.740 2671.840 105.045 2672.590 ;
        RECT 102.015 2665.385 105.045 2671.840 ;
        RECT 96.450 2631.735 98.035 2665.385 ;
        RECT 69.645 2631.215 98.035 2631.735 ;
        RECT 103.745 2635.300 105.045 2665.385 ;
        RECT 103.745 2631.215 107.065 2635.300 ;
      LAYER nwell ;
        RECT 112.260 2634.420 113.340 2634.495 ;
        RECT 111.720 2631.975 113.340 2634.420 ;
      LAYER pwell ;
        RECT 69.645 2625.785 107.065 2631.215 ;
      LAYER nwell ;
        RECT 108.180 2630.530 113.340 2631.975 ;
        RECT 108.180 2628.795 114.420 2630.530 ;
        RECT 107.600 2625.880 114.420 2628.795 ;
        RECT 118.765 2626.715 120.195 2650.815 ;
        RECT 138.980 2636.460 139.230 2639.535 ;
        RECT 138.980 2629.810 139.820 2636.460 ;
        RECT 137.660 2626.715 139.820 2629.810 ;
        RECT 141.980 2626.715 143.410 2649.515 ;
        RECT 176.920 2630.580 180.845 2690.830 ;
        RECT 107.600 2625.585 111.515 2625.880 ;
        RECT 118.765 2625.285 143.410 2626.715 ;
        RECT 190.675 2625.585 194.335 2629.110 ;
      LAYER pwell ;
        RECT 3388.935 2582.715 3411.790 2590.505 ;
      LAYER nwell ;
        RECT 3388.685 2523.035 3390.205 2582.140 ;
        RECT 197.795 2426.860 199.315 2485.965 ;
      LAYER pwell ;
        RECT 176.210 2418.495 199.065 2426.285 ;
      LAYER nwell ;
        RECT 3388.685 2082.035 3390.205 2141.140 ;
        RECT 29.770 2068.435 55.120 2068.440 ;
        RECT 21.025 2066.630 55.120 2068.435 ;
        RECT 21.025 2054.970 31.485 2066.630 ;
        RECT 21.025 1995.515 26.455 2054.970 ;
        RECT 29.525 1995.515 31.485 2054.970 ;
        RECT 21.025 1994.385 31.485 1995.515 ;
        RECT 53.310 1994.385 55.120 2066.630 ;
        RECT 21.025 1987.585 55.120 1994.385 ;
      LAYER pwell ;
        RECT 55.435 1987.710 59.315 2068.290 ;
      LAYER nwell ;
        RECT 59.615 2034.040 69.335 2068.440 ;
      LAYER pwell ;
        RECT 69.645 2065.865 104.025 2068.290 ;
        RECT 69.645 2054.910 74.865 2065.865 ;
      LAYER nwell ;
        RECT 59.620 1987.585 69.335 2034.040 ;
      LAYER pwell ;
        RECT 70.685 2028.245 74.865 2054.910 ;
        RECT 69.645 1993.735 74.865 2028.245 ;
        RECT 96.450 2064.770 104.025 2065.865 ;
        RECT 96.450 2040.880 100.480 2064.770 ;
        RECT 96.450 2027.385 99.180 2040.880 ;
        RECT 102.015 2033.840 104.025 2064.770 ;
      LAYER nwell ;
        RECT 104.835 2067.240 149.380 2068.670 ;
        RECT 104.835 2050.650 106.265 2067.240 ;
        RECT 104.835 2034.940 105.755 2050.650 ;
        RECT 115.655 2034.940 116.835 2067.240 ;
        RECT 126.225 2067.125 149.380 2067.240 ;
        RECT 126.225 2050.650 127.405 2067.125 ;
        RECT 133.955 2058.335 134.805 2067.125 ;
        RECT 147.950 2058.335 149.380 2067.125 ;
        RECT 126.735 2034.940 127.405 2050.650 ;
        RECT 163.945 2052.830 170.215 2068.450 ;
        RECT 174.655 2052.830 180.845 2068.450 ;
        RECT 163.945 2046.275 167.590 2052.830 ;
        RECT 163.945 2036.915 165.735 2046.275 ;
      LAYER pwell ;
        RECT 104.740 2033.840 105.045 2034.590 ;
        RECT 102.015 2027.385 105.045 2033.840 ;
        RECT 96.450 1993.735 98.035 2027.385 ;
        RECT 69.645 1993.215 98.035 1993.735 ;
        RECT 103.745 1997.300 105.045 2027.385 ;
        RECT 103.745 1993.215 107.065 1997.300 ;
      LAYER nwell ;
        RECT 112.260 1996.420 113.340 1996.495 ;
        RECT 111.720 1993.975 113.340 1996.420 ;
      LAYER pwell ;
        RECT 69.645 1987.785 107.065 1993.215 ;
      LAYER nwell ;
        RECT 108.180 1992.530 113.340 1993.975 ;
        RECT 108.180 1990.795 114.420 1992.530 ;
        RECT 107.600 1987.880 114.420 1990.795 ;
        RECT 118.765 1988.715 120.195 2012.815 ;
        RECT 138.980 1998.460 139.230 2001.535 ;
        RECT 138.980 1991.810 139.820 1998.460 ;
        RECT 137.660 1988.715 139.820 1991.810 ;
        RECT 141.980 1988.715 143.410 2011.515 ;
        RECT 176.920 1992.580 180.845 2052.830 ;
        RECT 107.600 1987.585 111.515 1987.880 ;
        RECT 118.765 1987.285 143.410 1988.715 ;
        RECT 190.675 1987.585 194.335 1991.110 ;
        RECT 3393.665 1929.890 3397.325 1933.415 ;
        RECT 3444.590 1932.285 3469.235 1933.715 ;
        RECT 3476.485 1933.120 3480.400 1933.415 ;
        RECT 3407.155 1868.170 3411.080 1928.420 ;
        RECT 3444.590 1909.485 3446.020 1932.285 ;
        RECT 3448.180 1929.190 3450.340 1932.285 ;
        RECT 3448.180 1922.540 3449.020 1929.190 ;
        RECT 3448.770 1919.465 3449.020 1922.540 ;
        RECT 3467.805 1908.185 3469.235 1932.285 ;
        RECT 3473.580 1930.205 3480.400 1933.120 ;
        RECT 3473.580 1928.470 3479.820 1930.205 ;
        RECT 3474.660 1927.025 3479.820 1928.470 ;
      LAYER pwell ;
        RECT 3480.935 1927.785 3518.355 1933.215 ;
      LAYER nwell ;
        RECT 3474.660 1924.580 3476.280 1927.025 ;
        RECT 3474.660 1924.505 3475.740 1924.580 ;
      LAYER pwell ;
        RECT 3480.935 1923.700 3484.255 1927.785 ;
        RECT 3482.955 1893.615 3484.255 1923.700 ;
        RECT 3489.965 1927.265 3518.355 1927.785 ;
        RECT 3489.965 1893.615 3491.550 1927.265 ;
        RECT 3482.955 1887.160 3485.985 1893.615 ;
        RECT 3482.955 1886.410 3483.260 1887.160 ;
      LAYER nwell ;
        RECT 3422.265 1874.725 3424.055 1884.085 ;
        RECT 3420.410 1868.170 3424.055 1874.725 ;
        RECT 29.770 1852.435 55.120 1852.440 ;
        RECT 21.025 1850.630 55.120 1852.435 ;
        RECT 21.025 1838.970 31.485 1850.630 ;
        RECT 21.025 1779.515 26.455 1838.970 ;
        RECT 29.525 1779.515 31.485 1838.970 ;
        RECT 21.025 1778.385 31.485 1779.515 ;
        RECT 53.310 1778.385 55.120 1850.630 ;
        RECT 21.025 1771.585 55.120 1778.385 ;
      LAYER pwell ;
        RECT 55.435 1771.710 59.315 1852.290 ;
      LAYER nwell ;
        RECT 59.615 1818.040 69.335 1852.440 ;
      LAYER pwell ;
        RECT 69.645 1849.865 104.025 1852.290 ;
        RECT 69.645 1838.910 74.865 1849.865 ;
      LAYER nwell ;
        RECT 59.620 1771.585 69.335 1818.040 ;
      LAYER pwell ;
        RECT 70.685 1812.245 74.865 1838.910 ;
        RECT 69.645 1777.735 74.865 1812.245 ;
        RECT 96.450 1848.770 104.025 1849.865 ;
        RECT 96.450 1824.880 100.480 1848.770 ;
        RECT 96.450 1811.385 99.180 1824.880 ;
        RECT 102.015 1817.840 104.025 1848.770 ;
      LAYER nwell ;
        RECT 104.835 1851.240 149.380 1852.670 ;
        RECT 3407.155 1852.550 3413.345 1868.170 ;
        RECT 3417.785 1852.550 3424.055 1868.170 ;
        RECT 3460.595 1870.350 3461.265 1886.060 ;
        RECT 3438.620 1853.875 3440.050 1862.665 ;
        RECT 3453.195 1853.875 3454.045 1862.665 ;
        RECT 3460.595 1853.875 3461.775 1870.350 ;
        RECT 3438.620 1853.760 3461.775 1853.875 ;
        RECT 3471.165 1853.760 3472.345 1886.060 ;
        RECT 3482.245 1870.350 3483.165 1886.060 ;
        RECT 3481.735 1853.760 3483.165 1870.350 ;
        RECT 104.835 1834.650 106.265 1851.240 ;
        RECT 104.835 1818.940 105.755 1834.650 ;
        RECT 115.655 1818.940 116.835 1851.240 ;
        RECT 126.225 1851.125 149.380 1851.240 ;
        RECT 126.225 1834.650 127.405 1851.125 ;
        RECT 133.955 1842.335 134.805 1851.125 ;
        RECT 147.950 1842.335 149.380 1851.125 ;
        RECT 126.735 1818.940 127.405 1834.650 ;
        RECT 163.945 1836.830 170.215 1852.450 ;
        RECT 174.655 1836.830 180.845 1852.450 ;
        RECT 3438.620 1852.330 3483.165 1853.760 ;
      LAYER pwell ;
        RECT 3483.975 1856.230 3485.985 1887.160 ;
        RECT 3488.820 1880.120 3491.550 1893.615 ;
        RECT 3487.520 1856.230 3491.550 1880.120 ;
        RECT 3483.975 1855.135 3491.550 1856.230 ;
        RECT 3513.135 1892.755 3518.355 1927.265 ;
        RECT 3513.135 1866.090 3517.315 1892.755 ;
      LAYER nwell ;
        RECT 3518.665 1886.960 3528.380 1933.415 ;
      LAYER pwell ;
        RECT 3513.135 1855.135 3518.355 1866.090 ;
        RECT 3483.975 1852.710 3518.355 1855.135 ;
      LAYER nwell ;
        RECT 3518.665 1852.560 3528.385 1886.960 ;
      LAYER pwell ;
        RECT 3528.685 1852.710 3532.565 1933.290 ;
      LAYER nwell ;
        RECT 3532.880 1926.615 3566.975 1933.415 ;
        RECT 3532.880 1854.370 3534.690 1926.615 ;
        RECT 3556.515 1925.485 3566.975 1926.615 ;
        RECT 3556.515 1866.030 3558.475 1925.485 ;
        RECT 3561.545 1866.030 3566.975 1925.485 ;
        RECT 3556.515 1854.370 3566.975 1866.030 ;
        RECT 3532.880 1852.565 3566.975 1854.370 ;
        RECT 3532.880 1852.560 3558.230 1852.565 ;
        RECT 163.945 1830.275 167.590 1836.830 ;
        RECT 163.945 1820.915 165.735 1830.275 ;
      LAYER pwell ;
        RECT 104.740 1817.840 105.045 1818.590 ;
        RECT 102.015 1811.385 105.045 1817.840 ;
        RECT 96.450 1777.735 98.035 1811.385 ;
        RECT 69.645 1777.215 98.035 1777.735 ;
        RECT 103.745 1781.300 105.045 1811.385 ;
        RECT 103.745 1777.215 107.065 1781.300 ;
      LAYER nwell ;
        RECT 112.260 1780.420 113.340 1780.495 ;
        RECT 111.720 1777.975 113.340 1780.420 ;
      LAYER pwell ;
        RECT 69.645 1771.785 107.065 1777.215 ;
      LAYER nwell ;
        RECT 108.180 1776.530 113.340 1777.975 ;
        RECT 108.180 1774.795 114.420 1776.530 ;
        RECT 107.600 1771.880 114.420 1774.795 ;
        RECT 118.765 1772.715 120.195 1796.815 ;
        RECT 138.980 1782.460 139.230 1785.535 ;
        RECT 138.980 1775.810 139.820 1782.460 ;
        RECT 137.660 1772.715 139.820 1775.810 ;
        RECT 141.980 1772.715 143.410 1795.515 ;
        RECT 176.920 1776.580 180.845 1836.830 ;
        RECT 107.600 1771.585 111.515 1771.880 ;
        RECT 118.765 1771.285 143.410 1772.715 ;
        RECT 190.675 1771.585 194.335 1775.110 ;
        RECT 3393.665 1703.890 3397.325 1707.415 ;
        RECT 3444.590 1706.285 3469.235 1707.715 ;
        RECT 3476.485 1707.120 3480.400 1707.415 ;
        RECT 3407.155 1642.170 3411.080 1702.420 ;
        RECT 3444.590 1683.485 3446.020 1706.285 ;
        RECT 3448.180 1703.190 3450.340 1706.285 ;
        RECT 3448.180 1696.540 3449.020 1703.190 ;
        RECT 3448.770 1693.465 3449.020 1696.540 ;
        RECT 3467.805 1682.185 3469.235 1706.285 ;
        RECT 3473.580 1704.205 3480.400 1707.120 ;
        RECT 3473.580 1702.470 3479.820 1704.205 ;
        RECT 3474.660 1701.025 3479.820 1702.470 ;
      LAYER pwell ;
        RECT 3480.935 1701.785 3518.355 1707.215 ;
      LAYER nwell ;
        RECT 3474.660 1698.580 3476.280 1701.025 ;
        RECT 3474.660 1698.505 3475.740 1698.580 ;
      LAYER pwell ;
        RECT 3480.935 1697.700 3484.255 1701.785 ;
        RECT 3482.955 1667.615 3484.255 1697.700 ;
        RECT 3489.965 1701.265 3518.355 1701.785 ;
        RECT 3489.965 1667.615 3491.550 1701.265 ;
        RECT 3482.955 1661.160 3485.985 1667.615 ;
        RECT 3482.955 1660.410 3483.260 1661.160 ;
      LAYER nwell ;
        RECT 3422.265 1648.725 3424.055 1658.085 ;
        RECT 3420.410 1642.170 3424.055 1648.725 ;
        RECT 29.770 1636.435 55.120 1636.440 ;
        RECT 21.025 1634.630 55.120 1636.435 ;
        RECT 21.025 1622.970 31.485 1634.630 ;
        RECT 21.025 1563.515 26.455 1622.970 ;
        RECT 29.525 1563.515 31.485 1622.970 ;
        RECT 21.025 1562.385 31.485 1563.515 ;
        RECT 53.310 1562.385 55.120 1634.630 ;
        RECT 21.025 1555.585 55.120 1562.385 ;
      LAYER pwell ;
        RECT 55.435 1555.710 59.315 1636.290 ;
      LAYER nwell ;
        RECT 59.615 1602.040 69.335 1636.440 ;
      LAYER pwell ;
        RECT 69.645 1633.865 104.025 1636.290 ;
        RECT 69.645 1622.910 74.865 1633.865 ;
      LAYER nwell ;
        RECT 59.620 1555.585 69.335 1602.040 ;
      LAYER pwell ;
        RECT 70.685 1596.245 74.865 1622.910 ;
        RECT 69.645 1561.735 74.865 1596.245 ;
        RECT 96.450 1632.770 104.025 1633.865 ;
        RECT 96.450 1608.880 100.480 1632.770 ;
        RECT 96.450 1595.385 99.180 1608.880 ;
        RECT 102.015 1601.840 104.025 1632.770 ;
      LAYER nwell ;
        RECT 104.835 1635.240 149.380 1636.670 ;
        RECT 104.835 1618.650 106.265 1635.240 ;
        RECT 104.835 1602.940 105.755 1618.650 ;
        RECT 115.655 1602.940 116.835 1635.240 ;
        RECT 126.225 1635.125 149.380 1635.240 ;
        RECT 126.225 1618.650 127.405 1635.125 ;
        RECT 133.955 1626.335 134.805 1635.125 ;
        RECT 147.950 1626.335 149.380 1635.125 ;
        RECT 126.735 1602.940 127.405 1618.650 ;
        RECT 163.945 1620.830 170.215 1636.450 ;
        RECT 174.655 1620.830 180.845 1636.450 ;
        RECT 3407.155 1626.550 3413.345 1642.170 ;
        RECT 3417.785 1626.550 3424.055 1642.170 ;
        RECT 3460.595 1644.350 3461.265 1660.060 ;
        RECT 3438.620 1627.875 3440.050 1636.665 ;
        RECT 3453.195 1627.875 3454.045 1636.665 ;
        RECT 3460.595 1627.875 3461.775 1644.350 ;
        RECT 3438.620 1627.760 3461.775 1627.875 ;
        RECT 3471.165 1627.760 3472.345 1660.060 ;
        RECT 3482.245 1644.350 3483.165 1660.060 ;
        RECT 3481.735 1627.760 3483.165 1644.350 ;
        RECT 3438.620 1626.330 3483.165 1627.760 ;
      LAYER pwell ;
        RECT 3483.975 1630.230 3485.985 1661.160 ;
        RECT 3488.820 1654.120 3491.550 1667.615 ;
        RECT 3487.520 1630.230 3491.550 1654.120 ;
        RECT 3483.975 1629.135 3491.550 1630.230 ;
        RECT 3513.135 1666.755 3518.355 1701.265 ;
        RECT 3513.135 1640.090 3517.315 1666.755 ;
      LAYER nwell ;
        RECT 3518.665 1660.960 3528.380 1707.415 ;
      LAYER pwell ;
        RECT 3513.135 1629.135 3518.355 1640.090 ;
        RECT 3483.975 1626.710 3518.355 1629.135 ;
      LAYER nwell ;
        RECT 3518.665 1626.560 3528.385 1660.960 ;
      LAYER pwell ;
        RECT 3528.685 1626.710 3532.565 1707.290 ;
      LAYER nwell ;
        RECT 3532.880 1700.615 3566.975 1707.415 ;
        RECT 3532.880 1628.370 3534.690 1700.615 ;
        RECT 3556.515 1699.485 3566.975 1700.615 ;
        RECT 3556.515 1640.030 3558.475 1699.485 ;
        RECT 3561.545 1640.030 3566.975 1699.485 ;
        RECT 3556.515 1628.370 3566.975 1640.030 ;
        RECT 3532.880 1626.565 3566.975 1628.370 ;
        RECT 3532.880 1626.560 3558.230 1626.565 ;
        RECT 163.945 1614.275 167.590 1620.830 ;
        RECT 163.945 1604.915 165.735 1614.275 ;
      LAYER pwell ;
        RECT 104.740 1601.840 105.045 1602.590 ;
        RECT 102.015 1595.385 105.045 1601.840 ;
        RECT 96.450 1561.735 98.035 1595.385 ;
        RECT 69.645 1561.215 98.035 1561.735 ;
        RECT 103.745 1565.300 105.045 1595.385 ;
        RECT 103.745 1561.215 107.065 1565.300 ;
      LAYER nwell ;
        RECT 112.260 1564.420 113.340 1564.495 ;
        RECT 111.720 1561.975 113.340 1564.420 ;
      LAYER pwell ;
        RECT 69.645 1555.785 107.065 1561.215 ;
      LAYER nwell ;
        RECT 108.180 1560.530 113.340 1561.975 ;
        RECT 108.180 1558.795 114.420 1560.530 ;
        RECT 107.600 1555.880 114.420 1558.795 ;
        RECT 118.765 1556.715 120.195 1580.815 ;
        RECT 138.980 1566.460 139.230 1569.535 ;
        RECT 138.980 1559.810 139.820 1566.460 ;
        RECT 137.660 1556.715 139.820 1559.810 ;
        RECT 141.980 1556.715 143.410 1579.515 ;
        RECT 176.920 1560.580 180.845 1620.830 ;
        RECT 107.600 1555.585 111.515 1555.880 ;
        RECT 118.765 1555.285 143.410 1556.715 ;
        RECT 190.675 1555.585 194.335 1559.110 ;
        RECT 3393.665 1478.890 3397.325 1482.415 ;
        RECT 3444.590 1481.285 3469.235 1482.715 ;
        RECT 3476.485 1482.120 3480.400 1482.415 ;
        RECT 29.770 1420.435 55.120 1420.440 ;
        RECT 21.025 1418.630 55.120 1420.435 ;
        RECT 21.025 1406.970 31.485 1418.630 ;
        RECT 21.025 1347.515 26.455 1406.970 ;
        RECT 29.525 1347.515 31.485 1406.970 ;
        RECT 21.025 1346.385 31.485 1347.515 ;
        RECT 53.310 1346.385 55.120 1418.630 ;
        RECT 21.025 1339.585 55.120 1346.385 ;
      LAYER pwell ;
        RECT 55.435 1339.710 59.315 1420.290 ;
      LAYER nwell ;
        RECT 59.615 1386.040 69.335 1420.440 ;
      LAYER pwell ;
        RECT 69.645 1417.865 104.025 1420.290 ;
        RECT 69.645 1406.910 74.865 1417.865 ;
      LAYER nwell ;
        RECT 59.620 1339.585 69.335 1386.040 ;
      LAYER pwell ;
        RECT 70.685 1380.245 74.865 1406.910 ;
        RECT 69.645 1345.735 74.865 1380.245 ;
        RECT 96.450 1416.770 104.025 1417.865 ;
        RECT 96.450 1392.880 100.480 1416.770 ;
        RECT 96.450 1379.385 99.180 1392.880 ;
        RECT 102.015 1385.840 104.025 1416.770 ;
      LAYER nwell ;
        RECT 104.835 1419.240 149.380 1420.670 ;
        RECT 104.835 1402.650 106.265 1419.240 ;
        RECT 104.835 1386.940 105.755 1402.650 ;
        RECT 115.655 1386.940 116.835 1419.240 ;
        RECT 126.225 1419.125 149.380 1419.240 ;
        RECT 126.225 1402.650 127.405 1419.125 ;
        RECT 133.955 1410.335 134.805 1419.125 ;
        RECT 147.950 1410.335 149.380 1419.125 ;
        RECT 126.735 1386.940 127.405 1402.650 ;
        RECT 163.945 1404.830 170.215 1420.450 ;
        RECT 174.655 1404.830 180.845 1420.450 ;
        RECT 163.945 1398.275 167.590 1404.830 ;
        RECT 163.945 1388.915 165.735 1398.275 ;
      LAYER pwell ;
        RECT 104.740 1385.840 105.045 1386.590 ;
        RECT 102.015 1379.385 105.045 1385.840 ;
        RECT 96.450 1345.735 98.035 1379.385 ;
        RECT 69.645 1345.215 98.035 1345.735 ;
        RECT 103.745 1349.300 105.045 1379.385 ;
        RECT 103.745 1345.215 107.065 1349.300 ;
      LAYER nwell ;
        RECT 112.260 1348.420 113.340 1348.495 ;
        RECT 111.720 1345.975 113.340 1348.420 ;
      LAYER pwell ;
        RECT 69.645 1339.785 107.065 1345.215 ;
      LAYER nwell ;
        RECT 108.180 1344.530 113.340 1345.975 ;
        RECT 108.180 1342.795 114.420 1344.530 ;
        RECT 107.600 1339.880 114.420 1342.795 ;
        RECT 118.765 1340.715 120.195 1364.815 ;
        RECT 138.980 1350.460 139.230 1353.535 ;
        RECT 138.980 1343.810 139.820 1350.460 ;
        RECT 137.660 1340.715 139.820 1343.810 ;
        RECT 141.980 1340.715 143.410 1363.515 ;
        RECT 176.920 1344.580 180.845 1404.830 ;
        RECT 3407.155 1417.170 3411.080 1477.420 ;
        RECT 3444.590 1458.485 3446.020 1481.285 ;
        RECT 3448.180 1478.190 3450.340 1481.285 ;
        RECT 3448.180 1471.540 3449.020 1478.190 ;
        RECT 3448.770 1468.465 3449.020 1471.540 ;
        RECT 3467.805 1457.185 3469.235 1481.285 ;
        RECT 3473.580 1479.205 3480.400 1482.120 ;
        RECT 3473.580 1477.470 3479.820 1479.205 ;
        RECT 3474.660 1476.025 3479.820 1477.470 ;
      LAYER pwell ;
        RECT 3480.935 1476.785 3518.355 1482.215 ;
      LAYER nwell ;
        RECT 3474.660 1473.580 3476.280 1476.025 ;
        RECT 3474.660 1473.505 3475.740 1473.580 ;
      LAYER pwell ;
        RECT 3480.935 1472.700 3484.255 1476.785 ;
        RECT 3482.955 1442.615 3484.255 1472.700 ;
        RECT 3489.965 1476.265 3518.355 1476.785 ;
        RECT 3489.965 1442.615 3491.550 1476.265 ;
        RECT 3482.955 1436.160 3485.985 1442.615 ;
        RECT 3482.955 1435.410 3483.260 1436.160 ;
      LAYER nwell ;
        RECT 3422.265 1423.725 3424.055 1433.085 ;
        RECT 3420.410 1417.170 3424.055 1423.725 ;
        RECT 3407.155 1401.550 3413.345 1417.170 ;
        RECT 3417.785 1401.550 3424.055 1417.170 ;
        RECT 3460.595 1419.350 3461.265 1435.060 ;
        RECT 3438.620 1402.875 3440.050 1411.665 ;
        RECT 3453.195 1402.875 3454.045 1411.665 ;
        RECT 3460.595 1402.875 3461.775 1419.350 ;
        RECT 3438.620 1402.760 3461.775 1402.875 ;
        RECT 3471.165 1402.760 3472.345 1435.060 ;
        RECT 3482.245 1419.350 3483.165 1435.060 ;
        RECT 3481.735 1402.760 3483.165 1419.350 ;
        RECT 3438.620 1401.330 3483.165 1402.760 ;
      LAYER pwell ;
        RECT 3483.975 1405.230 3485.985 1436.160 ;
        RECT 3488.820 1429.120 3491.550 1442.615 ;
        RECT 3487.520 1405.230 3491.550 1429.120 ;
        RECT 3483.975 1404.135 3491.550 1405.230 ;
        RECT 3513.135 1441.755 3518.355 1476.265 ;
        RECT 3513.135 1415.090 3517.315 1441.755 ;
      LAYER nwell ;
        RECT 3518.665 1435.960 3528.380 1482.415 ;
      LAYER pwell ;
        RECT 3513.135 1404.135 3518.355 1415.090 ;
        RECT 3483.975 1401.710 3518.355 1404.135 ;
      LAYER nwell ;
        RECT 3518.665 1401.560 3528.385 1435.960 ;
      LAYER pwell ;
        RECT 3528.685 1401.710 3532.565 1482.290 ;
      LAYER nwell ;
        RECT 3532.880 1475.615 3566.975 1482.415 ;
        RECT 3532.880 1403.370 3534.690 1475.615 ;
        RECT 3556.515 1474.485 3566.975 1475.615 ;
        RECT 3556.515 1415.030 3558.475 1474.485 ;
        RECT 3561.545 1415.030 3566.975 1474.485 ;
        RECT 3556.515 1403.370 3566.975 1415.030 ;
        RECT 3532.880 1401.565 3566.975 1403.370 ;
        RECT 3532.880 1401.560 3558.230 1401.565 ;
        RECT 107.600 1339.585 111.515 1339.880 ;
        RECT 118.765 1339.285 143.410 1340.715 ;
        RECT 190.675 1339.585 194.335 1343.110 ;
        RECT 3393.665 1253.890 3397.325 1257.415 ;
        RECT 3444.590 1256.285 3469.235 1257.715 ;
        RECT 3476.485 1257.120 3480.400 1257.415 ;
        RECT 29.770 1204.435 55.120 1204.440 ;
        RECT 21.025 1202.630 55.120 1204.435 ;
        RECT 21.025 1190.970 31.485 1202.630 ;
        RECT 21.025 1131.515 26.455 1190.970 ;
        RECT 29.525 1131.515 31.485 1190.970 ;
        RECT 21.025 1130.385 31.485 1131.515 ;
        RECT 53.310 1130.385 55.120 1202.630 ;
        RECT 21.025 1123.585 55.120 1130.385 ;
      LAYER pwell ;
        RECT 55.435 1123.710 59.315 1204.290 ;
      LAYER nwell ;
        RECT 59.615 1170.040 69.335 1204.440 ;
      LAYER pwell ;
        RECT 69.645 1201.865 104.025 1204.290 ;
        RECT 69.645 1190.910 74.865 1201.865 ;
      LAYER nwell ;
        RECT 59.620 1123.585 69.335 1170.040 ;
      LAYER pwell ;
        RECT 70.685 1164.245 74.865 1190.910 ;
        RECT 69.645 1129.735 74.865 1164.245 ;
        RECT 96.450 1200.770 104.025 1201.865 ;
        RECT 96.450 1176.880 100.480 1200.770 ;
        RECT 96.450 1163.385 99.180 1176.880 ;
        RECT 102.015 1169.840 104.025 1200.770 ;
      LAYER nwell ;
        RECT 104.835 1203.240 149.380 1204.670 ;
        RECT 104.835 1186.650 106.265 1203.240 ;
        RECT 104.835 1170.940 105.755 1186.650 ;
        RECT 115.655 1170.940 116.835 1203.240 ;
        RECT 126.225 1203.125 149.380 1203.240 ;
        RECT 126.225 1186.650 127.405 1203.125 ;
        RECT 133.955 1194.335 134.805 1203.125 ;
        RECT 147.950 1194.335 149.380 1203.125 ;
        RECT 126.735 1170.940 127.405 1186.650 ;
        RECT 163.945 1188.830 170.215 1204.450 ;
        RECT 174.655 1188.830 180.845 1204.450 ;
        RECT 163.945 1182.275 167.590 1188.830 ;
        RECT 163.945 1172.915 165.735 1182.275 ;
      LAYER pwell ;
        RECT 104.740 1169.840 105.045 1170.590 ;
        RECT 102.015 1163.385 105.045 1169.840 ;
        RECT 96.450 1129.735 98.035 1163.385 ;
        RECT 69.645 1129.215 98.035 1129.735 ;
        RECT 103.745 1133.300 105.045 1163.385 ;
        RECT 103.745 1129.215 107.065 1133.300 ;
      LAYER nwell ;
        RECT 112.260 1132.420 113.340 1132.495 ;
        RECT 111.720 1129.975 113.340 1132.420 ;
      LAYER pwell ;
        RECT 69.645 1123.785 107.065 1129.215 ;
      LAYER nwell ;
        RECT 108.180 1128.530 113.340 1129.975 ;
        RECT 108.180 1126.795 114.420 1128.530 ;
        RECT 107.600 1123.880 114.420 1126.795 ;
        RECT 118.765 1124.715 120.195 1148.815 ;
        RECT 138.980 1134.460 139.230 1137.535 ;
        RECT 138.980 1127.810 139.820 1134.460 ;
        RECT 137.660 1124.715 139.820 1127.810 ;
        RECT 141.980 1124.715 143.410 1147.515 ;
        RECT 176.920 1128.580 180.845 1188.830 ;
        RECT 3407.155 1192.170 3411.080 1252.420 ;
        RECT 3444.590 1233.485 3446.020 1256.285 ;
        RECT 3448.180 1253.190 3450.340 1256.285 ;
        RECT 3448.180 1246.540 3449.020 1253.190 ;
        RECT 3448.770 1243.465 3449.020 1246.540 ;
        RECT 3467.805 1232.185 3469.235 1256.285 ;
        RECT 3473.580 1254.205 3480.400 1257.120 ;
        RECT 3473.580 1252.470 3479.820 1254.205 ;
        RECT 3474.660 1251.025 3479.820 1252.470 ;
      LAYER pwell ;
        RECT 3480.935 1251.785 3518.355 1257.215 ;
      LAYER nwell ;
        RECT 3474.660 1248.580 3476.280 1251.025 ;
        RECT 3474.660 1248.505 3475.740 1248.580 ;
      LAYER pwell ;
        RECT 3480.935 1247.700 3484.255 1251.785 ;
        RECT 3482.955 1217.615 3484.255 1247.700 ;
        RECT 3489.965 1251.265 3518.355 1251.785 ;
        RECT 3489.965 1217.615 3491.550 1251.265 ;
        RECT 3482.955 1211.160 3485.985 1217.615 ;
        RECT 3482.955 1210.410 3483.260 1211.160 ;
      LAYER nwell ;
        RECT 3422.265 1198.725 3424.055 1208.085 ;
        RECT 3420.410 1192.170 3424.055 1198.725 ;
        RECT 3407.155 1176.550 3413.345 1192.170 ;
        RECT 3417.785 1176.550 3424.055 1192.170 ;
        RECT 3460.595 1194.350 3461.265 1210.060 ;
        RECT 3438.620 1177.875 3440.050 1186.665 ;
        RECT 3453.195 1177.875 3454.045 1186.665 ;
        RECT 3460.595 1177.875 3461.775 1194.350 ;
        RECT 3438.620 1177.760 3461.775 1177.875 ;
        RECT 3471.165 1177.760 3472.345 1210.060 ;
        RECT 3482.245 1194.350 3483.165 1210.060 ;
        RECT 3481.735 1177.760 3483.165 1194.350 ;
        RECT 3438.620 1176.330 3483.165 1177.760 ;
      LAYER pwell ;
        RECT 3483.975 1180.230 3485.985 1211.160 ;
        RECT 3488.820 1204.120 3491.550 1217.615 ;
        RECT 3487.520 1180.230 3491.550 1204.120 ;
        RECT 3483.975 1179.135 3491.550 1180.230 ;
        RECT 3513.135 1216.755 3518.355 1251.265 ;
        RECT 3513.135 1190.090 3517.315 1216.755 ;
      LAYER nwell ;
        RECT 3518.665 1210.960 3528.380 1257.415 ;
      LAYER pwell ;
        RECT 3513.135 1179.135 3518.355 1190.090 ;
        RECT 3483.975 1176.710 3518.355 1179.135 ;
      LAYER nwell ;
        RECT 3518.665 1176.560 3528.385 1210.960 ;
      LAYER pwell ;
        RECT 3528.685 1176.710 3532.565 1257.290 ;
      LAYER nwell ;
        RECT 3532.880 1250.615 3566.975 1257.415 ;
        RECT 3532.880 1178.370 3534.690 1250.615 ;
        RECT 3556.515 1249.485 3566.975 1250.615 ;
        RECT 3556.515 1190.030 3558.475 1249.485 ;
        RECT 3561.545 1190.030 3566.975 1249.485 ;
        RECT 3556.515 1178.370 3566.975 1190.030 ;
        RECT 3532.880 1176.565 3566.975 1178.370 ;
        RECT 3532.880 1176.560 3558.230 1176.565 ;
        RECT 107.600 1123.585 111.515 1123.880 ;
        RECT 118.765 1123.285 143.410 1124.715 ;
        RECT 190.675 1123.585 194.335 1127.110 ;
        RECT 3393.665 1027.890 3397.325 1031.415 ;
        RECT 3444.590 1030.285 3469.235 1031.715 ;
        RECT 3476.485 1031.120 3480.400 1031.415 ;
        RECT 29.770 988.435 55.120 988.440 ;
        RECT 21.025 986.630 55.120 988.435 ;
        RECT 21.025 974.970 31.485 986.630 ;
        RECT 21.025 915.515 26.455 974.970 ;
        RECT 29.525 915.515 31.485 974.970 ;
        RECT 21.025 914.385 31.485 915.515 ;
        RECT 53.310 914.385 55.120 986.630 ;
        RECT 21.025 907.585 55.120 914.385 ;
      LAYER pwell ;
        RECT 55.435 907.710 59.315 988.290 ;
      LAYER nwell ;
        RECT 59.615 954.040 69.335 988.440 ;
      LAYER pwell ;
        RECT 69.645 985.865 104.025 988.290 ;
        RECT 69.645 974.910 74.865 985.865 ;
      LAYER nwell ;
        RECT 59.620 907.585 69.335 954.040 ;
      LAYER pwell ;
        RECT 70.685 948.245 74.865 974.910 ;
        RECT 69.645 913.735 74.865 948.245 ;
        RECT 96.450 984.770 104.025 985.865 ;
        RECT 96.450 960.880 100.480 984.770 ;
        RECT 96.450 947.385 99.180 960.880 ;
        RECT 102.015 953.840 104.025 984.770 ;
      LAYER nwell ;
        RECT 104.835 987.240 149.380 988.670 ;
        RECT 104.835 970.650 106.265 987.240 ;
        RECT 104.835 954.940 105.755 970.650 ;
        RECT 115.655 954.940 116.835 987.240 ;
        RECT 126.225 987.125 149.380 987.240 ;
        RECT 126.225 970.650 127.405 987.125 ;
        RECT 133.955 978.335 134.805 987.125 ;
        RECT 147.950 978.335 149.380 987.125 ;
        RECT 126.735 954.940 127.405 970.650 ;
        RECT 163.945 972.830 170.215 988.450 ;
        RECT 174.655 972.830 180.845 988.450 ;
        RECT 163.945 966.275 167.590 972.830 ;
        RECT 163.945 956.915 165.735 966.275 ;
      LAYER pwell ;
        RECT 104.740 953.840 105.045 954.590 ;
        RECT 102.015 947.385 105.045 953.840 ;
        RECT 96.450 913.735 98.035 947.385 ;
        RECT 69.645 913.215 98.035 913.735 ;
        RECT 103.745 917.300 105.045 947.385 ;
        RECT 103.745 913.215 107.065 917.300 ;
      LAYER nwell ;
        RECT 112.260 916.420 113.340 916.495 ;
        RECT 111.720 913.975 113.340 916.420 ;
      LAYER pwell ;
        RECT 69.645 907.785 107.065 913.215 ;
      LAYER nwell ;
        RECT 108.180 912.530 113.340 913.975 ;
        RECT 108.180 910.795 114.420 912.530 ;
        RECT 107.600 907.880 114.420 910.795 ;
        RECT 118.765 908.715 120.195 932.815 ;
        RECT 138.980 918.460 139.230 921.535 ;
        RECT 138.980 911.810 139.820 918.460 ;
        RECT 137.660 908.715 139.820 911.810 ;
        RECT 141.980 908.715 143.410 931.515 ;
        RECT 176.920 912.580 180.845 972.830 ;
        RECT 3407.155 966.170 3411.080 1026.420 ;
        RECT 3444.590 1007.485 3446.020 1030.285 ;
        RECT 3448.180 1027.190 3450.340 1030.285 ;
        RECT 3448.180 1020.540 3449.020 1027.190 ;
        RECT 3448.770 1017.465 3449.020 1020.540 ;
        RECT 3467.805 1006.185 3469.235 1030.285 ;
        RECT 3473.580 1028.205 3480.400 1031.120 ;
        RECT 3473.580 1026.470 3479.820 1028.205 ;
        RECT 3474.660 1025.025 3479.820 1026.470 ;
      LAYER pwell ;
        RECT 3480.935 1025.785 3518.355 1031.215 ;
      LAYER nwell ;
        RECT 3474.660 1022.580 3476.280 1025.025 ;
        RECT 3474.660 1022.505 3475.740 1022.580 ;
      LAYER pwell ;
        RECT 3480.935 1021.700 3484.255 1025.785 ;
        RECT 3482.955 991.615 3484.255 1021.700 ;
        RECT 3489.965 1025.265 3518.355 1025.785 ;
        RECT 3489.965 991.615 3491.550 1025.265 ;
        RECT 3482.955 985.160 3485.985 991.615 ;
        RECT 3482.955 984.410 3483.260 985.160 ;
      LAYER nwell ;
        RECT 3422.265 972.725 3424.055 982.085 ;
        RECT 3420.410 966.170 3424.055 972.725 ;
        RECT 3407.155 950.550 3413.345 966.170 ;
        RECT 3417.785 950.550 3424.055 966.170 ;
        RECT 3460.595 968.350 3461.265 984.060 ;
        RECT 3438.620 951.875 3440.050 960.665 ;
        RECT 3453.195 951.875 3454.045 960.665 ;
        RECT 3460.595 951.875 3461.775 968.350 ;
        RECT 3438.620 951.760 3461.775 951.875 ;
        RECT 3471.165 951.760 3472.345 984.060 ;
        RECT 3482.245 968.350 3483.165 984.060 ;
        RECT 3481.735 951.760 3483.165 968.350 ;
        RECT 3438.620 950.330 3483.165 951.760 ;
      LAYER pwell ;
        RECT 3483.975 954.230 3485.985 985.160 ;
        RECT 3488.820 978.120 3491.550 991.615 ;
        RECT 3487.520 954.230 3491.550 978.120 ;
        RECT 3483.975 953.135 3491.550 954.230 ;
        RECT 3513.135 990.755 3518.355 1025.265 ;
        RECT 3513.135 964.090 3517.315 990.755 ;
      LAYER nwell ;
        RECT 3518.665 984.960 3528.380 1031.415 ;
      LAYER pwell ;
        RECT 3513.135 953.135 3518.355 964.090 ;
        RECT 3483.975 950.710 3518.355 953.135 ;
      LAYER nwell ;
        RECT 3518.665 950.560 3528.385 984.960 ;
      LAYER pwell ;
        RECT 3528.685 950.710 3532.565 1031.290 ;
      LAYER nwell ;
        RECT 3532.880 1024.615 3566.975 1031.415 ;
        RECT 3532.880 952.370 3534.690 1024.615 ;
        RECT 3556.515 1023.485 3566.975 1024.615 ;
        RECT 3556.515 964.030 3558.475 1023.485 ;
        RECT 3561.545 964.030 3566.975 1023.485 ;
        RECT 3556.515 952.370 3566.975 964.030 ;
        RECT 3532.880 950.565 3566.975 952.370 ;
        RECT 3532.880 950.560 3558.230 950.565 ;
        RECT 107.600 907.585 111.515 907.880 ;
        RECT 118.765 907.285 143.410 908.715 ;
        RECT 190.675 907.585 194.335 911.110 ;
        RECT 3393.665 802.890 3397.325 806.415 ;
        RECT 3444.590 805.285 3469.235 806.715 ;
        RECT 3476.485 806.120 3480.400 806.415 ;
        RECT 3407.155 741.170 3411.080 801.420 ;
        RECT 3444.590 782.485 3446.020 805.285 ;
        RECT 3448.180 802.190 3450.340 805.285 ;
        RECT 3448.180 795.540 3449.020 802.190 ;
        RECT 3448.770 792.465 3449.020 795.540 ;
        RECT 3467.805 781.185 3469.235 805.285 ;
        RECT 3473.580 803.205 3480.400 806.120 ;
        RECT 3473.580 801.470 3479.820 803.205 ;
        RECT 3474.660 800.025 3479.820 801.470 ;
      LAYER pwell ;
        RECT 3480.935 800.785 3518.355 806.215 ;
      LAYER nwell ;
        RECT 3474.660 797.580 3476.280 800.025 ;
        RECT 3474.660 797.505 3475.740 797.580 ;
      LAYER pwell ;
        RECT 3480.935 796.700 3484.255 800.785 ;
        RECT 3482.955 766.615 3484.255 796.700 ;
        RECT 3489.965 800.265 3518.355 800.785 ;
        RECT 3489.965 766.615 3491.550 800.265 ;
        RECT 3482.955 760.160 3485.985 766.615 ;
        RECT 3482.955 759.410 3483.260 760.160 ;
      LAYER nwell ;
        RECT 3422.265 747.725 3424.055 757.085 ;
        RECT 3420.410 741.170 3424.055 747.725 ;
        RECT 3407.155 725.550 3413.345 741.170 ;
        RECT 3417.785 725.550 3424.055 741.170 ;
        RECT 3460.595 743.350 3461.265 759.060 ;
        RECT 3438.620 726.875 3440.050 735.665 ;
        RECT 3453.195 726.875 3454.045 735.665 ;
        RECT 3460.595 726.875 3461.775 743.350 ;
        RECT 3438.620 726.760 3461.775 726.875 ;
        RECT 3471.165 726.760 3472.345 759.060 ;
        RECT 3482.245 743.350 3483.165 759.060 ;
        RECT 3481.735 726.760 3483.165 743.350 ;
        RECT 3438.620 725.330 3483.165 726.760 ;
      LAYER pwell ;
        RECT 3483.975 729.230 3485.985 760.160 ;
        RECT 3488.820 753.120 3491.550 766.615 ;
        RECT 3487.520 729.230 3491.550 753.120 ;
        RECT 3483.975 728.135 3491.550 729.230 ;
        RECT 3513.135 765.755 3518.355 800.265 ;
        RECT 3513.135 739.090 3517.315 765.755 ;
      LAYER nwell ;
        RECT 3518.665 759.960 3528.380 806.415 ;
      LAYER pwell ;
        RECT 3513.135 728.135 3518.355 739.090 ;
        RECT 3483.975 725.710 3518.355 728.135 ;
      LAYER nwell ;
        RECT 3518.665 725.560 3528.385 759.960 ;
      LAYER pwell ;
        RECT 3528.685 725.710 3532.565 806.290 ;
      LAYER nwell ;
        RECT 3532.880 799.615 3566.975 806.415 ;
        RECT 3532.880 727.370 3534.690 799.615 ;
        RECT 3556.515 798.485 3566.975 799.615 ;
        RECT 3556.515 739.030 3558.475 798.485 ;
        RECT 3561.545 739.030 3566.975 798.485 ;
        RECT 3556.515 727.370 3566.975 739.030 ;
        RECT 3532.880 725.565 3566.975 727.370 ;
        RECT 3532.880 725.560 3558.230 725.565 ;
        RECT 197.795 562.860 199.315 621.965 ;
        RECT 3393.665 576.890 3397.325 580.415 ;
        RECT 3444.590 579.285 3469.235 580.715 ;
        RECT 3476.485 580.120 3480.400 580.415 ;
      LAYER pwell ;
        RECT 176.210 554.495 199.065 562.285 ;
      LAYER nwell ;
        RECT 3407.155 515.170 3411.080 575.420 ;
        RECT 3444.590 556.485 3446.020 579.285 ;
        RECT 3448.180 576.190 3450.340 579.285 ;
        RECT 3448.180 569.540 3449.020 576.190 ;
        RECT 3448.770 566.465 3449.020 569.540 ;
        RECT 3467.805 555.185 3469.235 579.285 ;
        RECT 3473.580 577.205 3480.400 580.120 ;
        RECT 3473.580 575.470 3479.820 577.205 ;
        RECT 3474.660 574.025 3479.820 575.470 ;
      LAYER pwell ;
        RECT 3480.935 574.785 3518.355 580.215 ;
      LAYER nwell ;
        RECT 3474.660 571.580 3476.280 574.025 ;
        RECT 3474.660 571.505 3475.740 571.580 ;
      LAYER pwell ;
        RECT 3480.935 570.700 3484.255 574.785 ;
        RECT 3482.955 540.615 3484.255 570.700 ;
        RECT 3489.965 574.265 3518.355 574.785 ;
        RECT 3489.965 540.615 3491.550 574.265 ;
        RECT 3482.955 534.160 3485.985 540.615 ;
        RECT 3482.955 533.410 3483.260 534.160 ;
      LAYER nwell ;
        RECT 3422.265 521.725 3424.055 531.085 ;
        RECT 3420.410 515.170 3424.055 521.725 ;
        RECT 3407.155 499.550 3413.345 515.170 ;
        RECT 3417.785 499.550 3424.055 515.170 ;
        RECT 3460.595 517.350 3461.265 533.060 ;
        RECT 3438.620 500.875 3440.050 509.665 ;
        RECT 3453.195 500.875 3454.045 509.665 ;
        RECT 3460.595 500.875 3461.775 517.350 ;
        RECT 3438.620 500.760 3461.775 500.875 ;
        RECT 3471.165 500.760 3472.345 533.060 ;
        RECT 3482.245 517.350 3483.165 533.060 ;
        RECT 3481.735 500.760 3483.165 517.350 ;
        RECT 3438.620 499.330 3483.165 500.760 ;
      LAYER pwell ;
        RECT 3483.975 503.230 3485.985 534.160 ;
        RECT 3488.820 527.120 3491.550 540.615 ;
        RECT 3487.520 503.230 3491.550 527.120 ;
        RECT 3483.975 502.135 3491.550 503.230 ;
        RECT 3513.135 539.755 3518.355 574.265 ;
        RECT 3513.135 513.090 3517.315 539.755 ;
      LAYER nwell ;
        RECT 3518.665 533.960 3528.380 580.415 ;
      LAYER pwell ;
        RECT 3513.135 502.135 3518.355 513.090 ;
        RECT 3483.975 499.710 3518.355 502.135 ;
      LAYER nwell ;
        RECT 3518.665 499.560 3528.385 533.960 ;
      LAYER pwell ;
        RECT 3528.685 499.710 3532.565 580.290 ;
      LAYER nwell ;
        RECT 3532.880 573.615 3566.975 580.415 ;
        RECT 3532.880 501.370 3534.690 573.615 ;
        RECT 3556.515 572.485 3566.975 573.615 ;
        RECT 3556.515 513.030 3558.475 572.485 ;
        RECT 3561.545 513.030 3566.975 572.485 ;
        RECT 3556.515 501.370 3566.975 513.030 ;
        RECT 3532.880 499.565 3566.975 501.370 ;
        RECT 3532.880 499.560 3558.230 499.565 ;
        RECT 398.035 197.795 457.140 199.315 ;
        RECT 2849.035 197.795 2908.140 199.315 ;
        RECT 3118.035 197.795 3177.140 199.315 ;
        RECT 1008.890 190.675 1012.415 194.335 ;
        RECT 1551.890 190.675 1555.415 194.335 ;
        RECT 1825.890 190.675 1829.415 194.335 ;
        RECT 2099.890 190.675 2103.415 194.335 ;
        RECT 2373.890 190.675 2377.415 194.335 ;
        RECT 2647.890 190.675 2651.415 194.335 ;
        RECT 931.550 176.920 1007.420 180.845 ;
        RECT 1474.550 176.920 1550.420 180.845 ;
        RECT 1748.550 176.920 1824.420 180.845 ;
        RECT 2022.550 176.920 2098.420 180.845 ;
        RECT 2296.550 176.920 2372.420 180.845 ;
        RECT 2570.550 176.920 2646.420 180.845 ;
        RECT 931.550 174.655 947.170 176.920 ;
        RECT 1474.550 174.655 1490.170 176.920 ;
        RECT 1748.550 174.655 1764.170 176.920 ;
        RECT 2022.550 174.655 2038.170 176.920 ;
        RECT 2296.550 174.655 2312.170 176.920 ;
        RECT 2570.550 174.655 2586.170 176.920 ;
      LAYER pwell ;
        RECT 3177.715 176.210 3185.505 199.065 ;
      LAYER nwell ;
        RECT 931.550 167.590 947.170 170.215 ;
        RECT 1474.550 167.590 1490.170 170.215 ;
        RECT 1748.550 167.590 1764.170 170.215 ;
        RECT 2022.550 167.590 2038.170 170.215 ;
        RECT 2296.550 167.590 2312.170 170.215 ;
        RECT 2570.550 167.590 2586.170 170.215 ;
        RECT 931.550 165.735 953.725 167.590 ;
        RECT 1474.550 165.735 1496.725 167.590 ;
        RECT 1748.550 165.735 1770.725 167.590 ;
        RECT 2022.550 165.735 2044.725 167.590 ;
        RECT 2296.550 165.735 2318.725 167.590 ;
        RECT 2570.550 165.735 2592.725 167.590 ;
        RECT 931.550 163.945 963.085 165.735 ;
        RECT 1474.550 163.945 1506.085 165.735 ;
        RECT 1748.550 163.945 1780.085 165.735 ;
        RECT 2022.550 163.945 2054.085 165.735 ;
        RECT 2296.550 163.945 2328.085 165.735 ;
        RECT 2570.550 163.945 2602.085 165.735 ;
        RECT 931.330 147.950 941.665 149.380 ;
        RECT 1474.330 147.950 1484.665 149.380 ;
        RECT 1748.330 147.950 1758.665 149.380 ;
        RECT 2022.330 147.950 2032.665 149.380 ;
        RECT 2296.330 147.950 2306.665 149.380 ;
        RECT 2570.330 147.950 2580.665 149.380 ;
        RECT 931.330 134.805 932.875 147.950 ;
        RECT 988.485 141.980 1012.715 143.410 ;
        RECT 1011.285 139.820 1012.715 141.980 ;
        RECT 1001.540 139.230 1012.715 139.820 ;
        RECT 998.465 138.980 1012.715 139.230 ;
        RECT 1008.190 137.660 1012.715 138.980 ;
        RECT 931.330 133.955 941.665 134.805 ;
        RECT 931.330 127.405 932.875 133.955 ;
        RECT 931.330 126.735 965.060 127.405 ;
        RECT 931.330 126.225 949.350 126.735 ;
        RECT 931.330 116.835 932.760 126.225 ;
        RECT 1011.285 120.195 1012.715 137.660 ;
        RECT 987.185 118.765 1012.715 120.195 ;
        RECT 1474.330 134.805 1475.875 147.950 ;
        RECT 1531.485 141.980 1555.715 143.410 ;
        RECT 1554.285 139.820 1555.715 141.980 ;
        RECT 1544.540 139.230 1555.715 139.820 ;
        RECT 1541.465 138.980 1555.715 139.230 ;
        RECT 1551.190 137.660 1555.715 138.980 ;
        RECT 1474.330 133.955 1484.665 134.805 ;
        RECT 1474.330 127.405 1475.875 133.955 ;
        RECT 1474.330 126.735 1508.060 127.405 ;
        RECT 1474.330 126.225 1492.350 126.735 ;
        RECT 1474.330 116.835 1475.760 126.225 ;
        RECT 1554.285 120.195 1555.715 137.660 ;
        RECT 1530.185 118.765 1555.715 120.195 ;
        RECT 1748.330 134.805 1749.875 147.950 ;
        RECT 1805.485 141.980 1829.715 143.410 ;
        RECT 1828.285 139.820 1829.715 141.980 ;
        RECT 1818.540 139.230 1829.715 139.820 ;
        RECT 1815.465 138.980 1829.715 139.230 ;
        RECT 1825.190 137.660 1829.715 138.980 ;
        RECT 1748.330 133.955 1758.665 134.805 ;
        RECT 1748.330 127.405 1749.875 133.955 ;
        RECT 1748.330 126.735 1782.060 127.405 ;
        RECT 1748.330 126.225 1766.350 126.735 ;
        RECT 1748.330 116.835 1749.760 126.225 ;
        RECT 1828.285 120.195 1829.715 137.660 ;
        RECT 1804.185 118.765 1829.715 120.195 ;
        RECT 2022.330 134.805 2023.875 147.950 ;
        RECT 2079.485 141.980 2103.715 143.410 ;
        RECT 2102.285 139.820 2103.715 141.980 ;
        RECT 2092.540 139.230 2103.715 139.820 ;
        RECT 2089.465 138.980 2103.715 139.230 ;
        RECT 2099.190 137.660 2103.715 138.980 ;
        RECT 2022.330 133.955 2032.665 134.805 ;
        RECT 2022.330 127.405 2023.875 133.955 ;
        RECT 2022.330 126.735 2056.060 127.405 ;
        RECT 2022.330 126.225 2040.350 126.735 ;
        RECT 2022.330 116.835 2023.760 126.225 ;
        RECT 2102.285 120.195 2103.715 137.660 ;
        RECT 2078.185 118.765 2103.715 120.195 ;
        RECT 2296.330 134.805 2297.875 147.950 ;
        RECT 2353.485 141.980 2377.715 143.410 ;
        RECT 2376.285 139.820 2377.715 141.980 ;
        RECT 2366.540 139.230 2377.715 139.820 ;
        RECT 2363.465 138.980 2377.715 139.230 ;
        RECT 2373.190 137.660 2377.715 138.980 ;
        RECT 2296.330 133.955 2306.665 134.805 ;
        RECT 2296.330 127.405 2297.875 133.955 ;
        RECT 2296.330 126.735 2330.060 127.405 ;
        RECT 2296.330 126.225 2314.350 126.735 ;
        RECT 2296.330 116.835 2297.760 126.225 ;
        RECT 2376.285 120.195 2377.715 137.660 ;
        RECT 2352.185 118.765 2377.715 120.195 ;
        RECT 2570.330 134.805 2571.875 147.950 ;
        RECT 2627.485 141.980 2651.715 143.410 ;
        RECT 2650.285 139.820 2651.715 141.980 ;
        RECT 2640.540 139.230 2651.715 139.820 ;
        RECT 2637.465 138.980 2651.715 139.230 ;
        RECT 2647.190 137.660 2651.715 138.980 ;
        RECT 2570.330 133.955 2580.665 134.805 ;
        RECT 2570.330 127.405 2571.875 133.955 ;
        RECT 2570.330 126.735 2604.060 127.405 ;
        RECT 2570.330 126.225 2588.350 126.735 ;
        RECT 2570.330 116.835 2571.760 126.225 ;
        RECT 2650.285 120.195 2651.715 137.660 ;
        RECT 2626.185 118.765 2651.715 120.195 ;
        RECT 931.330 115.655 965.060 116.835 ;
        RECT 1474.330 115.655 1508.060 116.835 ;
        RECT 1748.330 115.655 1782.060 116.835 ;
        RECT 2022.330 115.655 2056.060 116.835 ;
        RECT 2296.330 115.655 2330.060 116.835 ;
        RECT 2570.330 115.655 2604.060 116.835 ;
        RECT 931.330 106.265 932.760 115.655 ;
        RECT 1007.470 113.340 1012.120 114.420 ;
        RECT 1003.505 112.260 1012.120 113.340 ;
        RECT 1003.580 111.720 1012.120 112.260 ;
        RECT 1006.025 111.515 1012.120 111.720 ;
        RECT 1006.025 108.180 1012.415 111.515 ;
        RECT 1009.205 107.600 1012.415 108.180 ;
        RECT 931.330 105.755 949.350 106.265 ;
        RECT 931.330 104.835 965.060 105.755 ;
      LAYER pwell ;
        RECT 1002.700 105.045 1012.215 107.065 ;
        RECT 965.410 104.740 1012.215 105.045 ;
      LAYER nwell ;
        RECT 1474.330 106.265 1475.760 115.655 ;
        RECT 1550.470 113.340 1555.120 114.420 ;
        RECT 1546.505 112.260 1555.120 113.340 ;
        RECT 1546.580 111.720 1555.120 112.260 ;
        RECT 1549.025 111.515 1555.120 111.720 ;
        RECT 1549.025 108.180 1555.415 111.515 ;
        RECT 1552.205 107.600 1555.415 108.180 ;
        RECT 1474.330 105.755 1492.350 106.265 ;
        RECT 1474.330 104.835 1508.060 105.755 ;
      LAYER pwell ;
        RECT 1545.700 105.045 1555.215 107.065 ;
        RECT 1508.410 104.740 1555.215 105.045 ;
      LAYER nwell ;
        RECT 1748.330 106.265 1749.760 115.655 ;
        RECT 1824.470 113.340 1829.120 114.420 ;
        RECT 1820.505 112.260 1829.120 113.340 ;
        RECT 1820.580 111.720 1829.120 112.260 ;
        RECT 1823.025 111.515 1829.120 111.720 ;
        RECT 1823.025 108.180 1829.415 111.515 ;
        RECT 1826.205 107.600 1829.415 108.180 ;
        RECT 1748.330 105.755 1766.350 106.265 ;
        RECT 1748.330 104.835 1782.060 105.755 ;
      LAYER pwell ;
        RECT 1819.700 105.045 1829.215 107.065 ;
        RECT 1782.410 104.740 1829.215 105.045 ;
      LAYER nwell ;
        RECT 2022.330 106.265 2023.760 115.655 ;
        RECT 2098.470 113.340 2103.120 114.420 ;
        RECT 2094.505 112.260 2103.120 113.340 ;
        RECT 2094.580 111.720 2103.120 112.260 ;
        RECT 2097.025 111.515 2103.120 111.720 ;
        RECT 2097.025 108.180 2103.415 111.515 ;
        RECT 2100.205 107.600 2103.415 108.180 ;
        RECT 2022.330 105.755 2040.350 106.265 ;
        RECT 2022.330 104.835 2056.060 105.755 ;
      LAYER pwell ;
        RECT 2093.700 105.045 2103.215 107.065 ;
        RECT 2056.410 104.740 2103.215 105.045 ;
      LAYER nwell ;
        RECT 2296.330 106.265 2297.760 115.655 ;
        RECT 2372.470 113.340 2377.120 114.420 ;
        RECT 2368.505 112.260 2377.120 113.340 ;
        RECT 2368.580 111.720 2377.120 112.260 ;
        RECT 2371.025 111.515 2377.120 111.720 ;
        RECT 2371.025 108.180 2377.415 111.515 ;
        RECT 2374.205 107.600 2377.415 108.180 ;
        RECT 2296.330 105.755 2314.350 106.265 ;
        RECT 2296.330 104.835 2330.060 105.755 ;
      LAYER pwell ;
        RECT 2367.700 105.045 2377.215 107.065 ;
        RECT 2330.410 104.740 2377.215 105.045 ;
      LAYER nwell ;
        RECT 2570.330 106.265 2571.760 115.655 ;
        RECT 2646.470 113.340 2651.120 114.420 ;
        RECT 2642.505 112.260 2651.120 113.340 ;
        RECT 2642.580 111.720 2651.120 112.260 ;
        RECT 2645.025 111.515 2651.120 111.720 ;
        RECT 2645.025 108.180 2651.415 111.515 ;
        RECT 2648.205 107.600 2651.415 108.180 ;
        RECT 2570.330 105.755 2588.350 106.265 ;
        RECT 2570.330 104.835 2604.060 105.755 ;
      LAYER pwell ;
        RECT 2641.700 105.045 2651.215 107.065 ;
        RECT 2604.410 104.740 2651.215 105.045 ;
        RECT 966.160 104.025 1012.215 104.740 ;
        RECT 1509.160 104.025 1555.215 104.740 ;
        RECT 1783.160 104.025 1829.215 104.740 ;
        RECT 2057.160 104.025 2103.215 104.740 ;
        RECT 2331.160 104.025 2377.215 104.740 ;
        RECT 2605.160 104.025 2651.215 104.740 ;
        RECT 931.710 103.745 1012.215 104.025 ;
        RECT 679.530 103.265 738.130 103.270 ;
        RECT 662.870 102.005 738.130 103.265 ;
        RECT 662.870 100.770 666.070 102.005 ;
        RECT 679.530 100.770 738.130 102.005 ;
        RECT 662.870 97.475 738.130 100.770 ;
        RECT 662.870 75.865 664.440 97.475 ;
        RECT 736.565 75.865 738.130 97.475 ;
        RECT 662.870 70.685 738.130 75.865 ;
        RECT 662.870 69.645 676.090 70.685 ;
        RECT 696.250 69.645 738.130 70.685 ;
        RECT 931.710 102.015 972.615 103.745 ;
        RECT 931.710 100.480 935.230 102.015 ;
        RECT 931.710 99.180 959.120 100.480 ;
        RECT 931.710 98.035 972.615 99.180 ;
        RECT 1006.785 98.035 1012.215 103.745 ;
        RECT 931.710 96.450 1012.215 98.035 ;
        RECT 931.710 74.865 934.135 96.450 ;
        RECT 1006.265 74.865 1012.215 96.450 ;
        RECT 931.710 70.685 1012.215 74.865 ;
        RECT 931.710 69.645 945.090 70.685 ;
        RECT 971.755 69.645 1012.215 70.685 ;
        RECT 1474.710 103.745 1555.215 104.025 ;
        RECT 1474.710 102.015 1515.615 103.745 ;
        RECT 1474.710 100.480 1478.230 102.015 ;
        RECT 1474.710 99.180 1502.120 100.480 ;
        RECT 1474.710 98.035 1515.615 99.180 ;
        RECT 1549.785 98.035 1555.215 103.745 ;
        RECT 1474.710 96.450 1555.215 98.035 ;
        RECT 1474.710 74.865 1477.135 96.450 ;
        RECT 1549.265 74.865 1555.215 96.450 ;
        RECT 1474.710 70.685 1555.215 74.865 ;
        RECT 1474.710 69.645 1488.090 70.685 ;
        RECT 1514.755 69.645 1555.215 70.685 ;
        RECT 1748.710 103.745 1829.215 104.025 ;
        RECT 1748.710 102.015 1789.615 103.745 ;
        RECT 1748.710 100.480 1752.230 102.015 ;
        RECT 1748.710 99.180 1776.120 100.480 ;
        RECT 1748.710 98.035 1789.615 99.180 ;
        RECT 1823.785 98.035 1829.215 103.745 ;
        RECT 1748.710 96.450 1829.215 98.035 ;
        RECT 1748.710 74.865 1751.135 96.450 ;
        RECT 1823.265 74.865 1829.215 96.450 ;
        RECT 1748.710 70.685 1829.215 74.865 ;
        RECT 1748.710 69.645 1762.090 70.685 ;
        RECT 1788.755 69.645 1829.215 70.685 ;
        RECT 2022.710 103.745 2103.215 104.025 ;
        RECT 2022.710 102.015 2063.615 103.745 ;
        RECT 2022.710 100.480 2026.230 102.015 ;
        RECT 2022.710 99.180 2050.120 100.480 ;
        RECT 2022.710 98.035 2063.615 99.180 ;
        RECT 2097.785 98.035 2103.215 103.745 ;
        RECT 2022.710 96.450 2103.215 98.035 ;
        RECT 2022.710 74.865 2025.135 96.450 ;
        RECT 2097.265 74.865 2103.215 96.450 ;
        RECT 2022.710 70.685 2103.215 74.865 ;
        RECT 2022.710 69.645 2036.090 70.685 ;
        RECT 2062.755 69.645 2103.215 70.685 ;
        RECT 2296.710 103.745 2377.215 104.025 ;
        RECT 2296.710 102.015 2337.615 103.745 ;
        RECT 2296.710 100.480 2300.230 102.015 ;
        RECT 2296.710 99.180 2324.120 100.480 ;
        RECT 2296.710 98.035 2337.615 99.180 ;
        RECT 2371.785 98.035 2377.215 103.745 ;
        RECT 2296.710 96.450 2377.215 98.035 ;
        RECT 2296.710 74.865 2299.135 96.450 ;
        RECT 2371.265 74.865 2377.215 96.450 ;
        RECT 2296.710 70.685 2377.215 74.865 ;
        RECT 2296.710 69.645 2310.090 70.685 ;
        RECT 2336.755 69.645 2377.215 70.685 ;
        RECT 2570.710 103.745 2651.215 104.025 ;
        RECT 2570.710 102.015 2611.615 103.745 ;
        RECT 2570.710 100.480 2574.230 102.015 ;
        RECT 2570.710 99.180 2598.120 100.480 ;
        RECT 2570.710 98.035 2611.615 99.180 ;
        RECT 2645.785 98.035 2651.215 103.745 ;
        RECT 2570.710 96.450 2651.215 98.035 ;
        RECT 2570.710 74.865 2573.135 96.450 ;
        RECT 2645.265 74.865 2651.215 96.450 ;
        RECT 2570.710 70.685 2651.215 74.865 ;
        RECT 2570.710 69.645 2584.090 70.685 ;
        RECT 2610.755 69.645 2651.215 70.685 ;
      LAYER nwell ;
        RECT 662.670 59.620 738.330 69.335 ;
        RECT 931.560 59.620 1012.415 69.335 ;
        RECT 1474.560 59.620 1555.415 69.335 ;
        RECT 1748.560 59.620 1829.415 69.335 ;
        RECT 2022.560 59.620 2103.415 69.335 ;
        RECT 2296.560 59.620 2377.415 69.335 ;
        RECT 2570.560 59.620 2651.415 69.335 ;
        RECT 931.560 59.615 965.960 59.620 ;
        RECT 1474.560 59.615 1508.960 59.620 ;
        RECT 1748.560 59.615 1782.960 59.620 ;
        RECT 2022.560 59.615 2056.960 59.620 ;
        RECT 2296.560 59.615 2330.960 59.620 ;
        RECT 2570.560 59.615 2604.960 59.620 ;
      LAYER pwell ;
        RECT 662.710 55.435 738.290 59.315 ;
        RECT 931.710 55.435 1012.290 59.315 ;
        RECT 1474.710 55.435 1555.290 59.315 ;
        RECT 1748.710 55.435 1829.290 59.315 ;
        RECT 2022.710 55.435 2103.290 59.315 ;
        RECT 2296.710 55.435 2377.290 59.315 ;
        RECT 2570.710 55.435 2651.290 59.315 ;
      LAYER nwell ;
        RECT 662.380 53.310 738.515 55.120 ;
        RECT 662.380 31.485 664.905 53.310 ;
        RECT 736.325 31.485 738.515 53.310 ;
        RECT 662.380 29.790 738.515 31.485 ;
        RECT 931.560 53.310 1012.415 55.120 ;
        RECT 931.560 31.485 933.370 53.310 ;
        RECT 1005.615 31.485 1012.415 53.310 ;
        RECT 931.560 29.770 1012.415 31.485 ;
        RECT 1474.560 53.310 1555.415 55.120 ;
        RECT 1474.560 31.485 1476.370 53.310 ;
        RECT 1548.615 31.485 1555.415 53.310 ;
        RECT 1474.560 29.770 1555.415 31.485 ;
        RECT 1748.560 53.310 1829.415 55.120 ;
        RECT 1748.560 31.485 1750.370 53.310 ;
        RECT 1822.615 31.485 1829.415 53.310 ;
        RECT 1748.560 29.770 1829.415 31.485 ;
        RECT 2022.560 53.310 2103.415 55.120 ;
        RECT 2022.560 31.485 2024.370 53.310 ;
        RECT 2096.615 31.485 2103.415 53.310 ;
        RECT 2022.560 29.770 2103.415 31.485 ;
        RECT 2296.560 53.310 2377.415 55.120 ;
        RECT 2296.560 31.485 2298.370 53.310 ;
        RECT 2370.615 31.485 2377.415 53.310 ;
        RECT 2296.560 29.770 2377.415 31.485 ;
        RECT 2570.560 53.310 2651.415 55.120 ;
        RECT 2570.560 31.485 2572.370 53.310 ;
        RECT 2644.615 31.485 2651.415 53.310 ;
        RECT 2570.560 29.770 2651.415 31.485 ;
        RECT 931.565 29.525 1012.415 29.770 ;
        RECT 931.565 26.455 945.030 29.525 ;
        RECT 1004.485 26.455 1012.415 29.525 ;
        RECT 931.565 21.025 1012.415 26.455 ;
        RECT 1474.565 29.525 1555.415 29.770 ;
        RECT 1474.565 26.455 1488.030 29.525 ;
        RECT 1547.485 26.455 1555.415 29.525 ;
        RECT 1474.565 21.025 1555.415 26.455 ;
        RECT 1748.565 29.525 1829.415 29.770 ;
        RECT 1748.565 26.455 1762.030 29.525 ;
        RECT 1821.485 26.455 1829.415 29.525 ;
        RECT 1748.565 21.025 1829.415 26.455 ;
        RECT 2022.565 29.525 2103.415 29.770 ;
        RECT 2022.565 26.455 2036.030 29.525 ;
        RECT 2095.485 26.455 2103.415 29.525 ;
        RECT 2022.565 21.025 2103.415 26.455 ;
        RECT 2296.565 29.525 2377.415 29.770 ;
        RECT 2296.565 26.455 2310.030 29.525 ;
        RECT 2369.485 26.455 2377.415 29.525 ;
        RECT 2296.565 21.025 2377.415 26.455 ;
        RECT 2570.565 29.525 2651.415 29.770 ;
        RECT 2570.565 26.455 2584.030 29.525 ;
        RECT 2643.485 26.455 2651.415 29.525 ;
        RECT 2570.565 21.025 2651.415 26.455 ;
      LAYER li1 ;
        RECT 381.000 5166.645 461.000 5187.705 ;
        RECT 638.000 5166.645 718.000 5187.705 ;
        RECT 895.000 5166.645 975.000 5187.705 ;
        RECT 1152.000 5166.645 1232.000 5187.705 ;
        RECT 1410.000 5166.645 1490.000 5187.705 ;
        RECT 380.915 5158.090 461.105 5166.645 ;
        RECT 637.915 5158.090 718.105 5166.645 ;
        RECT 894.915 5158.090 975.105 5166.645 ;
        RECT 1151.915 5158.090 1232.105 5166.645 ;
        RECT 1409.915 5158.090 1490.105 5166.645 ;
        RECT 380.885 5133.215 461.105 5158.090 ;
        RECT 637.885 5133.215 718.105 5158.090 ;
        RECT 894.885 5133.215 975.105 5158.090 ;
        RECT 1151.885 5133.215 1232.105 5158.090 ;
        RECT 1409.885 5133.215 1490.105 5158.090 ;
        RECT 380.885 5133.155 461.000 5133.215 ;
        RECT 637.885 5133.155 718.000 5133.215 ;
        RECT 894.885 5133.155 975.000 5133.215 ;
        RECT 1151.885 5133.155 1232.000 5133.215 ;
        RECT 1409.885 5133.155 1490.000 5133.215 ;
        RECT 381.000 5132.435 461.000 5133.155 ;
        RECT 638.000 5132.435 718.000 5133.155 ;
        RECT 895.000 5132.435 975.000 5133.155 ;
        RECT 1152.000 5132.435 1232.000 5133.155 ;
        RECT 1410.000 5132.435 1490.000 5133.155 ;
        RECT 380.840 5128.815 461.160 5132.435 ;
        RECT 637.840 5128.815 718.160 5132.435 ;
        RECT 894.840 5128.815 975.160 5132.435 ;
        RECT 1151.840 5128.815 1232.160 5132.435 ;
        RECT 1409.840 5128.815 1490.160 5132.435 ;
        RECT 381.000 5128.150 461.000 5128.815 ;
        RECT 638.000 5128.150 718.000 5128.815 ;
        RECT 895.000 5128.150 975.000 5128.815 ;
        RECT 1152.000 5128.150 1232.000 5128.815 ;
        RECT 1410.000 5128.150 1490.000 5128.815 ;
        RECT 380.885 5128.055 461.000 5128.150 ;
        RECT 637.885 5128.055 718.000 5128.150 ;
        RECT 894.885 5128.055 975.000 5128.150 ;
        RECT 1151.885 5128.055 1232.000 5128.150 ;
        RECT 1409.885 5128.055 1490.000 5128.150 ;
        RECT 380.885 5119.275 461.085 5128.055 ;
        RECT 637.885 5119.275 718.085 5128.055 ;
        RECT 894.885 5119.275 975.085 5128.055 ;
        RECT 1151.885 5119.275 1232.085 5128.055 ;
        RECT 1409.885 5119.275 1490.085 5128.055 ;
        RECT 380.915 5118.995 461.085 5119.275 ;
        RECT 637.915 5118.995 718.085 5119.275 ;
        RECT 894.915 5118.995 975.085 5119.275 ;
        RECT 1151.915 5118.995 1232.085 5119.275 ;
        RECT 1409.915 5118.995 1490.085 5119.275 ;
        RECT 381.000 5118.225 461.000 5118.995 ;
        RECT 638.000 5118.225 718.000 5118.995 ;
        RECT 895.000 5118.225 975.000 5118.995 ;
        RECT 1152.000 5118.225 1232.000 5118.995 ;
        RECT 1410.000 5118.225 1490.000 5118.995 ;
        RECT 380.915 5118.220 461.160 5118.225 ;
        RECT 637.915 5118.220 718.160 5118.225 ;
        RECT 894.915 5118.220 975.160 5118.225 ;
        RECT 1151.915 5118.220 1232.160 5118.225 ;
        RECT 1409.915 5118.220 1490.160 5118.225 ;
        RECT 380.885 5084.105 461.160 5118.220 ;
        RECT 637.885 5084.105 718.160 5118.220 ;
        RECT 894.885 5084.105 975.160 5118.220 ;
        RECT 1151.885 5084.105 1232.160 5118.220 ;
        RECT 1409.885 5084.105 1490.160 5118.220 ;
        RECT 380.885 5083.895 461.000 5084.105 ;
        RECT 637.885 5083.895 718.000 5084.105 ;
        RECT 894.885 5083.895 975.000 5084.105 ;
        RECT 1151.885 5083.895 1232.000 5084.105 ;
        RECT 1409.885 5083.895 1490.000 5084.105 ;
        RECT 380.915 5082.580 461.000 5083.895 ;
        RECT 637.915 5082.580 718.000 5083.895 ;
        RECT 894.915 5082.580 975.000 5083.895 ;
        RECT 1151.915 5082.580 1232.000 5083.895 ;
        RECT 1409.915 5082.580 1490.000 5083.895 ;
        RECT 380.915 5081.065 461.085 5082.580 ;
        RECT 637.915 5081.065 718.085 5082.580 ;
        RECT 894.915 5081.065 975.085 5082.580 ;
        RECT 1151.915 5081.065 1232.085 5082.580 ;
        RECT 1409.915 5081.065 1490.085 5082.580 ;
        RECT 381.000 5080.070 461.085 5081.065 ;
        RECT 638.000 5080.070 718.085 5081.065 ;
        RECT 895.000 5080.070 975.085 5081.065 ;
        RECT 1152.000 5080.070 1232.085 5081.065 ;
        RECT 1410.000 5080.070 1490.085 5081.065 ;
        RECT 380.915 5076.815 461.085 5080.070 ;
        RECT 637.915 5076.815 718.085 5080.070 ;
        RECT 894.915 5076.815 975.085 5080.070 ;
        RECT 1151.915 5076.815 1232.085 5080.070 ;
        RECT 1409.915 5076.815 1490.085 5080.070 ;
        RECT 381.000 5068.605 461.085 5076.815 ;
        RECT 638.000 5068.605 718.085 5076.815 ;
        RECT 895.000 5068.605 975.085 5076.815 ;
        RECT 1152.000 5068.605 1232.085 5076.815 ;
        RECT 1410.000 5068.605 1490.085 5076.815 ;
        RECT 380.915 5045.220 461.085 5068.605 ;
        RECT 637.915 5045.220 718.085 5068.605 ;
        RECT 894.915 5045.220 975.085 5068.605 ;
        RECT 1151.915 5045.220 1232.085 5068.605 ;
        RECT 1409.915 5045.220 1490.085 5068.605 ;
        RECT 381.000 5039.250 461.085 5045.220 ;
        RECT 638.000 5039.250 718.085 5045.220 ;
        RECT 895.000 5039.250 975.085 5045.220 ;
        RECT 1152.000 5039.250 1232.085 5045.220 ;
        RECT 1410.000 5039.250 1490.085 5045.220 ;
        RECT 381.000 5023.725 461.000 5039.250 ;
        RECT 638.000 5023.725 718.000 5039.250 ;
        RECT 895.000 5023.725 975.000 5039.250 ;
        RECT 1152.000 5023.725 1232.000 5039.250 ;
        RECT 1410.000 5023.725 1490.000 5039.250 ;
        RECT 381.000 5018.115 461.120 5023.725 ;
        RECT 638.000 5018.115 718.120 5023.725 ;
        RECT 895.000 5018.115 975.120 5023.725 ;
        RECT 1152.000 5018.115 1232.120 5023.725 ;
        RECT 1410.000 5018.115 1490.120 5023.725 ;
        RECT 381.000 5013.015 461.000 5018.115 ;
        RECT 638.000 5013.015 718.000 5018.115 ;
        RECT 895.000 5013.015 975.000 5018.115 ;
        RECT 1152.000 5013.015 1232.000 5018.115 ;
        RECT 1410.000 5013.015 1490.000 5018.115 ;
        RECT 381.000 5007.485 461.120 5013.015 ;
        RECT 638.000 5007.485 718.120 5013.015 ;
        RECT 895.000 5007.485 975.120 5013.015 ;
        RECT 1152.000 5007.485 1232.120 5013.015 ;
        RECT 1410.000 5007.485 1490.120 5013.015 ;
        RECT 381.000 4996.995 461.000 5007.485 ;
        RECT 638.000 4996.995 718.000 5007.485 ;
        RECT 895.000 4996.995 975.000 5007.485 ;
        RECT 1152.000 4996.995 1232.000 5007.485 ;
        RECT 1410.000 4996.995 1490.000 5007.485 ;
        RECT 380.915 4993.995 461.000 4996.995 ;
        RECT 637.915 4993.995 718.000 4996.995 ;
        RECT 894.915 4993.995 975.000 4996.995 ;
        RECT 1151.915 4993.995 1232.000 4996.995 ;
        RECT 1409.915 4993.995 1490.000 4996.995 ;
        RECT 381.000 4988.230 461.000 4993.995 ;
        RECT 638.000 4988.230 718.000 4993.995 ;
        RECT 895.000 4988.230 975.000 4993.995 ;
        RECT 1152.000 4988.230 1232.000 4993.995 ;
        RECT 1410.000 4988.230 1490.000 4993.995 ;
        RECT 1668.070 4990.035 1739.775 5187.695 ;
        RECT 1919.000 5166.645 1999.000 5187.705 ;
        RECT 2364.000 5166.645 2444.000 5187.705 ;
        RECT 2621.000 5166.645 2701.000 5187.705 ;
        RECT 1918.915 5158.090 1999.105 5166.645 ;
        RECT 2363.915 5158.090 2444.105 5166.645 ;
        RECT 2620.915 5158.090 2701.105 5166.645 ;
        RECT 1918.885 5133.215 1999.105 5158.090 ;
        RECT 2363.885 5133.215 2444.105 5158.090 ;
        RECT 2620.885 5133.215 2701.105 5158.090 ;
        RECT 1918.885 5133.155 1999.000 5133.215 ;
        RECT 2363.885 5133.155 2444.000 5133.215 ;
        RECT 2620.885 5133.155 2701.000 5133.215 ;
        RECT 1919.000 5132.435 1999.000 5133.155 ;
        RECT 2364.000 5132.435 2444.000 5133.155 ;
        RECT 2621.000 5132.435 2701.000 5133.155 ;
        RECT 1918.840 5128.815 1999.160 5132.435 ;
        RECT 2363.840 5128.815 2444.160 5132.435 ;
        RECT 2620.840 5128.815 2701.160 5132.435 ;
        RECT 1919.000 5128.150 1999.000 5128.815 ;
        RECT 2364.000 5128.150 2444.000 5128.815 ;
        RECT 2621.000 5128.150 2701.000 5128.815 ;
        RECT 1918.885 5128.055 1999.000 5128.150 ;
        RECT 2363.885 5128.055 2444.000 5128.150 ;
        RECT 2620.885 5128.055 2701.000 5128.150 ;
        RECT 1918.885 5119.275 1999.085 5128.055 ;
        RECT 2363.885 5119.275 2444.085 5128.055 ;
        RECT 2620.885 5119.275 2701.085 5128.055 ;
        RECT 1918.915 5118.995 1999.085 5119.275 ;
        RECT 2363.915 5118.995 2444.085 5119.275 ;
        RECT 2620.915 5118.995 2701.085 5119.275 ;
        RECT 1919.000 5118.225 1999.000 5118.995 ;
        RECT 2364.000 5118.225 2444.000 5118.995 ;
        RECT 2621.000 5118.225 2701.000 5118.995 ;
        RECT 1918.915 5118.220 1999.160 5118.225 ;
        RECT 2363.915 5118.220 2444.160 5118.225 ;
        RECT 2620.915 5118.220 2701.160 5118.225 ;
        RECT 1918.885 5084.105 1999.160 5118.220 ;
        RECT 2363.885 5084.105 2444.160 5118.220 ;
        RECT 2620.885 5084.105 2701.160 5118.220 ;
        RECT 1918.885 5083.895 1999.000 5084.105 ;
        RECT 2363.885 5083.895 2444.000 5084.105 ;
        RECT 2620.885 5083.895 2701.000 5084.105 ;
        RECT 1918.915 5082.580 1999.000 5083.895 ;
        RECT 2363.915 5082.580 2444.000 5083.895 ;
        RECT 2620.915 5082.580 2701.000 5083.895 ;
        RECT 1918.915 5081.065 1999.085 5082.580 ;
        RECT 2363.915 5081.065 2444.085 5082.580 ;
        RECT 2620.915 5081.065 2701.085 5082.580 ;
        RECT 1919.000 5080.070 1999.085 5081.065 ;
        RECT 2364.000 5080.070 2444.085 5081.065 ;
        RECT 2621.000 5080.070 2701.085 5081.065 ;
        RECT 1918.915 5076.815 1999.085 5080.070 ;
        RECT 2363.915 5076.815 2444.085 5080.070 ;
        RECT 2620.915 5076.815 2701.085 5080.070 ;
        RECT 1919.000 5068.605 1999.085 5076.815 ;
        RECT 2364.000 5068.605 2444.085 5076.815 ;
        RECT 2621.000 5068.605 2701.085 5076.815 ;
        RECT 1918.915 5045.220 1999.085 5068.605 ;
        RECT 2363.915 5045.220 2444.085 5068.605 ;
        RECT 2620.915 5045.220 2701.085 5068.605 ;
        RECT 1919.000 5039.250 1999.085 5045.220 ;
        RECT 2364.000 5039.250 2444.085 5045.220 ;
        RECT 2621.000 5039.250 2701.085 5045.220 ;
        RECT 1919.000 5023.725 1999.000 5039.250 ;
        RECT 2364.000 5023.725 2444.000 5039.250 ;
        RECT 2621.000 5023.725 2701.000 5039.250 ;
        RECT 1919.000 5018.115 1999.120 5023.725 ;
        RECT 2364.000 5018.115 2444.120 5023.725 ;
        RECT 2621.000 5018.115 2701.120 5023.725 ;
        RECT 1919.000 5013.015 1999.000 5018.115 ;
        RECT 2364.000 5013.015 2444.000 5018.115 ;
        RECT 2621.000 5013.015 2701.000 5018.115 ;
        RECT 1919.000 5007.485 1999.120 5013.015 ;
        RECT 2364.000 5007.485 2444.120 5013.015 ;
        RECT 2621.000 5007.485 2701.120 5013.015 ;
        RECT 1919.000 4996.995 1999.000 5007.485 ;
        RECT 2364.000 4996.995 2444.000 5007.485 ;
        RECT 2621.000 4996.995 2701.000 5007.485 ;
        RECT 1918.915 4993.995 1999.000 4996.995 ;
        RECT 2363.915 4993.995 2444.000 4996.995 ;
        RECT 2620.915 4993.995 2701.000 4996.995 ;
        RECT 1679.065 4989.890 1680.045 4990.035 ;
        RECT 1736.760 4989.890 1737.650 4990.035 ;
        RECT 1679.065 4989.000 1737.650 4989.890 ;
        RECT 1919.000 4988.230 1999.000 4993.995 ;
        RECT 2364.000 4988.230 2444.000 4993.995 ;
        RECT 2621.000 4988.230 2701.000 4993.995 ;
        RECT 2879.070 4990.035 2950.775 5187.695 ;
        RECT 3130.000 5166.645 3210.000 5187.705 ;
        RECT 3129.915 5158.090 3210.105 5166.645 ;
        RECT 3129.885 5133.215 3210.105 5158.090 ;
        RECT 3129.885 5133.155 3210.000 5133.215 ;
        RECT 3130.000 5132.435 3210.000 5133.155 ;
        RECT 3129.840 5128.815 3210.160 5132.435 ;
        RECT 3130.000 5128.150 3210.000 5128.815 ;
        RECT 3129.885 5128.055 3210.000 5128.150 ;
        RECT 3129.885 5119.275 3210.085 5128.055 ;
        RECT 3129.915 5118.995 3210.085 5119.275 ;
        RECT 3130.000 5118.225 3210.000 5118.995 ;
        RECT 3129.915 5118.220 3210.160 5118.225 ;
        RECT 3129.885 5084.105 3210.160 5118.220 ;
        RECT 3129.885 5083.895 3210.000 5084.105 ;
        RECT 3129.915 5082.580 3210.000 5083.895 ;
        RECT 3129.915 5081.065 3210.085 5082.580 ;
        RECT 3130.000 5080.070 3210.085 5081.065 ;
        RECT 3129.915 5076.815 3210.085 5080.070 ;
        RECT 3130.000 5068.605 3210.085 5076.815 ;
        RECT 3129.915 5045.220 3210.085 5068.605 ;
        RECT 3130.000 5039.250 3210.085 5045.220 ;
        RECT 3130.000 5023.725 3210.000 5039.250 ;
        RECT 3130.000 5018.115 3210.120 5023.725 ;
        RECT 3130.000 5013.015 3210.000 5018.115 ;
        RECT 3130.000 5007.485 3210.120 5013.015 ;
        RECT 3130.000 4996.995 3210.000 5007.485 ;
        RECT 3129.915 4993.995 3210.000 4996.995 ;
        RECT 2890.065 4989.890 2891.045 4990.035 ;
        RECT 2947.760 4989.890 2948.650 4990.035 ;
        RECT 2890.065 4989.000 2948.650 4989.890 ;
        RECT 3130.000 4988.230 3210.000 4993.995 ;
        RECT 21.355 4851.000 54.785 4851.105 ;
        RECT 55.565 4851.000 59.185 4851.160 ;
        RECT 59.945 4851.000 69.005 4851.085 ;
        RECT 69.775 4851.000 103.895 4851.160 ;
        RECT 105.420 4851.000 148.750 4851.085 ;
        RECT 164.275 4851.000 169.885 4851.120 ;
        RECT 174.985 4851.000 180.515 4851.120 ;
        RECT 0.295 4771.000 199.770 4851.000 ;
        RECT 3483.895 4838.085 3518.220 4838.115 ;
        RECT 3519.275 4838.085 3528.150 4838.115 ;
        RECT 3393.995 4838.000 3396.995 4838.085 ;
        RECT 3445.220 4838.000 3468.605 4838.085 ;
        RECT 3476.815 4838.000 3480.070 4838.085 ;
        RECT 3481.065 4838.000 3518.225 4838.085 ;
        RECT 3518.995 4838.000 3528.150 4838.085 ;
        RECT 3528.815 4838.000 3532.435 4838.160 ;
        RECT 3533.155 4838.085 3558.090 4838.115 ;
        RECT 3533.155 4838.000 3566.645 4838.085 ;
        RECT 21.355 4770.915 54.845 4771.000 ;
        RECT 29.910 4770.885 54.845 4770.915 ;
        RECT 55.565 4770.840 59.185 4771.000 ;
        RECT 59.850 4770.915 69.005 4771.000 ;
        RECT 69.775 4770.915 106.935 4771.000 ;
        RECT 107.930 4770.915 111.185 4771.000 ;
        RECT 119.395 4770.915 142.780 4771.000 ;
        RECT 191.005 4770.915 194.005 4771.000 ;
        RECT 59.850 4770.885 68.725 4770.915 ;
        RECT 69.780 4770.885 104.105 4770.915 ;
        RECT 3388.230 4758.000 3587.705 4838.000 ;
        RECT 3407.485 4757.880 3413.015 4758.000 ;
        RECT 3418.115 4757.880 3423.725 4758.000 ;
        RECT 3439.250 4757.915 3482.580 4758.000 ;
        RECT 3484.105 4757.840 3518.225 4758.000 ;
        RECT 3518.995 4757.915 3528.055 4758.000 ;
        RECT 3528.815 4757.840 3532.435 4758.000 ;
        RECT 3533.215 4757.895 3566.645 4758.000 ;
        RECT 0.220 4560.240 196.980 4634.755 ;
        RECT 3391.020 4538.245 3587.780 4612.760 ;
        RECT 0.305 4419.680 197.965 4421.855 ;
        RECT 0.305 4418.730 199.030 4419.680 ;
        RECT 0.305 4362.045 197.965 4418.730 ;
        RECT 198.080 4362.045 199.030 4418.730 ;
        RECT 3483.895 4392.085 3518.220 4392.115 ;
        RECT 3519.275 4392.085 3528.150 4392.115 ;
        RECT 3393.995 4392.000 3396.995 4392.085 ;
        RECT 3445.220 4392.000 3468.605 4392.085 ;
        RECT 3476.815 4392.000 3480.070 4392.085 ;
        RECT 3481.065 4392.000 3518.225 4392.085 ;
        RECT 3518.995 4392.000 3528.150 4392.085 ;
        RECT 3528.815 4392.000 3532.435 4392.160 ;
        RECT 3533.155 4392.085 3558.090 4392.115 ;
        RECT 3533.155 4392.000 3566.645 4392.085 ;
        RECT 0.305 4361.035 199.030 4362.045 ;
        RECT 0.305 4360.155 197.965 4361.035 ;
        RECT 0.305 4349.610 198.935 4360.155 ;
        RECT 3388.230 4312.000 3587.705 4392.000 ;
        RECT 3407.485 4311.880 3413.015 4312.000 ;
        RECT 3418.115 4311.880 3423.725 4312.000 ;
        RECT 3439.250 4311.915 3482.580 4312.000 ;
        RECT 3484.105 4311.840 3518.225 4312.000 ;
        RECT 3518.995 4311.915 3528.055 4312.000 ;
        RECT 3528.815 4311.840 3532.435 4312.000 ;
        RECT 3533.215 4311.895 3566.645 4312.000 ;
        RECT 0.305 4208.650 197.965 4210.775 ;
        RECT 0.305 4207.760 199.000 4208.650 ;
        RECT 0.305 4151.045 197.965 4207.760 ;
        RECT 198.110 4151.045 199.000 4207.760 ;
        RECT 3389.065 4155.845 3587.695 4166.390 ;
        RECT 3390.035 4154.965 3587.695 4155.845 ;
        RECT 0.305 4150.065 199.000 4151.045 ;
        RECT 3388.970 4153.955 3587.695 4154.965 ;
        RECT 0.305 4139.070 197.965 4150.065 ;
        RECT 3388.970 4097.270 3389.920 4153.955 ;
        RECT 3390.035 4097.270 3587.695 4153.955 ;
        RECT 3388.970 4096.320 3587.695 4097.270 ;
        RECT 3390.035 4094.145 3587.695 4096.320 ;
        RECT 21.355 4002.000 54.785 4002.105 ;
        RECT 55.565 4002.000 59.185 4002.160 ;
        RECT 59.945 4002.000 69.005 4002.085 ;
        RECT 69.775 4002.000 103.895 4002.160 ;
        RECT 105.420 4002.000 148.750 4002.085 ;
        RECT 164.275 4002.000 169.885 4002.120 ;
        RECT 174.985 4002.000 180.515 4002.120 ;
        RECT 0.295 3922.000 199.770 4002.000 ;
        RECT 3483.895 3946.085 3518.220 3946.115 ;
        RECT 3519.275 3946.085 3528.150 3946.115 ;
        RECT 3393.995 3946.000 3396.995 3946.085 ;
        RECT 3445.220 3946.000 3468.605 3946.085 ;
        RECT 3476.815 3946.000 3480.070 3946.085 ;
        RECT 3481.065 3946.000 3518.225 3946.085 ;
        RECT 3518.995 3946.000 3528.150 3946.085 ;
        RECT 3528.815 3946.000 3532.435 3946.160 ;
        RECT 3533.155 3946.085 3558.090 3946.115 ;
        RECT 3533.155 3946.000 3566.645 3946.085 ;
        RECT 21.355 3921.915 54.845 3922.000 ;
        RECT 29.910 3921.885 54.845 3921.915 ;
        RECT 55.565 3921.840 59.185 3922.000 ;
        RECT 59.850 3921.915 69.005 3922.000 ;
        RECT 69.775 3921.915 106.935 3922.000 ;
        RECT 107.930 3921.915 111.185 3922.000 ;
        RECT 119.395 3921.915 142.780 3922.000 ;
        RECT 191.005 3921.915 194.005 3922.000 ;
        RECT 59.850 3921.885 68.725 3921.915 ;
        RECT 69.780 3921.885 104.105 3921.915 ;
        RECT 3388.230 3866.000 3587.705 3946.000 ;
        RECT 3407.485 3865.880 3413.015 3866.000 ;
        RECT 3418.115 3865.880 3423.725 3866.000 ;
        RECT 3439.250 3865.915 3482.580 3866.000 ;
        RECT 3484.105 3865.840 3518.225 3866.000 ;
        RECT 3518.995 3865.915 3528.055 3866.000 ;
        RECT 3528.815 3865.840 3532.435 3866.000 ;
        RECT 3533.215 3865.895 3566.645 3866.000 ;
        RECT 21.355 3786.000 54.785 3786.105 ;
        RECT 55.565 3786.000 59.185 3786.160 ;
        RECT 59.945 3786.000 69.005 3786.085 ;
        RECT 69.775 3786.000 103.895 3786.160 ;
        RECT 105.420 3786.000 148.750 3786.085 ;
        RECT 164.275 3786.000 169.885 3786.120 ;
        RECT 174.985 3786.000 180.515 3786.120 ;
        RECT 0.295 3706.000 199.770 3786.000 ;
        RECT 3483.895 3721.085 3518.220 3721.115 ;
        RECT 3519.275 3721.085 3528.150 3721.115 ;
        RECT 3393.995 3721.000 3396.995 3721.085 ;
        RECT 3445.220 3721.000 3468.605 3721.085 ;
        RECT 3476.815 3721.000 3480.070 3721.085 ;
        RECT 3481.065 3721.000 3518.225 3721.085 ;
        RECT 3518.995 3721.000 3528.150 3721.085 ;
        RECT 3528.815 3721.000 3532.435 3721.160 ;
        RECT 3533.155 3721.085 3558.090 3721.115 ;
        RECT 3533.155 3721.000 3566.645 3721.085 ;
        RECT 21.355 3705.915 54.845 3706.000 ;
        RECT 29.910 3705.885 54.845 3705.915 ;
        RECT 55.565 3705.840 59.185 3706.000 ;
        RECT 59.850 3705.915 69.005 3706.000 ;
        RECT 69.775 3705.915 106.935 3706.000 ;
        RECT 107.930 3705.915 111.185 3706.000 ;
        RECT 119.395 3705.915 142.780 3706.000 ;
        RECT 191.005 3705.915 194.005 3706.000 ;
        RECT 59.850 3705.885 68.725 3705.915 ;
        RECT 69.780 3705.885 104.105 3705.915 ;
        RECT 3388.230 3641.000 3587.705 3721.000 ;
        RECT 3407.485 3640.880 3413.015 3641.000 ;
        RECT 3418.115 3640.880 3423.725 3641.000 ;
        RECT 3439.250 3640.915 3482.580 3641.000 ;
        RECT 3484.105 3640.840 3518.225 3641.000 ;
        RECT 3518.995 3640.915 3528.055 3641.000 ;
        RECT 3528.815 3640.840 3532.435 3641.000 ;
        RECT 3533.215 3640.895 3566.645 3641.000 ;
        RECT 21.355 3570.000 54.785 3570.105 ;
        RECT 55.565 3570.000 59.185 3570.160 ;
        RECT 59.945 3570.000 69.005 3570.085 ;
        RECT 69.775 3570.000 103.895 3570.160 ;
        RECT 105.420 3570.000 148.750 3570.085 ;
        RECT 164.275 3570.000 169.885 3570.120 ;
        RECT 174.985 3570.000 180.515 3570.120 ;
        RECT 0.295 3490.000 199.770 3570.000 ;
        RECT 3483.895 3496.085 3518.220 3496.115 ;
        RECT 3519.275 3496.085 3528.150 3496.115 ;
        RECT 3393.995 3496.000 3396.995 3496.085 ;
        RECT 3445.220 3496.000 3468.605 3496.085 ;
        RECT 3476.815 3496.000 3480.070 3496.085 ;
        RECT 3481.065 3496.000 3518.225 3496.085 ;
        RECT 3518.995 3496.000 3528.150 3496.085 ;
        RECT 3528.815 3496.000 3532.435 3496.160 ;
        RECT 3533.155 3496.085 3558.090 3496.115 ;
        RECT 3533.155 3496.000 3566.645 3496.085 ;
        RECT 21.355 3489.915 54.845 3490.000 ;
        RECT 29.910 3489.885 54.845 3489.915 ;
        RECT 55.565 3489.840 59.185 3490.000 ;
        RECT 59.850 3489.915 69.005 3490.000 ;
        RECT 69.775 3489.915 106.935 3490.000 ;
        RECT 107.930 3489.915 111.185 3490.000 ;
        RECT 119.395 3489.915 142.780 3490.000 ;
        RECT 191.005 3489.915 194.005 3490.000 ;
        RECT 59.850 3489.885 68.725 3489.915 ;
        RECT 69.780 3489.885 104.105 3489.915 ;
        RECT 3388.230 3416.000 3587.705 3496.000 ;
        RECT 3407.485 3415.880 3413.015 3416.000 ;
        RECT 3418.115 3415.880 3423.725 3416.000 ;
        RECT 3439.250 3415.915 3482.580 3416.000 ;
        RECT 3484.105 3415.840 3518.225 3416.000 ;
        RECT 3518.995 3415.915 3528.055 3416.000 ;
        RECT 3528.815 3415.840 3532.435 3416.000 ;
        RECT 3533.215 3415.895 3566.645 3416.000 ;
        RECT 21.355 3354.000 54.785 3354.105 ;
        RECT 55.565 3354.000 59.185 3354.160 ;
        RECT 59.945 3354.000 69.005 3354.085 ;
        RECT 69.775 3354.000 103.895 3354.160 ;
        RECT 105.420 3354.000 148.750 3354.085 ;
        RECT 164.275 3354.000 169.885 3354.120 ;
        RECT 174.985 3354.000 180.515 3354.120 ;
        RECT 0.295 3274.000 199.770 3354.000 ;
        RECT 21.355 3273.915 54.845 3274.000 ;
        RECT 29.910 3273.885 54.845 3273.915 ;
        RECT 55.565 3273.840 59.185 3274.000 ;
        RECT 59.850 3273.915 69.005 3274.000 ;
        RECT 69.775 3273.915 106.935 3274.000 ;
        RECT 107.930 3273.915 111.185 3274.000 ;
        RECT 119.395 3273.915 142.780 3274.000 ;
        RECT 191.005 3273.915 194.005 3274.000 ;
        RECT 59.850 3273.885 68.725 3273.915 ;
        RECT 69.780 3273.885 104.105 3273.915 ;
        RECT 3483.895 3270.085 3518.220 3270.115 ;
        RECT 3519.275 3270.085 3528.150 3270.115 ;
        RECT 3393.995 3270.000 3396.995 3270.085 ;
        RECT 3445.220 3270.000 3468.605 3270.085 ;
        RECT 3476.815 3270.000 3480.070 3270.085 ;
        RECT 3481.065 3270.000 3518.225 3270.085 ;
        RECT 3518.995 3270.000 3528.150 3270.085 ;
        RECT 3528.815 3270.000 3532.435 3270.160 ;
        RECT 3533.155 3270.085 3558.090 3270.115 ;
        RECT 3533.155 3270.000 3566.645 3270.085 ;
        RECT 3388.230 3190.000 3587.705 3270.000 ;
        RECT 3407.485 3189.880 3413.015 3190.000 ;
        RECT 3418.115 3189.880 3423.725 3190.000 ;
        RECT 3439.250 3189.915 3482.580 3190.000 ;
        RECT 3484.105 3189.840 3518.225 3190.000 ;
        RECT 3518.995 3189.915 3528.055 3190.000 ;
        RECT 3528.815 3189.840 3532.435 3190.000 ;
        RECT 3533.215 3189.895 3566.645 3190.000 ;
        RECT 21.355 3138.000 54.785 3138.105 ;
        RECT 55.565 3138.000 59.185 3138.160 ;
        RECT 59.945 3138.000 69.005 3138.085 ;
        RECT 69.775 3138.000 103.895 3138.160 ;
        RECT 105.420 3138.000 148.750 3138.085 ;
        RECT 164.275 3138.000 169.885 3138.120 ;
        RECT 174.985 3138.000 180.515 3138.120 ;
        RECT 0.295 3058.000 199.770 3138.000 ;
        RECT 21.355 3057.915 54.845 3058.000 ;
        RECT 29.910 3057.885 54.845 3057.915 ;
        RECT 55.565 3057.840 59.185 3058.000 ;
        RECT 59.850 3057.915 69.005 3058.000 ;
        RECT 69.775 3057.915 106.935 3058.000 ;
        RECT 107.930 3057.915 111.185 3058.000 ;
        RECT 119.395 3057.915 142.780 3058.000 ;
        RECT 191.005 3057.915 194.005 3058.000 ;
        RECT 59.850 3057.885 68.725 3057.915 ;
        RECT 69.780 3057.885 104.105 3057.915 ;
        RECT 3483.895 3045.085 3518.220 3045.115 ;
        RECT 3519.275 3045.085 3528.150 3045.115 ;
        RECT 3393.995 3045.000 3396.995 3045.085 ;
        RECT 3445.220 3045.000 3468.605 3045.085 ;
        RECT 3476.815 3045.000 3480.070 3045.085 ;
        RECT 3481.065 3045.000 3518.225 3045.085 ;
        RECT 3518.995 3045.000 3528.150 3045.085 ;
        RECT 3528.815 3045.000 3532.435 3045.160 ;
        RECT 3533.155 3045.085 3558.090 3045.115 ;
        RECT 3533.155 3045.000 3566.645 3045.085 ;
        RECT 3388.230 2965.000 3587.705 3045.000 ;
        RECT 3407.485 2964.880 3413.015 2965.000 ;
        RECT 3418.115 2964.880 3423.725 2965.000 ;
        RECT 3439.250 2964.915 3482.580 2965.000 ;
        RECT 3484.105 2964.840 3518.225 2965.000 ;
        RECT 3518.995 2964.915 3528.055 2965.000 ;
        RECT 3528.815 2964.840 3532.435 2965.000 ;
        RECT 3533.215 2964.895 3566.645 2965.000 ;
        RECT 21.355 2922.000 54.785 2922.105 ;
        RECT 55.565 2922.000 59.185 2922.160 ;
        RECT 59.945 2922.000 69.005 2922.085 ;
        RECT 69.775 2922.000 103.895 2922.160 ;
        RECT 105.420 2922.000 148.750 2922.085 ;
        RECT 164.275 2922.000 169.885 2922.120 ;
        RECT 174.985 2922.000 180.515 2922.120 ;
        RECT 0.295 2842.000 199.770 2922.000 ;
        RECT 21.355 2841.915 54.845 2842.000 ;
        RECT 29.910 2841.885 54.845 2841.915 ;
        RECT 55.565 2841.840 59.185 2842.000 ;
        RECT 59.850 2841.915 69.005 2842.000 ;
        RECT 69.775 2841.915 106.935 2842.000 ;
        RECT 107.930 2841.915 111.185 2842.000 ;
        RECT 119.395 2841.915 142.780 2842.000 ;
        RECT 191.005 2841.915 194.005 2842.000 ;
        RECT 59.850 2841.885 68.725 2841.915 ;
        RECT 69.780 2841.885 104.105 2841.915 ;
        RECT 3483.895 2819.085 3518.220 2819.115 ;
        RECT 3519.275 2819.085 3528.150 2819.115 ;
        RECT 3393.995 2819.000 3396.995 2819.085 ;
        RECT 3445.220 2819.000 3468.605 2819.085 ;
        RECT 3476.815 2819.000 3480.070 2819.085 ;
        RECT 3481.065 2819.000 3518.225 2819.085 ;
        RECT 3518.995 2819.000 3528.150 2819.085 ;
        RECT 3528.815 2819.000 3532.435 2819.160 ;
        RECT 3533.155 2819.085 3558.090 2819.115 ;
        RECT 3533.155 2819.000 3566.645 2819.085 ;
        RECT 3388.230 2739.000 3587.705 2819.000 ;
        RECT 3407.485 2738.880 3413.015 2739.000 ;
        RECT 3418.115 2738.880 3423.725 2739.000 ;
        RECT 3439.250 2738.915 3482.580 2739.000 ;
        RECT 3484.105 2738.840 3518.225 2739.000 ;
        RECT 3518.995 2738.915 3528.055 2739.000 ;
        RECT 3528.815 2738.840 3532.435 2739.000 ;
        RECT 3533.215 2738.895 3566.645 2739.000 ;
        RECT 21.355 2706.000 54.785 2706.105 ;
        RECT 55.565 2706.000 59.185 2706.160 ;
        RECT 59.945 2706.000 69.005 2706.085 ;
        RECT 69.775 2706.000 103.895 2706.160 ;
        RECT 105.420 2706.000 148.750 2706.085 ;
        RECT 164.275 2706.000 169.885 2706.120 ;
        RECT 174.985 2706.000 180.515 2706.120 ;
        RECT 0.295 2626.000 199.770 2706.000 ;
        RECT 21.355 2625.915 54.845 2626.000 ;
        RECT 29.910 2625.885 54.845 2625.915 ;
        RECT 55.565 2625.840 59.185 2626.000 ;
        RECT 59.850 2625.915 69.005 2626.000 ;
        RECT 69.775 2625.915 106.935 2626.000 ;
        RECT 107.930 2625.915 111.185 2626.000 ;
        RECT 119.395 2625.915 142.780 2626.000 ;
        RECT 191.005 2625.915 194.005 2626.000 ;
        RECT 59.850 2625.885 68.725 2625.915 ;
        RECT 69.780 2625.885 104.105 2625.915 ;
        RECT 3389.065 2582.845 3587.695 2593.390 ;
        RECT 3390.035 2581.965 3587.695 2582.845 ;
        RECT 3388.970 2580.955 3587.695 2581.965 ;
        RECT 3388.970 2524.270 3389.920 2580.955 ;
        RECT 3390.035 2524.270 3587.695 2580.955 ;
        RECT 3388.970 2523.320 3587.695 2524.270 ;
        RECT 3390.035 2521.145 3587.695 2523.320 ;
        RECT 0.305 2485.680 197.965 2487.855 ;
        RECT 0.305 2484.730 199.030 2485.680 ;
        RECT 0.305 2428.045 197.965 2484.730 ;
        RECT 198.080 2428.045 199.030 2484.730 ;
        RECT 0.305 2427.035 199.030 2428.045 ;
        RECT 0.305 2426.155 197.965 2427.035 ;
        RECT 0.305 2415.610 198.935 2426.155 ;
        RECT 3391.020 2299.245 3587.780 2373.760 ;
        RECT 0.220 2204.240 196.980 2278.755 ;
        RECT 3390.035 2140.935 3587.695 2151.930 ;
        RECT 3389.000 2139.955 3587.695 2140.935 ;
        RECT 3389.000 2083.240 3389.890 2139.955 ;
        RECT 3390.035 2083.240 3587.695 2139.955 ;
        RECT 3389.000 2082.350 3587.695 2083.240 ;
        RECT 3390.035 2080.225 3587.695 2082.350 ;
        RECT 21.355 2068.000 54.785 2068.105 ;
        RECT 55.565 2068.000 59.185 2068.160 ;
        RECT 59.945 2068.000 69.005 2068.085 ;
        RECT 69.775 2068.000 103.895 2068.160 ;
        RECT 105.420 2068.000 148.750 2068.085 ;
        RECT 164.275 2068.000 169.885 2068.120 ;
        RECT 174.985 2068.000 180.515 2068.120 ;
        RECT 0.295 1988.000 199.770 2068.000 ;
        RECT 21.355 1987.915 54.845 1988.000 ;
        RECT 29.910 1987.885 54.845 1987.915 ;
        RECT 55.565 1987.840 59.185 1988.000 ;
        RECT 59.850 1987.915 69.005 1988.000 ;
        RECT 69.775 1987.915 106.935 1988.000 ;
        RECT 107.930 1987.915 111.185 1988.000 ;
        RECT 119.395 1987.915 142.780 1988.000 ;
        RECT 191.005 1987.915 194.005 1988.000 ;
        RECT 59.850 1987.885 68.725 1987.915 ;
        RECT 69.780 1987.885 104.105 1987.915 ;
        RECT 3483.895 1933.085 3518.220 1933.115 ;
        RECT 3519.275 1933.085 3528.150 1933.115 ;
        RECT 3393.995 1933.000 3396.995 1933.085 ;
        RECT 3445.220 1933.000 3468.605 1933.085 ;
        RECT 3476.815 1933.000 3480.070 1933.085 ;
        RECT 3481.065 1933.000 3518.225 1933.085 ;
        RECT 3518.995 1933.000 3528.150 1933.085 ;
        RECT 3528.815 1933.000 3532.435 1933.160 ;
        RECT 3533.155 1933.085 3558.090 1933.115 ;
        RECT 3533.155 1933.000 3566.645 1933.085 ;
        RECT 3388.230 1853.000 3587.705 1933.000 ;
        RECT 3407.485 1852.880 3413.015 1853.000 ;
        RECT 3418.115 1852.880 3423.725 1853.000 ;
        RECT 3439.250 1852.915 3482.580 1853.000 ;
        RECT 3484.105 1852.840 3518.225 1853.000 ;
        RECT 3518.995 1852.915 3528.055 1853.000 ;
        RECT 3528.815 1852.840 3532.435 1853.000 ;
        RECT 3533.215 1852.895 3566.645 1853.000 ;
        RECT 21.355 1852.000 54.785 1852.105 ;
        RECT 55.565 1852.000 59.185 1852.160 ;
        RECT 59.945 1852.000 69.005 1852.085 ;
        RECT 69.775 1852.000 103.895 1852.160 ;
        RECT 105.420 1852.000 148.750 1852.085 ;
        RECT 164.275 1852.000 169.885 1852.120 ;
        RECT 174.985 1852.000 180.515 1852.120 ;
        RECT 0.295 1772.000 199.770 1852.000 ;
        RECT 21.355 1771.915 54.845 1772.000 ;
        RECT 29.910 1771.885 54.845 1771.915 ;
        RECT 55.565 1771.840 59.185 1772.000 ;
        RECT 59.850 1771.915 69.005 1772.000 ;
        RECT 69.775 1771.915 106.935 1772.000 ;
        RECT 107.930 1771.915 111.185 1772.000 ;
        RECT 119.395 1771.915 142.780 1772.000 ;
        RECT 191.005 1771.915 194.005 1772.000 ;
        RECT 59.850 1771.885 68.725 1771.915 ;
        RECT 69.780 1771.885 104.105 1771.915 ;
        RECT 3483.895 1707.085 3518.220 1707.115 ;
        RECT 3519.275 1707.085 3528.150 1707.115 ;
        RECT 3393.995 1707.000 3396.995 1707.085 ;
        RECT 3445.220 1707.000 3468.605 1707.085 ;
        RECT 3476.815 1707.000 3480.070 1707.085 ;
        RECT 3481.065 1707.000 3518.225 1707.085 ;
        RECT 3518.995 1707.000 3528.150 1707.085 ;
        RECT 3528.815 1707.000 3532.435 1707.160 ;
        RECT 3533.155 1707.085 3558.090 1707.115 ;
        RECT 3533.155 1707.000 3566.645 1707.085 ;
        RECT 21.355 1636.000 54.785 1636.105 ;
        RECT 55.565 1636.000 59.185 1636.160 ;
        RECT 59.945 1636.000 69.005 1636.085 ;
        RECT 69.775 1636.000 103.895 1636.160 ;
        RECT 105.420 1636.000 148.750 1636.085 ;
        RECT 164.275 1636.000 169.885 1636.120 ;
        RECT 174.985 1636.000 180.515 1636.120 ;
        RECT 0.295 1556.000 199.770 1636.000 ;
        RECT 3388.230 1627.000 3587.705 1707.000 ;
        RECT 3407.485 1626.880 3413.015 1627.000 ;
        RECT 3418.115 1626.880 3423.725 1627.000 ;
        RECT 3439.250 1626.915 3482.580 1627.000 ;
        RECT 3484.105 1626.840 3518.225 1627.000 ;
        RECT 3518.995 1626.915 3528.055 1627.000 ;
        RECT 3528.815 1626.840 3532.435 1627.000 ;
        RECT 3533.215 1626.895 3566.645 1627.000 ;
        RECT 21.355 1555.915 54.845 1556.000 ;
        RECT 29.910 1555.885 54.845 1555.915 ;
        RECT 55.565 1555.840 59.185 1556.000 ;
        RECT 59.850 1555.915 69.005 1556.000 ;
        RECT 69.775 1555.915 106.935 1556.000 ;
        RECT 107.930 1555.915 111.185 1556.000 ;
        RECT 119.395 1555.915 142.780 1556.000 ;
        RECT 191.005 1555.915 194.005 1556.000 ;
        RECT 59.850 1555.885 68.725 1555.915 ;
        RECT 69.780 1555.885 104.105 1555.915 ;
        RECT 3483.895 1482.085 3518.220 1482.115 ;
        RECT 3519.275 1482.085 3528.150 1482.115 ;
        RECT 3393.995 1482.000 3396.995 1482.085 ;
        RECT 3445.220 1482.000 3468.605 1482.085 ;
        RECT 3476.815 1482.000 3480.070 1482.085 ;
        RECT 3481.065 1482.000 3518.225 1482.085 ;
        RECT 3518.995 1482.000 3528.150 1482.085 ;
        RECT 3528.815 1482.000 3532.435 1482.160 ;
        RECT 3533.155 1482.085 3558.090 1482.115 ;
        RECT 3533.155 1482.000 3566.645 1482.085 ;
        RECT 21.355 1420.000 54.785 1420.105 ;
        RECT 55.565 1420.000 59.185 1420.160 ;
        RECT 59.945 1420.000 69.005 1420.085 ;
        RECT 69.775 1420.000 103.895 1420.160 ;
        RECT 105.420 1420.000 148.750 1420.085 ;
        RECT 164.275 1420.000 169.885 1420.120 ;
        RECT 174.985 1420.000 180.515 1420.120 ;
        RECT 0.295 1340.000 199.770 1420.000 ;
        RECT 3388.230 1402.000 3587.705 1482.000 ;
        RECT 3407.485 1401.880 3413.015 1402.000 ;
        RECT 3418.115 1401.880 3423.725 1402.000 ;
        RECT 3439.250 1401.915 3482.580 1402.000 ;
        RECT 3484.105 1401.840 3518.225 1402.000 ;
        RECT 3518.995 1401.915 3528.055 1402.000 ;
        RECT 3528.815 1401.840 3532.435 1402.000 ;
        RECT 3533.215 1401.895 3566.645 1402.000 ;
        RECT 21.355 1339.915 54.845 1340.000 ;
        RECT 29.910 1339.885 54.845 1339.915 ;
        RECT 55.565 1339.840 59.185 1340.000 ;
        RECT 59.850 1339.915 69.005 1340.000 ;
        RECT 69.775 1339.915 106.935 1340.000 ;
        RECT 107.930 1339.915 111.185 1340.000 ;
        RECT 119.395 1339.915 142.780 1340.000 ;
        RECT 191.005 1339.915 194.005 1340.000 ;
        RECT 59.850 1339.885 68.725 1339.915 ;
        RECT 69.780 1339.885 104.105 1339.915 ;
        RECT 3483.895 1257.085 3518.220 1257.115 ;
        RECT 3519.275 1257.085 3528.150 1257.115 ;
        RECT 3393.995 1257.000 3396.995 1257.085 ;
        RECT 3445.220 1257.000 3468.605 1257.085 ;
        RECT 3476.815 1257.000 3480.070 1257.085 ;
        RECT 3481.065 1257.000 3518.225 1257.085 ;
        RECT 3518.995 1257.000 3528.150 1257.085 ;
        RECT 3528.815 1257.000 3532.435 1257.160 ;
        RECT 3533.155 1257.085 3558.090 1257.115 ;
        RECT 3533.155 1257.000 3566.645 1257.085 ;
        RECT 21.355 1204.000 54.785 1204.105 ;
        RECT 55.565 1204.000 59.185 1204.160 ;
        RECT 59.945 1204.000 69.005 1204.085 ;
        RECT 69.775 1204.000 103.895 1204.160 ;
        RECT 105.420 1204.000 148.750 1204.085 ;
        RECT 164.275 1204.000 169.885 1204.120 ;
        RECT 174.985 1204.000 180.515 1204.120 ;
        RECT 0.295 1124.000 199.770 1204.000 ;
        RECT 3388.230 1177.000 3587.705 1257.000 ;
        RECT 3407.485 1176.880 3413.015 1177.000 ;
        RECT 3418.115 1176.880 3423.725 1177.000 ;
        RECT 3439.250 1176.915 3482.580 1177.000 ;
        RECT 3484.105 1176.840 3518.225 1177.000 ;
        RECT 3518.995 1176.915 3528.055 1177.000 ;
        RECT 3528.815 1176.840 3532.435 1177.000 ;
        RECT 3533.215 1176.895 3566.645 1177.000 ;
        RECT 21.355 1123.915 54.845 1124.000 ;
        RECT 29.910 1123.885 54.845 1123.915 ;
        RECT 55.565 1123.840 59.185 1124.000 ;
        RECT 59.850 1123.915 69.005 1124.000 ;
        RECT 69.775 1123.915 106.935 1124.000 ;
        RECT 107.930 1123.915 111.185 1124.000 ;
        RECT 119.395 1123.915 142.780 1124.000 ;
        RECT 191.005 1123.915 194.005 1124.000 ;
        RECT 59.850 1123.885 68.725 1123.915 ;
        RECT 69.780 1123.885 104.105 1123.915 ;
        RECT 3483.895 1031.085 3518.220 1031.115 ;
        RECT 3519.275 1031.085 3528.150 1031.115 ;
        RECT 3393.995 1031.000 3396.995 1031.085 ;
        RECT 3445.220 1031.000 3468.605 1031.085 ;
        RECT 3476.815 1031.000 3480.070 1031.085 ;
        RECT 3481.065 1031.000 3518.225 1031.085 ;
        RECT 3518.995 1031.000 3528.150 1031.085 ;
        RECT 3528.815 1031.000 3532.435 1031.160 ;
        RECT 3533.155 1031.085 3558.090 1031.115 ;
        RECT 3533.155 1031.000 3566.645 1031.085 ;
        RECT 21.355 988.000 54.785 988.105 ;
        RECT 55.565 988.000 59.185 988.160 ;
        RECT 59.945 988.000 69.005 988.085 ;
        RECT 69.775 988.000 103.895 988.160 ;
        RECT 105.420 988.000 148.750 988.085 ;
        RECT 164.275 988.000 169.885 988.120 ;
        RECT 174.985 988.000 180.515 988.120 ;
        RECT 0.295 908.000 199.770 988.000 ;
        RECT 3388.230 951.000 3587.705 1031.000 ;
        RECT 3407.485 950.880 3413.015 951.000 ;
        RECT 3418.115 950.880 3423.725 951.000 ;
        RECT 3439.250 950.915 3482.580 951.000 ;
        RECT 3484.105 950.840 3518.225 951.000 ;
        RECT 3518.995 950.915 3528.055 951.000 ;
        RECT 3528.815 950.840 3532.435 951.000 ;
        RECT 3533.215 950.895 3566.645 951.000 ;
        RECT 21.355 907.915 54.845 908.000 ;
        RECT 29.910 907.885 54.845 907.915 ;
        RECT 55.565 907.840 59.185 908.000 ;
        RECT 59.850 907.915 69.005 908.000 ;
        RECT 69.775 907.915 106.935 908.000 ;
        RECT 107.930 907.915 111.185 908.000 ;
        RECT 119.395 907.915 142.780 908.000 ;
        RECT 191.005 907.915 194.005 908.000 ;
        RECT 59.850 907.885 68.725 907.915 ;
        RECT 69.780 907.885 104.105 907.915 ;
        RECT 3483.895 806.085 3518.220 806.115 ;
        RECT 3519.275 806.085 3528.150 806.115 ;
        RECT 3393.995 806.000 3396.995 806.085 ;
        RECT 3445.220 806.000 3468.605 806.085 ;
        RECT 3476.815 806.000 3480.070 806.085 ;
        RECT 3481.065 806.000 3518.225 806.085 ;
        RECT 3518.995 806.000 3528.150 806.085 ;
        RECT 3528.815 806.000 3532.435 806.160 ;
        RECT 3533.155 806.085 3558.090 806.115 ;
        RECT 3533.155 806.000 3566.645 806.085 ;
        RECT 3388.230 726.000 3587.705 806.000 ;
        RECT 3407.485 725.880 3413.015 726.000 ;
        RECT 3418.115 725.880 3423.725 726.000 ;
        RECT 3439.250 725.915 3482.580 726.000 ;
        RECT 3484.105 725.840 3518.225 726.000 ;
        RECT 3518.995 725.915 3528.055 726.000 ;
        RECT 3528.815 725.840 3532.435 726.000 ;
        RECT 3533.215 725.895 3566.645 726.000 ;
        RECT 0.305 621.680 197.965 623.855 ;
        RECT 0.305 620.730 199.030 621.680 ;
        RECT 0.305 564.045 197.965 620.730 ;
        RECT 198.080 564.045 199.030 620.730 ;
        RECT 3483.895 580.085 3518.220 580.115 ;
        RECT 3519.275 580.085 3528.150 580.115 ;
        RECT 3393.995 580.000 3396.995 580.085 ;
        RECT 3445.220 580.000 3468.605 580.085 ;
        RECT 3476.815 580.000 3480.070 580.085 ;
        RECT 3481.065 580.000 3518.225 580.085 ;
        RECT 3518.995 580.000 3528.150 580.085 ;
        RECT 3528.815 580.000 3532.435 580.160 ;
        RECT 3533.155 580.085 3558.090 580.115 ;
        RECT 3533.155 580.000 3566.645 580.085 ;
        RECT 0.305 563.035 199.030 564.045 ;
        RECT 0.305 562.155 197.965 563.035 ;
        RECT 0.305 551.610 198.935 562.155 ;
        RECT 3388.230 500.000 3587.705 580.000 ;
        RECT 3407.485 499.880 3413.015 500.000 ;
        RECT 3418.115 499.880 3423.725 500.000 ;
        RECT 3439.250 499.915 3482.580 500.000 ;
        RECT 3484.105 499.840 3518.225 500.000 ;
        RECT 3518.995 499.915 3528.055 500.000 ;
        RECT 3528.815 499.840 3532.435 500.000 ;
        RECT 3533.215 499.895 3566.645 500.000 ;
        RECT 0.220 340.240 196.980 414.755 ;
        RECT 398.350 198.110 456.935 199.000 ;
        RECT 398.350 197.965 399.240 198.110 ;
        RECT 455.955 197.965 456.935 198.110 ;
        RECT 396.225 0.305 467.930 197.965 ;
        RECT 663.000 98.605 738.000 199.815 ;
        RECT 932.000 194.005 1012.000 199.770 ;
        RECT 932.000 191.005 1012.085 194.005 ;
        RECT 932.000 180.515 1012.000 191.005 ;
        RECT 931.880 174.985 1012.000 180.515 ;
        RECT 932.000 169.885 1012.000 174.985 ;
        RECT 931.880 164.275 1012.000 169.885 ;
        RECT 932.000 148.750 1012.000 164.275 ;
        RECT 931.915 142.780 1012.000 148.750 ;
        RECT 931.915 119.395 1012.085 142.780 ;
        RECT 931.915 111.185 1012.000 119.395 ;
        RECT 931.915 107.930 1012.085 111.185 ;
        RECT 931.915 106.935 1012.000 107.930 ;
        RECT 931.915 105.420 1012.085 106.935 ;
        RECT 932.000 104.105 1012.085 105.420 ;
        RECT 932.000 103.895 1012.115 104.105 ;
        RECT 663.000 69.775 738.265 98.605 ;
        RECT 931.840 69.780 1012.115 103.895 ;
        RECT 931.840 69.775 1012.085 69.780 ;
        RECT 663.000 59.185 738.000 69.775 ;
        RECT 932.000 69.005 1012.000 69.775 ;
        RECT 931.915 68.725 1012.085 69.005 ;
        RECT 931.915 59.945 1012.115 68.725 ;
        RECT 932.000 59.850 1012.115 59.945 ;
        RECT 932.000 59.185 1012.000 59.850 ;
        RECT 662.840 55.565 738.160 59.185 ;
        RECT 931.840 55.565 1012.160 59.185 ;
        RECT 663.000 0.780 738.000 55.565 ;
        RECT 932.000 54.845 1012.000 55.565 ;
        RECT 932.000 54.785 1012.115 54.845 ;
        RECT 931.895 29.910 1012.115 54.785 ;
        RECT 931.895 21.355 1012.085 29.910 ;
        RECT 932.000 0.295 1012.000 21.355 ;
        RECT 1206.245 0.220 1280.760 196.980 ;
        RECT 1475.000 194.005 1555.000 199.770 ;
        RECT 1749.000 194.005 1829.000 199.770 ;
        RECT 2023.000 194.005 2103.000 199.770 ;
        RECT 2297.000 194.005 2377.000 199.770 ;
        RECT 2571.000 194.005 2651.000 199.770 ;
        RECT 2849.350 198.110 2907.935 199.000 ;
        RECT 2849.350 197.965 2850.240 198.110 ;
        RECT 2906.955 197.965 2907.935 198.110 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.270 198.080 ;
        RECT 3175.955 197.965 3176.965 198.080 ;
        RECT 3177.845 197.965 3188.390 198.935 ;
        RECT 1475.000 191.005 1555.085 194.005 ;
        RECT 1749.000 191.005 1829.085 194.005 ;
        RECT 2023.000 191.005 2103.085 194.005 ;
        RECT 2297.000 191.005 2377.085 194.005 ;
        RECT 2571.000 191.005 2651.085 194.005 ;
        RECT 1475.000 180.515 1555.000 191.005 ;
        RECT 1749.000 180.515 1829.000 191.005 ;
        RECT 2023.000 180.515 2103.000 191.005 ;
        RECT 2297.000 180.515 2377.000 191.005 ;
        RECT 2571.000 180.515 2651.000 191.005 ;
        RECT 1474.880 174.985 1555.000 180.515 ;
        RECT 1748.880 174.985 1829.000 180.515 ;
        RECT 2022.880 174.985 2103.000 180.515 ;
        RECT 2296.880 174.985 2377.000 180.515 ;
        RECT 2570.880 174.985 2651.000 180.515 ;
        RECT 1475.000 169.885 1555.000 174.985 ;
        RECT 1749.000 169.885 1829.000 174.985 ;
        RECT 2023.000 169.885 2103.000 174.985 ;
        RECT 2297.000 169.885 2377.000 174.985 ;
        RECT 2571.000 169.885 2651.000 174.985 ;
        RECT 1474.880 164.275 1555.000 169.885 ;
        RECT 1748.880 164.275 1829.000 169.885 ;
        RECT 2022.880 164.275 2103.000 169.885 ;
        RECT 2296.880 164.275 2377.000 169.885 ;
        RECT 2570.880 164.275 2651.000 169.885 ;
        RECT 1475.000 148.750 1555.000 164.275 ;
        RECT 1749.000 148.750 1829.000 164.275 ;
        RECT 2023.000 148.750 2103.000 164.275 ;
        RECT 2297.000 148.750 2377.000 164.275 ;
        RECT 2571.000 148.750 2651.000 164.275 ;
        RECT 1474.915 142.780 1555.000 148.750 ;
        RECT 1748.915 142.780 1829.000 148.750 ;
        RECT 2022.915 142.780 2103.000 148.750 ;
        RECT 2296.915 142.780 2377.000 148.750 ;
        RECT 2570.915 142.780 2651.000 148.750 ;
        RECT 1474.915 119.395 1555.085 142.780 ;
        RECT 1748.915 119.395 1829.085 142.780 ;
        RECT 2022.915 119.395 2103.085 142.780 ;
        RECT 2296.915 119.395 2377.085 142.780 ;
        RECT 2570.915 119.395 2651.085 142.780 ;
        RECT 1474.915 111.185 1555.000 119.395 ;
        RECT 1748.915 111.185 1829.000 119.395 ;
        RECT 2022.915 111.185 2103.000 119.395 ;
        RECT 2296.915 111.185 2377.000 119.395 ;
        RECT 2570.915 111.185 2651.000 119.395 ;
        RECT 1474.915 107.930 1555.085 111.185 ;
        RECT 1748.915 107.930 1829.085 111.185 ;
        RECT 2022.915 107.930 2103.085 111.185 ;
        RECT 2296.915 107.930 2377.085 111.185 ;
        RECT 2570.915 107.930 2651.085 111.185 ;
        RECT 1474.915 106.935 1555.000 107.930 ;
        RECT 1748.915 106.935 1829.000 107.930 ;
        RECT 2022.915 106.935 2103.000 107.930 ;
        RECT 2296.915 106.935 2377.000 107.930 ;
        RECT 2570.915 106.935 2651.000 107.930 ;
        RECT 1474.915 105.420 1555.085 106.935 ;
        RECT 1748.915 105.420 1829.085 106.935 ;
        RECT 2022.915 105.420 2103.085 106.935 ;
        RECT 2296.915 105.420 2377.085 106.935 ;
        RECT 2570.915 105.420 2651.085 106.935 ;
        RECT 1475.000 104.105 1555.085 105.420 ;
        RECT 1749.000 104.105 1829.085 105.420 ;
        RECT 2023.000 104.105 2103.085 105.420 ;
        RECT 2297.000 104.105 2377.085 105.420 ;
        RECT 2571.000 104.105 2651.085 105.420 ;
        RECT 1475.000 103.895 1555.115 104.105 ;
        RECT 1749.000 103.895 1829.115 104.105 ;
        RECT 2023.000 103.895 2103.115 104.105 ;
        RECT 2297.000 103.895 2377.115 104.105 ;
        RECT 2571.000 103.895 2651.115 104.105 ;
        RECT 1474.840 69.780 1555.115 103.895 ;
        RECT 1748.840 69.780 1829.115 103.895 ;
        RECT 2022.840 69.780 2103.115 103.895 ;
        RECT 2296.840 69.780 2377.115 103.895 ;
        RECT 2570.840 69.780 2651.115 103.895 ;
        RECT 1474.840 69.775 1555.085 69.780 ;
        RECT 1748.840 69.775 1829.085 69.780 ;
        RECT 2022.840 69.775 2103.085 69.780 ;
        RECT 2296.840 69.775 2377.085 69.780 ;
        RECT 2570.840 69.775 2651.085 69.780 ;
        RECT 1475.000 69.005 1555.000 69.775 ;
        RECT 1749.000 69.005 1829.000 69.775 ;
        RECT 2023.000 69.005 2103.000 69.775 ;
        RECT 2297.000 69.005 2377.000 69.775 ;
        RECT 2571.000 69.005 2651.000 69.775 ;
        RECT 1474.915 68.725 1555.085 69.005 ;
        RECT 1748.915 68.725 1829.085 69.005 ;
        RECT 2022.915 68.725 2103.085 69.005 ;
        RECT 2296.915 68.725 2377.085 69.005 ;
        RECT 2570.915 68.725 2651.085 69.005 ;
        RECT 1474.915 59.945 1555.115 68.725 ;
        RECT 1748.915 59.945 1829.115 68.725 ;
        RECT 2022.915 59.945 2103.115 68.725 ;
        RECT 2296.915 59.945 2377.115 68.725 ;
        RECT 2570.915 59.945 2651.115 68.725 ;
        RECT 1475.000 59.850 1555.115 59.945 ;
        RECT 1749.000 59.850 1829.115 59.945 ;
        RECT 2023.000 59.850 2103.115 59.945 ;
        RECT 2297.000 59.850 2377.115 59.945 ;
        RECT 2571.000 59.850 2651.115 59.945 ;
        RECT 1475.000 59.185 1555.000 59.850 ;
        RECT 1749.000 59.185 1829.000 59.850 ;
        RECT 2023.000 59.185 2103.000 59.850 ;
        RECT 2297.000 59.185 2377.000 59.850 ;
        RECT 2571.000 59.185 2651.000 59.850 ;
        RECT 1474.840 55.565 1555.160 59.185 ;
        RECT 1748.840 55.565 1829.160 59.185 ;
        RECT 2022.840 55.565 2103.160 59.185 ;
        RECT 2296.840 55.565 2377.160 59.185 ;
        RECT 2570.840 55.565 2651.160 59.185 ;
        RECT 1475.000 54.845 1555.000 55.565 ;
        RECT 1749.000 54.845 1829.000 55.565 ;
        RECT 2023.000 54.845 2103.000 55.565 ;
        RECT 2297.000 54.845 2377.000 55.565 ;
        RECT 2571.000 54.845 2651.000 55.565 ;
        RECT 1475.000 54.785 1555.115 54.845 ;
        RECT 1749.000 54.785 1829.115 54.845 ;
        RECT 2023.000 54.785 2103.115 54.845 ;
        RECT 2297.000 54.785 2377.115 54.845 ;
        RECT 2571.000 54.785 2651.115 54.845 ;
        RECT 1474.895 29.910 1555.115 54.785 ;
        RECT 1748.895 29.910 1829.115 54.785 ;
        RECT 2022.895 29.910 2103.115 54.785 ;
        RECT 2296.895 29.910 2377.115 54.785 ;
        RECT 2570.895 29.910 2651.115 54.785 ;
        RECT 1474.895 21.355 1555.085 29.910 ;
        RECT 1748.895 21.355 1829.085 29.910 ;
        RECT 2022.895 21.355 2103.085 29.910 ;
        RECT 2296.895 21.355 2377.085 29.910 ;
        RECT 2570.895 21.355 2651.085 29.910 ;
        RECT 1475.000 0.295 1555.000 21.355 ;
        RECT 1749.000 0.295 1829.000 21.355 ;
        RECT 2023.000 0.295 2103.000 21.355 ;
        RECT 2297.000 0.295 2377.000 21.355 ;
        RECT 2571.000 0.295 2651.000 21.355 ;
        RECT 2847.225 0.305 2918.930 197.965 ;
        RECT 3116.145 0.305 3188.390 197.965 ;
      LAYER met1 ;
        RECT 381.000 5168.975 461.000 5188.000 ;
        RECT 638.000 5168.975 718.000 5188.000 ;
        RECT 895.000 5168.975 975.000 5188.000 ;
        RECT 1152.000 5168.975 1232.000 5188.000 ;
        RECT 1410.000 5168.975 1490.000 5188.000 ;
        RECT 381.000 5166.900 461.020 5168.975 ;
        RECT 638.000 5166.900 718.020 5168.975 ;
        RECT 895.000 5166.900 975.020 5168.975 ;
        RECT 1152.000 5166.900 1232.020 5168.975 ;
        RECT 1410.000 5166.900 1490.020 5168.975 ;
        RECT 381.000 5158.090 461.000 5166.900 ;
        RECT 638.000 5158.090 718.000 5166.900 ;
        RECT 895.000 5158.090 975.000 5166.900 ;
        RECT 1152.000 5158.090 1232.000 5166.900 ;
        RECT 1410.000 5158.090 1490.000 5166.900 ;
        RECT 380.885 5119.275 461.145 5158.090 ;
        RECT 637.885 5119.275 718.145 5158.090 ;
        RECT 894.885 5119.275 975.145 5158.090 ;
        RECT 1151.885 5119.275 1232.145 5158.090 ;
        RECT 1409.885 5119.275 1490.145 5158.090 ;
        RECT 381.000 5118.220 461.000 5119.275 ;
        RECT 638.000 5118.220 718.000 5119.275 ;
        RECT 895.000 5118.220 975.000 5119.275 ;
        RECT 1152.000 5118.220 1232.000 5119.275 ;
        RECT 1410.000 5118.220 1490.000 5119.275 ;
        RECT 380.885 5083.895 461.145 5118.220 ;
        RECT 637.885 5083.895 718.145 5118.220 ;
        RECT 894.885 5083.895 975.145 5118.220 ;
        RECT 1151.885 5083.895 1232.145 5118.220 ;
        RECT 1409.885 5083.895 1490.145 5118.220 ;
        RECT 381.000 5082.580 461.000 5083.895 ;
        RECT 638.000 5082.580 718.000 5083.895 ;
        RECT 895.000 5082.580 975.000 5083.895 ;
        RECT 1152.000 5082.580 1232.000 5083.895 ;
        RECT 1410.000 5082.580 1490.000 5083.895 ;
        RECT 381.000 5079.480 461.060 5082.580 ;
        RECT 638.000 5079.480 718.060 5082.580 ;
        RECT 895.000 5079.480 975.060 5082.580 ;
        RECT 1152.000 5079.480 1232.060 5082.580 ;
        RECT 1410.000 5079.480 1490.060 5082.580 ;
        RECT 380.855 5077.750 461.060 5079.480 ;
        RECT 637.855 5077.750 718.060 5079.480 ;
        RECT 894.855 5077.750 975.060 5079.480 ;
        RECT 1151.855 5077.750 1232.060 5079.480 ;
        RECT 1409.855 5077.750 1490.060 5079.480 ;
        RECT 381.000 5068.635 461.060 5077.750 ;
        RECT 638.000 5068.635 718.060 5077.750 ;
        RECT 895.000 5068.635 975.060 5077.750 ;
        RECT 1152.000 5068.635 1232.060 5077.750 ;
        RECT 1410.000 5068.635 1490.060 5077.750 ;
        RECT 380.885 5060.930 461.060 5068.635 ;
        POLYGON 461.060 5060.985 461.115 5060.930 461.060 5060.930 ;
        RECT 380.885 5045.190 461.115 5060.930 ;
        RECT 637.885 5060.930 718.060 5068.635 ;
        POLYGON 718.060 5060.985 718.115 5060.930 718.060 5060.930 ;
        RECT 637.885 5045.190 718.115 5060.930 ;
        RECT 894.885 5060.930 975.060 5068.635 ;
        POLYGON 975.060 5060.985 975.115 5060.930 975.060 5060.930 ;
        RECT 894.885 5045.190 975.115 5060.930 ;
        RECT 1151.885 5060.930 1232.060 5068.635 ;
        POLYGON 1232.060 5060.985 1232.115 5060.930 1232.060 5060.930 ;
        RECT 1151.885 5045.190 1232.115 5060.930 ;
        RECT 1409.885 5060.930 1490.060 5068.635 ;
        POLYGON 1490.060 5060.985 1490.115 5060.930 1490.060 5060.930 ;
        RECT 1409.885 5045.190 1490.115 5060.930 ;
        RECT 381.000 5039.220 461.115 5045.190 ;
        RECT 638.000 5039.220 718.115 5045.190 ;
        RECT 895.000 5039.220 975.115 5045.190 ;
        RECT 1152.000 5039.220 1232.115 5045.190 ;
        RECT 1410.000 5039.220 1490.115 5045.190 ;
        RECT 381.000 5023.725 461.000 5039.220 ;
        RECT 638.000 5023.725 718.000 5039.220 ;
        RECT 895.000 5023.725 975.000 5039.220 ;
        RECT 1152.000 5023.725 1232.000 5039.220 ;
        RECT 1410.000 5023.725 1490.000 5039.220 ;
        RECT 381.000 5018.120 461.115 5023.725 ;
        RECT 638.000 5018.120 718.115 5023.725 ;
        RECT 895.000 5018.120 975.115 5023.725 ;
        RECT 1152.000 5018.120 1232.115 5023.725 ;
        RECT 1410.000 5018.120 1490.115 5023.725 ;
        RECT 381.000 5013.015 461.000 5018.120 ;
        RECT 638.000 5013.015 718.000 5018.120 ;
        RECT 895.000 5013.015 975.000 5018.120 ;
        RECT 1152.000 5013.015 1232.000 5018.120 ;
        RECT 1410.000 5013.015 1490.000 5018.120 ;
        RECT 381.000 5007.485 461.115 5013.015 ;
        RECT 638.000 5007.485 718.115 5013.015 ;
        RECT 895.000 5007.485 975.115 5013.015 ;
        RECT 1152.000 5007.485 1232.115 5013.015 ;
        RECT 1410.000 5007.485 1490.115 5013.015 ;
        RECT 381.000 4981.155 461.000 5007.485 ;
        RECT 638.000 4981.155 718.000 5007.485 ;
        RECT 895.000 4981.155 975.000 5007.485 ;
        RECT 1152.000 4981.155 1232.000 5007.485 ;
        RECT 1410.000 4981.155 1490.000 5007.485 ;
        RECT 1667.185 4990.035 1740.620 5187.725 ;
        RECT 1919.000 5168.975 1999.000 5188.000 ;
        RECT 2364.000 5168.975 2444.000 5188.000 ;
        RECT 2621.000 5168.975 2701.000 5188.000 ;
        RECT 1919.000 5166.900 1999.020 5168.975 ;
        RECT 2364.000 5166.900 2444.020 5168.975 ;
        RECT 2621.000 5166.900 2701.020 5168.975 ;
        RECT 1919.000 5158.090 1999.000 5166.900 ;
        RECT 2364.000 5158.090 2444.000 5166.900 ;
        RECT 2621.000 5158.090 2701.000 5166.900 ;
        RECT 1918.885 5119.275 1999.145 5158.090 ;
        RECT 2363.885 5119.275 2444.145 5158.090 ;
        RECT 2620.885 5119.275 2701.145 5158.090 ;
        RECT 1919.000 5118.220 1999.000 5119.275 ;
        RECT 2364.000 5118.220 2444.000 5119.275 ;
        RECT 2621.000 5118.220 2701.000 5119.275 ;
        RECT 1918.885 5083.895 1999.145 5118.220 ;
        RECT 2363.885 5083.895 2444.145 5118.220 ;
        RECT 2620.885 5083.895 2701.145 5118.220 ;
        RECT 1919.000 5082.580 1999.000 5083.895 ;
        RECT 2364.000 5082.580 2444.000 5083.895 ;
        RECT 2621.000 5082.580 2701.000 5083.895 ;
        RECT 1919.000 5079.480 1999.060 5082.580 ;
        RECT 2364.000 5079.480 2444.060 5082.580 ;
        RECT 2621.000 5079.480 2701.060 5082.580 ;
        RECT 1918.855 5077.750 1999.060 5079.480 ;
        RECT 2363.855 5077.750 2444.060 5079.480 ;
        RECT 2620.855 5077.750 2701.060 5079.480 ;
        RECT 1919.000 5068.635 1999.060 5077.750 ;
        RECT 2364.000 5068.635 2444.060 5077.750 ;
        RECT 2621.000 5068.635 2701.060 5077.750 ;
        RECT 1918.885 5060.930 1999.060 5068.635 ;
        POLYGON 1999.060 5060.985 1999.115 5060.930 1999.060 5060.930 ;
        RECT 1918.885 5045.190 1999.115 5060.930 ;
        RECT 2363.885 5060.930 2444.060 5068.635 ;
        POLYGON 2444.060 5060.985 2444.115 5060.930 2444.060 5060.930 ;
        RECT 2363.885 5045.190 2444.115 5060.930 ;
        RECT 2620.885 5060.930 2701.060 5068.635 ;
        POLYGON 2701.060 5060.985 2701.115 5060.930 2701.060 5060.930 ;
        RECT 2620.885 5045.190 2701.115 5060.930 ;
        RECT 1919.000 5039.220 1999.115 5045.190 ;
        RECT 2364.000 5039.220 2444.115 5045.190 ;
        RECT 2621.000 5039.220 2701.115 5045.190 ;
        RECT 1919.000 5023.725 1999.000 5039.220 ;
        RECT 2364.000 5023.725 2444.000 5039.220 ;
        RECT 2621.000 5023.725 2701.000 5039.220 ;
        RECT 1919.000 5018.120 1999.115 5023.725 ;
        RECT 2364.000 5018.120 2444.115 5023.725 ;
        RECT 2621.000 5018.120 2701.115 5023.725 ;
        RECT 1919.000 5013.015 1999.000 5018.120 ;
        RECT 2364.000 5013.015 2444.000 5018.120 ;
        RECT 2621.000 5013.015 2701.000 5018.120 ;
        RECT 1919.000 5007.485 1999.115 5013.015 ;
        RECT 2364.000 5007.485 2444.115 5013.015 ;
        RECT 2621.000 5007.485 2701.115 5013.015 ;
        RECT 1679.035 4989.920 1680.350 4990.035 ;
        POLYGON 1680.350 4990.035 1680.465 4989.920 1680.350 4989.920 ;
        POLYGON 1736.540 4990.035 1736.540 4989.920 1736.425 4989.920 ;
        RECT 1736.540 4989.920 1737.680 4990.035 ;
        RECT 1679.035 4988.970 1737.680 4989.920 ;
        RECT 1919.000 4981.155 1999.000 5007.485 ;
        RECT 2364.000 4981.155 2444.000 5007.485 ;
        RECT 2621.000 4981.155 2701.000 5007.485 ;
        RECT 2878.185 4990.035 2951.620 5187.725 ;
        RECT 3130.000 5168.975 3210.000 5188.000 ;
        RECT 3130.000 5166.900 3210.020 5168.975 ;
        RECT 3130.000 5158.090 3210.000 5166.900 ;
        RECT 3129.885 5119.275 3210.145 5158.090 ;
        RECT 3130.000 5118.220 3210.000 5119.275 ;
        RECT 3129.885 5083.895 3210.145 5118.220 ;
        RECT 3130.000 5082.580 3210.000 5083.895 ;
        RECT 3130.000 5079.480 3210.060 5082.580 ;
        RECT 3129.855 5077.750 3210.060 5079.480 ;
        RECT 3130.000 5068.635 3210.060 5077.750 ;
        RECT 3129.885 5060.930 3210.060 5068.635 ;
        POLYGON 3210.060 5060.985 3210.115 5060.930 3210.060 5060.930 ;
        RECT 3129.885 5045.190 3210.115 5060.930 ;
        RECT 3130.000 5039.220 3210.115 5045.190 ;
        RECT 3130.000 5023.725 3210.000 5039.220 ;
        RECT 3130.000 5018.120 3210.115 5023.725 ;
        RECT 3130.000 5013.015 3210.000 5018.120 ;
        RECT 3130.000 5007.485 3210.115 5013.015 ;
        RECT 2890.035 4989.920 2891.350 4990.035 ;
        POLYGON 2891.350 4990.035 2891.465 4989.920 2891.350 4989.920 ;
        POLYGON 2947.540 4990.035 2947.540 4989.920 2947.425 4989.920 ;
        RECT 2947.540 4989.920 2948.680 4990.035 ;
        RECT 2890.035 4988.970 2948.680 4989.920 ;
        RECT 3130.000 4981.155 3210.000 5007.485 ;
      LAYER met1 ;
        RECT 2690.610 4976.480 2690.930 4976.540 ;
        RECT 2699.350 4976.480 2699.670 4976.540 ;
        RECT 2690.610 4976.340 2699.670 4976.480 ;
        RECT 2690.610 4976.280 2690.930 4976.340 ;
        RECT 2699.350 4976.280 2699.670 4976.340 ;
        RECT 710.310 4975.120 710.630 4975.180 ;
        RECT 716.290 4975.120 716.610 4975.180 ;
        RECT 710.310 4974.980 716.610 4975.120 ;
        RECT 710.310 4974.920 710.630 4974.980 ;
        RECT 716.290 4974.920 716.610 4974.980 ;
        RECT 1953.780 4968.180 1954.840 4968.320 ;
        RECT 416.370 4967.980 416.690 4968.040 ;
        RECT 669.830 4967.980 670.150 4968.040 ;
        RECT 675.810 4967.980 676.130 4968.040 ;
        RECT 416.370 4967.840 676.130 4967.980 ;
        RECT 416.370 4967.780 416.690 4967.840 ;
        RECT 669.830 4967.780 670.150 4967.840 ;
        RECT 675.810 4967.780 676.130 4967.840 ;
        RECT 676.270 4967.980 676.590 4968.040 ;
        RECT 710.310 4967.980 710.630 4968.040 ;
        RECT 676.270 4967.840 710.630 4967.980 ;
        RECT 676.270 4967.780 676.590 4967.840 ;
        RECT 710.310 4967.780 710.630 4967.840 ;
        RECT 933.410 4967.980 933.730 4968.040 ;
        RECT 973.430 4967.980 973.750 4968.040 ;
        RECT 933.410 4967.840 973.750 4967.980 ;
        RECT 933.410 4967.780 933.730 4967.840 ;
        RECT 973.430 4967.780 973.750 4967.840 ;
        RECT 1168.470 4967.980 1168.790 4968.040 ;
        RECT 1187.330 4967.980 1187.650 4968.040 ;
        RECT 1441.710 4967.980 1442.030 4968.040 ;
        RECT 1168.470 4967.840 1187.650 4967.980 ;
        RECT 1168.470 4967.780 1168.790 4967.840 ;
        RECT 1187.330 4967.780 1187.650 4967.840 ;
        RECT 1193.630 4967.840 1442.030 4967.980 ;
        RECT 397.510 4967.640 397.830 4967.700 ;
        RECT 654.650 4967.640 654.970 4967.700 ;
        RECT 911.790 4967.640 912.110 4967.700 ;
        RECT 917.310 4967.640 917.630 4967.700 ;
        RECT 397.510 4967.500 917.630 4967.640 ;
        RECT 397.510 4967.440 397.830 4967.500 ;
        RECT 654.650 4967.440 654.970 4967.500 ;
        RECT 911.790 4967.440 912.110 4967.500 ;
        RECT 917.310 4967.440 917.630 4967.500 ;
        RECT 926.970 4967.640 927.290 4967.700 ;
        RECT 1183.650 4967.640 1183.970 4967.700 ;
        RECT 1193.630 4967.640 1193.770 4967.840 ;
        RECT 1441.710 4967.780 1442.030 4967.840 ;
        RECT 1448.150 4967.980 1448.470 4968.040 ;
        RECT 1488.170 4967.980 1488.490 4968.040 ;
        RECT 1448.150 4967.840 1488.490 4967.980 ;
        RECT 1448.150 4967.780 1448.470 4967.840 ;
        RECT 1488.170 4967.780 1488.490 4967.840 ;
        RECT 1478.970 4967.640 1479.290 4967.700 ;
        RECT 1953.780 4967.640 1953.920 4968.180 ;
        RECT 1954.700 4967.980 1954.840 4968.180 ;
        RECT 1957.370 4967.980 1957.690 4968.040 ;
        RECT 1997.390 4967.980 1997.710 4968.040 ;
        RECT 1954.700 4967.840 1955.300 4967.980 ;
        RECT 926.970 4967.500 1193.770 4967.640 ;
        RECT 1241.930 4967.500 1953.920 4967.640 ;
        RECT 1955.160 4967.640 1955.300 4967.840 ;
        RECT 1957.370 4967.840 1997.710 4967.980 ;
        RECT 1957.370 4967.780 1957.690 4967.840 ;
        RECT 1997.390 4967.780 1997.710 4967.840 ;
        RECT 2402.190 4967.980 2402.510 4968.040 ;
        RECT 2442.210 4967.980 2442.530 4968.040 ;
        RECT 2402.190 4967.840 2442.530 4967.980 ;
        RECT 2402.190 4967.780 2402.510 4967.840 ;
        RECT 2442.210 4967.780 2442.530 4967.840 ;
        RECT 2659.330 4967.980 2659.650 4968.040 ;
        RECT 2690.610 4967.980 2690.930 4968.040 ;
        RECT 2659.330 4967.840 2690.930 4967.980 ;
        RECT 2659.330 4967.780 2659.650 4967.840 ;
        RECT 2690.610 4967.780 2690.930 4967.840 ;
        RECT 3168.090 4967.980 3168.410 4968.040 ;
        RECT 3208.110 4967.980 3208.430 4968.040 ;
        RECT 3168.090 4967.840 3208.430 4967.980 ;
        RECT 3168.090 4967.780 3168.410 4967.840 ;
        RECT 3208.110 4967.780 3208.430 4967.840 ;
        RECT 1988.190 4967.640 1988.510 4967.700 ;
        RECT 2433.010 4967.640 2433.330 4967.700 ;
        RECT 2690.150 4967.640 2690.470 4967.700 ;
        RECT 3198.910 4967.640 3199.230 4967.700 ;
        RECT 1955.160 4967.500 3199.230 4967.640 ;
        RECT 926.970 4967.440 927.290 4967.500 ;
        RECT 1183.650 4967.440 1183.970 4967.500 ;
        RECT 449.950 4967.300 450.270 4967.360 ;
        RECT 707.090 4967.300 707.410 4967.360 ;
        RECT 964.230 4967.300 964.550 4967.360 ;
        RECT 1220.910 4967.300 1221.230 4967.360 ;
        RECT 1241.930 4967.300 1242.070 4967.500 ;
        RECT 1478.970 4967.440 1479.290 4967.500 ;
        RECT 1988.190 4967.440 1988.510 4967.500 ;
        RECT 2433.010 4967.440 2433.330 4967.500 ;
        RECT 2690.150 4967.440 2690.470 4967.500 ;
        RECT 3198.910 4967.440 3199.230 4967.500 ;
        RECT 2380.570 4967.300 2380.890 4967.360 ;
        RECT 2637.710 4967.300 2638.030 4967.360 ;
        RECT 2641.390 4967.300 2641.710 4967.360 ;
        RECT 449.950 4967.160 1242.070 4967.300 ;
        RECT 1954.240 4967.160 2641.710 4967.300 ;
        RECT 449.950 4967.100 450.270 4967.160 ;
        RECT 707.090 4967.100 707.410 4967.160 ;
        RECT 964.230 4967.100 964.550 4967.160 ;
        RECT 1220.910 4967.100 1221.230 4967.160 ;
        RECT 1187.330 4966.960 1187.650 4967.020 ;
        RECT 1426.530 4966.960 1426.850 4967.020 ;
        RECT 1666.190 4966.960 1666.510 4967.020 ;
        RECT 1935.750 4966.960 1936.070 4967.020 ;
        RECT 1954.240 4966.960 1954.380 4967.160 ;
        RECT 2380.570 4967.100 2380.890 4967.160 ;
        RECT 2637.710 4967.100 2638.030 4967.160 ;
        RECT 2641.390 4967.100 2641.710 4967.160 ;
        RECT 2656.110 4967.300 2656.430 4967.360 ;
        RECT 3161.650 4967.300 3161.970 4967.360 ;
        RECT 2656.110 4967.160 3161.970 4967.300 ;
        RECT 2656.110 4967.100 2656.430 4967.160 ;
        RECT 3161.650 4967.100 3161.970 4967.160 ;
        RECT 1187.330 4966.820 1954.380 4966.960 ;
        RECT 1187.330 4966.760 1187.650 4966.820 ;
        RECT 1426.530 4966.760 1426.850 4966.820 ;
        RECT 1666.190 4966.760 1666.510 4966.820 ;
        RECT 1935.750 4966.760 1936.070 4966.820 ;
        RECT 419.130 4966.620 419.450 4966.680 ;
        RECT 459.150 4966.620 459.470 4966.680 ;
        RECT 419.130 4966.480 459.470 4966.620 ;
        RECT 419.130 4966.420 419.450 4966.480 ;
        RECT 459.150 4966.420 459.470 4966.480 ;
        RECT 917.310 4966.620 917.630 4966.680 ;
        RECT 1168.470 4966.620 1168.790 4966.680 ;
        RECT 1950.930 4966.620 1951.250 4966.680 ;
        RECT 2395.750 4966.620 2396.070 4966.680 ;
        RECT 2641.390 4966.620 2641.710 4966.680 ;
        RECT 3146.470 4966.620 3146.790 4966.680 ;
        RECT 917.310 4966.480 1168.790 4966.620 ;
        RECT 917.310 4966.420 917.630 4966.480 ;
        RECT 1168.470 4966.420 1168.790 4966.480 ;
        RECT 1483.430 4966.480 2401.270 4966.620 ;
        RECT 675.810 4966.280 676.130 4966.340 ;
        RECT 926.970 4966.280 927.290 4966.340 ;
        RECT 675.810 4966.140 927.290 4966.280 ;
        RECT 675.810 4966.080 676.130 4966.140 ;
        RECT 926.970 4966.080 927.290 4966.140 ;
        RECT 1190.090 4966.280 1190.410 4966.340 ;
        RECT 1230.110 4966.280 1230.430 4966.340 ;
        RECT 1190.090 4966.140 1230.430 4966.280 ;
        RECT 1190.090 4966.080 1190.410 4966.140 ;
        RECT 1230.110 4966.080 1230.430 4966.140 ;
        RECT 1441.710 4966.280 1442.030 4966.340 ;
        RECT 1483.430 4966.280 1483.570 4966.480 ;
        RECT 1950.930 4966.420 1951.250 4966.480 ;
        RECT 2395.750 4966.420 2396.070 4966.480 ;
        RECT 1441.710 4966.140 1483.570 4966.280 ;
        RECT 2401.130 4966.280 2401.270 4966.480 ;
        RECT 2641.390 4966.480 3146.790 4966.620 ;
        RECT 2641.390 4966.420 2641.710 4966.480 ;
        RECT 3146.470 4966.420 3146.790 4966.480 ;
        RECT 2652.890 4966.280 2653.210 4966.340 ;
        RECT 2656.110 4966.280 2656.430 4966.340 ;
        RECT 2401.130 4966.140 2656.430 4966.280 ;
        RECT 1441.710 4966.080 1442.030 4966.140 ;
        RECT 2652.890 4966.080 2653.210 4966.140 ;
        RECT 2656.110 4966.080 2656.430 4966.140 ;
        RECT 3198.910 4965.600 3199.230 4965.660 ;
        RECT 3370.950 4965.600 3371.270 4965.660 ;
        RECT 3198.910 4965.460 3371.270 4965.600 ;
        RECT 3198.910 4965.400 3199.230 4965.460 ;
        RECT 3370.950 4965.400 3371.270 4965.460 ;
        RECT 217.190 4965.260 217.510 4965.320 ;
        RECT 397.510 4965.260 397.830 4965.320 ;
        RECT 217.190 4965.120 397.830 4965.260 ;
        RECT 217.190 4965.060 217.510 4965.120 ;
        RECT 397.510 4965.060 397.830 4965.120 ;
        RECT 3161.650 4965.260 3161.970 4965.320 ;
        RECT 3371.410 4965.260 3371.730 4965.320 ;
        RECT 3161.650 4965.120 3371.730 4965.260 ;
        RECT 3161.650 4965.060 3161.970 4965.120 ;
        RECT 3371.410 4965.060 3371.730 4965.120 ;
        RECT 217.650 4964.920 217.970 4964.980 ;
        RECT 412.690 4964.920 413.010 4964.980 ;
        RECT 416.370 4964.920 416.690 4964.980 ;
        RECT 217.650 4964.780 416.690 4964.920 ;
        RECT 217.650 4964.720 217.970 4964.780 ;
        RECT 412.690 4964.720 413.010 4964.780 ;
        RECT 416.370 4964.720 416.690 4964.780 ;
        RECT 211.670 4964.580 211.990 4964.640 ;
        RECT 449.950 4964.580 450.270 4964.640 ;
        RECT 211.670 4964.440 450.270 4964.580 ;
        RECT 211.670 4964.380 211.990 4964.440 ;
        RECT 449.950 4964.380 450.270 4964.440 ;
        RECT 3146.470 4964.580 3146.790 4964.640 ;
        RECT 3375.550 4964.580 3375.870 4964.640 ;
        RECT 3146.470 4964.440 3375.870 4964.580 ;
        RECT 3146.470 4964.380 3146.790 4964.440 ;
        RECT 3375.550 4964.380 3375.870 4964.440 ;
        RECT 2902.670 4950.640 2902.990 4950.700 ;
        RECT 3370.490 4950.640 3370.810 4950.700 ;
        RECT 2902.670 4950.500 3370.810 4950.640 ;
        RECT 2902.670 4950.440 2902.990 4950.500 ;
        RECT 3370.490 4950.440 3370.810 4950.500 ;
      LAYER met1 ;
        RECT 19.025 4851.000 21.100 4851.020 ;
        RECT 29.910 4851.000 68.725 4851.145 ;
        RECT 69.780 4851.000 104.105 4851.145 ;
        POLYGON 127.070 4851.115 127.070 4851.060 127.015 4851.060 ;
        RECT 127.070 4851.060 148.780 4851.115 ;
        RECT 105.420 4851.000 148.780 4851.060 ;
        RECT 164.275 4851.000 169.880 4851.115 ;
        RECT 174.985 4851.000 180.515 4851.115 ;
        RECT 0.000 4771.000 206.845 4851.000 ;
      LAYER met1 ;
        RECT 208.910 4839.800 209.230 4839.860 ;
        RECT 212.130 4839.800 212.450 4839.860 ;
        RECT 208.910 4839.660 212.450 4839.800 ;
        RECT 208.910 4839.600 209.230 4839.660 ;
        RECT 212.130 4839.600 212.450 4839.660 ;
      LAYER met1 ;
        RECT 3445.190 4838.000 3468.635 4838.115 ;
        RECT 3477.750 4838.000 3479.480 4838.145 ;
        RECT 3483.895 4838.000 3518.220 4838.115 ;
        RECT 3519.275 4838.000 3558.090 4838.115 ;
      LAYER met1 ;
        RECT 3371.410 4820.760 3371.730 4820.820 ;
        RECT 3376.470 4820.760 3376.790 4820.820 ;
        RECT 3371.410 4820.620 3376.790 4820.760 ;
        RECT 3371.410 4820.560 3371.730 4820.620 ;
        RECT 3376.470 4820.560 3376.790 4820.620 ;
        RECT 3374.630 4803.420 3374.950 4803.480 ;
        RECT 3376.930 4803.420 3377.250 4803.480 ;
        RECT 3374.630 4803.280 3377.250 4803.420 ;
        RECT 3374.630 4803.220 3374.950 4803.280 ;
        RECT 3376.930 4803.220 3377.250 4803.280 ;
        RECT 3376.010 4800.840 3376.330 4801.100 ;
        RECT 3376.100 4800.080 3376.240 4800.840 ;
        RECT 3376.010 4799.820 3376.330 4800.080 ;
        RECT 211.210 4795.260 211.530 4795.320 ;
        RECT 213.050 4795.260 213.370 4795.320 ;
        RECT 217.650 4795.260 217.970 4795.320 ;
        RECT 211.210 4795.120 217.970 4795.260 ;
        RECT 211.210 4795.060 211.530 4795.120 ;
        RECT 213.050 4795.060 213.370 4795.120 ;
        RECT 217.650 4795.060 217.970 4795.120 ;
        RECT 208.910 4788.460 209.230 4788.520 ;
        RECT 217.190 4788.460 217.510 4788.520 ;
        RECT 208.910 4788.320 217.510 4788.460 ;
        RECT 208.910 4788.260 209.230 4788.320 ;
        RECT 217.190 4788.260 217.510 4788.320 ;
        RECT 212.130 4787.240 212.450 4787.500 ;
        RECT 212.220 4786.480 212.360 4787.240 ;
        RECT 212.130 4786.220 212.450 4786.480 ;
      LAYER met1 ;
        RECT 29.910 4770.885 68.725 4771.000 ;
        RECT 69.780 4770.885 104.105 4771.000 ;
        RECT 108.520 4770.855 110.250 4771.000 ;
        RECT 119.365 4770.885 142.810 4771.000 ;
      LAYER met1 ;
        RECT 3370.950 4766.700 3371.270 4766.760 ;
        RECT 3375.550 4766.700 3375.870 4766.760 ;
        RECT 3377.850 4766.700 3378.170 4766.760 ;
        RECT 3370.950 4766.560 3378.170 4766.700 ;
        RECT 3370.950 4766.500 3371.270 4766.560 ;
        RECT 3375.550 4766.500 3375.870 4766.560 ;
        RECT 3377.850 4766.500 3378.170 4766.560 ;
      LAYER met1 ;
        RECT 3381.155 4758.000 3588.000 4838.000 ;
        RECT 3407.485 4757.885 3413.015 4758.000 ;
        RECT 3418.120 4757.885 3423.725 4758.000 ;
        RECT 3439.220 4757.940 3482.580 4758.000 ;
        RECT 3439.220 4757.885 3460.930 4757.940 ;
        POLYGON 3460.930 4757.940 3460.985 4757.940 3460.930 4757.885 ;
        RECT 3483.895 4757.855 3518.220 4758.000 ;
        RECT 3519.275 4757.855 3558.090 4758.000 ;
        RECT 3566.900 4757.980 3568.975 4758.000 ;
        RECT 122.615 4641.935 204.885 4645.935 ;
        POLYGON 204.885 4645.935 208.885 4641.935 204.885 4641.935 ;
        RECT 122.615 4636.200 208.885 4641.935 ;
        RECT 0.160 4616.565 197.965 4635.000 ;
        RECT 198.780 4616.565 208.885 4636.200 ;
        RECT 0.160 4580.925 208.885 4616.565 ;
        RECT 3390.035 4596.345 3587.840 4612.880 ;
        RECT 3390.000 4592.075 3587.840 4596.345 ;
        RECT 0.160 4576.655 198.000 4580.925 ;
        RECT 0.160 4560.120 197.965 4576.655 ;
        RECT 3379.115 4556.435 3587.840 4592.075 ;
        RECT 3379.115 4536.800 3389.220 4556.435 ;
        RECT 3390.035 4538.000 3587.840 4556.435 ;
        RECT 3379.115 4531.065 3465.385 4536.800 ;
        POLYGON 3379.115 4531.065 3383.115 4531.065 3383.115 4527.065 ;
        RECT 3383.115 4527.065 3465.385 4531.065 ;
        RECT 0.275 4419.680 197.965 4421.915 ;
        RECT 0.275 4418.540 199.030 4419.680 ;
        RECT 0.275 4362.350 197.965 4418.540 ;
        POLYGON 197.965 4418.540 198.080 4418.540 198.080 4418.425 ;
        POLYGON 198.080 4362.465 198.080 4362.350 197.965 4362.350 ;
        RECT 198.080 4362.350 199.030 4418.540 ;
        RECT 3445.190 4392.000 3468.635 4392.115 ;
        RECT 3477.750 4392.000 3479.480 4392.145 ;
        RECT 3483.895 4392.000 3518.220 4392.115 ;
        RECT 3519.275 4392.000 3558.090 4392.115 ;
      LAYER met1 ;
        RECT 3374.170 4372.640 3374.490 4372.700 ;
        RECT 3376.010 4372.640 3376.330 4372.700 ;
        RECT 3376.930 4372.640 3377.250 4372.700 ;
        RECT 3374.170 4372.500 3377.250 4372.640 ;
        RECT 3374.170 4372.440 3374.490 4372.500 ;
        RECT 3376.010 4372.440 3376.330 4372.500 ;
        RECT 3376.930 4372.440 3377.250 4372.500 ;
      LAYER met1 ;
        RECT 0.275 4361.035 199.030 4362.350 ;
        RECT 0.275 4357.855 197.965 4361.035 ;
      LAYER met1 ;
        RECT 3375.090 4358.360 3375.410 4358.420 ;
        RECT 3376.930 4358.360 3377.250 4358.420 ;
        RECT 3375.090 4358.220 3377.250 4358.360 ;
        RECT 3375.090 4358.160 3375.410 4358.220 ;
        RECT 3376.930 4358.160 3377.250 4358.220 ;
      LAYER met1 ;
        RECT 0.275 4352.625 198.870 4357.855 ;
        RECT 0.275 4349.185 197.965 4352.625 ;
      LAYER met1 ;
        RECT 3374.630 4320.620 3374.950 4320.680 ;
        RECT 3375.550 4320.620 3375.870 4320.680 ;
        RECT 3376.930 4320.620 3377.250 4320.680 ;
        RECT 3374.630 4320.480 3377.250 4320.620 ;
        RECT 3374.630 4320.420 3374.950 4320.480 ;
        RECT 3375.550 4320.420 3375.870 4320.480 ;
        RECT 3376.930 4320.420 3377.250 4320.480 ;
      LAYER met1 ;
        RECT 3381.155 4312.000 3588.000 4392.000 ;
        RECT 3407.485 4311.885 3413.015 4312.000 ;
        RECT 3418.120 4311.885 3423.725 4312.000 ;
        RECT 3439.220 4311.940 3482.580 4312.000 ;
        RECT 3439.220 4311.885 3460.930 4311.940 ;
        POLYGON 3460.930 4311.940 3460.985 4311.940 3460.930 4311.885 ;
        RECT 3483.895 4311.855 3518.220 4312.000 ;
        RECT 3519.275 4311.855 3558.090 4312.000 ;
        RECT 3566.900 4311.980 3568.975 4312.000 ;
        RECT 0.275 4208.680 197.965 4211.620 ;
        RECT 0.275 4207.540 199.030 4208.680 ;
        RECT 0.275 4151.350 197.965 4207.540 ;
        POLYGON 197.965 4207.540 198.080 4207.540 198.080 4207.425 ;
        POLYGON 198.080 4151.465 198.080 4151.350 197.965 4151.350 ;
        RECT 198.080 4151.350 199.030 4207.540 ;
        RECT 3390.035 4163.375 3587.725 4166.815 ;
        RECT 3389.130 4158.145 3587.725 4163.375 ;
        RECT 3390.035 4154.965 3587.725 4158.145 ;
        RECT 0.275 4150.035 199.030 4151.350 ;
        RECT 3388.970 4153.650 3587.725 4154.965 ;
        RECT 0.275 4138.185 197.965 4150.035 ;
        RECT 3388.970 4097.460 3389.920 4153.650 ;
        POLYGON 3389.920 4153.650 3390.035 4153.650 3389.920 4153.535 ;
        POLYGON 3389.920 4097.575 3390.035 4097.460 3389.920 4097.460 ;
        RECT 3390.035 4097.460 3587.725 4153.650 ;
        RECT 3388.970 4096.320 3587.725 4097.460 ;
        RECT 3390.035 4094.085 3587.725 4096.320 ;
      LAYER met1 ;
        RECT 3376.470 4091.800 3376.790 4091.860 ;
        RECT 3387.510 4091.800 3387.830 4091.860 ;
        RECT 3376.470 4091.660 3387.830 4091.800 ;
        RECT 3376.470 4091.600 3376.790 4091.660 ;
        RECT 3387.510 4091.600 3387.830 4091.660 ;
      LAYER met1 ;
        RECT 19.025 4002.000 21.100 4002.020 ;
        RECT 29.910 4002.000 68.725 4002.145 ;
        RECT 69.780 4002.000 104.105 4002.145 ;
        POLYGON 127.070 4002.115 127.070 4002.060 127.015 4002.060 ;
        RECT 127.070 4002.060 148.780 4002.115 ;
        RECT 105.420 4002.000 148.780 4002.060 ;
        RECT 164.275 4002.000 169.880 4002.115 ;
        RECT 174.985 4002.000 180.515 4002.115 ;
        RECT 0.000 3922.000 206.845 4002.000 ;
      LAYER met1 ;
        RECT 208.910 3997.960 209.230 3998.020 ;
        RECT 211.670 3997.960 211.990 3998.020 ;
        RECT 208.910 3997.820 211.990 3997.960 ;
        RECT 208.910 3997.760 209.230 3997.820 ;
        RECT 211.670 3997.760 211.990 3997.820 ;
        RECT 208.910 3988.780 209.230 3988.840 ;
        RECT 212.130 3988.780 212.450 3988.840 ;
        RECT 213.050 3988.780 213.370 3988.840 ;
        RECT 208.910 3988.640 213.370 3988.780 ;
        RECT 208.910 3988.580 209.230 3988.640 ;
        RECT 212.130 3988.580 212.450 3988.640 ;
        RECT 213.050 3988.580 213.370 3988.640 ;
        RECT 208.910 3962.940 209.230 3963.000 ;
        RECT 211.670 3962.940 211.990 3963.000 ;
        RECT 208.910 3962.800 211.990 3962.940 ;
        RECT 208.910 3962.740 209.230 3962.800 ;
        RECT 211.670 3962.740 211.990 3962.800 ;
      LAYER met1 ;
        RECT 3445.190 3946.000 3468.635 3946.115 ;
        RECT 3477.750 3946.000 3479.480 3946.145 ;
        RECT 3483.895 3946.000 3518.220 3946.115 ;
        RECT 3519.275 3946.000 3558.090 3946.115 ;
      LAYER met1 ;
        RECT 208.910 3936.420 209.230 3936.480 ;
        RECT 212.590 3936.420 212.910 3936.480 ;
        RECT 208.910 3936.280 212.910 3936.420 ;
        RECT 208.910 3936.220 209.230 3936.280 ;
        RECT 212.590 3936.220 212.910 3936.280 ;
        RECT 3374.170 3926.560 3374.490 3926.620 ;
        RECT 3376.930 3926.560 3377.250 3926.620 ;
        RECT 3374.170 3926.420 3377.250 3926.560 ;
        RECT 3374.170 3926.360 3374.490 3926.420 ;
        RECT 3376.930 3926.360 3377.250 3926.420 ;
      LAYER met1 ;
        RECT 29.910 3921.885 68.725 3922.000 ;
        RECT 69.780 3921.885 104.105 3922.000 ;
        RECT 108.520 3921.855 110.250 3922.000 ;
        RECT 119.365 3921.885 142.810 3922.000 ;
      LAYER met1 ;
        RECT 3375.090 3916.360 3375.410 3916.420 ;
        RECT 3376.930 3916.360 3377.250 3916.420 ;
        RECT 3375.090 3916.220 3377.250 3916.360 ;
        RECT 3375.090 3916.160 3375.410 3916.220 ;
        RECT 3376.930 3916.160 3377.250 3916.220 ;
        RECT 3376.010 3905.140 3376.330 3905.200 ;
        RECT 3376.930 3905.140 3377.250 3905.200 ;
        RECT 3376.010 3905.000 3377.250 3905.140 ;
        RECT 3376.010 3904.940 3376.330 3905.000 ;
        RECT 3376.930 3904.940 3377.250 3905.000 ;
        RECT 3374.630 3875.220 3374.950 3875.280 ;
        RECT 3376.930 3875.220 3377.250 3875.280 ;
        RECT 3374.630 3875.080 3377.250 3875.220 ;
        RECT 3374.630 3875.020 3374.950 3875.080 ;
        RECT 3376.930 3875.020 3377.250 3875.080 ;
        RECT 3376.010 3870.120 3376.330 3870.180 ;
        RECT 3376.930 3870.120 3377.250 3870.180 ;
        RECT 3376.010 3869.980 3377.250 3870.120 ;
        RECT 3376.010 3869.920 3376.330 3869.980 ;
        RECT 3376.930 3869.920 3377.250 3869.980 ;
      LAYER met1 ;
        RECT 3381.155 3866.000 3588.000 3946.000 ;
        RECT 3407.485 3865.885 3413.015 3866.000 ;
        RECT 3418.120 3865.885 3423.725 3866.000 ;
        RECT 3439.220 3865.940 3482.580 3866.000 ;
        RECT 3439.220 3865.885 3460.930 3865.940 ;
        POLYGON 3460.930 3865.940 3460.985 3865.940 3460.930 3865.885 ;
        RECT 3483.895 3865.855 3518.220 3866.000 ;
        RECT 3519.275 3865.855 3558.090 3866.000 ;
        RECT 3566.900 3865.980 3568.975 3866.000 ;
        RECT 19.025 3786.000 21.100 3786.020 ;
        RECT 29.910 3786.000 68.725 3786.145 ;
        RECT 69.780 3786.000 104.105 3786.145 ;
        POLYGON 127.070 3786.115 127.070 3786.060 127.015 3786.060 ;
        RECT 127.070 3786.060 148.780 3786.115 ;
        RECT 105.420 3786.000 148.780 3786.060 ;
        RECT 164.275 3786.000 169.880 3786.115 ;
        RECT 174.985 3786.000 180.515 3786.115 ;
        RECT 0.000 3706.000 206.845 3786.000 ;
      LAYER met1 ;
        RECT 208.910 3782.060 209.230 3782.120 ;
        RECT 213.510 3782.060 213.830 3782.120 ;
        RECT 208.910 3781.920 213.830 3782.060 ;
        RECT 208.910 3781.860 209.230 3781.920 ;
        RECT 213.510 3781.860 213.830 3781.920 ;
        RECT 208.910 3776.960 209.230 3777.020 ;
        RECT 212.130 3776.960 212.450 3777.020 ;
        RECT 213.050 3776.960 213.370 3777.020 ;
        RECT 208.910 3776.820 213.370 3776.960 ;
        RECT 208.910 3776.760 209.230 3776.820 ;
        RECT 212.130 3776.760 212.450 3776.820 ;
        RECT 213.050 3776.760 213.370 3776.820 ;
        RECT 208.910 3747.040 209.230 3747.100 ;
        RECT 213.510 3747.040 213.830 3747.100 ;
        RECT 208.910 3746.900 213.830 3747.040 ;
        RECT 208.910 3746.840 209.230 3746.900 ;
        RECT 213.510 3746.840 213.830 3746.900 ;
        RECT 208.910 3725.620 209.230 3725.680 ;
        RECT 212.590 3725.620 212.910 3725.680 ;
        RECT 208.910 3725.480 212.910 3725.620 ;
        RECT 208.910 3725.420 209.230 3725.480 ;
        RECT 212.590 3725.420 212.910 3725.480 ;
      LAYER met1 ;
        RECT 3445.190 3721.000 3468.635 3721.115 ;
        RECT 3477.750 3721.000 3479.480 3721.145 ;
        RECT 3483.895 3721.000 3518.220 3721.115 ;
        RECT 3519.275 3721.000 3558.090 3721.115 ;
        RECT 29.910 3705.885 68.725 3706.000 ;
        RECT 69.780 3705.885 104.105 3706.000 ;
        RECT 108.520 3705.855 110.250 3706.000 ;
        RECT 119.365 3705.885 142.810 3706.000 ;
      LAYER met1 ;
        RECT 3374.170 3701.820 3374.490 3701.880 ;
        RECT 3376.010 3701.820 3376.330 3701.880 ;
        RECT 3376.930 3701.820 3377.250 3701.880 ;
        RECT 3374.170 3701.680 3377.250 3701.820 ;
        RECT 3374.170 3701.620 3374.490 3701.680 ;
        RECT 3376.010 3701.620 3376.330 3701.680 ;
        RECT 3376.930 3701.620 3377.250 3701.680 ;
        RECT 3375.090 3686.520 3375.410 3686.580 ;
        RECT 3376.930 3686.520 3377.250 3686.580 ;
        RECT 3375.090 3686.380 3377.250 3686.520 ;
        RECT 3375.090 3686.320 3375.410 3686.380 ;
        RECT 3376.930 3686.320 3377.250 3686.380 ;
        RECT 3374.170 3680.060 3374.490 3680.120 ;
        RECT 3376.930 3680.060 3377.250 3680.120 ;
        RECT 3374.170 3679.920 3377.250 3680.060 ;
        RECT 3374.170 3679.860 3374.490 3679.920 ;
        RECT 3376.930 3679.860 3377.250 3679.920 ;
        RECT 3374.630 3649.800 3374.950 3649.860 ;
        RECT 3376.930 3649.800 3377.250 3649.860 ;
        RECT 3374.630 3649.660 3377.250 3649.800 ;
        RECT 3374.630 3649.600 3374.950 3649.660 ;
        RECT 3376.930 3649.600 3377.250 3649.660 ;
        RECT 3374.170 3645.380 3374.490 3645.440 ;
        RECT 3376.930 3645.380 3377.250 3645.440 ;
        RECT 3374.170 3645.240 3377.250 3645.380 ;
        RECT 3374.170 3645.180 3374.490 3645.240 ;
        RECT 3376.930 3645.180 3377.250 3645.240 ;
      LAYER met1 ;
        RECT 3381.155 3641.000 3588.000 3721.000 ;
        RECT 3407.485 3640.885 3413.015 3641.000 ;
        RECT 3418.120 3640.885 3423.725 3641.000 ;
        RECT 3439.220 3640.940 3482.580 3641.000 ;
        RECT 3439.220 3640.885 3460.930 3640.940 ;
        POLYGON 3460.930 3640.940 3460.985 3640.940 3460.930 3640.885 ;
        RECT 3483.895 3640.855 3518.220 3641.000 ;
        RECT 3519.275 3640.855 3558.090 3641.000 ;
        RECT 3566.900 3640.980 3568.975 3641.000 ;
      LAYER met1 ;
        RECT 3376.470 3633.280 3376.790 3633.540 ;
        RECT 3376.560 3632.520 3376.700 3633.280 ;
        RECT 3374.630 3632.460 3374.950 3632.520 ;
        RECT 3376.010 3632.460 3376.330 3632.520 ;
        RECT 3374.630 3632.320 3376.330 3632.460 ;
        RECT 3374.630 3632.260 3374.950 3632.320 ;
        RECT 3376.010 3632.260 3376.330 3632.320 ;
        RECT 3376.470 3632.260 3376.790 3632.520 ;
      LAYER met1 ;
        RECT 19.025 3570.000 21.100 3570.020 ;
        RECT 29.910 3570.000 68.725 3570.145 ;
        RECT 69.780 3570.000 104.105 3570.145 ;
        POLYGON 127.070 3570.115 127.070 3570.060 127.015 3570.060 ;
        RECT 127.070 3570.060 148.780 3570.115 ;
        RECT 105.420 3570.000 148.780 3570.060 ;
        RECT 164.275 3570.000 169.880 3570.115 ;
        RECT 174.985 3570.000 180.515 3570.115 ;
        RECT 0.000 3490.000 206.845 3570.000 ;
      LAYER met1 ;
        RECT 208.910 3565.820 209.230 3565.880 ;
        RECT 212.130 3565.820 212.450 3565.880 ;
        RECT 208.910 3565.680 212.450 3565.820 ;
        RECT 208.910 3565.620 209.230 3565.680 ;
        RECT 212.130 3565.620 212.450 3565.680 ;
        RECT 208.910 3558.680 209.230 3558.740 ;
        RECT 213.050 3558.680 213.370 3558.740 ;
        RECT 208.910 3558.540 213.370 3558.680 ;
        RECT 208.910 3558.480 209.230 3558.540 ;
        RECT 213.050 3558.480 213.370 3558.540 ;
        RECT 208.910 3531.140 209.230 3531.200 ;
        RECT 212.130 3531.140 212.450 3531.200 ;
        RECT 208.910 3531.000 212.450 3531.140 ;
        RECT 208.910 3530.940 209.230 3531.000 ;
        RECT 212.130 3530.940 212.450 3531.000 ;
        RECT 211.210 3525.840 211.530 3526.100 ;
        RECT 208.910 3524.680 209.230 3524.740 ;
        RECT 211.300 3524.680 211.440 3525.840 ;
        RECT 212.590 3524.680 212.910 3524.740 ;
        RECT 208.910 3524.540 212.910 3524.680 ;
        RECT 208.910 3524.480 209.230 3524.540 ;
        RECT 212.590 3524.480 212.910 3524.540 ;
        RECT 208.910 3504.280 209.230 3504.340 ;
        RECT 213.510 3504.280 213.830 3504.340 ;
        RECT 208.910 3504.140 213.830 3504.280 ;
        RECT 208.910 3504.080 209.230 3504.140 ;
        RECT 211.300 3502.640 211.440 3504.140 ;
        RECT 213.510 3504.080 213.830 3504.140 ;
        RECT 211.210 3502.380 211.530 3502.640 ;
      LAYER met1 ;
        RECT 3445.190 3496.000 3468.635 3496.115 ;
        RECT 3477.750 3496.000 3479.480 3496.145 ;
        RECT 3483.895 3496.000 3518.220 3496.115 ;
        RECT 3519.275 3496.000 3558.090 3496.115 ;
      LAYER met1 ;
        RECT 3374.630 3495.100 3374.950 3495.160 ;
        RECT 3376.930 3495.100 3377.250 3495.160 ;
        RECT 3374.630 3494.960 3377.250 3495.100 ;
        RECT 3374.630 3494.900 3374.950 3494.960 ;
        RECT 3376.930 3494.900 3377.250 3494.960 ;
      LAYER met1 ;
        RECT 29.910 3489.885 68.725 3490.000 ;
        RECT 69.780 3489.885 104.105 3490.000 ;
        RECT 108.520 3489.855 110.250 3490.000 ;
        RECT 119.365 3489.885 142.810 3490.000 ;
      LAYER met1 ;
        RECT 3374.630 3480.960 3374.950 3481.220 ;
        RECT 3374.720 3480.200 3374.860 3480.960 ;
        RECT 3374.630 3479.940 3374.950 3480.200 ;
        RECT 3374.630 3476.740 3374.950 3476.800 ;
        RECT 3376.930 3476.740 3377.250 3476.800 ;
        RECT 3374.630 3476.600 3377.250 3476.740 ;
        RECT 3374.630 3476.540 3374.950 3476.600 ;
        RECT 3376.930 3476.540 3377.250 3476.600 ;
        RECT 3374.170 3466.200 3374.490 3466.260 ;
        RECT 3376.930 3466.200 3377.250 3466.260 ;
        RECT 3374.170 3466.060 3377.250 3466.200 ;
        RECT 3374.170 3466.000 3374.490 3466.060 ;
        RECT 3376.930 3466.000 3377.250 3466.060 ;
        RECT 3376.010 3458.380 3376.330 3458.440 ;
        RECT 3376.930 3458.380 3377.250 3458.440 ;
        RECT 3376.010 3458.240 3377.250 3458.380 ;
        RECT 3376.010 3458.180 3376.330 3458.240 ;
        RECT 3376.930 3458.180 3377.250 3458.240 ;
        RECT 3376.470 3457.840 3376.790 3458.100 ;
        RECT 3376.560 3457.080 3376.700 3457.840 ;
        RECT 3376.470 3456.820 3376.790 3457.080 ;
        RECT 3375.550 3426.080 3375.870 3426.140 ;
        RECT 3376.930 3426.080 3377.250 3426.140 ;
        RECT 3375.550 3425.940 3377.250 3426.080 ;
        RECT 3375.550 3425.880 3375.870 3425.940 ;
        RECT 3376.930 3425.880 3377.250 3425.940 ;
        RECT 3376.010 3420.300 3376.330 3420.360 ;
        RECT 3376.930 3420.300 3377.250 3420.360 ;
        RECT 3376.010 3420.160 3377.250 3420.300 ;
        RECT 3376.010 3420.100 3376.330 3420.160 ;
        RECT 3376.930 3420.100 3377.250 3420.160 ;
      LAYER met1 ;
        RECT 3381.155 3416.000 3588.000 3496.000 ;
        RECT 3407.485 3415.885 3413.015 3416.000 ;
        RECT 3418.120 3415.885 3423.725 3416.000 ;
        RECT 3439.220 3415.940 3482.580 3416.000 ;
        RECT 3439.220 3415.885 3460.930 3415.940 ;
        POLYGON 3460.930 3415.940 3460.985 3415.940 3460.930 3415.885 ;
        RECT 3483.895 3415.855 3518.220 3416.000 ;
        RECT 3519.275 3415.855 3558.090 3416.000 ;
        RECT 3566.900 3415.980 3568.975 3416.000 ;
      LAYER met1 ;
        RECT 3375.090 3357.060 3375.410 3357.120 ;
        RECT 3376.010 3357.060 3376.330 3357.120 ;
        RECT 3375.090 3356.920 3376.330 3357.060 ;
        RECT 3375.090 3356.860 3375.410 3356.920 ;
        RECT 3376.010 3356.860 3376.330 3356.920 ;
      LAYER met1 ;
        RECT 19.025 3354.000 21.100 3354.020 ;
        RECT 29.910 3354.000 68.725 3354.145 ;
        RECT 69.780 3354.000 104.105 3354.145 ;
        POLYGON 127.070 3354.115 127.070 3354.060 127.015 3354.060 ;
        RECT 127.070 3354.060 148.780 3354.115 ;
        RECT 105.420 3354.000 148.780 3354.060 ;
        RECT 164.275 3354.000 169.880 3354.115 ;
        RECT 174.985 3354.000 180.515 3354.115 ;
        RECT 0.000 3274.000 206.845 3354.000 ;
      LAYER met1 ;
        RECT 208.910 3349.920 209.230 3349.980 ;
        RECT 212.130 3349.920 212.450 3349.980 ;
        RECT 208.910 3349.780 212.450 3349.920 ;
        RECT 208.910 3349.720 209.230 3349.780 ;
        RECT 212.130 3349.720 212.450 3349.780 ;
        RECT 208.910 3342.780 209.230 3342.840 ;
        RECT 213.050 3342.780 213.370 3342.840 ;
        RECT 208.910 3342.640 213.370 3342.780 ;
        RECT 208.910 3342.580 209.230 3342.640 ;
        RECT 213.050 3342.580 213.370 3342.640 ;
        RECT 212.130 3315.580 212.450 3315.640 ;
        RECT 209.000 3315.440 212.450 3315.580 ;
        RECT 209.000 3315.300 209.140 3315.440 ;
        RECT 212.130 3315.380 212.450 3315.440 ;
        RECT 208.910 3315.040 209.230 3315.300 ;
        RECT 211.210 3315.240 211.530 3315.300 ;
        RECT 211.210 3315.100 212.360 3315.240 ;
        RECT 211.210 3315.040 211.530 3315.100 ;
        RECT 212.220 3314.280 212.360 3315.100 ;
        RECT 212.130 3314.020 212.450 3314.280 ;
        RECT 208.910 3304.020 209.230 3304.080 ;
        RECT 212.130 3304.020 212.450 3304.080 ;
        RECT 208.910 3303.880 212.450 3304.020 ;
        RECT 208.910 3303.820 209.230 3303.880 ;
        RECT 212.130 3303.820 212.450 3303.880 ;
        RECT 208.910 3293.480 209.230 3293.540 ;
        RECT 211.670 3293.480 211.990 3293.540 ;
        RECT 213.510 3293.480 213.830 3293.540 ;
        RECT 208.910 3293.340 213.830 3293.480 ;
        RECT 208.910 3293.280 209.230 3293.340 ;
        RECT 211.670 3293.280 211.990 3293.340 ;
        RECT 213.510 3293.280 213.830 3293.340 ;
      LAYER met1 ;
        RECT 29.910 3273.885 68.725 3274.000 ;
        RECT 69.780 3273.885 104.105 3274.000 ;
        RECT 108.520 3273.855 110.250 3274.000 ;
        RECT 119.365 3273.885 142.810 3274.000 ;
        RECT 3445.190 3270.000 3468.635 3270.115 ;
        RECT 3477.750 3270.000 3479.480 3270.145 ;
        RECT 3483.895 3270.000 3518.220 3270.115 ;
        RECT 3519.275 3270.000 3558.090 3270.115 ;
      LAYER met1 ;
        RECT 3374.630 3250.640 3374.950 3250.700 ;
        RECT 3376.930 3250.640 3377.250 3250.700 ;
        RECT 3374.630 3250.500 3377.250 3250.640 ;
        RECT 3374.630 3250.440 3374.950 3250.500 ;
        RECT 3376.930 3250.440 3377.250 3250.500 ;
        RECT 3374.170 3240.100 3374.490 3240.160 ;
        RECT 3376.930 3240.100 3377.250 3240.160 ;
        RECT 3374.170 3239.960 3377.250 3240.100 ;
        RECT 3374.170 3239.900 3374.490 3239.960 ;
        RECT 3376.930 3239.900 3377.250 3239.960 ;
        RECT 3376.010 3228.880 3376.330 3228.940 ;
        RECT 3376.930 3228.880 3377.250 3228.940 ;
        RECT 3376.010 3228.740 3377.250 3228.880 ;
        RECT 3376.010 3228.680 3376.330 3228.740 ;
        RECT 3376.930 3228.680 3377.250 3228.740 ;
        RECT 3375.090 3198.960 3375.410 3199.020 ;
        RECT 3376.930 3198.960 3377.250 3199.020 ;
        RECT 3375.090 3198.820 3377.250 3198.960 ;
        RECT 3375.090 3198.760 3375.410 3198.820 ;
        RECT 3376.930 3198.760 3377.250 3198.820 ;
        RECT 3376.010 3194.200 3376.330 3194.260 ;
        RECT 3376.930 3194.200 3377.250 3194.260 ;
        RECT 3376.010 3194.060 3377.250 3194.200 ;
        RECT 3376.010 3194.000 3376.330 3194.060 ;
        RECT 3376.930 3194.000 3377.250 3194.060 ;
      LAYER met1 ;
        RECT 3381.155 3190.000 3588.000 3270.000 ;
        RECT 3407.485 3189.885 3413.015 3190.000 ;
        RECT 3418.120 3189.885 3423.725 3190.000 ;
        RECT 3439.220 3189.940 3482.580 3190.000 ;
        RECT 3439.220 3189.885 3460.930 3189.940 ;
        POLYGON 3460.930 3189.940 3460.985 3189.940 3460.930 3189.885 ;
        RECT 3483.895 3189.855 3518.220 3190.000 ;
        RECT 3519.275 3189.855 3558.090 3190.000 ;
        RECT 3566.900 3189.980 3568.975 3190.000 ;
        RECT 19.025 3138.000 21.100 3138.020 ;
        RECT 29.910 3138.000 68.725 3138.145 ;
        RECT 69.780 3138.000 104.105 3138.145 ;
        POLYGON 127.070 3138.115 127.070 3138.060 127.015 3138.060 ;
        RECT 127.070 3138.060 148.780 3138.115 ;
        RECT 105.420 3138.000 148.780 3138.060 ;
        RECT 164.275 3138.000 169.880 3138.115 ;
        RECT 174.985 3138.000 180.515 3138.115 ;
        RECT 0.000 3058.000 206.845 3138.000 ;
      LAYER met1 ;
        RECT 209.830 3125.520 210.150 3125.580 ;
        RECT 213.050 3125.520 213.370 3125.580 ;
        RECT 209.830 3125.380 213.370 3125.520 ;
        RECT 209.830 3125.320 210.150 3125.380 ;
        RECT 213.050 3125.320 213.370 3125.380 ;
        RECT 208.910 3092.540 209.230 3092.600 ;
        RECT 212.130 3092.540 212.450 3092.600 ;
        RECT 208.910 3092.400 212.450 3092.540 ;
        RECT 208.910 3092.340 209.230 3092.400 ;
        RECT 212.130 3092.340 212.450 3092.400 ;
        RECT 211.210 3074.860 211.530 3074.920 ;
        RECT 213.510 3074.860 213.830 3074.920 ;
        RECT 211.210 3074.720 213.830 3074.860 ;
        RECT 211.210 3074.660 211.530 3074.720 ;
        RECT 213.510 3074.660 213.830 3074.720 ;
      LAYER met1 ;
        RECT 29.910 3057.885 68.725 3058.000 ;
        RECT 69.780 3057.885 104.105 3058.000 ;
        RECT 108.520 3057.855 110.250 3058.000 ;
        RECT 119.365 3057.885 142.810 3058.000 ;
        RECT 3445.190 3045.000 3468.635 3045.115 ;
        RECT 3477.750 3045.000 3479.480 3045.145 ;
        RECT 3483.895 3045.000 3518.220 3045.115 ;
        RECT 3519.275 3045.000 3558.090 3045.115 ;
      LAYER met1 ;
        RECT 212.590 3029.300 212.910 3029.360 ;
        RECT 213.510 3029.300 213.830 3029.360 ;
        RECT 212.590 3029.160 213.830 3029.300 ;
        RECT 212.590 3029.100 212.910 3029.160 ;
        RECT 213.510 3029.100 213.830 3029.160 ;
        RECT 3374.630 3027.600 3374.950 3027.660 ;
        RECT 3376.930 3027.600 3377.250 3027.660 ;
        RECT 3374.630 3027.460 3377.250 3027.600 ;
        RECT 3374.630 3027.400 3374.950 3027.460 ;
        RECT 3376.930 3027.400 3377.250 3027.460 ;
        RECT 3374.170 3011.960 3374.490 3012.020 ;
        RECT 3374.170 3011.820 3374.860 3011.960 ;
        RECT 3374.170 3011.760 3374.490 3011.820 ;
        RECT 3374.720 3010.660 3374.860 3011.820 ;
        RECT 3374.630 3010.600 3374.950 3010.660 ;
        RECT 3376.930 3010.600 3377.250 3010.660 ;
        RECT 3374.630 3010.460 3377.250 3010.600 ;
        RECT 3374.630 3010.400 3374.950 3010.460 ;
        RECT 3376.930 3010.400 3377.250 3010.460 ;
        RECT 3376.010 3004.140 3376.330 3004.200 ;
        RECT 3376.930 3004.140 3377.250 3004.200 ;
        RECT 3376.010 3004.000 3377.250 3004.140 ;
        RECT 3376.010 3003.940 3376.330 3004.000 ;
        RECT 3376.930 3003.940 3377.250 3004.000 ;
        RECT 3375.090 2973.540 3375.410 2973.600 ;
        RECT 3376.930 2973.540 3377.250 2973.600 ;
        RECT 3375.090 2973.400 3377.250 2973.540 ;
        RECT 3375.090 2973.340 3375.410 2973.400 ;
        RECT 3376.930 2973.340 3377.250 2973.400 ;
        RECT 3376.010 2969.120 3376.330 2969.180 ;
        RECT 3376.930 2969.120 3377.250 2969.180 ;
        RECT 3376.010 2968.980 3377.250 2969.120 ;
        RECT 3376.010 2968.920 3376.330 2968.980 ;
        RECT 3376.930 2968.920 3377.250 2968.980 ;
      LAYER met1 ;
        RECT 3381.155 2965.000 3588.000 3045.000 ;
        RECT 3407.485 2964.885 3413.015 2965.000 ;
        RECT 3418.120 2964.885 3423.725 2965.000 ;
        RECT 3439.220 2964.940 3482.580 2965.000 ;
        RECT 3439.220 2964.885 3460.930 2964.940 ;
        POLYGON 3460.930 2964.940 3460.985 2964.940 3460.930 2964.885 ;
        RECT 3483.895 2964.855 3518.220 2965.000 ;
        RECT 3519.275 2964.855 3558.090 2965.000 ;
        RECT 3566.900 2964.980 3568.975 2965.000 ;
        RECT 19.025 2922.000 21.100 2922.020 ;
        RECT 29.910 2922.000 68.725 2922.145 ;
        RECT 69.780 2922.000 104.105 2922.145 ;
        POLYGON 127.070 2922.115 127.070 2922.060 127.015 2922.060 ;
        RECT 127.070 2922.060 148.780 2922.115 ;
        RECT 105.420 2922.000 148.780 2922.060 ;
        RECT 164.275 2922.000 169.880 2922.115 ;
        RECT 174.985 2922.000 180.515 2922.115 ;
        RECT 0.000 2842.000 206.845 2922.000 ;
      LAYER met1 ;
        RECT 208.910 2917.780 209.230 2917.840 ;
        RECT 212.130 2917.780 212.450 2917.840 ;
        RECT 208.910 2917.640 212.450 2917.780 ;
        RECT 208.910 2917.580 209.230 2917.640 ;
        RECT 212.130 2917.580 212.450 2917.640 ;
        RECT 208.910 2909.280 209.230 2909.340 ;
        RECT 212.590 2909.280 212.910 2909.340 ;
        RECT 208.910 2909.140 212.910 2909.280 ;
        RECT 208.910 2909.080 209.230 2909.140 ;
        RECT 212.590 2909.080 212.910 2909.140 ;
        RECT 208.910 2882.420 209.230 2882.480 ;
        RECT 212.130 2882.420 212.450 2882.480 ;
        RECT 208.910 2882.280 212.450 2882.420 ;
        RECT 208.910 2882.220 209.230 2882.280 ;
        RECT 212.130 2882.220 212.450 2882.280 ;
        RECT 211.210 2881.400 211.530 2881.460 ;
        RECT 213.510 2881.400 213.830 2881.460 ;
        RECT 211.210 2881.260 213.830 2881.400 ;
        RECT 211.210 2881.200 211.530 2881.260 ;
        RECT 213.510 2881.200 213.830 2881.260 ;
        RECT 208.910 2871.880 209.230 2871.940 ;
        RECT 212.130 2871.880 212.450 2871.940 ;
        RECT 213.050 2871.880 213.370 2871.940 ;
        RECT 208.910 2871.740 213.370 2871.880 ;
        RECT 208.910 2871.680 209.230 2871.740 ;
        RECT 212.130 2871.680 212.450 2871.740 ;
        RECT 213.050 2871.680 213.370 2871.740 ;
        RECT 208.910 2858.280 209.230 2858.340 ;
        RECT 213.050 2858.280 213.370 2858.340 ;
        RECT 208.910 2858.140 213.370 2858.280 ;
        RECT 208.910 2858.080 209.230 2858.140 ;
        RECT 213.050 2858.080 213.370 2858.140 ;
      LAYER met1 ;
        RECT 29.910 2841.885 68.725 2842.000 ;
        RECT 69.780 2841.885 104.105 2842.000 ;
        RECT 108.520 2841.855 110.250 2842.000 ;
        RECT 119.365 2841.885 142.810 2842.000 ;
        RECT 3445.190 2819.000 3468.635 2819.115 ;
        RECT 3477.750 2819.000 3479.480 2819.145 ;
        RECT 3483.895 2819.000 3518.220 2819.115 ;
        RECT 3519.275 2819.000 3558.090 2819.115 ;
      LAYER met1 ;
        RECT 3374.170 2804.900 3374.490 2804.960 ;
        RECT 3376.930 2804.900 3377.250 2804.960 ;
        RECT 3374.170 2804.760 3377.250 2804.900 ;
        RECT 3374.170 2804.700 3374.490 2804.760 ;
        RECT 3376.930 2804.700 3377.250 2804.760 ;
        RECT 3374.630 2789.260 3374.950 2789.320 ;
        RECT 3376.930 2789.260 3377.250 2789.320 ;
        RECT 3374.630 2789.120 3377.250 2789.260 ;
        RECT 3374.630 2789.060 3374.950 2789.120 ;
        RECT 3376.930 2789.060 3377.250 2789.120 ;
        RECT 3376.010 2778.040 3376.330 2778.100 ;
        RECT 3376.930 2778.040 3377.250 2778.100 ;
        RECT 3376.010 2777.900 3377.250 2778.040 ;
        RECT 3376.010 2777.840 3376.330 2777.900 ;
        RECT 3376.930 2777.840 3377.250 2777.900 ;
        RECT 3375.090 2752.540 3375.410 2752.600 ;
        RECT 3376.930 2752.540 3377.250 2752.600 ;
        RECT 3375.090 2752.400 3377.250 2752.540 ;
        RECT 3375.090 2752.340 3375.410 2752.400 ;
        RECT 3376.930 2752.340 3377.250 2752.400 ;
      LAYER met1 ;
        RECT 3381.155 2739.000 3588.000 2819.000 ;
        RECT 3407.485 2738.885 3413.015 2739.000 ;
        RECT 3418.120 2738.885 3423.725 2739.000 ;
        RECT 3439.220 2738.940 3482.580 2739.000 ;
        RECT 3439.220 2738.885 3460.930 2738.940 ;
        POLYGON 3460.930 2738.940 3460.985 2738.940 3460.930 2738.885 ;
        RECT 3483.895 2738.855 3518.220 2739.000 ;
        RECT 3519.275 2738.855 3558.090 2739.000 ;
        RECT 3566.900 2738.980 3568.975 2739.000 ;
        RECT 19.025 2706.000 21.100 2706.020 ;
        RECT 29.910 2706.000 68.725 2706.145 ;
        RECT 69.780 2706.000 104.105 2706.145 ;
        POLYGON 127.070 2706.115 127.070 2706.060 127.015 2706.060 ;
        RECT 127.070 2706.060 148.780 2706.115 ;
        RECT 105.420 2706.000 148.780 2706.060 ;
        RECT 164.275 2706.000 169.880 2706.115 ;
        RECT 174.985 2706.000 180.515 2706.115 ;
        RECT 0.000 2626.000 206.845 2706.000 ;
      LAYER met1 ;
        RECT 208.910 2695.760 209.230 2695.820 ;
        RECT 212.590 2695.760 212.910 2695.820 ;
        RECT 208.910 2695.620 212.910 2695.760 ;
        RECT 208.910 2695.560 209.230 2695.620 ;
        RECT 212.590 2695.560 212.910 2695.620 ;
        RECT 208.910 2660.740 209.230 2660.800 ;
        RECT 212.130 2660.740 212.450 2660.800 ;
        RECT 208.910 2660.600 212.450 2660.740 ;
        RECT 208.910 2660.540 209.230 2660.600 ;
        RECT 212.130 2660.540 212.450 2660.600 ;
        RECT 209.830 2642.380 210.150 2642.440 ;
        RECT 213.510 2642.380 213.830 2642.440 ;
        RECT 209.830 2642.240 213.830 2642.380 ;
        RECT 209.830 2642.180 210.150 2642.240 ;
        RECT 213.510 2642.180 213.830 2642.240 ;
      LAYER met1 ;
        RECT 29.910 2625.885 68.725 2626.000 ;
        RECT 69.780 2625.885 104.105 2626.000 ;
        RECT 108.520 2625.855 110.250 2626.000 ;
        RECT 119.365 2625.885 142.810 2626.000 ;
        RECT 3390.035 2590.375 3587.725 2593.815 ;
        RECT 3389.130 2585.145 3587.725 2590.375 ;
        RECT 3390.035 2581.965 3587.725 2585.145 ;
        RECT 3388.970 2580.650 3587.725 2581.965 ;
        RECT 3388.970 2524.460 3389.920 2580.650 ;
        POLYGON 3389.920 2580.650 3390.035 2580.650 3389.920 2580.535 ;
        POLYGON 3389.920 2524.575 3390.035 2524.460 3389.920 2524.460 ;
        RECT 3390.035 2524.460 3587.725 2580.650 ;
        RECT 3388.970 2523.320 3587.725 2524.460 ;
        RECT 3390.035 2521.085 3587.725 2523.320 ;
      LAYER met1 ;
        RECT 3376.470 2519.640 3376.790 2519.700 ;
        RECT 3387.510 2519.640 3387.830 2519.700 ;
        RECT 3376.470 2519.500 3387.830 2519.640 ;
        RECT 3376.470 2519.440 3376.790 2519.500 ;
        RECT 3387.510 2519.440 3387.830 2519.500 ;
      LAYER met1 ;
        RECT 0.275 2485.680 197.965 2487.915 ;
        RECT 0.275 2484.540 199.030 2485.680 ;
        RECT 0.275 2428.350 197.965 2484.540 ;
        POLYGON 197.965 2484.540 198.080 2484.540 198.080 2484.425 ;
        POLYGON 198.080 2428.465 198.080 2428.350 197.965 2428.350 ;
        RECT 198.080 2428.350 199.030 2484.540 ;
        RECT 0.275 2427.035 199.030 2428.350 ;
        RECT 0.275 2423.855 197.965 2427.035 ;
        RECT 0.275 2418.625 198.870 2423.855 ;
        RECT 0.275 2415.185 197.965 2418.625 ;
        RECT 3390.035 2357.345 3587.840 2373.880 ;
        RECT 3390.000 2353.075 3587.840 2357.345 ;
        RECT 3379.115 2317.435 3587.840 2353.075 ;
        RECT 3379.115 2297.800 3389.220 2317.435 ;
        RECT 3390.035 2299.000 3587.840 2317.435 ;
        RECT 3379.115 2292.065 3465.385 2297.800 ;
        POLYGON 3379.115 2292.065 3381.245 2292.065 3381.245 2289.935 ;
        RECT 3381.245 2289.935 3465.385 2292.065 ;
        RECT 122.615 2285.935 204.885 2289.935 ;
        POLYGON 204.885 2289.935 208.885 2285.935 204.885 2285.935 ;
        POLYGON 3381.245 2289.935 3383.115 2289.935 3383.115 2288.065 ;
        RECT 3383.115 2288.065 3465.385 2289.935 ;
        RECT 122.615 2280.200 208.885 2285.935 ;
        RECT 0.160 2260.565 197.965 2279.000 ;
        RECT 198.780 2260.565 208.885 2280.200 ;
        RECT 0.160 2224.925 208.885 2260.565 ;
        RECT 0.160 2220.655 198.000 2224.925 ;
        RECT 0.160 2204.120 197.965 2220.655 ;
        RECT 3390.035 2140.965 3587.725 2152.815 ;
        RECT 3388.970 2139.650 3587.725 2140.965 ;
      LAYER met1 ;
        RECT 3370.490 2139.180 3370.810 2139.240 ;
        RECT 3387.510 2139.180 3387.830 2139.240 ;
        RECT 3370.490 2139.040 3387.830 2139.180 ;
        RECT 3370.490 2138.980 3370.810 2139.040 ;
        RECT 3387.510 2138.980 3387.830 2139.040 ;
      LAYER met1 ;
        RECT 3388.970 2083.460 3389.920 2139.650 ;
        POLYGON 3389.920 2139.650 3390.035 2139.650 3389.920 2139.535 ;
        POLYGON 3389.920 2083.575 3390.035 2083.460 3389.920 2083.460 ;
        RECT 3390.035 2083.460 3587.725 2139.650 ;
        RECT 3388.970 2082.320 3587.725 2083.460 ;
        RECT 3390.035 2079.380 3587.725 2082.320 ;
        RECT 19.025 2068.000 21.100 2068.020 ;
        RECT 29.910 2068.000 68.725 2068.145 ;
        RECT 69.780 2068.000 104.105 2068.145 ;
        POLYGON 127.070 2068.115 127.070 2068.060 127.015 2068.060 ;
        RECT 127.070 2068.060 148.780 2068.115 ;
        RECT 105.420 2068.000 148.780 2068.060 ;
        RECT 164.275 2068.000 169.880 2068.115 ;
        RECT 174.985 2068.000 180.515 2068.115 ;
        RECT 0.000 1988.000 206.845 2068.000 ;
      LAYER met1 ;
        RECT 208.910 2064.720 209.230 2064.780 ;
        RECT 211.670 2064.720 211.990 2064.780 ;
        RECT 208.910 2064.580 211.990 2064.720 ;
        RECT 208.910 2064.520 209.230 2064.580 ;
        RECT 211.670 2064.520 211.990 2064.580 ;
        RECT 208.910 2054.860 209.230 2054.920 ;
        RECT 213.050 2054.860 213.370 2054.920 ;
        RECT 208.910 2054.720 213.370 2054.860 ;
        RECT 208.910 2054.660 209.230 2054.720 ;
        RECT 213.050 2054.660 213.370 2054.720 ;
        RECT 208.910 2029.020 209.230 2029.080 ;
        RECT 211.670 2029.020 211.990 2029.080 ;
        RECT 208.910 2028.880 211.990 2029.020 ;
        RECT 208.910 2028.820 209.230 2028.880 ;
        RECT 211.670 2028.820 211.990 2028.880 ;
        RECT 208.910 2022.560 209.230 2022.620 ;
        RECT 212.130 2022.560 212.450 2022.620 ;
        RECT 208.910 2022.420 212.450 2022.560 ;
        RECT 208.910 2022.360 209.230 2022.420 ;
        RECT 212.130 2022.360 212.450 2022.420 ;
        RECT 208.910 2002.160 209.230 2002.220 ;
        RECT 212.130 2002.160 212.450 2002.220 ;
        RECT 213.510 2002.160 213.830 2002.220 ;
        RECT 208.910 2002.020 213.830 2002.160 ;
        RECT 208.910 2001.960 209.230 2002.020 ;
        RECT 212.130 2001.960 212.450 2002.020 ;
        RECT 213.510 2001.960 213.830 2002.020 ;
      LAYER met1 ;
        RECT 29.910 1987.885 68.725 1988.000 ;
        RECT 69.780 1987.885 104.105 1988.000 ;
        RECT 108.520 1987.855 110.250 1988.000 ;
        RECT 119.365 1987.885 142.810 1988.000 ;
        RECT 3445.190 1933.000 3468.635 1933.115 ;
        RECT 3477.750 1933.000 3479.480 1933.145 ;
        RECT 3483.895 1933.000 3518.220 1933.115 ;
        RECT 3519.275 1933.000 3558.090 1933.115 ;
      LAYER met1 ;
        RECT 3374.170 1918.860 3374.490 1918.920 ;
        RECT 3376.930 1918.860 3377.250 1918.920 ;
        RECT 3374.170 1918.720 3377.250 1918.860 ;
        RECT 3374.170 1918.660 3374.490 1918.720 ;
        RECT 3376.930 1918.660 3377.250 1918.720 ;
        RECT 3375.090 1899.140 3375.410 1899.200 ;
        RECT 3376.930 1899.140 3377.250 1899.200 ;
        RECT 3375.090 1899.000 3377.250 1899.140 ;
        RECT 3375.090 1898.940 3375.410 1899.000 ;
        RECT 3376.930 1898.940 3377.250 1899.000 ;
        RECT 3374.170 1892.000 3374.490 1892.060 ;
        RECT 3376.930 1892.000 3377.250 1892.060 ;
        RECT 3374.170 1891.860 3377.250 1892.000 ;
        RECT 3374.170 1891.800 3374.490 1891.860 ;
        RECT 3376.930 1891.800 3377.250 1891.860 ;
        RECT 3374.170 1857.320 3374.490 1857.380 ;
        RECT 3376.930 1857.320 3377.250 1857.380 ;
        RECT 3374.170 1857.180 3377.250 1857.320 ;
        RECT 3374.170 1857.120 3374.490 1857.180 ;
        RECT 3376.930 1857.120 3377.250 1857.180 ;
      LAYER met1 ;
        RECT 3381.155 1853.000 3588.000 1933.000 ;
        RECT 3407.485 1852.885 3413.015 1853.000 ;
        RECT 3418.120 1852.885 3423.725 1853.000 ;
        RECT 3439.220 1852.940 3482.580 1853.000 ;
        RECT 3439.220 1852.885 3460.930 1852.940 ;
        POLYGON 3460.930 1852.940 3460.985 1852.940 3460.930 1852.885 ;
        RECT 3483.895 1852.855 3518.220 1853.000 ;
        RECT 3519.275 1852.855 3558.090 1853.000 ;
        RECT 3566.900 1852.980 3568.975 1853.000 ;
        RECT 19.025 1852.000 21.100 1852.020 ;
        RECT 29.910 1852.000 68.725 1852.145 ;
        RECT 69.780 1852.000 104.105 1852.145 ;
        POLYGON 127.070 1852.115 127.070 1852.060 127.015 1852.060 ;
        RECT 127.070 1852.060 148.780 1852.115 ;
        RECT 105.420 1852.000 148.780 1852.060 ;
        RECT 164.275 1852.000 169.880 1852.115 ;
        RECT 174.985 1852.000 180.515 1852.115 ;
        RECT 0.000 1772.000 206.845 1852.000 ;
      LAYER met1 ;
        RECT 208.910 1847.800 209.230 1847.860 ;
        RECT 211.670 1847.800 211.990 1847.860 ;
        RECT 208.910 1847.660 211.990 1847.800 ;
        RECT 208.910 1847.600 209.230 1847.660 ;
        RECT 211.670 1847.600 211.990 1847.660 ;
        RECT 208.910 1843.380 209.230 1843.440 ;
        RECT 213.050 1843.380 213.370 1843.440 ;
        RECT 208.910 1843.240 213.370 1843.380 ;
        RECT 208.910 1843.180 209.230 1843.240 ;
        RECT 213.050 1843.180 213.370 1843.240 ;
        RECT 208.910 1813.120 209.230 1813.180 ;
        RECT 211.670 1813.120 211.990 1813.180 ;
        RECT 208.910 1812.980 211.990 1813.120 ;
        RECT 208.910 1812.920 209.230 1812.980 ;
        RECT 211.670 1812.920 211.990 1812.980 ;
        RECT 208.910 1801.900 209.230 1801.960 ;
        RECT 212.590 1801.900 212.910 1801.960 ;
        RECT 213.510 1801.900 213.830 1801.960 ;
        RECT 208.910 1801.760 213.830 1801.900 ;
        RECT 208.910 1801.700 209.230 1801.760 ;
        RECT 212.590 1801.700 212.910 1801.760 ;
        RECT 213.510 1801.700 213.830 1801.760 ;
        RECT 208.910 1786.260 209.230 1786.320 ;
        RECT 212.130 1786.260 212.450 1786.320 ;
        RECT 208.910 1786.120 212.450 1786.260 ;
        RECT 208.910 1786.060 209.230 1786.120 ;
        RECT 211.300 1785.300 211.440 1786.120 ;
        RECT 212.130 1786.060 212.450 1786.120 ;
        RECT 211.210 1785.040 211.530 1785.300 ;
      LAYER met1 ;
        RECT 29.910 1771.885 68.725 1772.000 ;
        RECT 69.780 1771.885 104.105 1772.000 ;
        RECT 108.520 1771.855 110.250 1772.000 ;
        RECT 119.365 1771.885 142.810 1772.000 ;
        RECT 3445.190 1707.000 3468.635 1707.115 ;
        RECT 3477.750 1707.000 3479.480 1707.145 ;
        RECT 3483.895 1707.000 3518.220 1707.115 ;
        RECT 3519.275 1707.000 3558.090 1707.115 ;
      LAYER met1 ;
        RECT 3374.630 1687.660 3374.950 1687.720 ;
        RECT 3376.930 1687.660 3377.250 1687.720 ;
        RECT 3374.630 1687.520 3377.250 1687.660 ;
        RECT 3374.630 1687.460 3374.950 1687.520 ;
        RECT 3376.930 1687.460 3377.250 1687.520 ;
        RECT 3375.090 1677.120 3375.410 1677.180 ;
        RECT 3376.010 1677.120 3376.330 1677.180 ;
        RECT 3376.930 1677.120 3377.250 1677.180 ;
        RECT 3375.090 1676.980 3377.250 1677.120 ;
        RECT 3375.090 1676.920 3375.410 1676.980 ;
        RECT 3376.010 1676.920 3376.330 1676.980 ;
        RECT 3376.930 1676.920 3377.250 1676.980 ;
        RECT 3374.170 1640.400 3374.490 1640.460 ;
        RECT 3375.550 1640.400 3375.870 1640.460 ;
        RECT 3376.930 1640.400 3377.250 1640.460 ;
        RECT 3374.170 1640.260 3377.250 1640.400 ;
        RECT 3374.170 1640.200 3374.490 1640.260 ;
        RECT 3375.550 1640.200 3375.870 1640.260 ;
        RECT 3376.930 1640.200 3377.250 1640.260 ;
      LAYER met1 ;
        RECT 19.025 1636.000 21.100 1636.020 ;
        RECT 29.910 1636.000 68.725 1636.145 ;
        RECT 69.780 1636.000 104.105 1636.145 ;
        POLYGON 127.070 1636.115 127.070 1636.060 127.015 1636.060 ;
        RECT 127.070 1636.060 148.780 1636.115 ;
        RECT 105.420 1636.000 148.780 1636.060 ;
        RECT 164.275 1636.000 169.880 1636.115 ;
        RECT 174.985 1636.000 180.515 1636.115 ;
        RECT 0.000 1556.000 206.845 1636.000 ;
      LAYER met1 ;
        RECT 208.910 1631.900 209.230 1631.960 ;
        RECT 212.130 1631.900 212.450 1631.960 ;
        RECT 208.910 1631.760 212.450 1631.900 ;
        RECT 208.910 1631.700 209.230 1631.760 ;
        RECT 212.130 1631.700 212.450 1631.760 ;
      LAYER met1 ;
        RECT 3381.155 1627.000 3588.000 1707.000 ;
        RECT 3407.485 1626.885 3413.015 1627.000 ;
        RECT 3418.120 1626.885 3423.725 1627.000 ;
        RECT 3439.220 1626.940 3482.580 1627.000 ;
        RECT 3439.220 1626.885 3460.930 1626.940 ;
        POLYGON 3460.930 1626.940 3460.985 1626.940 3460.930 1626.885 ;
        RECT 3483.895 1626.855 3518.220 1627.000 ;
        RECT 3519.275 1626.855 3558.090 1627.000 ;
        RECT 3566.900 1626.980 3568.975 1627.000 ;
      LAYER met1 ;
        RECT 208.910 1625.780 209.230 1625.840 ;
        RECT 212.590 1625.780 212.910 1625.840 ;
        RECT 208.910 1625.640 212.910 1625.780 ;
        RECT 208.910 1625.580 209.230 1625.640 ;
        RECT 212.590 1625.580 212.910 1625.640 ;
        RECT 208.910 1597.220 209.230 1597.280 ;
        RECT 212.130 1597.220 212.450 1597.280 ;
        RECT 208.910 1597.080 212.450 1597.220 ;
        RECT 208.910 1597.020 209.230 1597.080 ;
        RECT 212.130 1597.020 212.450 1597.080 ;
        RECT 208.910 1590.760 209.230 1590.820 ;
        RECT 213.510 1590.760 213.830 1590.820 ;
        RECT 208.910 1590.620 213.830 1590.760 ;
        RECT 208.910 1590.560 209.230 1590.620 ;
        RECT 213.510 1590.560 213.830 1590.620 ;
      LAYER met1 ;
        RECT 29.910 1555.885 68.725 1556.000 ;
        RECT 69.780 1555.885 104.105 1556.000 ;
        RECT 108.520 1555.855 110.250 1556.000 ;
        RECT 119.365 1555.885 142.810 1556.000 ;
        RECT 3445.190 1482.000 3468.635 1482.115 ;
        RECT 3477.750 1482.000 3479.480 1482.145 ;
        RECT 3483.895 1482.000 3518.220 1482.115 ;
        RECT 3519.275 1482.000 3558.090 1482.115 ;
      LAYER met1 ;
        RECT 3374.630 1466.320 3374.950 1466.380 ;
        RECT 3376.930 1466.320 3377.250 1466.380 ;
        RECT 3374.630 1466.180 3377.250 1466.320 ;
        RECT 3374.630 1466.120 3374.950 1466.180 ;
        RECT 3376.930 1466.120 3377.250 1466.180 ;
        RECT 3374.630 1447.620 3374.950 1447.680 ;
        RECT 3375.550 1447.620 3375.870 1447.680 ;
        RECT 3376.930 1447.620 3377.250 1447.680 ;
        RECT 3374.630 1447.480 3377.250 1447.620 ;
        RECT 3374.630 1447.420 3374.950 1447.480 ;
        RECT 3375.550 1447.420 3375.870 1447.480 ;
        RECT 3376.930 1447.420 3377.250 1447.480 ;
        RECT 3375.090 1443.200 3375.410 1443.260 ;
        RECT 3376.470 1443.200 3376.790 1443.260 ;
        RECT 3375.090 1443.060 3376.790 1443.200 ;
        RECT 3375.090 1443.000 3375.410 1443.060 ;
        RECT 3376.470 1443.000 3376.790 1443.060 ;
      LAYER met1 ;
        RECT 19.025 1420.000 21.100 1420.020 ;
        RECT 29.910 1420.000 68.725 1420.145 ;
        RECT 69.780 1420.000 104.105 1420.145 ;
        POLYGON 127.070 1420.115 127.070 1420.060 127.015 1420.060 ;
        RECT 127.070 1420.060 148.780 1420.115 ;
        RECT 105.420 1420.000 148.780 1420.060 ;
        RECT 164.275 1420.000 169.880 1420.115 ;
        RECT 174.985 1420.000 180.515 1420.115 ;
        RECT 0.000 1340.000 206.845 1420.000 ;
      LAYER met1 ;
        RECT 208.910 1416.000 209.230 1416.060 ;
        RECT 212.130 1416.000 212.450 1416.060 ;
        RECT 208.910 1415.860 212.450 1416.000 ;
        RECT 208.910 1415.800 209.230 1415.860 ;
        RECT 212.130 1415.800 212.450 1415.860 ;
        RECT 3374.170 1411.580 3374.490 1411.640 ;
        RECT 3376.930 1411.580 3377.250 1411.640 ;
        RECT 3374.170 1411.440 3377.250 1411.580 ;
        RECT 3374.170 1411.380 3374.490 1411.440 ;
        RECT 3376.930 1411.380 3377.250 1411.440 ;
        RECT 208.910 1410.560 209.230 1410.620 ;
        RECT 212.590 1410.560 212.910 1410.620 ;
        RECT 208.910 1410.420 212.910 1410.560 ;
        RECT 208.910 1410.360 209.230 1410.420 ;
        RECT 212.590 1410.360 212.910 1410.420 ;
        RECT 3376.010 1406.140 3376.330 1406.200 ;
        RECT 3376.930 1406.140 3377.250 1406.200 ;
        RECT 3376.010 1406.000 3377.250 1406.140 ;
        RECT 3376.010 1405.940 3376.330 1406.000 ;
        RECT 3376.930 1405.940 3377.250 1406.000 ;
      LAYER met1 ;
        RECT 3381.155 1402.000 3588.000 1482.000 ;
        RECT 3407.485 1401.885 3413.015 1402.000 ;
        RECT 3418.120 1401.885 3423.725 1402.000 ;
        RECT 3439.220 1401.940 3482.580 1402.000 ;
        RECT 3439.220 1401.885 3460.930 1401.940 ;
        POLYGON 3460.930 1401.940 3460.985 1401.940 3460.930 1401.885 ;
        RECT 3483.895 1401.855 3518.220 1402.000 ;
        RECT 3519.275 1401.855 3558.090 1402.000 ;
        RECT 3566.900 1401.980 3568.975 1402.000 ;
      LAYER met1 ;
        RECT 208.910 1380.980 209.230 1381.040 ;
        RECT 212.130 1380.980 212.450 1381.040 ;
        RECT 208.910 1380.840 212.450 1380.980 ;
        RECT 208.910 1380.780 209.230 1380.840 ;
        RECT 212.130 1380.780 212.450 1380.840 ;
        RECT 208.910 1369.760 209.230 1369.820 ;
        RECT 213.050 1369.760 213.370 1369.820 ;
        RECT 208.910 1369.620 213.370 1369.760 ;
        RECT 208.910 1369.560 209.230 1369.620 ;
        RECT 213.050 1369.560 213.370 1369.620 ;
      LAYER met1 ;
        RECT 29.910 1339.885 68.725 1340.000 ;
        RECT 69.780 1339.885 104.105 1340.000 ;
        RECT 108.520 1339.855 110.250 1340.000 ;
        RECT 119.365 1339.885 142.810 1340.000 ;
        RECT 3445.190 1257.000 3468.635 1257.115 ;
        RECT 3477.750 1257.000 3479.480 1257.145 ;
        RECT 3483.895 1257.000 3518.220 1257.115 ;
        RECT 3519.275 1257.000 3558.090 1257.115 ;
      LAYER met1 ;
        RECT 3375.090 1237.500 3375.410 1237.560 ;
        RECT 3376.930 1237.500 3377.250 1237.560 ;
        RECT 3375.090 1237.360 3377.250 1237.500 ;
        RECT 3375.090 1237.300 3375.410 1237.360 ;
        RECT 3376.930 1237.300 3377.250 1237.360 ;
        RECT 3374.630 1222.540 3374.950 1222.600 ;
        RECT 3376.930 1222.540 3377.250 1222.600 ;
        RECT 3374.630 1222.400 3377.250 1222.540 ;
        RECT 3374.630 1222.340 3374.950 1222.400 ;
        RECT 3376.930 1222.340 3377.250 1222.400 ;
      LAYER met1 ;
        RECT 19.025 1204.000 21.100 1204.020 ;
        RECT 29.910 1204.000 68.725 1204.145 ;
        RECT 69.780 1204.000 104.105 1204.145 ;
        POLYGON 127.070 1204.115 127.070 1204.060 127.015 1204.060 ;
        RECT 127.070 1204.060 148.780 1204.115 ;
        RECT 105.420 1204.000 148.780 1204.060 ;
        RECT 164.275 1204.000 169.880 1204.115 ;
        RECT 174.985 1204.000 180.515 1204.115 ;
        RECT 0.000 1124.000 206.845 1204.000 ;
      LAYER met1 ;
        RECT 208.910 1199.760 209.230 1199.820 ;
        RECT 212.130 1199.760 212.450 1199.820 ;
        RECT 208.910 1199.620 212.450 1199.760 ;
        RECT 208.910 1199.560 209.230 1199.620 ;
        RECT 212.130 1199.560 212.450 1199.620 ;
        RECT 208.910 1192.620 209.230 1192.680 ;
        RECT 212.590 1192.620 212.910 1192.680 ;
        RECT 208.910 1192.480 212.910 1192.620 ;
        RECT 208.910 1192.420 209.230 1192.480 ;
        RECT 212.590 1192.420 212.910 1192.480 ;
        RECT 3374.170 1188.540 3374.490 1188.600 ;
        RECT 3376.930 1188.540 3377.250 1188.600 ;
        RECT 3374.170 1188.400 3377.250 1188.540 ;
        RECT 3374.170 1188.340 3374.490 1188.400 ;
        RECT 3376.930 1188.340 3377.250 1188.400 ;
        RECT 3376.010 1181.400 3376.330 1181.460 ;
        RECT 3376.930 1181.400 3377.250 1181.460 ;
        RECT 3376.010 1181.260 3377.250 1181.400 ;
        RECT 3376.010 1181.200 3376.330 1181.260 ;
        RECT 3376.930 1181.200 3377.250 1181.260 ;
      LAYER met1 ;
        RECT 3381.155 1177.000 3588.000 1257.000 ;
        RECT 3407.485 1176.885 3413.015 1177.000 ;
        RECT 3418.120 1176.885 3423.725 1177.000 ;
        RECT 3439.220 1176.940 3482.580 1177.000 ;
        RECT 3439.220 1176.885 3460.930 1176.940 ;
        POLYGON 3460.930 1176.940 3460.985 1176.940 3460.930 1176.885 ;
        RECT 3483.895 1176.855 3518.220 1177.000 ;
        RECT 3519.275 1176.855 3558.090 1177.000 ;
        RECT 3566.900 1176.980 3568.975 1177.000 ;
      LAYER met1 ;
        RECT 208.910 1165.080 209.230 1165.140 ;
        RECT 212.130 1165.080 212.450 1165.140 ;
        RECT 208.910 1164.940 212.450 1165.080 ;
        RECT 208.910 1164.880 209.230 1164.940 ;
        RECT 212.130 1164.880 212.450 1164.940 ;
        RECT 208.910 1158.620 209.230 1158.680 ;
        RECT 213.050 1158.620 213.370 1158.680 ;
        RECT 208.910 1158.480 213.370 1158.620 ;
        RECT 208.910 1158.420 209.230 1158.480 ;
        RECT 213.050 1158.420 213.370 1158.480 ;
      LAYER met1 ;
        RECT 29.910 1123.885 68.725 1124.000 ;
        RECT 69.780 1123.885 104.105 1124.000 ;
        RECT 108.520 1123.855 110.250 1124.000 ;
        RECT 119.365 1123.885 142.810 1124.000 ;
        RECT 3445.190 1031.000 3468.635 1031.115 ;
        RECT 3477.750 1031.000 3479.480 1031.145 ;
        RECT 3483.895 1031.000 3518.220 1031.115 ;
        RECT 3519.275 1031.000 3558.090 1031.115 ;
      LAYER met1 ;
        RECT 3375.090 1011.740 3375.410 1011.800 ;
        RECT 3376.930 1011.740 3377.250 1011.800 ;
        RECT 3375.090 1011.600 3377.250 1011.740 ;
        RECT 3375.090 1011.540 3375.410 1011.600 ;
        RECT 3376.930 1011.540 3377.250 1011.600 ;
        RECT 3374.630 1001.200 3374.950 1001.260 ;
        RECT 3376.930 1001.200 3377.250 1001.260 ;
        RECT 3374.630 1001.060 3377.250 1001.200 ;
        RECT 3374.630 1001.000 3374.950 1001.060 ;
        RECT 3376.930 1001.000 3377.250 1001.060 ;
        RECT 3376.010 996.240 3376.330 996.500 ;
        RECT 3376.100 995.480 3376.240 996.240 ;
        RECT 3376.010 995.220 3376.330 995.480 ;
      LAYER met1 ;
        RECT 19.025 988.000 21.100 988.020 ;
        RECT 29.910 988.000 68.725 988.145 ;
        RECT 69.780 988.000 104.105 988.145 ;
        POLYGON 127.070 988.115 127.070 988.060 127.015 988.060 ;
        RECT 127.070 988.060 148.780 988.115 ;
        RECT 105.420 988.000 148.780 988.060 ;
        RECT 164.275 988.000 169.880 988.115 ;
        RECT 174.985 988.000 180.515 988.115 ;
        RECT 0.000 908.000 206.845 988.000 ;
      LAYER met1 ;
        RECT 208.910 983.860 209.230 983.920 ;
        RECT 213.510 983.860 213.830 983.920 ;
        RECT 208.910 983.720 213.830 983.860 ;
        RECT 208.910 983.660 209.230 983.720 ;
        RECT 213.510 983.660 213.830 983.720 ;
        RECT 208.910 976.720 209.230 976.780 ;
        RECT 212.130 976.720 212.450 976.780 ;
        RECT 208.910 976.580 212.450 976.720 ;
        RECT 208.910 976.520 209.230 976.580 ;
        RECT 212.130 976.520 212.450 976.580 ;
        RECT 3376.010 959.720 3376.330 959.780 ;
        RECT 3376.930 959.720 3377.250 959.780 ;
        RECT 3376.010 959.580 3377.250 959.720 ;
        RECT 3376.010 959.520 3376.330 959.580 ;
        RECT 3376.930 959.520 3377.250 959.580 ;
      LAYER met1 ;
        RECT 3381.155 951.000 3588.000 1031.000 ;
        RECT 3407.485 950.885 3413.015 951.000 ;
        RECT 3418.120 950.885 3423.725 951.000 ;
        RECT 3439.220 950.940 3482.580 951.000 ;
        RECT 3439.220 950.885 3460.930 950.940 ;
        POLYGON 3460.930 950.940 3460.985 950.940 3460.930 950.885 ;
        RECT 3483.895 950.855 3518.220 951.000 ;
        RECT 3519.275 950.855 3558.090 951.000 ;
        RECT 3566.900 950.980 3568.975 951.000 ;
      LAYER met1 ;
        RECT 208.910 949.180 209.230 949.240 ;
        RECT 213.510 949.180 213.830 949.240 ;
        RECT 208.910 949.040 213.830 949.180 ;
        RECT 208.910 948.980 209.230 949.040 ;
        RECT 213.510 948.980 213.830 949.040 ;
        RECT 208.910 937.960 209.230 938.020 ;
        RECT 212.590 937.960 212.910 938.020 ;
        RECT 208.910 937.820 212.910 937.960 ;
        RECT 208.910 937.760 209.230 937.820 ;
        RECT 212.590 937.760 212.910 937.820 ;
      LAYER met1 ;
        RECT 29.910 907.885 68.725 908.000 ;
        RECT 69.780 907.885 104.105 908.000 ;
        RECT 108.520 907.855 110.250 908.000 ;
        RECT 119.365 907.885 142.810 908.000 ;
        RECT 3445.190 806.000 3468.635 806.115 ;
        RECT 3477.750 806.000 3479.480 806.145 ;
        RECT 3483.895 806.000 3518.220 806.115 ;
        RECT 3519.275 806.000 3558.090 806.115 ;
      LAYER met1 ;
        RECT 3376.470 793.600 3376.790 793.860 ;
        RECT 3375.550 792.780 3375.870 792.840 ;
        RECT 3376.560 792.780 3376.700 793.600 ;
        RECT 3375.550 792.640 3376.700 792.780 ;
        RECT 3375.550 792.580 3375.870 792.640 ;
        RECT 3374.170 786.660 3374.490 786.720 ;
        RECT 3375.090 786.660 3375.410 786.720 ;
        RECT 3376.930 786.660 3377.250 786.720 ;
        RECT 3374.170 786.520 3377.250 786.660 ;
        RECT 3374.170 786.460 3374.490 786.520 ;
        RECT 3375.090 786.460 3375.410 786.520 ;
        RECT 3376.930 786.460 3377.250 786.520 ;
        RECT 3374.630 776.120 3374.950 776.180 ;
        RECT 3376.930 776.120 3377.250 776.180 ;
        RECT 3374.630 775.980 3377.250 776.120 ;
        RECT 3374.630 775.920 3374.950 775.980 ;
        RECT 3376.930 775.920 3377.250 775.980 ;
        RECT 3375.090 735.660 3375.410 735.720 ;
        RECT 3376.010 735.660 3376.330 735.720 ;
        RECT 3376.930 735.660 3377.250 735.720 ;
        RECT 3375.090 735.520 3377.250 735.660 ;
        RECT 3375.090 735.460 3375.410 735.520 ;
        RECT 3376.010 735.460 3376.330 735.520 ;
        RECT 3376.930 735.460 3377.250 735.520 ;
      LAYER met1 ;
        RECT 3381.155 726.000 3588.000 806.000 ;
        RECT 3407.485 725.885 3413.015 726.000 ;
        RECT 3418.120 725.885 3423.725 726.000 ;
        RECT 3439.220 725.940 3482.580 726.000 ;
        RECT 3439.220 725.885 3460.930 725.940 ;
        POLYGON 3460.930 725.940 3460.985 725.940 3460.930 725.885 ;
        RECT 3483.895 725.855 3518.220 726.000 ;
        RECT 3519.275 725.855 3558.090 726.000 ;
        RECT 3566.900 725.980 3568.975 726.000 ;
        RECT 0.275 621.680 197.965 623.915 ;
        RECT 0.275 620.540 199.030 621.680 ;
        RECT 0.275 564.350 197.965 620.540 ;
        POLYGON 197.965 620.540 198.080 620.540 198.080 620.425 ;
        POLYGON 198.080 564.465 198.080 564.350 197.965 564.350 ;
        RECT 198.080 564.350 199.030 620.540 ;
        RECT 3445.190 580.000 3468.635 580.115 ;
        RECT 3477.750 580.000 3479.480 580.145 ;
        RECT 3483.895 580.000 3518.220 580.115 ;
        RECT 3519.275 580.000 3558.090 580.115 ;
        RECT 0.275 563.035 199.030 564.350 ;
        RECT 0.275 559.855 197.965 563.035 ;
      LAYER met1 ;
        RECT 3374.170 562.600 3374.490 562.660 ;
        RECT 3376.930 562.600 3377.250 562.660 ;
        RECT 3374.170 562.460 3377.250 562.600 ;
        RECT 3374.170 562.400 3374.490 562.460 ;
        RECT 3376.930 562.400 3377.250 562.460 ;
      LAYER met1 ;
        RECT 0.275 554.625 198.870 559.855 ;
        RECT 0.275 551.185 197.965 554.625 ;
      LAYER met1 ;
        RECT 3374.630 545.600 3374.950 545.660 ;
        RECT 3376.930 545.600 3377.250 545.660 ;
        RECT 3374.630 545.460 3377.250 545.600 ;
        RECT 3374.630 545.400 3374.950 545.460 ;
        RECT 3376.930 545.400 3377.250 545.460 ;
        RECT 3376.010 539.140 3376.330 539.200 ;
        RECT 3376.930 539.140 3377.250 539.200 ;
        RECT 3376.010 539.000 3377.250 539.140 ;
        RECT 3376.010 538.940 3376.330 539.000 ;
        RECT 3376.930 538.940 3377.250 539.000 ;
        RECT 3376.010 510.040 3376.330 510.300 ;
        RECT 3376.100 509.220 3376.240 510.040 ;
        RECT 3376.470 509.220 3376.790 509.280 ;
        RECT 3376.100 509.080 3376.790 509.220 ;
        RECT 3376.470 509.020 3376.790 509.080 ;
      LAYER met1 ;
        RECT 3381.155 500.000 3588.000 580.000 ;
        RECT 3407.485 499.885 3413.015 500.000 ;
        RECT 3418.120 499.885 3423.725 500.000 ;
        RECT 3439.220 499.940 3482.580 500.000 ;
        RECT 3439.220 499.885 3460.930 499.940 ;
        POLYGON 3460.930 499.940 3460.985 499.940 3460.930 499.885 ;
        RECT 3483.895 499.855 3518.220 500.000 ;
        RECT 3519.275 499.855 3558.090 500.000 ;
        RECT 3566.900 499.980 3568.975 500.000 ;
        RECT 159.640 425.935 163.510 426.195 ;
        RECT 159.640 421.935 204.500 425.935 ;
        POLYGON 204.500 425.935 208.500 421.935 204.500 421.935 ;
        RECT 159.640 416.200 208.500 421.935 ;
        RECT 159.640 415.245 163.510 416.200 ;
        RECT 0.160 396.565 197.965 415.000 ;
        RECT 198.780 396.565 208.500 416.200 ;
        RECT 0.160 360.495 208.500 396.565 ;
        RECT 0.160 356.655 198.000 360.495 ;
        RECT 198.980 358.655 208.500 360.495 ;
        POLYGON 198.980 358.655 200.980 358.655 200.980 356.655 ;
        RECT 200.980 356.655 206.500 358.655 ;
        POLYGON 206.500 358.655 208.500 358.655 206.500 356.655 ;
        RECT 0.160 340.120 197.965 356.655 ;
      LAYER met1 ;
        RECT 210.750 224.640 211.070 224.700 ;
        RECT 738.370 224.640 738.690 224.700 ;
        RECT 210.750 224.500 738.690 224.640 ;
        RECT 210.750 224.440 211.070 224.500 ;
        RECT 738.370 224.440 738.690 224.500 ;
        RECT 2618.850 224.640 2619.170 224.700 ;
        RECT 3374.630 224.640 3374.950 224.700 ;
        RECT 2618.850 224.500 3374.950 224.640 ;
        RECT 2618.850 224.440 2619.170 224.500 ;
        RECT 3374.630 224.440 3374.950 224.500 ;
        RECT 210.290 224.300 210.610 224.360 ;
        RECT 979.870 224.300 980.190 224.360 ;
        RECT 210.290 224.160 980.190 224.300 ;
        RECT 210.290 224.100 210.610 224.160 ;
        RECT 979.870 224.100 980.190 224.160 ;
        RECT 2580.670 224.300 2580.990 224.360 ;
        RECT 3375.550 224.300 3375.870 224.360 ;
        RECT 2580.670 224.160 3375.870 224.300 ;
        RECT 2580.670 224.100 2580.990 224.160 ;
        RECT 3375.550 224.100 3375.870 224.160 ;
        RECT 2298.230 223.960 2298.550 224.020 ;
        RECT 2338.250 223.960 2338.570 224.020 ;
        RECT 2298.230 223.820 2338.570 223.960 ;
        RECT 2298.230 223.760 2298.550 223.820 ;
        RECT 2338.250 223.760 2338.570 223.820 ;
        RECT 2076.510 223.620 2076.830 223.680 ;
        RECT 2339.170 223.620 2339.490 223.680 ;
        RECT 2076.510 223.480 2339.490 223.620 ;
        RECT 2076.510 223.420 2076.830 223.480 ;
        RECT 2339.170 223.420 2339.490 223.480 ;
        RECT 2366.310 223.620 2366.630 223.680 ;
        RECT 2634.030 223.620 2634.350 223.680 ;
        RECT 2366.310 223.480 2634.350 223.620 ;
        RECT 2366.310 223.420 2366.630 223.480 ;
        RECT 2634.030 223.420 2634.350 223.480 ;
        RECT 2307.430 223.280 2307.750 223.340 ;
        RECT 2580.670 223.280 2580.990 223.340 ;
        RECT 2256.230 223.140 2580.990 223.280 ;
        RECT 1476.210 222.940 1476.530 223.000 ;
        RECT 1516.230 222.940 1516.550 223.000 ;
        RECT 1476.210 222.800 1516.550 222.940 ;
        RECT 1476.210 222.740 1476.530 222.800 ;
        RECT 1516.230 222.740 1516.550 222.800 ;
        RECT 1750.370 222.940 1750.690 223.000 ;
        RECT 1790.390 222.940 1790.710 223.000 ;
        RECT 1750.370 222.800 1790.710 222.940 ;
        RECT 1750.370 222.740 1750.690 222.800 ;
        RECT 1790.390 222.740 1790.710 222.800 ;
        RECT 1802.810 222.940 1803.130 223.000 ;
        RECT 2033.730 222.940 2034.050 223.000 ;
        RECT 2256.230 222.940 2256.370 223.140 ;
        RECT 2307.430 223.080 2307.750 223.140 ;
        RECT 2580.670 223.080 2580.990 223.140 ;
        RECT 1802.810 222.800 2256.370 222.940 ;
        RECT 2339.170 222.940 2339.490 223.000 ;
        RECT 2344.690 222.940 2345.010 223.000 ;
        RECT 2618.850 222.940 2619.170 223.000 ;
        RECT 2339.170 222.800 2619.170 222.940 ;
        RECT 1802.810 222.740 1803.130 222.800 ;
        RECT 2033.730 222.740 2034.050 222.800 ;
        RECT 2339.170 222.740 2339.490 222.800 ;
        RECT 2344.690 222.740 2345.010 222.800 ;
        RECT 2618.850 222.740 2619.170 222.800 ;
        RECT 1537.850 222.600 1538.170 222.660 ;
        RECT 1812.010 222.600 1812.330 222.660 ;
        RECT 2086.170 222.600 2086.490 222.660 ;
        RECT 2359.870 222.600 2360.190 222.660 ;
        RECT 2366.310 222.600 2366.630 222.660 ;
        RECT 1000.430 222.460 2366.630 222.600 ;
        RECT 443.970 222.260 444.290 222.320 ;
        RECT 995.050 222.260 995.370 222.320 ;
        RECT 1000.430 222.260 1000.570 222.460 ;
        RECT 1537.850 222.400 1538.170 222.460 ;
        RECT 1812.010 222.400 1812.330 222.460 ;
        RECT 2086.170 222.400 2086.490 222.460 ;
        RECT 2359.870 222.400 2360.190 222.460 ;
        RECT 2366.310 222.400 2366.630 222.460 ;
        RECT 2572.390 222.600 2572.710 222.660 ;
        RECT 2612.410 222.600 2612.730 222.660 ;
        RECT 2572.390 222.460 2612.730 222.600 ;
        RECT 2572.390 222.400 2572.710 222.460 ;
        RECT 2612.410 222.400 2612.730 222.460 ;
        RECT 443.970 222.120 1000.570 222.260 ;
        RECT 1004.250 222.260 1004.570 222.320 ;
        RECT 1206.650 222.260 1206.970 222.320 ;
        RECT 1488.630 222.260 1488.950 222.320 ;
        RECT 1503.810 222.260 1504.130 222.320 ;
        RECT 1525.430 222.260 1525.750 222.320 ;
        RECT 1004.250 222.120 1525.750 222.260 ;
        RECT 443.970 222.060 444.290 222.120 ;
        RECT 995.050 222.060 995.370 222.120 ;
        RECT 1004.250 222.060 1004.570 222.120 ;
        RECT 1206.650 222.060 1206.970 222.120 ;
        RECT 1488.630 222.060 1488.950 222.120 ;
        RECT 1503.810 222.060 1504.130 222.120 ;
        RECT 1525.430 222.060 1525.750 222.120 ;
        RECT 1547.050 222.260 1547.370 222.320 ;
        RECT 1762.790 222.260 1763.110 222.320 ;
        RECT 1777.970 222.260 1778.290 222.320 ;
        RECT 1799.590 222.260 1799.910 222.320 ;
        RECT 1547.050 222.120 1799.910 222.260 ;
        RECT 1547.050 222.060 1547.370 222.120 ;
        RECT 1762.790 222.060 1763.110 222.120 ;
        RECT 1777.970 222.060 1778.290 222.120 ;
        RECT 1799.590 222.060 1799.910 222.120 ;
        RECT 1821.210 222.260 1821.530 222.320 ;
        RECT 2036.950 222.260 2037.270 222.320 ;
        RECT 2052.130 222.260 2052.450 222.320 ;
        RECT 1821.210 222.120 2052.450 222.260 ;
        RECT 1821.210 222.060 1821.530 222.120 ;
        RECT 2036.950 222.060 2037.270 222.120 ;
        RECT 2052.130 222.060 2052.450 222.120 ;
        RECT 2080.190 222.260 2080.510 222.320 ;
        RECT 2095.370 222.260 2095.690 222.320 ;
        RECT 2310.650 222.260 2310.970 222.320 ;
        RECT 2325.830 222.260 2326.150 222.320 ;
        RECT 2080.190 222.120 2326.150 222.260 ;
        RECT 2080.190 222.060 2080.510 222.120 ;
        RECT 2095.370 222.060 2095.690 222.120 ;
        RECT 2310.650 222.060 2310.970 222.120 ;
        RECT 2325.830 222.060 2326.150 222.120 ;
        RECT 2353.890 222.260 2354.210 222.320 ;
        RECT 2369.070 222.260 2369.390 222.320 ;
        RECT 2584.810 222.260 2585.130 222.320 ;
        RECT 2599.990 222.260 2600.310 222.320 ;
        RECT 2353.890 222.120 2600.310 222.260 ;
        RECT 2353.890 222.060 2354.210 222.120 ;
        RECT 2369.070 222.060 2369.390 222.120 ;
        RECT 2584.810 222.060 2585.130 222.120 ;
        RECT 2599.990 222.060 2600.310 222.120 ;
        RECT 942.610 221.920 942.930 221.980 ;
        RECT 964.230 221.920 964.550 221.980 ;
        RECT 1007.470 221.920 1007.790 221.980 ;
        RECT 1485.410 221.920 1485.730 221.980 ;
        RECT 1497.830 221.920 1498.150 221.980 ;
        RECT 1528.650 221.920 1528.970 221.980 ;
        RECT 1759.570 221.920 1759.890 221.980 ;
        RECT 1771.990 221.920 1772.310 221.980 ;
        RECT 1802.810 221.920 1803.130 221.980 ;
        RECT 942.610 221.780 1803.130 221.920 ;
        RECT 942.610 221.720 942.930 221.780 ;
        RECT 964.230 221.720 964.550 221.780 ;
        RECT 1007.470 221.720 1007.790 221.780 ;
        RECT 1485.410 221.720 1485.730 221.780 ;
        RECT 1497.830 221.720 1498.150 221.780 ;
        RECT 1528.650 221.720 1528.970 221.780 ;
        RECT 1759.570 221.720 1759.890 221.780 ;
        RECT 1771.990 221.720 1772.310 221.780 ;
        RECT 1802.810 221.720 1803.130 221.780 ;
        RECT 2024.530 221.920 2024.850 221.980 ;
        RECT 2064.550 221.920 2064.870 221.980 ;
        RECT 2024.530 221.780 2064.870 221.920 ;
        RECT 2024.530 221.720 2024.850 221.780 ;
        RECT 2064.550 221.720 2064.870 221.780 ;
        RECT 738.370 221.240 738.690 221.300 ;
        RECT 942.610 221.240 942.930 221.300 ;
        RECT 738.370 221.100 942.930 221.240 ;
        RECT 738.370 221.040 738.690 221.100 ;
        RECT 942.610 221.040 942.930 221.100 ;
        RECT 979.870 221.240 980.190 221.300 ;
        RECT 1522.670 221.240 1522.990 221.300 ;
        RECT 1796.830 221.240 1797.150 221.300 ;
        RECT 2070.990 221.240 2071.310 221.300 ;
        RECT 2076.510 221.240 2076.830 221.300 ;
        RECT 979.870 221.100 2076.830 221.240 ;
        RECT 979.870 221.040 980.190 221.100 ;
        RECT 1522.670 221.040 1522.990 221.100 ;
        RECT 1796.830 221.040 1797.150 221.100 ;
        RECT 2070.990 221.040 2071.310 221.100 ;
        RECT 2076.510 221.040 2076.830 221.100 ;
        RECT 933.410 220.900 933.730 220.960 ;
        RECT 973.430 220.900 973.750 220.960 ;
        RECT 933.410 220.760 973.750 220.900 ;
        RECT 933.410 220.700 933.730 220.760 ;
        RECT 973.430 220.700 973.750 220.760 ;
        RECT 211.210 210.700 211.530 210.760 ;
        RECT 704.790 210.700 705.110 210.760 ;
        RECT 211.210 210.560 705.110 210.700 ;
        RECT 211.210 210.500 211.530 210.560 ;
        RECT 704.790 210.500 705.110 210.560 ;
        RECT 2348.370 210.020 2348.690 210.080 ;
        RECT 2353.430 210.020 2353.750 210.080 ;
        RECT 2348.370 209.880 2353.750 210.020 ;
        RECT 2348.370 209.820 2348.690 209.880 ;
        RECT 2353.430 209.820 2353.750 209.880 ;
        RECT 992.290 209.680 992.610 209.740 ;
        RECT 1000.570 209.680 1000.890 209.740 ;
        RECT 992.290 209.540 1000.890 209.680 ;
        RECT 992.290 209.480 992.610 209.540 ;
        RECT 1000.570 209.480 1000.890 209.540 ;
        RECT 1526.350 209.680 1526.670 209.740 ;
        RECT 1531.410 209.680 1531.730 209.740 ;
        RECT 1543.370 209.680 1543.690 209.740 ;
        RECT 1526.350 209.540 1543.690 209.680 ;
        RECT 1526.350 209.480 1526.670 209.540 ;
        RECT 1531.410 209.480 1531.730 209.540 ;
        RECT 1543.370 209.480 1543.690 209.540 ;
        RECT 946.290 209.000 946.610 209.060 ;
        RECT 955.490 209.000 955.810 209.060 ;
        RECT 961.470 209.000 961.790 209.060 ;
        RECT 967.910 209.000 968.230 209.060 ;
        RECT 982.170 209.000 982.490 209.060 ;
        RECT 946.290 208.860 982.490 209.000 ;
        RECT 946.290 208.800 946.610 208.860 ;
        RECT 955.490 208.800 955.810 208.860 ;
        RECT 961.470 208.800 961.790 208.860 ;
        RECT 967.910 208.800 968.230 208.860 ;
        RECT 982.170 208.800 982.490 208.860 ;
        RECT 1800.050 209.000 1800.370 209.060 ;
        RECT 1805.570 209.000 1805.890 209.060 ;
        RECT 1817.530 209.000 1817.850 209.060 ;
        RECT 1800.050 208.860 1817.850 209.000 ;
        RECT 1800.050 208.800 1800.370 208.860 ;
        RECT 1805.570 208.800 1805.890 208.860 ;
        RECT 1817.530 208.800 1817.850 208.860 ;
        RECT 2052.590 209.000 2052.910 209.060 ;
        RECT 2057.650 209.000 2057.970 209.060 ;
        RECT 2074.210 209.000 2074.530 209.060 ;
        RECT 2079.270 209.000 2079.590 209.060 ;
        RECT 2052.590 208.860 2079.590 209.000 ;
        RECT 2052.590 208.800 2052.910 208.860 ;
        RECT 2057.650 208.800 2057.970 208.860 ;
        RECT 2074.210 208.800 2074.530 208.860 ;
        RECT 2079.270 208.800 2079.590 208.860 ;
        RECT 2326.750 209.000 2327.070 209.060 ;
        RECT 2331.810 209.000 2332.130 209.060 ;
        RECT 2346.990 209.000 2347.310 209.060 ;
        RECT 2326.750 208.860 2347.310 209.000 ;
        RECT 2326.750 208.800 2327.070 208.860 ;
        RECT 2331.810 208.800 2332.130 208.860 ;
        RECT 2346.990 208.800 2347.310 208.860 ;
        RECT 2600.450 209.000 2600.770 209.060 ;
        RECT 2605.970 209.000 2606.290 209.060 ;
        RECT 2621.150 209.000 2621.470 209.060 ;
        RECT 2627.590 209.000 2627.910 209.060 ;
        RECT 2639.550 209.000 2639.870 209.060 ;
        RECT 2600.450 208.860 2639.870 209.000 ;
        RECT 2600.450 208.800 2600.770 208.860 ;
        RECT 2605.970 208.800 2606.290 208.860 ;
        RECT 2621.150 208.800 2621.470 208.860 ;
        RECT 2627.590 208.800 2627.910 208.860 ;
        RECT 2639.550 208.800 2639.870 208.860 ;
      LAYER met1 ;
        POLYGON 1199.065 208.500 1199.065 207.360 1197.925 207.360 ;
        RECT 1199.065 207.360 1262.345 208.500 ;
      LAYER met1 ;
        RECT 715.370 207.300 715.690 207.360 ;
      LAYER met1 ;
        POLYGON 1197.925 207.360 1197.925 207.300 1197.865 207.300 ;
        RECT 1197.925 207.300 1262.345 207.360 ;
      LAYER met1 ;
        RECT 715.370 207.160 723.420 207.300 ;
        RECT 715.370 207.100 715.690 207.160 ;
        RECT 723.280 207.020 723.420 207.160 ;
        RECT 931.430 207.160 1012.760 207.300 ;
        RECT 723.190 206.960 723.510 207.020 ;
        RECT 931.430 206.960 931.570 207.160 ;
        RECT 723.190 206.820 931.570 206.960 ;
        RECT 1012.620 206.960 1012.760 207.160 ;
      LAYER met1 ;
        POLYGON 1197.865 207.300 1197.865 206.960 1197.525 206.960 ;
        RECT 1197.865 206.960 1262.345 207.300 ;
        POLYGON 1262.345 208.500 1263.885 206.960 1262.345 206.960 ;
      LAYER met1 ;
        RECT 1474.460 207.160 1555.560 207.300 ;
        RECT 1474.460 206.960 1474.600 207.160 ;
        RECT 723.190 206.760 723.510 206.820 ;
        RECT 704.950 200.500 705.270 200.560 ;
        RECT 715.370 200.500 715.690 200.560 ;
        RECT 704.950 200.360 715.690 200.500 ;
        RECT 704.950 200.300 705.270 200.360 ;
        RECT 712.930 200.000 713.070 200.360 ;
        RECT 715.370 200.300 715.690 200.360 ;
      LAYER met1 ;
        RECT 663.000 199.390 704.700 199.815 ;
      LAYER met1 ;
        RECT 704.980 199.670 705.240 200.000 ;
      LAYER met1 ;
        RECT 705.520 199.390 706.565 199.815 ;
      LAYER met1 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met1 ;
        RECT 707.775 199.390 709.490 199.815 ;
      LAYER met1 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met1 ;
        RECT 710.700 199.390 712.585 199.815 ;
        RECT 398.320 198.080 456.965 199.030 ;
        RECT 398.320 197.965 399.460 198.080 ;
        POLYGON 399.460 198.080 399.575 198.080 399.460 197.965 ;
        POLYGON 455.535 198.080 455.650 198.080 455.650 197.965 ;
        RECT 455.650 197.965 456.965 198.080 ;
        RECT 395.380 0.275 468.815 197.965 ;
        RECT 663.000 189.745 712.585 199.390 ;
      LAYER met1 ;
        RECT 712.865 190.025 713.095 200.000 ;
      LAYER met1 ;
        RECT 713.375 199.390 715.060 199.815 ;
      LAYER met1 ;
        RECT 715.340 199.670 715.640 200.000 ;
      LAYER met1 ;
        RECT 715.920 199.390 722.585 199.815 ;
      LAYER met1 ;
        RECT 722.865 199.670 723.445 200.000 ;
      LAYER met1 ;
        RECT 723.725 199.390 725.175 199.815 ;
      LAYER met1 ;
        RECT 725.455 199.670 725.715 200.000 ;
      LAYER met1 ;
        RECT 725.995 199.390 738.000 199.815 ;
        RECT 713.375 189.745 738.000 199.390 ;
        RECT 663.000 104.105 738.000 189.745 ;
        RECT 932.000 180.515 1012.000 206.845 ;
      LAYER met1 ;
        RECT 1012.620 206.820 1197.385 206.960 ;
        POLYGON 1197.385 206.960 1197.525 206.960 1197.385 206.820 ;
      LAYER met1 ;
        RECT 1197.525 206.820 1263.885 206.960 ;
        POLYGON 1263.885 206.960 1264.025 206.820 1263.885 206.820 ;
      LAYER met1 ;
        RECT 1264.025 206.820 1474.600 206.960 ;
        RECT 1555.420 206.960 1555.560 207.160 ;
        RECT 1748.160 207.160 1829.720 207.300 ;
        RECT 1748.160 206.960 1748.300 207.160 ;
      LAYER met1 ;
        RECT 931.885 174.985 1012.000 180.515 ;
        RECT 932.000 169.880 1012.000 174.985 ;
        RECT 931.885 164.275 1012.000 169.880 ;
        RECT 932.000 148.780 1012.000 164.275 ;
        POLYGON 1197.385 206.820 1197.385 204.500 1195.065 204.500 ;
        RECT 1197.385 206.500 1264.025 206.820 ;
        POLYGON 1264.025 206.820 1264.345 206.500 1264.025 206.500 ;
        RECT 1197.385 204.500 1264.345 206.500 ;
        RECT 1195.065 200.980 1264.345 204.500 ;
        RECT 1195.065 198.980 1262.345 200.980 ;
        POLYGON 1262.345 200.980 1264.345 200.980 1262.345 198.980 ;
        RECT 1195.065 198.780 1260.505 198.980 ;
        RECT 1195.065 163.510 1204.800 198.780 ;
        RECT 1224.435 198.000 1260.505 198.780 ;
        RECT 1224.435 197.965 1264.345 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 931.885 142.810 1012.000 148.780 ;
        RECT 931.885 127.070 1012.115 142.810 ;
        POLYGON 931.885 127.070 931.940 127.070 931.940 127.015 ;
        RECT 931.940 119.365 1012.115 127.070 ;
        RECT 931.940 110.250 1012.000 119.365 ;
        RECT 931.940 108.520 1012.145 110.250 ;
        RECT 931.940 105.420 1012.000 108.520 ;
        RECT 932.000 104.105 1012.000 105.420 ;
        RECT 662.855 69.780 738.145 104.105 ;
        RECT 931.855 69.780 1012.115 104.105 ;
        RECT 663.000 68.725 738.000 69.780 ;
        RECT 932.000 68.725 1012.000 69.780 ;
        RECT 662.855 29.910 738.145 68.725 ;
        RECT 931.855 29.910 1012.115 68.725 ;
        RECT 663.000 0.790 738.000 29.910 ;
        RECT 932.000 21.100 1012.000 29.910 ;
        RECT 931.980 19.025 1012.000 21.100 ;
        RECT 932.000 0.000 1012.000 19.025 ;
        RECT 1206.000 0.160 1280.880 197.965 ;
        RECT 1475.000 180.515 1555.000 206.845 ;
      LAYER met1 ;
        RECT 1555.420 206.820 1748.300 206.960 ;
        RECT 1829.580 206.960 1829.720 207.160 ;
        RECT 2022.320 207.160 2103.880 207.300 ;
        RECT 2022.320 206.960 2022.460 207.160 ;
      LAYER met1 ;
        RECT 1749.000 180.515 1829.000 206.845 ;
      LAYER met1 ;
        RECT 1829.580 206.820 2022.460 206.960 ;
        RECT 2103.740 206.960 2103.880 207.160 ;
        RECT 2296.480 207.160 2377.580 207.300 ;
        RECT 2296.480 206.960 2296.620 207.160 ;
      LAYER met1 ;
        RECT 2023.000 180.515 2103.000 206.845 ;
      LAYER met1 ;
        RECT 2103.740 206.820 2296.620 206.960 ;
        RECT 2377.440 206.960 2377.580 207.160 ;
        RECT 2570.180 207.160 2651.740 207.300 ;
        RECT 2570.180 206.960 2570.320 207.160 ;
      LAYER met1 ;
        RECT 2297.000 180.515 2377.000 206.845 ;
      LAYER met1 ;
        RECT 2377.440 206.820 2570.320 206.960 ;
        RECT 2651.600 206.960 2651.740 207.160 ;
        RECT 2863.570 206.960 2863.890 207.020 ;
      LAYER met1 ;
        RECT 2571.000 180.515 2651.000 206.845 ;
      LAYER met1 ;
        RECT 2651.600 206.820 2863.890 206.960 ;
        RECT 2863.570 206.760 2863.890 206.820 ;
        RECT 2863.570 203.560 2863.890 203.620 ;
        RECT 3374.170 203.560 3374.490 203.620 ;
        RECT 2863.570 203.420 3374.490 203.560 ;
        RECT 2863.570 203.360 2863.890 203.420 ;
        RECT 3374.170 203.360 3374.490 203.420 ;
      LAYER met1 ;
        RECT 2849.320 198.080 2907.965 199.030 ;
        RECT 2849.320 197.965 2850.460 198.080 ;
        POLYGON 2850.460 198.080 2850.575 198.080 2850.460 197.965 ;
        POLYGON 2906.535 198.080 2906.650 198.080 2906.650 197.965 ;
        RECT 2906.650 197.965 2907.965 198.080 ;
        RECT 3118.320 198.080 3176.965 199.030 ;
        RECT 3118.320 197.965 3119.460 198.080 ;
        POLYGON 3119.460 198.080 3119.575 198.080 3119.460 197.965 ;
        POLYGON 3175.535 198.080 3175.650 198.080 3175.650 197.965 ;
        RECT 3175.650 197.965 3176.965 198.080 ;
        RECT 3180.145 197.965 3185.375 198.870 ;
        RECT 1474.885 174.985 1555.000 180.515 ;
        RECT 1748.885 174.985 1829.000 180.515 ;
        RECT 2022.885 174.985 2103.000 180.515 ;
        RECT 2296.885 174.985 2377.000 180.515 ;
        RECT 2570.885 174.985 2651.000 180.515 ;
        RECT 1475.000 169.880 1555.000 174.985 ;
        RECT 1749.000 169.880 1829.000 174.985 ;
        RECT 2023.000 169.880 2103.000 174.985 ;
        RECT 2297.000 169.880 2377.000 174.985 ;
        RECT 2571.000 169.880 2651.000 174.985 ;
        RECT 1474.885 164.275 1555.000 169.880 ;
        RECT 1748.885 164.275 1829.000 169.880 ;
        RECT 2022.885 164.275 2103.000 169.880 ;
        RECT 2296.885 164.275 2377.000 169.880 ;
        RECT 2570.885 164.275 2651.000 169.880 ;
        RECT 1475.000 148.780 1555.000 164.275 ;
        RECT 1749.000 148.780 1829.000 164.275 ;
        RECT 2023.000 148.780 2103.000 164.275 ;
        RECT 2297.000 148.780 2377.000 164.275 ;
        RECT 2571.000 148.780 2651.000 164.275 ;
        RECT 1474.885 142.810 1555.000 148.780 ;
        RECT 1748.885 142.810 1829.000 148.780 ;
        RECT 2022.885 142.810 2103.000 148.780 ;
        RECT 2296.885 142.810 2377.000 148.780 ;
        RECT 2570.885 142.810 2651.000 148.780 ;
        RECT 1474.885 127.070 1555.115 142.810 ;
        POLYGON 1474.885 127.070 1474.940 127.070 1474.940 127.015 ;
        RECT 1474.940 119.365 1555.115 127.070 ;
        RECT 1748.885 127.070 1829.115 142.810 ;
        POLYGON 1748.885 127.070 1748.940 127.070 1748.940 127.015 ;
        RECT 1748.940 119.365 1829.115 127.070 ;
        RECT 2022.885 127.070 2103.115 142.810 ;
        POLYGON 2022.885 127.070 2022.940 127.070 2022.940 127.015 ;
        RECT 2022.940 119.365 2103.115 127.070 ;
        RECT 2296.885 127.070 2377.115 142.810 ;
        POLYGON 2296.885 127.070 2296.940 127.070 2296.940 127.015 ;
        RECT 2296.940 119.365 2377.115 127.070 ;
        RECT 2570.885 127.070 2651.115 142.810 ;
        POLYGON 2570.885 127.070 2570.940 127.070 2570.940 127.015 ;
        RECT 2570.940 119.365 2651.115 127.070 ;
        RECT 1474.940 110.250 1555.000 119.365 ;
        RECT 1748.940 110.250 1829.000 119.365 ;
        RECT 2022.940 110.250 2103.000 119.365 ;
        RECT 2296.940 110.250 2377.000 119.365 ;
        RECT 2570.940 110.250 2651.000 119.365 ;
        RECT 1474.940 108.520 1555.145 110.250 ;
        RECT 1748.940 108.520 1829.145 110.250 ;
        RECT 2022.940 108.520 2103.145 110.250 ;
        RECT 2296.940 108.520 2377.145 110.250 ;
        RECT 2570.940 108.520 2651.145 110.250 ;
        RECT 1474.940 105.420 1555.000 108.520 ;
        RECT 1748.940 105.420 1829.000 108.520 ;
        RECT 2022.940 105.420 2103.000 108.520 ;
        RECT 2296.940 105.420 2377.000 108.520 ;
        RECT 2570.940 105.420 2651.000 108.520 ;
        RECT 1475.000 104.105 1555.000 105.420 ;
        RECT 1749.000 104.105 1829.000 105.420 ;
        RECT 2023.000 104.105 2103.000 105.420 ;
        RECT 2297.000 104.105 2377.000 105.420 ;
        RECT 2571.000 104.105 2651.000 105.420 ;
        RECT 1474.855 69.780 1555.115 104.105 ;
        RECT 1748.855 69.780 1829.115 104.105 ;
        RECT 2022.855 69.780 2103.115 104.105 ;
        RECT 2296.855 69.780 2377.115 104.105 ;
        RECT 2570.855 69.780 2651.115 104.105 ;
        RECT 1475.000 68.725 1555.000 69.780 ;
        RECT 1749.000 68.725 1829.000 69.780 ;
        RECT 2023.000 68.725 2103.000 69.780 ;
        RECT 2297.000 68.725 2377.000 69.780 ;
        RECT 2571.000 68.725 2651.000 69.780 ;
        RECT 1474.855 29.910 1555.115 68.725 ;
        RECT 1748.855 29.910 1829.115 68.725 ;
        RECT 2022.855 29.910 2103.115 68.725 ;
        RECT 2296.855 29.910 2377.115 68.725 ;
        RECT 2570.855 29.910 2651.115 68.725 ;
        RECT 1475.000 21.100 1555.000 29.910 ;
        RECT 1749.000 21.100 1829.000 29.910 ;
        RECT 2023.000 21.100 2103.000 29.910 ;
        RECT 2297.000 21.100 2377.000 29.910 ;
        RECT 2571.000 21.100 2651.000 29.910 ;
        RECT 1474.980 19.025 1555.000 21.100 ;
        RECT 1748.980 19.025 1829.000 21.100 ;
        RECT 2022.980 19.025 2103.000 21.100 ;
        RECT 2296.980 19.025 2377.000 21.100 ;
        RECT 2570.980 19.025 2651.000 21.100 ;
        RECT 1475.000 0.000 1555.000 19.025 ;
        RECT 1749.000 0.000 1829.000 19.025 ;
        RECT 2023.000 0.000 2103.000 19.025 ;
        RECT 2297.000 0.000 2377.000 19.025 ;
        RECT 2571.000 0.000 2651.000 19.025 ;
        RECT 2846.380 0.275 2919.815 197.965 ;
        RECT 3116.085 0.275 3188.815 197.965 ;
      LAYER via ;
        RECT 2690.640 4976.280 2690.900 4976.540 ;
        RECT 2699.380 4976.280 2699.640 4976.540 ;
        RECT 710.340 4974.920 710.600 4975.180 ;
        RECT 716.320 4974.920 716.580 4975.180 ;
        RECT 416.400 4967.780 416.660 4968.040 ;
        RECT 669.860 4967.780 670.120 4968.040 ;
        RECT 675.840 4967.780 676.100 4968.040 ;
        RECT 676.300 4967.780 676.560 4968.040 ;
        RECT 710.340 4967.780 710.600 4968.040 ;
        RECT 933.440 4967.780 933.700 4968.040 ;
        RECT 973.460 4967.780 973.720 4968.040 ;
        RECT 1168.500 4967.780 1168.760 4968.040 ;
        RECT 1187.360 4967.780 1187.620 4968.040 ;
        RECT 397.540 4967.440 397.800 4967.700 ;
        RECT 654.680 4967.440 654.940 4967.700 ;
        RECT 911.820 4967.440 912.080 4967.700 ;
        RECT 917.340 4967.440 917.600 4967.700 ;
        RECT 927.000 4967.440 927.260 4967.700 ;
        RECT 1183.680 4967.440 1183.940 4967.700 ;
        RECT 1441.740 4967.780 1442.000 4968.040 ;
        RECT 1448.180 4967.780 1448.440 4968.040 ;
        RECT 1488.200 4967.780 1488.460 4968.040 ;
        RECT 449.980 4967.100 450.240 4967.360 ;
        RECT 707.120 4967.100 707.380 4967.360 ;
        RECT 964.260 4967.100 964.520 4967.360 ;
        RECT 1220.940 4967.100 1221.200 4967.360 ;
        RECT 1479.000 4967.440 1479.260 4967.700 ;
        RECT 1957.400 4967.780 1957.660 4968.040 ;
        RECT 1997.420 4967.780 1997.680 4968.040 ;
        RECT 2402.220 4967.780 2402.480 4968.040 ;
        RECT 2442.240 4967.780 2442.500 4968.040 ;
        RECT 2659.360 4967.780 2659.620 4968.040 ;
        RECT 2690.640 4967.780 2690.900 4968.040 ;
        RECT 3168.120 4967.780 3168.380 4968.040 ;
        RECT 3208.140 4967.780 3208.400 4968.040 ;
        RECT 1988.220 4967.440 1988.480 4967.700 ;
        RECT 2433.040 4967.440 2433.300 4967.700 ;
        RECT 2690.180 4967.440 2690.440 4967.700 ;
        RECT 3198.940 4967.440 3199.200 4967.700 ;
        RECT 1187.360 4966.760 1187.620 4967.020 ;
        RECT 1426.560 4966.760 1426.820 4967.020 ;
        RECT 1666.220 4966.760 1666.480 4967.020 ;
        RECT 1935.780 4966.760 1936.040 4967.020 ;
        RECT 2380.600 4967.100 2380.860 4967.360 ;
        RECT 2637.740 4967.100 2638.000 4967.360 ;
        RECT 2641.420 4967.100 2641.680 4967.360 ;
        RECT 2656.140 4967.100 2656.400 4967.360 ;
        RECT 3161.680 4967.100 3161.940 4967.360 ;
        RECT 419.160 4966.420 419.420 4966.680 ;
        RECT 459.180 4966.420 459.440 4966.680 ;
        RECT 917.340 4966.420 917.600 4966.680 ;
        RECT 1168.500 4966.420 1168.760 4966.680 ;
        RECT 675.840 4966.080 676.100 4966.340 ;
        RECT 927.000 4966.080 927.260 4966.340 ;
        RECT 1190.120 4966.080 1190.380 4966.340 ;
        RECT 1230.140 4966.080 1230.400 4966.340 ;
        RECT 1441.740 4966.080 1442.000 4966.340 ;
        RECT 1950.960 4966.420 1951.220 4966.680 ;
        RECT 2395.780 4966.420 2396.040 4966.680 ;
        RECT 2641.420 4966.420 2641.680 4966.680 ;
        RECT 3146.500 4966.420 3146.760 4966.680 ;
        RECT 2652.920 4966.080 2653.180 4966.340 ;
        RECT 2656.140 4966.080 2656.400 4966.340 ;
        RECT 3198.940 4965.400 3199.200 4965.660 ;
        RECT 3370.980 4965.400 3371.240 4965.660 ;
        RECT 217.220 4965.060 217.480 4965.320 ;
        RECT 397.540 4965.060 397.800 4965.320 ;
        RECT 3161.680 4965.060 3161.940 4965.320 ;
        RECT 3371.440 4965.060 3371.700 4965.320 ;
        RECT 217.680 4964.720 217.940 4964.980 ;
        RECT 412.720 4964.720 412.980 4964.980 ;
        RECT 416.400 4964.720 416.660 4964.980 ;
        RECT 211.700 4964.380 211.960 4964.640 ;
        RECT 449.980 4964.380 450.240 4964.640 ;
        RECT 3146.500 4964.380 3146.760 4964.640 ;
        RECT 3375.580 4964.380 3375.840 4964.640 ;
        RECT 2902.700 4950.440 2902.960 4950.700 ;
        RECT 3370.520 4950.440 3370.780 4950.700 ;
        RECT 208.940 4839.600 209.200 4839.860 ;
        RECT 212.160 4839.600 212.420 4839.860 ;
        RECT 3371.440 4820.560 3371.700 4820.820 ;
        RECT 3376.500 4820.560 3376.760 4820.820 ;
        RECT 3374.660 4803.220 3374.920 4803.480 ;
        RECT 3376.960 4803.220 3377.220 4803.480 ;
        RECT 3376.040 4800.840 3376.300 4801.100 ;
        RECT 3376.040 4799.820 3376.300 4800.080 ;
        RECT 211.240 4795.060 211.500 4795.320 ;
        RECT 213.080 4795.060 213.340 4795.320 ;
        RECT 217.680 4795.060 217.940 4795.320 ;
        RECT 208.940 4788.260 209.200 4788.520 ;
        RECT 217.220 4788.260 217.480 4788.520 ;
        RECT 212.160 4787.240 212.420 4787.500 ;
        RECT 212.160 4786.220 212.420 4786.480 ;
        RECT 3370.980 4766.500 3371.240 4766.760 ;
        RECT 3375.580 4766.500 3375.840 4766.760 ;
        RECT 3377.880 4766.500 3378.140 4766.760 ;
        RECT 3374.200 4372.440 3374.460 4372.700 ;
        RECT 3376.040 4372.440 3376.300 4372.700 ;
        RECT 3376.960 4372.440 3377.220 4372.700 ;
        RECT 3375.120 4358.160 3375.380 4358.420 ;
        RECT 3376.960 4358.160 3377.220 4358.420 ;
        RECT 3374.660 4320.420 3374.920 4320.680 ;
        RECT 3375.580 4320.420 3375.840 4320.680 ;
        RECT 3376.960 4320.420 3377.220 4320.680 ;
        RECT 3376.500 4091.600 3376.760 4091.860 ;
        RECT 3387.540 4091.600 3387.800 4091.860 ;
        RECT 208.940 3997.760 209.200 3998.020 ;
        RECT 211.700 3997.760 211.960 3998.020 ;
        RECT 208.940 3988.580 209.200 3988.840 ;
        RECT 212.160 3988.580 212.420 3988.840 ;
        RECT 213.080 3988.580 213.340 3988.840 ;
        RECT 208.940 3962.740 209.200 3963.000 ;
        RECT 211.700 3962.740 211.960 3963.000 ;
        RECT 208.940 3936.220 209.200 3936.480 ;
        RECT 212.620 3936.220 212.880 3936.480 ;
        RECT 3374.200 3926.360 3374.460 3926.620 ;
        RECT 3376.960 3926.360 3377.220 3926.620 ;
        RECT 3375.120 3916.160 3375.380 3916.420 ;
        RECT 3376.960 3916.160 3377.220 3916.420 ;
        RECT 3376.040 3904.940 3376.300 3905.200 ;
        RECT 3376.960 3904.940 3377.220 3905.200 ;
        RECT 3374.660 3875.020 3374.920 3875.280 ;
        RECT 3376.960 3875.020 3377.220 3875.280 ;
        RECT 3376.040 3869.920 3376.300 3870.180 ;
        RECT 3376.960 3869.920 3377.220 3870.180 ;
        RECT 208.940 3781.860 209.200 3782.120 ;
        RECT 213.540 3781.860 213.800 3782.120 ;
        RECT 208.940 3776.760 209.200 3777.020 ;
        RECT 212.160 3776.760 212.420 3777.020 ;
        RECT 213.080 3776.760 213.340 3777.020 ;
        RECT 208.940 3746.840 209.200 3747.100 ;
        RECT 213.540 3746.840 213.800 3747.100 ;
        RECT 208.940 3725.420 209.200 3725.680 ;
        RECT 212.620 3725.420 212.880 3725.680 ;
        RECT 3374.200 3701.620 3374.460 3701.880 ;
        RECT 3376.040 3701.620 3376.300 3701.880 ;
        RECT 3376.960 3701.620 3377.220 3701.880 ;
        RECT 3375.120 3686.320 3375.380 3686.580 ;
        RECT 3376.960 3686.320 3377.220 3686.580 ;
        RECT 3374.200 3679.860 3374.460 3680.120 ;
        RECT 3376.960 3679.860 3377.220 3680.120 ;
        RECT 3374.660 3649.600 3374.920 3649.860 ;
        RECT 3376.960 3649.600 3377.220 3649.860 ;
        RECT 3374.200 3645.180 3374.460 3645.440 ;
        RECT 3376.960 3645.180 3377.220 3645.440 ;
        RECT 3376.500 3633.280 3376.760 3633.540 ;
        RECT 3374.660 3632.260 3374.920 3632.520 ;
        RECT 3376.040 3632.260 3376.300 3632.520 ;
        RECT 3376.500 3632.260 3376.760 3632.520 ;
        RECT 208.940 3565.620 209.200 3565.880 ;
        RECT 212.160 3565.620 212.420 3565.880 ;
        RECT 208.940 3558.480 209.200 3558.740 ;
        RECT 213.080 3558.480 213.340 3558.740 ;
        RECT 208.940 3530.940 209.200 3531.200 ;
        RECT 212.160 3530.940 212.420 3531.200 ;
        RECT 211.240 3525.840 211.500 3526.100 ;
        RECT 208.940 3524.480 209.200 3524.740 ;
        RECT 212.620 3524.480 212.880 3524.740 ;
        RECT 208.940 3504.080 209.200 3504.340 ;
        RECT 213.540 3504.080 213.800 3504.340 ;
        RECT 211.240 3502.380 211.500 3502.640 ;
        RECT 3374.660 3494.900 3374.920 3495.160 ;
        RECT 3376.960 3494.900 3377.220 3495.160 ;
        RECT 3374.660 3480.960 3374.920 3481.220 ;
        RECT 3374.660 3479.940 3374.920 3480.200 ;
        RECT 3374.660 3476.540 3374.920 3476.800 ;
        RECT 3376.960 3476.540 3377.220 3476.800 ;
        RECT 3374.200 3466.000 3374.460 3466.260 ;
        RECT 3376.960 3466.000 3377.220 3466.260 ;
        RECT 3376.040 3458.180 3376.300 3458.440 ;
        RECT 3376.960 3458.180 3377.220 3458.440 ;
        RECT 3376.500 3457.840 3376.760 3458.100 ;
        RECT 3376.500 3456.820 3376.760 3457.080 ;
        RECT 3375.580 3425.880 3375.840 3426.140 ;
        RECT 3376.960 3425.880 3377.220 3426.140 ;
        RECT 3376.040 3420.100 3376.300 3420.360 ;
        RECT 3376.960 3420.100 3377.220 3420.360 ;
        RECT 3375.120 3356.860 3375.380 3357.120 ;
        RECT 3376.040 3356.860 3376.300 3357.120 ;
        RECT 208.940 3349.720 209.200 3349.980 ;
        RECT 212.160 3349.720 212.420 3349.980 ;
        RECT 208.940 3342.580 209.200 3342.840 ;
        RECT 213.080 3342.580 213.340 3342.840 ;
        RECT 212.160 3315.380 212.420 3315.640 ;
        RECT 208.940 3315.040 209.200 3315.300 ;
        RECT 211.240 3315.040 211.500 3315.300 ;
        RECT 212.160 3314.020 212.420 3314.280 ;
        RECT 208.940 3303.820 209.200 3304.080 ;
        RECT 212.160 3303.820 212.420 3304.080 ;
        RECT 208.940 3293.280 209.200 3293.540 ;
        RECT 211.700 3293.280 211.960 3293.540 ;
        RECT 213.540 3293.280 213.800 3293.540 ;
        RECT 3374.660 3250.440 3374.920 3250.700 ;
        RECT 3376.960 3250.440 3377.220 3250.700 ;
        RECT 3374.200 3239.900 3374.460 3240.160 ;
        RECT 3376.960 3239.900 3377.220 3240.160 ;
        RECT 3376.040 3228.680 3376.300 3228.940 ;
        RECT 3376.960 3228.680 3377.220 3228.940 ;
        RECT 3375.120 3198.760 3375.380 3199.020 ;
        RECT 3376.960 3198.760 3377.220 3199.020 ;
        RECT 3376.040 3194.000 3376.300 3194.260 ;
        RECT 3376.960 3194.000 3377.220 3194.260 ;
        RECT 209.860 3125.320 210.120 3125.580 ;
        RECT 213.080 3125.320 213.340 3125.580 ;
        RECT 208.940 3092.340 209.200 3092.600 ;
        RECT 212.160 3092.340 212.420 3092.600 ;
        RECT 211.240 3074.660 211.500 3074.920 ;
        RECT 213.540 3074.660 213.800 3074.920 ;
        RECT 212.620 3029.100 212.880 3029.360 ;
        RECT 213.540 3029.100 213.800 3029.360 ;
        RECT 3374.660 3027.400 3374.920 3027.660 ;
        RECT 3376.960 3027.400 3377.220 3027.660 ;
        RECT 3374.200 3011.760 3374.460 3012.020 ;
        RECT 3374.660 3010.400 3374.920 3010.660 ;
        RECT 3376.960 3010.400 3377.220 3010.660 ;
        RECT 3376.040 3003.940 3376.300 3004.200 ;
        RECT 3376.960 3003.940 3377.220 3004.200 ;
        RECT 3375.120 2973.340 3375.380 2973.600 ;
        RECT 3376.960 2973.340 3377.220 2973.600 ;
        RECT 3376.040 2968.920 3376.300 2969.180 ;
        RECT 3376.960 2968.920 3377.220 2969.180 ;
        RECT 208.940 2917.580 209.200 2917.840 ;
        RECT 212.160 2917.580 212.420 2917.840 ;
        RECT 208.940 2909.080 209.200 2909.340 ;
        RECT 212.620 2909.080 212.880 2909.340 ;
        RECT 208.940 2882.220 209.200 2882.480 ;
        RECT 212.160 2882.220 212.420 2882.480 ;
        RECT 211.240 2881.200 211.500 2881.460 ;
        RECT 213.540 2881.200 213.800 2881.460 ;
        RECT 208.940 2871.680 209.200 2871.940 ;
        RECT 212.160 2871.680 212.420 2871.940 ;
        RECT 213.080 2871.680 213.340 2871.940 ;
        RECT 208.940 2858.080 209.200 2858.340 ;
        RECT 213.080 2858.080 213.340 2858.340 ;
        RECT 3374.200 2804.700 3374.460 2804.960 ;
        RECT 3376.960 2804.700 3377.220 2804.960 ;
        RECT 3374.660 2789.060 3374.920 2789.320 ;
        RECT 3376.960 2789.060 3377.220 2789.320 ;
        RECT 3376.040 2777.840 3376.300 2778.100 ;
        RECT 3376.960 2777.840 3377.220 2778.100 ;
        RECT 3375.120 2752.340 3375.380 2752.600 ;
        RECT 3376.960 2752.340 3377.220 2752.600 ;
        RECT 208.940 2695.560 209.200 2695.820 ;
        RECT 212.620 2695.560 212.880 2695.820 ;
        RECT 208.940 2660.540 209.200 2660.800 ;
        RECT 212.160 2660.540 212.420 2660.800 ;
        RECT 209.860 2642.180 210.120 2642.440 ;
        RECT 213.540 2642.180 213.800 2642.440 ;
        RECT 3376.500 2519.440 3376.760 2519.700 ;
        RECT 3387.540 2519.440 3387.800 2519.700 ;
        RECT 3370.520 2138.980 3370.780 2139.240 ;
        RECT 3387.540 2138.980 3387.800 2139.240 ;
        RECT 208.940 2064.520 209.200 2064.780 ;
        RECT 211.700 2064.520 211.960 2064.780 ;
        RECT 208.940 2054.660 209.200 2054.920 ;
        RECT 213.080 2054.660 213.340 2054.920 ;
        RECT 208.940 2028.820 209.200 2029.080 ;
        RECT 211.700 2028.820 211.960 2029.080 ;
        RECT 208.940 2022.360 209.200 2022.620 ;
        RECT 212.160 2022.360 212.420 2022.620 ;
        RECT 208.940 2001.960 209.200 2002.220 ;
        RECT 212.160 2001.960 212.420 2002.220 ;
        RECT 213.540 2001.960 213.800 2002.220 ;
        RECT 3374.200 1918.660 3374.460 1918.920 ;
        RECT 3376.960 1918.660 3377.220 1918.920 ;
        RECT 3375.120 1898.940 3375.380 1899.200 ;
        RECT 3376.960 1898.940 3377.220 1899.200 ;
        RECT 3374.200 1891.800 3374.460 1892.060 ;
        RECT 3376.960 1891.800 3377.220 1892.060 ;
        RECT 3374.200 1857.120 3374.460 1857.380 ;
        RECT 3376.960 1857.120 3377.220 1857.380 ;
        RECT 208.940 1847.600 209.200 1847.860 ;
        RECT 211.700 1847.600 211.960 1847.860 ;
        RECT 208.940 1843.180 209.200 1843.440 ;
        RECT 213.080 1843.180 213.340 1843.440 ;
        RECT 208.940 1812.920 209.200 1813.180 ;
        RECT 211.700 1812.920 211.960 1813.180 ;
        RECT 208.940 1801.700 209.200 1801.960 ;
        RECT 212.620 1801.700 212.880 1801.960 ;
        RECT 213.540 1801.700 213.800 1801.960 ;
        RECT 208.940 1786.060 209.200 1786.320 ;
        RECT 212.160 1786.060 212.420 1786.320 ;
        RECT 211.240 1785.040 211.500 1785.300 ;
        RECT 3374.660 1687.460 3374.920 1687.720 ;
        RECT 3376.960 1687.460 3377.220 1687.720 ;
        RECT 3375.120 1676.920 3375.380 1677.180 ;
        RECT 3376.040 1676.920 3376.300 1677.180 ;
        RECT 3376.960 1676.920 3377.220 1677.180 ;
        RECT 3374.200 1640.200 3374.460 1640.460 ;
        RECT 3375.580 1640.200 3375.840 1640.460 ;
        RECT 3376.960 1640.200 3377.220 1640.460 ;
        RECT 208.940 1631.700 209.200 1631.960 ;
        RECT 212.160 1631.700 212.420 1631.960 ;
        RECT 208.940 1625.580 209.200 1625.840 ;
        RECT 212.620 1625.580 212.880 1625.840 ;
        RECT 208.940 1597.020 209.200 1597.280 ;
        RECT 212.160 1597.020 212.420 1597.280 ;
        RECT 208.940 1590.560 209.200 1590.820 ;
        RECT 213.540 1590.560 213.800 1590.820 ;
        RECT 3374.660 1466.120 3374.920 1466.380 ;
        RECT 3376.960 1466.120 3377.220 1466.380 ;
        RECT 3374.660 1447.420 3374.920 1447.680 ;
        RECT 3375.580 1447.420 3375.840 1447.680 ;
        RECT 3376.960 1447.420 3377.220 1447.680 ;
        RECT 3375.120 1443.000 3375.380 1443.260 ;
        RECT 3376.500 1443.000 3376.760 1443.260 ;
        RECT 208.940 1415.800 209.200 1416.060 ;
        RECT 212.160 1415.800 212.420 1416.060 ;
        RECT 3374.200 1411.380 3374.460 1411.640 ;
        RECT 3376.960 1411.380 3377.220 1411.640 ;
        RECT 208.940 1410.360 209.200 1410.620 ;
        RECT 212.620 1410.360 212.880 1410.620 ;
        RECT 3376.040 1405.940 3376.300 1406.200 ;
        RECT 3376.960 1405.940 3377.220 1406.200 ;
        RECT 208.940 1380.780 209.200 1381.040 ;
        RECT 212.160 1380.780 212.420 1381.040 ;
        RECT 208.940 1369.560 209.200 1369.820 ;
        RECT 213.080 1369.560 213.340 1369.820 ;
        RECT 3375.120 1237.300 3375.380 1237.560 ;
        RECT 3376.960 1237.300 3377.220 1237.560 ;
        RECT 3374.660 1222.340 3374.920 1222.600 ;
        RECT 3376.960 1222.340 3377.220 1222.600 ;
        RECT 208.940 1199.560 209.200 1199.820 ;
        RECT 212.160 1199.560 212.420 1199.820 ;
        RECT 208.940 1192.420 209.200 1192.680 ;
        RECT 212.620 1192.420 212.880 1192.680 ;
        RECT 3374.200 1188.340 3374.460 1188.600 ;
        RECT 3376.960 1188.340 3377.220 1188.600 ;
        RECT 3376.040 1181.200 3376.300 1181.460 ;
        RECT 3376.960 1181.200 3377.220 1181.460 ;
        RECT 208.940 1164.880 209.200 1165.140 ;
        RECT 212.160 1164.880 212.420 1165.140 ;
        RECT 208.940 1158.420 209.200 1158.680 ;
        RECT 213.080 1158.420 213.340 1158.680 ;
        RECT 3375.120 1011.540 3375.380 1011.800 ;
        RECT 3376.960 1011.540 3377.220 1011.800 ;
        RECT 3374.660 1001.000 3374.920 1001.260 ;
        RECT 3376.960 1001.000 3377.220 1001.260 ;
        RECT 3376.040 996.240 3376.300 996.500 ;
        RECT 3376.040 995.220 3376.300 995.480 ;
        RECT 208.940 983.660 209.200 983.920 ;
        RECT 213.540 983.660 213.800 983.920 ;
        RECT 208.940 976.520 209.200 976.780 ;
        RECT 212.160 976.520 212.420 976.780 ;
        RECT 3376.040 959.520 3376.300 959.780 ;
        RECT 3376.960 959.520 3377.220 959.780 ;
        RECT 208.940 948.980 209.200 949.240 ;
        RECT 213.540 948.980 213.800 949.240 ;
        RECT 208.940 937.760 209.200 938.020 ;
        RECT 212.620 937.760 212.880 938.020 ;
        RECT 3376.500 793.600 3376.760 793.860 ;
        RECT 3375.580 792.580 3375.840 792.840 ;
        RECT 3374.200 786.460 3374.460 786.720 ;
        RECT 3375.120 786.460 3375.380 786.720 ;
        RECT 3376.960 786.460 3377.220 786.720 ;
        RECT 3374.660 775.920 3374.920 776.180 ;
        RECT 3376.960 775.920 3377.220 776.180 ;
        RECT 3375.120 735.460 3375.380 735.720 ;
        RECT 3376.040 735.460 3376.300 735.720 ;
        RECT 3376.960 735.460 3377.220 735.720 ;
        RECT 3374.200 562.400 3374.460 562.660 ;
        RECT 3376.960 562.400 3377.220 562.660 ;
        RECT 3374.660 545.400 3374.920 545.660 ;
        RECT 3376.960 545.400 3377.220 545.660 ;
        RECT 3376.040 538.940 3376.300 539.200 ;
        RECT 3376.960 538.940 3377.220 539.200 ;
        RECT 3376.040 510.040 3376.300 510.300 ;
        RECT 3376.500 509.020 3376.760 509.280 ;
        RECT 210.780 224.440 211.040 224.700 ;
        RECT 738.400 224.440 738.660 224.700 ;
        RECT 2618.880 224.440 2619.140 224.700 ;
        RECT 3374.660 224.440 3374.920 224.700 ;
        RECT 210.320 224.100 210.580 224.360 ;
        RECT 979.900 224.100 980.160 224.360 ;
        RECT 2580.700 224.100 2580.960 224.360 ;
        RECT 3375.580 224.100 3375.840 224.360 ;
        RECT 2298.260 223.760 2298.520 224.020 ;
        RECT 2338.280 223.760 2338.540 224.020 ;
        RECT 2076.540 223.420 2076.800 223.680 ;
        RECT 2339.200 223.420 2339.460 223.680 ;
        RECT 2366.340 223.420 2366.600 223.680 ;
        RECT 2634.060 223.420 2634.320 223.680 ;
        RECT 1476.240 222.740 1476.500 223.000 ;
        RECT 1516.260 222.740 1516.520 223.000 ;
        RECT 1750.400 222.740 1750.660 223.000 ;
        RECT 1790.420 222.740 1790.680 223.000 ;
        RECT 1802.840 222.740 1803.100 223.000 ;
        RECT 2033.760 222.740 2034.020 223.000 ;
        RECT 2307.460 223.080 2307.720 223.340 ;
        RECT 2580.700 223.080 2580.960 223.340 ;
        RECT 2339.200 222.740 2339.460 223.000 ;
        RECT 2344.720 222.740 2344.980 223.000 ;
        RECT 2618.880 222.740 2619.140 223.000 ;
        RECT 444.000 222.060 444.260 222.320 ;
        RECT 995.080 222.060 995.340 222.320 ;
        RECT 1537.880 222.400 1538.140 222.660 ;
        RECT 1812.040 222.400 1812.300 222.660 ;
        RECT 2086.200 222.400 2086.460 222.660 ;
        RECT 2359.900 222.400 2360.160 222.660 ;
        RECT 2366.340 222.400 2366.600 222.660 ;
        RECT 2572.420 222.400 2572.680 222.660 ;
        RECT 2612.440 222.400 2612.700 222.660 ;
        RECT 1004.280 222.060 1004.540 222.320 ;
        RECT 1206.680 222.060 1206.940 222.320 ;
        RECT 1488.660 222.060 1488.920 222.320 ;
        RECT 1503.840 222.060 1504.100 222.320 ;
        RECT 1525.460 222.060 1525.720 222.320 ;
        RECT 1547.080 222.060 1547.340 222.320 ;
        RECT 1762.820 222.060 1763.080 222.320 ;
        RECT 1778.000 222.060 1778.260 222.320 ;
        RECT 1799.620 222.060 1799.880 222.320 ;
        RECT 1821.240 222.060 1821.500 222.320 ;
        RECT 2036.980 222.060 2037.240 222.320 ;
        RECT 2052.160 222.060 2052.420 222.320 ;
        RECT 2080.220 222.060 2080.480 222.320 ;
        RECT 2095.400 222.060 2095.660 222.320 ;
        RECT 2310.680 222.060 2310.940 222.320 ;
        RECT 2325.860 222.060 2326.120 222.320 ;
        RECT 2353.920 222.060 2354.180 222.320 ;
        RECT 2369.100 222.060 2369.360 222.320 ;
        RECT 2584.840 222.060 2585.100 222.320 ;
        RECT 2600.020 222.060 2600.280 222.320 ;
        RECT 942.640 221.720 942.900 221.980 ;
        RECT 964.260 221.720 964.520 221.980 ;
        RECT 1007.500 221.720 1007.760 221.980 ;
        RECT 1485.440 221.720 1485.700 221.980 ;
        RECT 1497.860 221.720 1498.120 221.980 ;
        RECT 1528.680 221.720 1528.940 221.980 ;
        RECT 1759.600 221.720 1759.860 221.980 ;
        RECT 1772.020 221.720 1772.280 221.980 ;
        RECT 1802.840 221.720 1803.100 221.980 ;
        RECT 2024.560 221.720 2024.820 221.980 ;
        RECT 2064.580 221.720 2064.840 221.980 ;
        RECT 738.400 221.040 738.660 221.300 ;
        RECT 942.640 221.040 942.900 221.300 ;
        RECT 979.900 221.040 980.160 221.300 ;
        RECT 1522.700 221.040 1522.960 221.300 ;
        RECT 1796.860 221.040 1797.120 221.300 ;
        RECT 2071.020 221.040 2071.280 221.300 ;
        RECT 2076.540 221.040 2076.800 221.300 ;
        RECT 933.440 220.700 933.700 220.960 ;
        RECT 973.460 220.700 973.720 220.960 ;
        RECT 211.240 210.500 211.500 210.760 ;
        RECT 704.820 210.500 705.080 210.760 ;
        RECT 2348.400 209.820 2348.660 210.080 ;
        RECT 2353.460 209.820 2353.720 210.080 ;
        RECT 992.320 209.480 992.580 209.740 ;
        RECT 1000.600 209.480 1000.860 209.740 ;
        RECT 1526.380 209.480 1526.640 209.740 ;
        RECT 1531.440 209.480 1531.700 209.740 ;
        RECT 1543.400 209.480 1543.660 209.740 ;
        RECT 946.320 208.800 946.580 209.060 ;
        RECT 955.520 208.800 955.780 209.060 ;
        RECT 961.500 208.800 961.760 209.060 ;
        RECT 967.940 208.800 968.200 209.060 ;
        RECT 982.200 208.800 982.460 209.060 ;
        RECT 1800.080 208.800 1800.340 209.060 ;
        RECT 1805.600 208.800 1805.860 209.060 ;
        RECT 1817.560 208.800 1817.820 209.060 ;
        RECT 2052.620 208.800 2052.880 209.060 ;
        RECT 2057.680 208.800 2057.940 209.060 ;
        RECT 2074.240 208.800 2074.500 209.060 ;
        RECT 2079.300 208.800 2079.560 209.060 ;
        RECT 2326.780 208.800 2327.040 209.060 ;
        RECT 2331.840 208.800 2332.100 209.060 ;
        RECT 2347.020 208.800 2347.280 209.060 ;
        RECT 2600.480 208.800 2600.740 209.060 ;
        RECT 2606.000 208.800 2606.260 209.060 ;
        RECT 2621.180 208.800 2621.440 209.060 ;
        RECT 2627.620 208.800 2627.880 209.060 ;
        RECT 2639.580 208.800 2639.840 209.060 ;
        RECT 715.400 207.100 715.660 207.360 ;
        RECT 723.220 206.760 723.480 207.020 ;
        RECT 704.980 200.300 705.240 200.560 ;
        RECT 715.400 200.300 715.660 200.560 ;
        RECT 2863.600 206.760 2863.860 207.020 ;
        RECT 2863.600 203.360 2863.860 203.620 ;
        RECT 3374.200 203.360 3374.460 203.620 ;
      LAYER met2 ;
        RECT 381.210 4979.715 460.915 5188.000 ;
        RECT 381.210 4979.435 382.205 4979.715 ;
        RECT 383.045 4979.435 384.965 4979.715 ;
        RECT 385.805 4979.435 388.185 4979.715 ;
        RECT 389.025 4979.435 391.405 4979.715 ;
        RECT 392.245 4979.435 394.165 4979.715 ;
        RECT 395.005 4979.435 397.385 4979.715 ;
        RECT 398.225 4979.435 400.605 4979.715 ;
        RECT 401.445 4979.435 403.365 4979.715 ;
        RECT 404.205 4979.435 406.585 4979.715 ;
        RECT 407.425 4979.435 409.805 4979.715 ;
        RECT 410.645 4979.435 412.565 4979.715 ;
        RECT 413.405 4979.435 415.785 4979.715 ;
        RECT 416.625 4979.435 419.005 4979.715 ;
        RECT 419.845 4979.435 422.225 4979.715 ;
        RECT 423.065 4979.435 424.985 4979.715 ;
        RECT 425.825 4979.435 428.205 4979.715 ;
        RECT 429.045 4979.435 431.425 4979.715 ;
        RECT 432.265 4979.435 434.185 4979.715 ;
        RECT 435.025 4979.435 437.405 4979.715 ;
        RECT 438.245 4979.435 440.625 4979.715 ;
        RECT 441.465 4979.435 443.385 4979.715 ;
        RECT 444.225 4979.435 446.605 4979.715 ;
        RECT 447.445 4979.435 449.825 4979.715 ;
        RECT 450.665 4979.435 452.585 4979.715 ;
        RECT 453.425 4979.435 455.805 4979.715 ;
        RECT 456.645 4979.435 459.025 4979.715 ;
        RECT 459.865 4979.435 460.915 4979.715 ;
        RECT 638.210 4979.715 717.915 5188.000 ;
        RECT 638.210 4979.435 639.205 4979.715 ;
        RECT 640.045 4979.435 641.965 4979.715 ;
        RECT 642.805 4979.435 645.185 4979.715 ;
        RECT 646.025 4979.435 648.405 4979.715 ;
        RECT 649.245 4979.435 651.165 4979.715 ;
        RECT 652.005 4979.435 654.385 4979.715 ;
        RECT 655.225 4979.435 657.605 4979.715 ;
        RECT 658.445 4979.435 660.365 4979.715 ;
        RECT 661.205 4979.435 663.585 4979.715 ;
        RECT 664.425 4979.435 666.805 4979.715 ;
        RECT 667.645 4979.435 669.565 4979.715 ;
        RECT 670.405 4979.435 672.785 4979.715 ;
        RECT 673.625 4979.435 676.005 4979.715 ;
        RECT 676.845 4979.435 679.225 4979.715 ;
        RECT 680.065 4979.435 681.985 4979.715 ;
        RECT 682.825 4979.435 685.205 4979.715 ;
        RECT 686.045 4979.435 688.425 4979.715 ;
        RECT 689.265 4979.435 691.185 4979.715 ;
        RECT 692.025 4979.435 694.405 4979.715 ;
        RECT 695.245 4979.435 697.625 4979.715 ;
        RECT 698.465 4979.435 700.385 4979.715 ;
        RECT 701.225 4979.435 703.605 4979.715 ;
        RECT 704.445 4979.435 706.825 4979.715 ;
        RECT 707.665 4979.435 709.585 4979.715 ;
        RECT 710.425 4979.435 712.805 4979.715 ;
        RECT 713.645 4979.435 716.025 4979.715 ;
        RECT 716.865 4979.435 717.915 4979.715 ;
        RECT 895.210 4979.715 974.915 5188.000 ;
        RECT 895.210 4979.435 896.205 4979.715 ;
        RECT 897.045 4979.435 898.965 4979.715 ;
        RECT 899.805 4979.435 902.185 4979.715 ;
        RECT 903.025 4979.435 905.405 4979.715 ;
        RECT 906.245 4979.435 908.165 4979.715 ;
        RECT 909.005 4979.435 911.385 4979.715 ;
        RECT 912.225 4979.435 914.605 4979.715 ;
        RECT 915.445 4979.435 917.365 4979.715 ;
        RECT 918.205 4979.435 920.585 4979.715 ;
        RECT 921.425 4979.435 923.805 4979.715 ;
        RECT 924.645 4979.435 926.565 4979.715 ;
        RECT 927.405 4979.435 929.785 4979.715 ;
        RECT 930.625 4979.435 933.005 4979.715 ;
        RECT 933.845 4979.435 936.225 4979.715 ;
        RECT 937.065 4979.435 938.985 4979.715 ;
        RECT 939.825 4979.435 942.205 4979.715 ;
        RECT 943.045 4979.435 945.425 4979.715 ;
        RECT 946.265 4979.435 948.185 4979.715 ;
        RECT 949.025 4979.435 951.405 4979.715 ;
        RECT 952.245 4979.435 954.625 4979.715 ;
        RECT 955.465 4979.435 957.385 4979.715 ;
        RECT 958.225 4979.435 960.605 4979.715 ;
        RECT 961.445 4979.435 963.825 4979.715 ;
        RECT 964.665 4979.435 966.585 4979.715 ;
        RECT 967.425 4979.435 969.805 4979.715 ;
        RECT 970.645 4979.435 973.025 4979.715 ;
        RECT 973.865 4979.435 974.915 4979.715 ;
        RECT 1152.210 4979.715 1231.915 5188.000 ;
        RECT 1152.210 4979.435 1153.205 4979.715 ;
        RECT 1154.045 4979.435 1155.965 4979.715 ;
        RECT 1156.805 4979.435 1159.185 4979.715 ;
        RECT 1160.025 4979.435 1162.405 4979.715 ;
        RECT 1163.245 4979.435 1165.165 4979.715 ;
        RECT 1166.005 4979.435 1168.385 4979.715 ;
        RECT 1169.225 4979.435 1171.605 4979.715 ;
        RECT 1172.445 4979.435 1174.365 4979.715 ;
        RECT 1175.205 4979.435 1177.585 4979.715 ;
        RECT 1178.425 4979.435 1180.805 4979.715 ;
        RECT 1181.645 4979.435 1183.565 4979.715 ;
        RECT 1184.405 4979.435 1186.785 4979.715 ;
        RECT 1187.625 4979.435 1190.005 4979.715 ;
        RECT 1190.845 4979.435 1193.225 4979.715 ;
        RECT 1194.065 4979.435 1195.985 4979.715 ;
        RECT 1196.825 4979.435 1199.205 4979.715 ;
        RECT 1200.045 4979.435 1202.425 4979.715 ;
        RECT 1203.265 4979.435 1205.185 4979.715 ;
        RECT 1206.025 4979.435 1208.405 4979.715 ;
        RECT 1209.245 4979.435 1211.625 4979.715 ;
        RECT 1212.465 4979.435 1214.385 4979.715 ;
        RECT 1215.225 4979.435 1217.605 4979.715 ;
        RECT 1218.445 4979.435 1220.825 4979.715 ;
        RECT 1221.665 4979.435 1223.585 4979.715 ;
        RECT 1224.425 4979.435 1226.805 4979.715 ;
        RECT 1227.645 4979.435 1230.025 4979.715 ;
        RECT 1230.865 4979.435 1231.915 4979.715 ;
        RECT 1410.210 4979.715 1489.915 5188.000 ;
        RECT 1667.265 4990.035 1741.290 5183.075 ;
      LAYER met2 ;
        RECT 1666.210 4989.315 1666.490 4989.685 ;
      LAYER met2 ;
        RECT 1410.210 4979.435 1411.205 4979.715 ;
        RECT 1412.045 4979.435 1413.965 4979.715 ;
        RECT 1414.805 4979.435 1417.185 4979.715 ;
        RECT 1418.025 4979.435 1420.405 4979.715 ;
        RECT 1421.245 4979.435 1423.165 4979.715 ;
        RECT 1424.005 4979.435 1426.385 4979.715 ;
        RECT 1427.225 4979.435 1429.605 4979.715 ;
        RECT 1430.445 4979.435 1432.365 4979.715 ;
        RECT 1433.205 4979.435 1435.585 4979.715 ;
        RECT 1436.425 4979.435 1438.805 4979.715 ;
        RECT 1439.645 4979.435 1441.565 4979.715 ;
        RECT 1442.405 4979.435 1444.785 4979.715 ;
        RECT 1445.625 4979.435 1448.005 4979.715 ;
        RECT 1448.845 4979.435 1451.225 4979.715 ;
        RECT 1452.065 4979.435 1453.985 4979.715 ;
        RECT 1454.825 4979.435 1457.205 4979.715 ;
        RECT 1458.045 4979.435 1460.425 4979.715 ;
        RECT 1461.265 4979.435 1463.185 4979.715 ;
        RECT 1464.025 4979.435 1466.405 4979.715 ;
        RECT 1467.245 4979.435 1469.625 4979.715 ;
        RECT 1470.465 4979.435 1472.385 4979.715 ;
        RECT 1473.225 4979.435 1475.605 4979.715 ;
        RECT 1476.445 4979.435 1478.825 4979.715 ;
        RECT 1479.665 4979.435 1481.585 4979.715 ;
        RECT 1482.425 4979.435 1484.805 4979.715 ;
        RECT 1485.645 4979.435 1488.025 4979.715 ;
        RECT 1488.865 4979.435 1489.915 4979.715 ;
      LAYER met2 ;
        RECT 382.485 4977.035 382.765 4979.435 ;
        RECT 397.665 4977.260 397.945 4979.435 ;
        RECT 412.845 4977.260 413.125 4979.435 ;
        RECT 419.285 4977.260 419.565 4979.435 ;
        RECT 397.600 4977.035 397.945 4977.260 ;
        RECT 412.780 4977.035 413.125 4977.260 ;
        RECT 419.220 4977.035 419.565 4977.260 ;
        RECT 434.465 4977.035 434.745 4979.435 ;
        RECT 440.905 4977.035 441.185 4979.435 ;
        RECT 450.105 4977.260 450.385 4979.435 ;
        RECT 450.040 4977.035 450.385 4977.260 ;
        RECT 452.865 4977.035 453.145 4979.435 ;
        RECT 459.305 4977.260 459.585 4979.435 ;
        RECT 459.240 4977.035 459.585 4977.260 ;
        RECT 639.485 4977.035 639.765 4979.435 ;
        RECT 654.665 4977.035 654.945 4979.435 ;
        RECT 669.845 4977.035 670.125 4979.435 ;
        RECT 676.285 4977.035 676.565 4979.435 ;
        RECT 691.465 4977.035 691.745 4979.435 ;
        RECT 697.905 4977.035 698.185 4979.435 ;
        RECT 707.105 4977.035 707.385 4979.435 ;
        RECT 709.865 4977.035 710.145 4979.435 ;
        RECT 716.305 4977.035 716.585 4979.435 ;
        RECT 896.485 4977.035 896.765 4979.435 ;
        RECT 911.665 4977.330 911.945 4979.435 ;
        RECT 926.845 4977.330 927.125 4979.435 ;
        RECT 933.285 4977.330 933.565 4979.435 ;
        RECT 911.665 4977.035 912.020 4977.330 ;
        RECT 926.845 4977.035 927.200 4977.330 ;
        RECT 933.285 4977.035 933.640 4977.330 ;
        RECT 948.465 4977.035 948.745 4979.435 ;
        RECT 954.905 4977.035 955.185 4979.435 ;
        RECT 964.105 4977.330 964.385 4979.435 ;
        RECT 964.105 4977.035 964.460 4977.330 ;
        RECT 966.865 4977.035 967.145 4979.435 ;
        RECT 973.305 4977.330 973.585 4979.435 ;
        RECT 973.305 4977.035 973.660 4977.330 ;
        RECT 1153.485 4977.035 1153.765 4979.435 ;
        RECT 1168.665 4977.330 1168.945 4979.435 ;
        RECT 1183.845 4977.330 1184.125 4979.435 ;
        RECT 1190.285 4977.330 1190.565 4979.435 ;
        RECT 1168.560 4977.035 1168.945 4977.330 ;
        RECT 1183.740 4977.035 1184.125 4977.330 ;
        RECT 1190.180 4977.035 1190.565 4977.330 ;
        RECT 1205.465 4977.035 1205.745 4979.435 ;
        RECT 1211.905 4977.035 1212.185 4979.435 ;
        RECT 1221.105 4977.330 1221.385 4979.435 ;
        RECT 1221.000 4977.035 1221.385 4977.330 ;
        RECT 1223.865 4977.035 1224.145 4979.435 ;
        RECT 1230.305 4977.330 1230.585 4979.435 ;
        RECT 1230.200 4977.035 1230.585 4977.330 ;
        RECT 1411.485 4977.035 1411.765 4979.435 ;
        RECT 1426.665 4977.260 1426.945 4979.435 ;
        RECT 1441.845 4977.260 1442.125 4979.435 ;
        RECT 1448.285 4977.260 1448.565 4979.435 ;
        RECT 1426.620 4977.035 1426.945 4977.260 ;
        RECT 1441.800 4977.035 1442.125 4977.260 ;
        RECT 1448.240 4977.035 1448.565 4977.260 ;
        RECT 1463.465 4977.035 1463.745 4979.435 ;
        RECT 1469.905 4977.035 1470.185 4979.435 ;
        RECT 1479.105 4977.260 1479.385 4979.435 ;
        RECT 1479.060 4977.035 1479.385 4977.260 ;
        RECT 1481.865 4977.035 1482.145 4979.435 ;
        RECT 1488.305 4977.260 1488.585 4979.435 ;
        RECT 1488.260 4977.035 1488.585 4977.260 ;
        RECT 397.600 4967.730 397.740 4977.035 ;
        RECT 397.540 4967.410 397.800 4967.730 ;
        RECT 397.600 4965.350 397.740 4967.410 ;
        RECT 217.220 4965.030 217.480 4965.350 ;
        RECT 397.540 4965.030 397.800 4965.350 ;
        RECT 211.700 4964.350 211.960 4964.670 ;
        RECT 211.760 4912.870 211.900 4964.350 ;
        RECT 211.760 4912.730 212.360 4912.870 ;
      LAYER met2 ;
        RECT 0.000 4849.865 208.565 4850.915 ;
        RECT 0.000 4849.025 208.285 4849.865 ;
      LAYER met2 ;
        RECT 208.565 4849.305 210.965 4849.585 ;
      LAYER met2 ;
        RECT 0.000 4846.645 208.565 4849.025 ;
      LAYER met2 ;
        RECT 209.460 4846.770 209.600 4849.305 ;
      LAYER met2 ;
        RECT 0.000 4845.805 208.285 4846.645 ;
      LAYER met2 ;
        RECT 209.460 4846.630 211.440 4846.770 ;
      LAYER met2 ;
        RECT 0.000 4843.425 208.565 4845.805 ;
        RECT 0.000 4842.585 208.285 4843.425 ;
      LAYER met2 ;
        RECT 208.565 4842.865 210.965 4843.145 ;
      LAYER met2 ;
        RECT 0.000 4840.665 208.565 4842.585 ;
        RECT 0.000 4839.825 208.285 4840.665 ;
      LAYER met2 ;
        RECT 208.565 4840.105 210.965 4840.385 ;
        RECT 209.000 4839.890 209.140 4840.105 ;
      LAYER met2 ;
        RECT 0.000 4837.445 208.565 4839.825 ;
      LAYER met2 ;
        RECT 208.940 4839.570 209.200 4839.890 ;
      LAYER met2 ;
        RECT 0.000 4836.605 208.285 4837.445 ;
        RECT 0.000 4834.225 208.565 4836.605 ;
        RECT 0.000 4833.385 208.285 4834.225 ;
        RECT 0.000 4831.465 208.565 4833.385 ;
        RECT 0.000 4830.625 208.285 4831.465 ;
      LAYER met2 ;
        RECT 208.565 4830.905 210.965 4831.185 ;
      LAYER met2 ;
        RECT 0.000 4828.245 208.565 4830.625 ;
        RECT 0.000 4827.405 208.285 4828.245 ;
        RECT 0.000 4825.025 208.565 4827.405 ;
        RECT 0.000 4824.185 208.285 4825.025 ;
      LAYER met2 ;
        RECT 208.565 4824.465 210.965 4824.745 ;
      LAYER met2 ;
        RECT 0.000 4822.265 208.565 4824.185 ;
        RECT 0.000 4821.425 208.285 4822.265 ;
        RECT 0.000 4819.045 208.565 4821.425 ;
        RECT 0.000 4818.205 208.285 4819.045 ;
        RECT 0.000 4815.825 208.565 4818.205 ;
        RECT 0.000 4814.985 208.285 4815.825 ;
        RECT 0.000 4813.065 208.565 4814.985 ;
        RECT 0.000 4812.225 208.285 4813.065 ;
        RECT 0.000 4809.845 208.565 4812.225 ;
      LAYER met2 ;
        RECT 211.300 4810.050 211.440 4846.630 ;
        RECT 212.220 4839.890 212.360 4912.730 ;
        RECT 212.160 4839.570 212.420 4839.890 ;
        RECT 209.000 4809.910 211.440 4810.050 ;
      LAYER met2 ;
        RECT 0.000 4809.005 208.285 4809.845 ;
      LAYER met2 ;
        RECT 209.000 4809.565 209.140 4809.910 ;
        RECT 208.565 4809.285 210.965 4809.565 ;
        RECT 208.610 4809.230 209.140 4809.285 ;
      LAYER met2 ;
        RECT 0.000 4806.625 208.565 4809.005 ;
        RECT 0.000 4805.785 208.285 4806.625 ;
        RECT 0.000 4803.405 208.565 4805.785 ;
        RECT 0.000 4802.565 208.285 4803.405 ;
      LAYER met2 ;
        RECT 208.565 4802.845 210.965 4803.125 ;
        RECT 209.460 4802.570 209.600 4802.845 ;
      LAYER met2 ;
        RECT 0.000 4800.645 208.565 4802.565 ;
      LAYER met2 ;
        RECT 209.460 4802.430 211.440 4802.570 ;
      LAYER met2 ;
        RECT 0.000 4799.805 208.285 4800.645 ;
        RECT 0.000 4797.425 208.565 4799.805 ;
        RECT 0.000 4796.585 208.285 4797.425 ;
        RECT 0.000 4794.205 208.565 4796.585 ;
      LAYER met2 ;
        RECT 211.300 4795.350 211.440 4802.430 ;
        RECT 211.240 4795.030 211.500 4795.350 ;
      LAYER met2 ;
        RECT 0.000 4793.365 208.285 4794.205 ;
        RECT 0.000 4791.445 208.565 4793.365 ;
        RECT 0.000 4790.605 208.285 4791.445 ;
        RECT 0.000 4788.225 208.565 4790.605 ;
      LAYER met2 ;
        RECT 208.940 4788.230 209.200 4788.550 ;
      LAYER met2 ;
        RECT 0.000 4787.385 208.285 4788.225 ;
      LAYER met2 ;
        RECT 209.000 4787.945 209.140 4788.230 ;
        RECT 208.565 4787.665 210.965 4787.945 ;
        RECT 212.220 4787.530 212.360 4839.570 ;
        RECT 213.080 4795.030 213.340 4795.350 ;
      LAYER met2 ;
        RECT 0.000 4785.005 208.565 4787.385 ;
      LAYER met2 ;
        RECT 212.160 4787.210 212.420 4787.530 ;
        RECT 212.160 4786.190 212.420 4786.510 ;
      LAYER met2 ;
        RECT 0.000 4784.165 208.285 4785.005 ;
        RECT 0.000 4782.245 208.565 4784.165 ;
        RECT 0.000 4781.405 208.285 4782.245 ;
        RECT 0.000 4779.025 208.565 4781.405 ;
        RECT 0.000 4778.185 208.285 4779.025 ;
        RECT 0.000 4775.805 208.565 4778.185 ;
        RECT 0.000 4774.965 208.285 4775.805 ;
        RECT 0.000 4773.045 208.565 4774.965 ;
        RECT 0.000 4772.205 208.285 4773.045 ;
      LAYER met2 ;
        RECT 208.565 4772.485 210.965 4772.765 ;
      LAYER met2 ;
        RECT 0.000 4771.210 208.565 4772.205 ;
        RECT 0.035 4636.200 151.405 4645.935 ;
        RECT 153.765 4635.000 158.415 4646.140 ;
        RECT 160.165 4636.200 174.575 4645.935 ;
        RECT 0.035 4634.700 197.965 4635.000 ;
        RECT 0.035 4614.095 198.000 4634.700 ;
        RECT 0.035 4613.535 197.965 4614.095 ;
        RECT 0.035 4580.925 198.000 4613.535 ;
        RECT 0.035 4580.495 197.965 4580.925 ;
        RECT 0.035 4560.500 198.000 4580.495 ;
        RECT 0.035 4560.000 197.965 4560.500 ;
        RECT 153.800 4549.025 158.450 4560.000 ;
        RECT 4.925 4399.390 200.000 4423.290 ;
      LAYER met2 ;
        RECT 207.090 4409.275 207.370 4409.645 ;
        RECT 207.160 4400.125 207.300 4409.275 ;
        RECT 207.090 4399.755 207.370 4400.125 ;
        RECT 211.230 4399.755 211.510 4400.125 ;
      LAYER met2 ;
        RECT 4.925 4373.395 197.965 4399.390 ;
        RECT 198.080 4374.895 200.000 4376.895 ;
        RECT 4.925 4349.495 200.000 4373.395 ;
        RECT 4.925 4349.265 197.965 4349.495 ;
        RECT 4.925 4188.390 200.000 4212.290 ;
        RECT 4.925 4162.395 197.965 4188.390 ;
        RECT 198.080 4163.895 200.000 4165.895 ;
        RECT 4.925 4138.495 200.000 4162.395 ;
        RECT 4.925 4138.265 197.965 4138.495 ;
        RECT 0.000 4000.865 208.565 4001.915 ;
        RECT 0.000 4000.025 208.285 4000.865 ;
      LAYER met2 ;
        RECT 208.565 4000.305 210.965 4000.585 ;
      LAYER met2 ;
        RECT 0.000 3997.645 208.565 4000.025 ;
      LAYER met2 ;
        RECT 209.000 3998.050 209.140 4000.305 ;
        RECT 208.940 3997.730 209.200 3998.050 ;
      LAYER met2 ;
        RECT 0.000 3996.805 208.285 3997.645 ;
        RECT 0.000 3994.425 208.565 3996.805 ;
        RECT 0.000 3993.585 208.285 3994.425 ;
      LAYER met2 ;
        RECT 208.565 3993.865 210.965 3994.145 ;
      LAYER met2 ;
        RECT 0.000 3991.665 208.565 3993.585 ;
        RECT 0.000 3990.825 208.285 3991.665 ;
      LAYER met2 ;
        RECT 208.565 3991.105 210.965 3991.385 ;
      LAYER met2 ;
        RECT 0.000 3988.445 208.565 3990.825 ;
      LAYER met2 ;
        RECT 209.000 3988.870 209.140 3991.105 ;
        RECT 208.940 3988.550 209.200 3988.870 ;
      LAYER met2 ;
        RECT 0.000 3987.605 208.285 3988.445 ;
        RECT 0.000 3985.225 208.565 3987.605 ;
        RECT 0.000 3984.385 208.285 3985.225 ;
        RECT 0.000 3982.465 208.565 3984.385 ;
        RECT 0.000 3981.625 208.285 3982.465 ;
      LAYER met2 ;
        RECT 208.565 3981.905 210.965 3982.185 ;
      LAYER met2 ;
        RECT 0.000 3979.245 208.565 3981.625 ;
        RECT 0.000 3978.405 208.285 3979.245 ;
        RECT 0.000 3976.025 208.565 3978.405 ;
        RECT 0.000 3975.185 208.285 3976.025 ;
      LAYER met2 ;
        RECT 208.565 3975.465 210.965 3975.745 ;
      LAYER met2 ;
        RECT 0.000 3973.265 208.565 3975.185 ;
        RECT 0.000 3972.425 208.285 3973.265 ;
        RECT 0.000 3970.045 208.565 3972.425 ;
        RECT 0.000 3969.205 208.285 3970.045 ;
        RECT 0.000 3966.825 208.565 3969.205 ;
        RECT 0.000 3965.985 208.285 3966.825 ;
        RECT 0.000 3964.065 208.565 3965.985 ;
        RECT 0.000 3963.225 208.285 3964.065 ;
        RECT 0.000 3960.845 208.565 3963.225 ;
      LAYER met2 ;
        RECT 208.940 3962.710 209.200 3963.030 ;
      LAYER met2 ;
        RECT 0.000 3960.005 208.285 3960.845 ;
      LAYER met2 ;
        RECT 209.000 3960.565 209.140 3962.710 ;
        RECT 208.565 3960.285 210.965 3960.565 ;
      LAYER met2 ;
        RECT 0.000 3957.625 208.565 3960.005 ;
        RECT 0.000 3956.785 208.285 3957.625 ;
        RECT 0.000 3954.405 208.565 3956.785 ;
      LAYER met2 ;
        RECT 211.300 3954.610 211.440 4399.755 ;
        RECT 211.700 3997.730 211.960 3998.050 ;
        RECT 211.760 3963.030 211.900 3997.730 ;
        RECT 212.220 3988.870 212.360 4786.190 ;
        RECT 213.140 4409.645 213.280 4795.030 ;
        RECT 217.280 4788.550 217.420 4965.030 ;
        RECT 412.780 4965.010 412.920 4977.035 ;
        RECT 416.400 4967.750 416.660 4968.070 ;
        RECT 416.460 4965.010 416.600 4967.750 ;
        RECT 419.220 4966.710 419.360 4977.035 ;
        RECT 450.040 4967.390 450.180 4977.035 ;
        RECT 449.980 4967.070 450.240 4967.390 ;
        RECT 419.160 4966.390 419.420 4966.710 ;
        RECT 217.680 4964.690 217.940 4965.010 ;
        RECT 412.720 4964.690 412.980 4965.010 ;
        RECT 416.400 4964.690 416.660 4965.010 ;
        RECT 217.740 4795.350 217.880 4964.690 ;
        RECT 450.040 4964.670 450.180 4967.070 ;
        RECT 459.240 4966.710 459.380 4977.035 ;
        RECT 654.740 4967.730 654.880 4977.035 ;
        RECT 669.920 4968.070 670.060 4977.035 ;
        RECT 676.360 4968.070 676.500 4977.035 ;
        RECT 669.860 4967.750 670.120 4968.070 ;
        RECT 675.840 4967.750 676.100 4968.070 ;
        RECT 676.300 4967.750 676.560 4968.070 ;
        RECT 654.680 4967.410 654.940 4967.730 ;
        RECT 459.180 4966.390 459.440 4966.710 ;
        RECT 675.900 4966.370 676.040 4967.750 ;
        RECT 707.180 4967.390 707.320 4977.035 ;
        RECT 716.380 4975.210 716.520 4977.035 ;
        RECT 710.340 4974.890 710.600 4975.210 ;
        RECT 716.320 4974.890 716.580 4975.210 ;
        RECT 710.400 4968.070 710.540 4974.890 ;
        RECT 710.340 4967.750 710.600 4968.070 ;
        RECT 911.880 4967.730 912.020 4977.035 ;
        RECT 927.060 4967.730 927.200 4977.035 ;
        RECT 933.500 4968.070 933.640 4977.035 ;
        RECT 933.440 4967.750 933.700 4968.070 ;
        RECT 911.820 4967.410 912.080 4967.730 ;
        RECT 917.340 4967.410 917.600 4967.730 ;
        RECT 927.000 4967.410 927.260 4967.730 ;
        RECT 707.120 4967.070 707.380 4967.390 ;
        RECT 917.400 4966.710 917.540 4967.410 ;
        RECT 917.340 4966.390 917.600 4966.710 ;
        RECT 927.060 4966.370 927.200 4967.410 ;
        RECT 964.320 4967.390 964.460 4977.035 ;
        RECT 973.520 4968.070 973.660 4977.035 ;
        RECT 1168.560 4968.070 1168.700 4977.035 ;
        RECT 973.460 4967.750 973.720 4968.070 ;
        RECT 1168.500 4967.750 1168.760 4968.070 ;
        RECT 964.260 4967.070 964.520 4967.390 ;
        RECT 1168.560 4966.710 1168.700 4967.750 ;
        RECT 1183.740 4967.730 1183.880 4977.035 ;
        RECT 1187.360 4967.750 1187.620 4968.070 ;
        RECT 1183.680 4967.410 1183.940 4967.730 ;
        RECT 1187.420 4967.050 1187.560 4967.750 ;
        RECT 1187.360 4966.730 1187.620 4967.050 ;
        RECT 1168.500 4966.390 1168.760 4966.710 ;
        RECT 1190.180 4966.370 1190.320 4977.035 ;
        RECT 1221.000 4967.390 1221.140 4977.035 ;
        RECT 1220.940 4967.070 1221.200 4967.390 ;
        RECT 1230.200 4966.370 1230.340 4977.035 ;
        RECT 1426.620 4967.050 1426.760 4977.035 ;
        RECT 1441.800 4968.070 1441.940 4977.035 ;
        RECT 1448.240 4968.070 1448.380 4977.035 ;
        RECT 1441.740 4967.750 1442.000 4968.070 ;
        RECT 1448.180 4967.750 1448.440 4968.070 ;
        RECT 1426.560 4966.730 1426.820 4967.050 ;
        RECT 1441.800 4966.370 1441.940 4967.750 ;
        RECT 1479.060 4967.730 1479.200 4977.035 ;
        RECT 1488.260 4968.070 1488.400 4977.035 ;
        RECT 1488.200 4967.750 1488.460 4968.070 ;
        RECT 1479.000 4967.410 1479.260 4967.730 ;
        RECT 1666.280 4967.050 1666.420 4989.315 ;
      LAYER met2 ;
        RECT 1667.495 4988.000 1691.395 4990.035 ;
        RECT 1692.895 4988.000 1694.895 4989.920 ;
        RECT 1717.390 4988.000 1741.290 4990.035 ;
        RECT 1919.210 4979.715 1998.915 5188.000 ;
        RECT 1919.210 4979.435 1920.205 4979.715 ;
        RECT 1921.045 4979.435 1922.965 4979.715 ;
        RECT 1923.805 4979.435 1926.185 4979.715 ;
        RECT 1927.025 4979.435 1929.405 4979.715 ;
        RECT 1930.245 4979.435 1932.165 4979.715 ;
        RECT 1933.005 4979.435 1935.385 4979.715 ;
        RECT 1936.225 4979.435 1938.605 4979.715 ;
        RECT 1939.445 4979.435 1941.365 4979.715 ;
        RECT 1942.205 4979.435 1944.585 4979.715 ;
        RECT 1945.425 4979.435 1947.805 4979.715 ;
        RECT 1948.645 4979.435 1950.565 4979.715 ;
        RECT 1951.405 4979.435 1953.785 4979.715 ;
        RECT 1954.625 4979.435 1957.005 4979.715 ;
        RECT 1957.845 4979.435 1960.225 4979.715 ;
        RECT 1961.065 4979.435 1962.985 4979.715 ;
        RECT 1963.825 4979.435 1966.205 4979.715 ;
        RECT 1967.045 4979.435 1969.425 4979.715 ;
        RECT 1970.265 4979.435 1972.185 4979.715 ;
        RECT 1973.025 4979.435 1975.405 4979.715 ;
        RECT 1976.245 4979.435 1978.625 4979.715 ;
        RECT 1979.465 4979.435 1981.385 4979.715 ;
        RECT 1982.225 4979.435 1984.605 4979.715 ;
        RECT 1985.445 4979.435 1987.825 4979.715 ;
        RECT 1988.665 4979.435 1990.585 4979.715 ;
        RECT 1991.425 4979.435 1993.805 4979.715 ;
        RECT 1994.645 4979.435 1997.025 4979.715 ;
        RECT 1997.865 4979.435 1998.915 4979.715 ;
        RECT 2364.210 4979.715 2443.915 5188.000 ;
        RECT 2364.210 4979.435 2365.205 4979.715 ;
        RECT 2366.045 4979.435 2367.965 4979.715 ;
        RECT 2368.805 4979.435 2371.185 4979.715 ;
        RECT 2372.025 4979.435 2374.405 4979.715 ;
        RECT 2375.245 4979.435 2377.165 4979.715 ;
        RECT 2378.005 4979.435 2380.385 4979.715 ;
        RECT 2381.225 4979.435 2383.605 4979.715 ;
        RECT 2384.445 4979.435 2386.365 4979.715 ;
        RECT 2387.205 4979.435 2389.585 4979.715 ;
        RECT 2390.425 4979.435 2392.805 4979.715 ;
        RECT 2393.645 4979.435 2395.565 4979.715 ;
        RECT 2396.405 4979.435 2398.785 4979.715 ;
        RECT 2399.625 4979.435 2402.005 4979.715 ;
        RECT 2402.845 4979.435 2405.225 4979.715 ;
        RECT 2406.065 4979.435 2407.985 4979.715 ;
        RECT 2408.825 4979.435 2411.205 4979.715 ;
        RECT 2412.045 4979.435 2414.425 4979.715 ;
        RECT 2415.265 4979.435 2417.185 4979.715 ;
        RECT 2418.025 4979.435 2420.405 4979.715 ;
        RECT 2421.245 4979.435 2423.625 4979.715 ;
        RECT 2424.465 4979.435 2426.385 4979.715 ;
        RECT 2427.225 4979.435 2429.605 4979.715 ;
        RECT 2430.445 4979.435 2432.825 4979.715 ;
        RECT 2433.665 4979.435 2435.585 4979.715 ;
        RECT 2436.425 4979.435 2438.805 4979.715 ;
        RECT 2439.645 4979.435 2442.025 4979.715 ;
        RECT 2442.865 4979.435 2443.915 4979.715 ;
        RECT 2621.210 4979.715 2700.915 5188.000 ;
        RECT 2878.265 4990.035 2952.290 5183.075 ;
        RECT 2878.495 4988.000 2902.395 4990.035 ;
      LAYER met2 ;
        RECT 2903.150 4989.315 2903.430 4989.685 ;
      LAYER met2 ;
        RECT 2621.210 4979.435 2622.205 4979.715 ;
        RECT 2623.045 4979.435 2624.965 4979.715 ;
        RECT 2625.805 4979.435 2628.185 4979.715 ;
        RECT 2629.025 4979.435 2631.405 4979.715 ;
        RECT 2632.245 4979.435 2634.165 4979.715 ;
        RECT 2635.005 4979.435 2637.385 4979.715 ;
        RECT 2638.225 4979.435 2640.605 4979.715 ;
        RECT 2641.445 4979.435 2643.365 4979.715 ;
        RECT 2644.205 4979.435 2646.585 4979.715 ;
        RECT 2647.425 4979.435 2649.805 4979.715 ;
        RECT 2650.645 4979.435 2652.565 4979.715 ;
        RECT 2653.405 4979.435 2655.785 4979.715 ;
        RECT 2656.625 4979.435 2659.005 4979.715 ;
        RECT 2659.845 4979.435 2662.225 4979.715 ;
        RECT 2663.065 4979.435 2664.985 4979.715 ;
        RECT 2665.825 4979.435 2668.205 4979.715 ;
        RECT 2669.045 4979.435 2671.425 4979.715 ;
        RECT 2672.265 4979.435 2674.185 4979.715 ;
        RECT 2675.025 4979.435 2677.405 4979.715 ;
        RECT 2678.245 4979.435 2680.625 4979.715 ;
        RECT 2681.465 4979.435 2683.385 4979.715 ;
        RECT 2684.225 4979.435 2686.605 4979.715 ;
        RECT 2687.445 4979.435 2689.825 4979.715 ;
        RECT 2690.665 4979.435 2692.585 4979.715 ;
        RECT 2693.425 4979.435 2695.805 4979.715 ;
        RECT 2696.645 4979.435 2699.025 4979.715 ;
        RECT 2699.865 4979.435 2700.915 4979.715 ;
      LAYER met2 ;
        RECT 1920.485 4977.035 1920.765 4979.435 ;
        RECT 1935.665 4977.260 1935.945 4979.435 ;
        RECT 1950.845 4977.260 1951.125 4979.435 ;
        RECT 1957.285 4977.260 1957.565 4979.435 ;
        RECT 1935.665 4977.035 1935.980 4977.260 ;
        RECT 1950.845 4977.035 1951.160 4977.260 ;
        RECT 1957.285 4977.035 1957.600 4977.260 ;
        RECT 1972.465 4977.035 1972.745 4979.435 ;
        RECT 1978.905 4977.035 1979.185 4979.435 ;
        RECT 1988.105 4977.260 1988.385 4979.435 ;
        RECT 1988.105 4977.035 1988.420 4977.260 ;
        RECT 1990.865 4977.035 1991.145 4979.435 ;
        RECT 1997.305 4977.260 1997.585 4979.435 ;
        RECT 1997.305 4977.035 1997.620 4977.260 ;
        RECT 2365.485 4977.035 2365.765 4979.435 ;
        RECT 2380.665 4977.260 2380.945 4979.435 ;
        RECT 2395.845 4977.260 2396.125 4979.435 ;
        RECT 2402.285 4977.260 2402.565 4979.435 ;
        RECT 2380.660 4977.035 2380.945 4977.260 ;
        RECT 2395.840 4977.035 2396.125 4977.260 ;
        RECT 2402.280 4977.035 2402.565 4977.260 ;
        RECT 2417.465 4977.035 2417.745 4979.435 ;
        RECT 2423.905 4977.035 2424.185 4979.435 ;
        RECT 2433.105 4977.260 2433.385 4979.435 ;
        RECT 2433.100 4977.035 2433.385 4977.260 ;
        RECT 2435.865 4977.035 2436.145 4979.435 ;
        RECT 2442.305 4977.260 2442.585 4979.435 ;
        RECT 2442.300 4977.035 2442.585 4977.260 ;
        RECT 2622.485 4977.035 2622.765 4979.435 ;
        RECT 2637.665 4977.035 2637.945 4979.435 ;
        RECT 2652.845 4977.035 2653.125 4979.435 ;
        RECT 2659.285 4977.035 2659.565 4979.435 ;
        RECT 2674.465 4977.035 2674.745 4979.435 ;
        RECT 2680.905 4977.035 2681.185 4979.435 ;
        RECT 2690.105 4977.035 2690.385 4979.435 ;
        RECT 2692.865 4977.035 2693.145 4979.435 ;
        RECT 2699.305 4977.035 2699.585 4979.435 ;
        RECT 1935.840 4967.050 1935.980 4977.035 ;
        RECT 1666.220 4966.730 1666.480 4967.050 ;
        RECT 1935.780 4966.730 1936.040 4967.050 ;
        RECT 1951.020 4966.710 1951.160 4977.035 ;
        RECT 1957.460 4968.070 1957.600 4977.035 ;
        RECT 1957.400 4967.750 1957.660 4968.070 ;
        RECT 1988.280 4967.730 1988.420 4977.035 ;
        RECT 1997.480 4968.070 1997.620 4977.035 ;
        RECT 1997.420 4967.750 1997.680 4968.070 ;
        RECT 1988.220 4967.410 1988.480 4967.730 ;
        RECT 2380.660 4967.390 2380.800 4977.035 ;
        RECT 2380.600 4967.070 2380.860 4967.390 ;
        RECT 2395.840 4966.710 2395.980 4977.035 ;
        RECT 2402.280 4968.070 2402.420 4977.035 ;
        RECT 2402.220 4967.750 2402.480 4968.070 ;
        RECT 2433.100 4967.730 2433.240 4977.035 ;
        RECT 2442.300 4968.070 2442.440 4977.035 ;
        RECT 2442.240 4967.750 2442.500 4968.070 ;
        RECT 2433.040 4967.410 2433.300 4967.730 ;
        RECT 2637.800 4967.390 2637.940 4977.035 ;
        RECT 2637.740 4967.070 2638.000 4967.390 ;
        RECT 2641.420 4967.070 2641.680 4967.390 ;
        RECT 2641.480 4966.710 2641.620 4967.070 ;
        RECT 1950.960 4966.390 1951.220 4966.710 ;
        RECT 2395.780 4966.390 2396.040 4966.710 ;
        RECT 2641.420 4966.390 2641.680 4966.710 ;
        RECT 2652.980 4966.370 2653.120 4977.035 ;
        RECT 2659.420 4968.070 2659.560 4977.035 ;
        RECT 2659.360 4967.750 2659.620 4968.070 ;
        RECT 2690.240 4967.730 2690.380 4977.035 ;
        RECT 2699.440 4976.570 2699.580 4977.035 ;
        RECT 2690.640 4976.250 2690.900 4976.570 ;
        RECT 2699.380 4976.250 2699.640 4976.570 ;
        RECT 2690.700 4968.070 2690.840 4976.250 ;
        RECT 2690.640 4967.750 2690.900 4968.070 ;
        RECT 2690.180 4967.410 2690.440 4967.730 ;
        RECT 2656.140 4967.070 2656.400 4967.390 ;
        RECT 2656.200 4966.370 2656.340 4967.070 ;
        RECT 675.840 4966.050 676.100 4966.370 ;
        RECT 927.000 4966.050 927.260 4966.370 ;
        RECT 1190.120 4966.050 1190.380 4966.370 ;
        RECT 1230.140 4966.050 1230.400 4966.370 ;
        RECT 1441.740 4966.050 1442.000 4966.370 ;
        RECT 2652.920 4966.050 2653.180 4966.370 ;
        RECT 2656.140 4966.050 2656.400 4966.370 ;
        RECT 449.980 4964.350 450.240 4964.670 ;
        RECT 2903.220 4961.170 2903.360 4989.315 ;
      LAYER met2 ;
        RECT 2903.895 4988.000 2905.895 4989.920 ;
        RECT 2928.390 4988.000 2952.290 4990.035 ;
        RECT 3130.210 4979.715 3209.915 5188.000 ;
        RECT 3130.210 4979.435 3131.205 4979.715 ;
        RECT 3132.045 4979.435 3133.965 4979.715 ;
        RECT 3134.805 4979.435 3137.185 4979.715 ;
        RECT 3138.025 4979.435 3140.405 4979.715 ;
        RECT 3141.245 4979.435 3143.165 4979.715 ;
        RECT 3144.005 4979.435 3146.385 4979.715 ;
        RECT 3147.225 4979.435 3149.605 4979.715 ;
        RECT 3150.445 4979.435 3152.365 4979.715 ;
        RECT 3153.205 4979.435 3155.585 4979.715 ;
        RECT 3156.425 4979.435 3158.805 4979.715 ;
        RECT 3159.645 4979.435 3161.565 4979.715 ;
        RECT 3162.405 4979.435 3164.785 4979.715 ;
        RECT 3165.625 4979.435 3168.005 4979.715 ;
        RECT 3168.845 4979.435 3171.225 4979.715 ;
        RECT 3172.065 4979.435 3173.985 4979.715 ;
        RECT 3174.825 4979.435 3177.205 4979.715 ;
        RECT 3178.045 4979.435 3180.425 4979.715 ;
        RECT 3181.265 4979.435 3183.185 4979.715 ;
        RECT 3184.025 4979.435 3186.405 4979.715 ;
        RECT 3187.245 4979.435 3189.625 4979.715 ;
        RECT 3190.465 4979.435 3192.385 4979.715 ;
        RECT 3193.225 4979.435 3195.605 4979.715 ;
        RECT 3196.445 4979.435 3198.825 4979.715 ;
        RECT 3199.665 4979.435 3201.585 4979.715 ;
        RECT 3202.425 4979.435 3204.805 4979.715 ;
        RECT 3205.645 4979.435 3208.025 4979.715 ;
        RECT 3208.865 4979.435 3209.915 4979.715 ;
      LAYER met2 ;
        RECT 3131.485 4977.035 3131.765 4979.435 ;
        RECT 3146.665 4977.330 3146.945 4979.435 ;
        RECT 3161.845 4977.330 3162.125 4979.435 ;
        RECT 3168.285 4977.330 3168.565 4979.435 ;
        RECT 3146.560 4977.035 3146.945 4977.330 ;
        RECT 3161.740 4977.035 3162.125 4977.330 ;
        RECT 3168.180 4977.035 3168.565 4977.330 ;
        RECT 3183.465 4977.035 3183.745 4979.435 ;
        RECT 3189.905 4977.035 3190.185 4979.435 ;
        RECT 3199.105 4977.330 3199.385 4979.435 ;
        RECT 3199.000 4977.035 3199.385 4977.330 ;
        RECT 3201.865 4977.035 3202.145 4979.435 ;
        RECT 3208.305 4977.330 3208.585 4979.435 ;
        RECT 3208.200 4977.035 3208.585 4977.330 ;
        RECT 3146.560 4966.710 3146.700 4977.035 ;
        RECT 3161.740 4967.390 3161.880 4977.035 ;
        RECT 3168.180 4968.070 3168.320 4977.035 ;
        RECT 3168.120 4967.750 3168.380 4968.070 ;
        RECT 3199.000 4967.730 3199.140 4977.035 ;
        RECT 3208.200 4968.070 3208.340 4977.035 ;
        RECT 3208.140 4967.750 3208.400 4968.070 ;
        RECT 3198.940 4967.410 3199.200 4967.730 ;
        RECT 3161.680 4967.070 3161.940 4967.390 ;
        RECT 3146.500 4966.390 3146.760 4966.710 ;
        RECT 3146.560 4964.670 3146.700 4966.390 ;
        RECT 3161.740 4965.350 3161.880 4967.070 ;
        RECT 3199.000 4965.690 3199.140 4967.410 ;
        RECT 3198.940 4965.370 3199.200 4965.690 ;
        RECT 3370.980 4965.370 3371.240 4965.690 ;
        RECT 3161.680 4965.030 3161.940 4965.350 ;
        RECT 3146.500 4964.350 3146.760 4964.670 ;
        RECT 2902.760 4961.030 2903.360 4961.170 ;
        RECT 2902.760 4950.730 2902.900 4961.030 ;
        RECT 2902.700 4950.410 2902.960 4950.730 ;
        RECT 3370.520 4950.410 3370.780 4950.730 ;
        RECT 217.680 4795.030 217.940 4795.350 ;
        RECT 217.220 4788.230 217.480 4788.550 ;
        RECT 213.070 4409.275 213.350 4409.645 ;
        RECT 212.160 3988.550 212.420 3988.870 ;
        RECT 213.080 3988.550 213.340 3988.870 ;
        RECT 211.700 3962.710 211.960 3963.030 ;
        RECT 209.460 3954.470 211.440 3954.610 ;
      LAYER met2 ;
        RECT 0.000 3953.565 208.285 3954.405 ;
      LAYER met2 ;
        RECT 209.460 3954.125 209.600 3954.470 ;
        RECT 208.565 3953.845 210.965 3954.125 ;
        RECT 208.610 3953.790 209.600 3953.845 ;
      LAYER met2 ;
        RECT 0.000 3951.645 208.565 3953.565 ;
        RECT 0.000 3950.805 208.285 3951.645 ;
        RECT 0.000 3948.425 208.565 3950.805 ;
        RECT 0.000 3947.585 208.285 3948.425 ;
        RECT 0.000 3945.205 208.565 3947.585 ;
        RECT 0.000 3944.365 208.285 3945.205 ;
        RECT 0.000 3942.445 208.565 3944.365 ;
        RECT 0.000 3941.605 208.285 3942.445 ;
        RECT 0.000 3939.225 208.565 3941.605 ;
        RECT 0.000 3938.385 208.285 3939.225 ;
      LAYER met2 ;
        RECT 208.610 3938.945 209.140 3938.970 ;
        RECT 208.565 3938.665 210.965 3938.945 ;
      LAYER met2 ;
        RECT 0.000 3936.005 208.565 3938.385 ;
      LAYER met2 ;
        RECT 209.000 3936.510 209.140 3938.665 ;
        RECT 208.940 3936.190 209.200 3936.510 ;
      LAYER met2 ;
        RECT 0.000 3935.165 208.285 3936.005 ;
        RECT 0.000 3933.245 208.565 3935.165 ;
        RECT 0.000 3932.405 208.285 3933.245 ;
        RECT 0.000 3930.025 208.565 3932.405 ;
        RECT 0.000 3929.185 208.285 3930.025 ;
        RECT 0.000 3926.805 208.565 3929.185 ;
        RECT 0.000 3925.965 208.285 3926.805 ;
        RECT 0.000 3924.045 208.565 3925.965 ;
        RECT 0.000 3923.205 208.285 3924.045 ;
      LAYER met2 ;
        RECT 208.565 3923.485 210.965 3923.765 ;
      LAYER met2 ;
        RECT 0.000 3922.210 208.565 3923.205 ;
        RECT 0.000 3784.865 208.565 3785.915 ;
        RECT 0.000 3784.025 208.285 3784.865 ;
      LAYER met2 ;
        RECT 208.610 3784.585 209.140 3784.610 ;
        RECT 208.565 3784.305 210.965 3784.585 ;
      LAYER met2 ;
        RECT 0.000 3781.645 208.565 3784.025 ;
      LAYER met2 ;
        RECT 209.000 3782.150 209.140 3784.305 ;
        RECT 208.940 3781.830 209.200 3782.150 ;
      LAYER met2 ;
        RECT 0.000 3780.805 208.285 3781.645 ;
        RECT 0.000 3778.425 208.565 3780.805 ;
        RECT 0.000 3777.585 208.285 3778.425 ;
      LAYER met2 ;
        RECT 208.565 3777.865 210.965 3778.145 ;
      LAYER met2 ;
        RECT 0.000 3775.665 208.565 3777.585 ;
      LAYER met2 ;
        RECT 208.940 3776.730 209.200 3777.050 ;
      LAYER met2 ;
        RECT 0.000 3774.825 208.285 3775.665 ;
      LAYER met2 ;
        RECT 209.000 3775.385 209.140 3776.730 ;
        RECT 208.565 3775.105 210.965 3775.385 ;
      LAYER met2 ;
        RECT 0.000 3772.445 208.565 3774.825 ;
        RECT 0.000 3771.605 208.285 3772.445 ;
        RECT 0.000 3769.225 208.565 3771.605 ;
        RECT 0.000 3768.385 208.285 3769.225 ;
        RECT 0.000 3766.465 208.565 3768.385 ;
        RECT 0.000 3765.625 208.285 3766.465 ;
      LAYER met2 ;
        RECT 208.565 3765.905 210.965 3766.185 ;
      LAYER met2 ;
        RECT 0.000 3763.245 208.565 3765.625 ;
        RECT 0.000 3762.405 208.285 3763.245 ;
        RECT 0.000 3760.025 208.565 3762.405 ;
        RECT 0.000 3759.185 208.285 3760.025 ;
      LAYER met2 ;
        RECT 208.565 3759.465 210.965 3759.745 ;
      LAYER met2 ;
        RECT 0.000 3757.265 208.565 3759.185 ;
        RECT 0.000 3756.425 208.285 3757.265 ;
        RECT 0.000 3754.045 208.565 3756.425 ;
        RECT 0.000 3753.205 208.285 3754.045 ;
        RECT 0.000 3750.825 208.565 3753.205 ;
        RECT 0.000 3749.985 208.285 3750.825 ;
        RECT 0.000 3748.065 208.565 3749.985 ;
        RECT 0.000 3747.225 208.285 3748.065 ;
        RECT 0.000 3744.845 208.565 3747.225 ;
      LAYER met2 ;
        RECT 208.940 3746.810 209.200 3747.130 ;
      LAYER met2 ;
        RECT 0.000 3744.005 208.285 3744.845 ;
      LAYER met2 ;
        RECT 209.000 3744.565 209.140 3746.810 ;
        RECT 208.565 3744.285 210.965 3744.565 ;
      LAYER met2 ;
        RECT 0.000 3741.625 208.565 3744.005 ;
        RECT 0.000 3740.785 208.285 3741.625 ;
        RECT 0.000 3738.405 208.565 3740.785 ;
        RECT 0.000 3737.565 208.285 3738.405 ;
      LAYER met2 ;
        RECT 208.565 3737.845 210.965 3738.125 ;
      LAYER met2 ;
        RECT 0.000 3735.645 208.565 3737.565 ;
      LAYER met2 ;
        RECT 209.000 3735.650 209.140 3737.845 ;
        RECT 211.300 3735.650 211.440 3954.470 ;
        RECT 212.620 3936.190 212.880 3936.510 ;
        RECT 212.160 3776.730 212.420 3777.050 ;
      LAYER met2 ;
        RECT 0.000 3734.805 208.285 3735.645 ;
      LAYER met2 ;
        RECT 209.000 3735.510 211.440 3735.650 ;
      LAYER met2 ;
        RECT 0.000 3732.425 208.565 3734.805 ;
        RECT 0.000 3731.585 208.285 3732.425 ;
        RECT 0.000 3729.205 208.565 3731.585 ;
        RECT 0.000 3728.365 208.285 3729.205 ;
        RECT 0.000 3726.445 208.565 3728.365 ;
        RECT 0.000 3725.605 208.285 3726.445 ;
        RECT 0.000 3723.225 208.565 3725.605 ;
      LAYER met2 ;
        RECT 208.940 3725.390 209.200 3725.710 ;
      LAYER met2 ;
        RECT 0.000 3722.385 208.285 3723.225 ;
      LAYER met2 ;
        RECT 209.000 3722.945 209.140 3725.390 ;
        RECT 208.565 3722.665 210.965 3722.945 ;
      LAYER met2 ;
        RECT 0.000 3720.005 208.565 3722.385 ;
        RECT 0.000 3719.165 208.285 3720.005 ;
        RECT 0.000 3717.245 208.565 3719.165 ;
        RECT 0.000 3716.405 208.285 3717.245 ;
        RECT 0.000 3714.025 208.565 3716.405 ;
        RECT 0.000 3713.185 208.285 3714.025 ;
        RECT 0.000 3710.805 208.565 3713.185 ;
        RECT 0.000 3709.965 208.285 3710.805 ;
        RECT 0.000 3708.045 208.565 3709.965 ;
        RECT 0.000 3707.205 208.285 3708.045 ;
      LAYER met2 ;
        RECT 208.565 3707.485 210.965 3707.765 ;
      LAYER met2 ;
        RECT 0.000 3706.210 208.565 3707.205 ;
        RECT 0.000 3568.865 208.565 3569.915 ;
        RECT 0.000 3568.025 208.285 3568.865 ;
      LAYER met2 ;
        RECT 208.565 3568.305 210.965 3568.585 ;
      LAYER met2 ;
        RECT 0.000 3565.645 208.565 3568.025 ;
      LAYER met2 ;
        RECT 209.000 3565.910 209.140 3568.305 ;
      LAYER met2 ;
        RECT 0.000 3564.805 208.285 3565.645 ;
      LAYER met2 ;
        RECT 208.940 3565.590 209.200 3565.910 ;
      LAYER met2 ;
        RECT 0.000 3562.425 208.565 3564.805 ;
        RECT 0.000 3561.585 208.285 3562.425 ;
      LAYER met2 ;
        RECT 208.565 3561.865 210.965 3562.145 ;
      LAYER met2 ;
        RECT 0.000 3559.665 208.565 3561.585 ;
        RECT 0.000 3558.825 208.285 3559.665 ;
      LAYER met2 ;
        RECT 208.565 3559.105 210.965 3559.385 ;
      LAYER met2 ;
        RECT 0.000 3556.445 208.565 3558.825 ;
      LAYER met2 ;
        RECT 209.000 3558.770 209.140 3559.105 ;
        RECT 208.940 3558.450 209.200 3558.770 ;
      LAYER met2 ;
        RECT 0.000 3555.605 208.285 3556.445 ;
        RECT 0.000 3553.225 208.565 3555.605 ;
        RECT 0.000 3552.385 208.285 3553.225 ;
        RECT 0.000 3550.465 208.565 3552.385 ;
        RECT 0.000 3549.625 208.285 3550.465 ;
      LAYER met2 ;
        RECT 208.565 3549.905 210.965 3550.185 ;
      LAYER met2 ;
        RECT 0.000 3547.245 208.565 3549.625 ;
        RECT 0.000 3546.405 208.285 3547.245 ;
        RECT 0.000 3544.025 208.565 3546.405 ;
        RECT 0.000 3543.185 208.285 3544.025 ;
      LAYER met2 ;
        RECT 208.565 3543.465 210.965 3543.745 ;
      LAYER met2 ;
        RECT 0.000 3541.265 208.565 3543.185 ;
        RECT 0.000 3540.425 208.285 3541.265 ;
        RECT 0.000 3538.045 208.565 3540.425 ;
        RECT 0.000 3537.205 208.285 3538.045 ;
        RECT 0.000 3534.825 208.565 3537.205 ;
        RECT 0.000 3533.985 208.285 3534.825 ;
        RECT 0.000 3532.065 208.565 3533.985 ;
        RECT 0.000 3531.225 208.285 3532.065 ;
        RECT 0.000 3528.845 208.565 3531.225 ;
      LAYER met2 ;
        RECT 208.940 3530.910 209.200 3531.230 ;
      LAYER met2 ;
        RECT 0.000 3528.005 208.285 3528.845 ;
      LAYER met2 ;
        RECT 209.000 3528.565 209.140 3530.910 ;
        RECT 208.565 3528.285 210.965 3528.565 ;
      LAYER met2 ;
        RECT 0.000 3525.625 208.565 3528.005 ;
      LAYER met2 ;
        RECT 211.300 3526.130 211.440 3735.510 ;
        RECT 212.220 3657.070 212.360 3776.730 ;
        RECT 212.680 3725.710 212.820 3936.190 ;
        RECT 213.140 3777.050 213.280 3988.550 ;
        RECT 213.540 3781.830 213.800 3782.150 ;
        RECT 213.080 3776.730 213.340 3777.050 ;
        RECT 213.600 3747.130 213.740 3781.830 ;
        RECT 213.540 3746.810 213.800 3747.130 ;
        RECT 212.620 3725.390 212.880 3725.710 ;
        RECT 212.680 3705.370 212.820 3725.390 ;
        RECT 212.680 3705.230 213.740 3705.370 ;
        RECT 212.220 3656.930 213.280 3657.070 ;
        RECT 212.160 3565.590 212.420 3565.910 ;
        RECT 212.220 3531.230 212.360 3565.590 ;
        RECT 213.140 3558.770 213.280 3656.930 ;
        RECT 213.080 3558.450 213.340 3558.770 ;
        RECT 212.160 3530.910 212.420 3531.230 ;
        RECT 211.240 3525.810 211.500 3526.130 ;
      LAYER met2 ;
        RECT 0.000 3524.785 208.285 3525.625 ;
        RECT 0.000 3522.405 208.565 3524.785 ;
      LAYER met2 ;
        RECT 208.940 3524.450 209.200 3524.770 ;
        RECT 212.620 3524.450 212.880 3524.770 ;
      LAYER met2 ;
        RECT 0.000 3521.565 208.285 3522.405 ;
      LAYER met2 ;
        RECT 209.000 3522.130 209.140 3524.450 ;
        RECT 208.610 3522.125 209.140 3522.130 ;
        RECT 208.565 3521.845 210.965 3522.125 ;
      LAYER met2 ;
        RECT 0.000 3519.645 208.565 3521.565 ;
        RECT 0.000 3518.805 208.285 3519.645 ;
        RECT 0.000 3516.425 208.565 3518.805 ;
        RECT 0.000 3515.585 208.285 3516.425 ;
        RECT 0.000 3513.205 208.565 3515.585 ;
        RECT 0.000 3512.365 208.285 3513.205 ;
        RECT 0.000 3510.445 208.565 3512.365 ;
        RECT 0.000 3509.605 208.285 3510.445 ;
        RECT 0.000 3507.225 208.565 3509.605 ;
        RECT 0.000 3506.385 208.285 3507.225 ;
      LAYER met2 ;
        RECT 208.565 3506.665 210.965 3506.945 ;
      LAYER met2 ;
        RECT 0.000 3504.005 208.565 3506.385 ;
      LAYER met2 ;
        RECT 209.000 3504.370 209.140 3506.665 ;
        RECT 208.940 3504.050 209.200 3504.370 ;
      LAYER met2 ;
        RECT 0.000 3503.165 208.285 3504.005 ;
        RECT 0.000 3501.245 208.565 3503.165 ;
      LAYER met2 ;
        RECT 211.240 3502.350 211.500 3502.670 ;
      LAYER met2 ;
        RECT 0.000 3500.405 208.285 3501.245 ;
        RECT 0.000 3498.025 208.565 3500.405 ;
        RECT 0.000 3497.185 208.285 3498.025 ;
        RECT 0.000 3494.805 208.565 3497.185 ;
        RECT 0.000 3493.965 208.285 3494.805 ;
        RECT 0.000 3492.045 208.565 3493.965 ;
        RECT 0.000 3491.205 208.285 3492.045 ;
      LAYER met2 ;
        RECT 208.565 3491.485 210.965 3491.765 ;
      LAYER met2 ;
        RECT 0.000 3490.210 208.565 3491.205 ;
        RECT 0.000 3352.865 208.565 3353.915 ;
        RECT 0.000 3352.025 208.285 3352.865 ;
      LAYER met2 ;
        RECT 208.565 3352.305 210.965 3352.585 ;
      LAYER met2 ;
        RECT 0.000 3349.645 208.565 3352.025 ;
      LAYER met2 ;
        RECT 209.000 3350.010 209.140 3352.305 ;
        RECT 208.940 3349.690 209.200 3350.010 ;
      LAYER met2 ;
        RECT 0.000 3348.805 208.285 3349.645 ;
        RECT 0.000 3346.425 208.565 3348.805 ;
        RECT 0.000 3345.585 208.285 3346.425 ;
      LAYER met2 ;
        RECT 208.565 3345.865 210.965 3346.145 ;
      LAYER met2 ;
        RECT 0.000 3343.665 208.565 3345.585 ;
        RECT 0.000 3342.825 208.285 3343.665 ;
      LAYER met2 ;
        RECT 208.565 3343.105 210.965 3343.385 ;
        RECT 209.000 3342.870 209.140 3343.105 ;
      LAYER met2 ;
        RECT 0.000 3340.445 208.565 3342.825 ;
      LAYER met2 ;
        RECT 208.940 3342.550 209.200 3342.870 ;
      LAYER met2 ;
        RECT 0.000 3339.605 208.285 3340.445 ;
        RECT 0.000 3337.225 208.565 3339.605 ;
        RECT 0.000 3336.385 208.285 3337.225 ;
        RECT 0.000 3334.465 208.565 3336.385 ;
        RECT 0.000 3333.625 208.285 3334.465 ;
      LAYER met2 ;
        RECT 208.565 3333.905 210.965 3334.185 ;
      LAYER met2 ;
        RECT 0.000 3331.245 208.565 3333.625 ;
        RECT 0.000 3330.405 208.285 3331.245 ;
        RECT 0.000 3328.025 208.565 3330.405 ;
        RECT 0.000 3327.185 208.285 3328.025 ;
      LAYER met2 ;
        RECT 208.565 3327.465 210.965 3327.745 ;
      LAYER met2 ;
        RECT 0.000 3325.265 208.565 3327.185 ;
        RECT 0.000 3324.425 208.285 3325.265 ;
        RECT 0.000 3322.045 208.565 3324.425 ;
        RECT 0.000 3321.205 208.285 3322.045 ;
        RECT 0.000 3318.825 208.565 3321.205 ;
        RECT 0.000 3317.985 208.285 3318.825 ;
        RECT 0.000 3316.065 208.565 3317.985 ;
        RECT 0.000 3315.225 208.285 3316.065 ;
      LAYER met2 ;
        RECT 211.300 3315.330 211.440 3502.350 ;
        RECT 212.160 3349.690 212.420 3350.010 ;
        RECT 212.220 3315.670 212.360 3349.690 ;
        RECT 212.160 3315.350 212.420 3315.670 ;
      LAYER met2 ;
        RECT 0.000 3312.845 208.565 3315.225 ;
      LAYER met2 ;
        RECT 208.940 3315.010 209.200 3315.330 ;
        RECT 211.240 3315.010 211.500 3315.330 ;
      LAYER met2 ;
        RECT 0.000 3312.005 208.285 3312.845 ;
      LAYER met2 ;
        RECT 209.000 3312.565 209.140 3315.010 ;
        RECT 212.160 3313.990 212.420 3314.310 ;
        RECT 208.565 3312.285 210.965 3312.565 ;
      LAYER met2 ;
        RECT 0.000 3309.625 208.565 3312.005 ;
        RECT 0.000 3308.785 208.285 3309.625 ;
        RECT 0.000 3306.405 208.565 3308.785 ;
        RECT 0.000 3305.565 208.285 3306.405 ;
      LAYER met2 ;
        RECT 208.565 3305.845 210.965 3306.125 ;
      LAYER met2 ;
        RECT 0.000 3303.645 208.565 3305.565 ;
      LAYER met2 ;
        RECT 209.000 3304.110 209.140 3305.845 ;
        RECT 212.220 3305.210 212.360 3313.990 ;
        RECT 211.760 3305.070 212.360 3305.210 ;
        RECT 208.940 3303.790 209.200 3304.110 ;
      LAYER met2 ;
        RECT 0.000 3302.805 208.285 3303.645 ;
        RECT 0.000 3300.425 208.565 3302.805 ;
        RECT 0.000 3299.585 208.285 3300.425 ;
        RECT 0.000 3297.205 208.565 3299.585 ;
        RECT 0.000 3296.365 208.285 3297.205 ;
        RECT 0.000 3294.445 208.565 3296.365 ;
        RECT 0.000 3293.605 208.285 3294.445 ;
        RECT 0.000 3291.225 208.565 3293.605 ;
      LAYER met2 ;
        RECT 211.760 3293.570 211.900 3305.070 ;
        RECT 212.680 3304.530 212.820 3524.450 ;
        RECT 213.140 3342.870 213.280 3558.450 ;
        RECT 213.600 3504.370 213.740 3705.230 ;
        RECT 213.540 3504.050 213.800 3504.370 ;
        RECT 213.080 3342.550 213.340 3342.870 ;
        RECT 212.220 3304.390 212.820 3304.530 ;
        RECT 212.220 3304.110 212.360 3304.390 ;
        RECT 212.160 3303.790 212.420 3304.110 ;
        RECT 208.940 3293.250 209.200 3293.570 ;
        RECT 211.700 3293.250 211.960 3293.570 ;
      LAYER met2 ;
        RECT 0.000 3290.385 208.285 3291.225 ;
      LAYER met2 ;
        RECT 209.000 3290.945 209.140 3293.250 ;
        RECT 208.565 3290.665 210.965 3290.945 ;
      LAYER met2 ;
        RECT 0.000 3288.005 208.565 3290.385 ;
        RECT 0.000 3287.165 208.285 3288.005 ;
        RECT 0.000 3285.245 208.565 3287.165 ;
        RECT 0.000 3284.405 208.285 3285.245 ;
        RECT 0.000 3282.025 208.565 3284.405 ;
        RECT 0.000 3281.185 208.285 3282.025 ;
        RECT 0.000 3278.805 208.565 3281.185 ;
        RECT 0.000 3277.965 208.285 3278.805 ;
        RECT 0.000 3276.045 208.565 3277.965 ;
        RECT 0.000 3275.205 208.285 3276.045 ;
      LAYER met2 ;
        RECT 208.565 3275.485 210.965 3275.765 ;
      LAYER met2 ;
        RECT 0.000 3274.210 208.565 3275.205 ;
        RECT 0.000 3136.865 208.565 3137.915 ;
        RECT 0.000 3136.025 208.285 3136.865 ;
      LAYER met2 ;
        RECT 208.565 3136.305 210.965 3136.585 ;
      LAYER met2 ;
        RECT 0.000 3133.645 208.565 3136.025 ;
      LAYER met2 ;
        RECT 209.000 3135.890 209.140 3136.305 ;
        RECT 209.000 3135.750 211.440 3135.890 ;
      LAYER met2 ;
        RECT 0.000 3132.805 208.285 3133.645 ;
        RECT 0.000 3130.425 208.565 3132.805 ;
        RECT 0.000 3129.585 208.285 3130.425 ;
      LAYER met2 ;
        RECT 208.565 3129.865 210.965 3130.145 ;
      LAYER met2 ;
        RECT 0.000 3127.665 208.565 3129.585 ;
        RECT 0.000 3126.825 208.285 3127.665 ;
      LAYER met2 ;
        RECT 208.565 3127.105 210.965 3127.385 ;
      LAYER met2 ;
        RECT 0.000 3124.445 208.565 3126.825 ;
      LAYER met2 ;
        RECT 209.920 3125.610 210.060 3127.105 ;
        RECT 209.860 3125.290 210.120 3125.610 ;
      LAYER met2 ;
        RECT 0.000 3123.605 208.285 3124.445 ;
        RECT 0.000 3121.225 208.565 3123.605 ;
        RECT 0.000 3120.385 208.285 3121.225 ;
        RECT 0.000 3118.465 208.565 3120.385 ;
        RECT 0.000 3117.625 208.285 3118.465 ;
      LAYER met2 ;
        RECT 208.565 3117.905 210.965 3118.185 ;
      LAYER met2 ;
        RECT 0.000 3115.245 208.565 3117.625 ;
        RECT 0.000 3114.405 208.285 3115.245 ;
        RECT 0.000 3112.025 208.565 3114.405 ;
        RECT 0.000 3111.185 208.285 3112.025 ;
      LAYER met2 ;
        RECT 208.565 3111.465 210.965 3111.745 ;
      LAYER met2 ;
        RECT 0.000 3109.265 208.565 3111.185 ;
        RECT 0.000 3108.425 208.285 3109.265 ;
        RECT 0.000 3106.045 208.565 3108.425 ;
        RECT 0.000 3105.205 208.285 3106.045 ;
        RECT 0.000 3102.825 208.565 3105.205 ;
        RECT 0.000 3101.985 208.285 3102.825 ;
        RECT 0.000 3100.065 208.565 3101.985 ;
        RECT 0.000 3099.225 208.285 3100.065 ;
        RECT 0.000 3096.845 208.565 3099.225 ;
      LAYER met2 ;
        RECT 211.300 3097.130 211.440 3135.750 ;
        RECT 209.000 3096.990 211.440 3097.130 ;
      LAYER met2 ;
        RECT 0.000 3096.005 208.285 3096.845 ;
      LAYER met2 ;
        RECT 209.000 3096.565 209.140 3096.990 ;
        RECT 208.565 3096.285 210.965 3096.565 ;
      LAYER met2 ;
        RECT 0.000 3093.625 208.565 3096.005 ;
        RECT 0.000 3092.785 208.285 3093.625 ;
        RECT 0.000 3090.405 208.565 3092.785 ;
      LAYER met2 ;
        RECT 212.220 3092.630 212.360 3303.790 ;
        RECT 213.140 3125.610 213.280 3342.550 ;
        RECT 213.540 3293.250 213.800 3293.570 ;
        RECT 213.080 3125.290 213.340 3125.610 ;
        RECT 208.940 3092.310 209.200 3092.630 ;
        RECT 212.160 3092.310 212.420 3092.630 ;
      LAYER met2 ;
        RECT 0.000 3089.565 208.285 3090.405 ;
      LAYER met2 ;
        RECT 209.000 3090.125 209.140 3092.310 ;
        RECT 208.565 3089.845 210.965 3090.125 ;
      LAYER met2 ;
        RECT 0.000 3087.645 208.565 3089.565 ;
        RECT 0.000 3086.805 208.285 3087.645 ;
        RECT 0.000 3084.425 208.565 3086.805 ;
        RECT 0.000 3083.585 208.285 3084.425 ;
        RECT 0.000 3081.205 208.565 3083.585 ;
        RECT 0.000 3080.365 208.285 3081.205 ;
        RECT 0.000 3078.445 208.565 3080.365 ;
        RECT 0.000 3077.605 208.285 3078.445 ;
        RECT 0.000 3075.225 208.565 3077.605 ;
        RECT 0.000 3074.385 208.285 3075.225 ;
      LAYER met2 ;
        RECT 211.300 3074.950 211.440 3075.105 ;
        RECT 208.565 3074.805 210.965 3074.945 ;
        RECT 208.540 3074.690 210.965 3074.805 ;
        RECT 211.240 3074.690 211.500 3074.950 ;
        RECT 208.540 3074.630 211.500 3074.690 ;
        RECT 208.540 3074.550 211.440 3074.630 ;
      LAYER met2 ;
        RECT 0.000 3072.005 208.565 3074.385 ;
        RECT 0.000 3071.165 208.285 3072.005 ;
        RECT 0.000 3069.245 208.565 3071.165 ;
        RECT 0.000 3068.405 208.285 3069.245 ;
        RECT 0.000 3066.025 208.565 3068.405 ;
        RECT 0.000 3065.185 208.285 3066.025 ;
        RECT 0.000 3062.805 208.565 3065.185 ;
        RECT 0.000 3061.965 208.285 3062.805 ;
        RECT 0.000 3060.045 208.565 3061.965 ;
        RECT 0.000 3059.205 208.285 3060.045 ;
      LAYER met2 ;
        RECT 208.565 3059.485 210.965 3059.765 ;
      LAYER met2 ;
        RECT 0.000 3058.210 208.565 3059.205 ;
        RECT 0.000 2920.865 208.565 2921.915 ;
        RECT 0.000 2920.025 208.285 2920.865 ;
      LAYER met2 ;
        RECT 208.565 2920.305 210.965 2920.585 ;
      LAYER met2 ;
        RECT 0.000 2917.645 208.565 2920.025 ;
      LAYER met2 ;
        RECT 209.000 2917.870 209.140 2920.305 ;
      LAYER met2 ;
        RECT 0.000 2916.805 208.285 2917.645 ;
      LAYER met2 ;
        RECT 208.940 2917.550 209.200 2917.870 ;
      LAYER met2 ;
        RECT 0.000 2914.425 208.565 2916.805 ;
        RECT 0.000 2913.585 208.285 2914.425 ;
      LAYER met2 ;
        RECT 208.565 2913.865 210.965 2914.145 ;
      LAYER met2 ;
        RECT 0.000 2911.665 208.565 2913.585 ;
        RECT 0.000 2910.825 208.285 2911.665 ;
      LAYER met2 ;
        RECT 208.565 2911.105 210.965 2911.385 ;
      LAYER met2 ;
        RECT 0.000 2908.445 208.565 2910.825 ;
      LAYER met2 ;
        RECT 209.000 2909.370 209.140 2911.105 ;
        RECT 208.940 2909.050 209.200 2909.370 ;
      LAYER met2 ;
        RECT 0.000 2907.605 208.285 2908.445 ;
        RECT 0.000 2905.225 208.565 2907.605 ;
        RECT 0.000 2904.385 208.285 2905.225 ;
        RECT 0.000 2902.465 208.565 2904.385 ;
        RECT 0.000 2901.625 208.285 2902.465 ;
      LAYER met2 ;
        RECT 208.565 2901.905 210.965 2902.185 ;
      LAYER met2 ;
        RECT 0.000 2899.245 208.565 2901.625 ;
        RECT 0.000 2898.405 208.285 2899.245 ;
        RECT 0.000 2896.025 208.565 2898.405 ;
        RECT 0.000 2895.185 208.285 2896.025 ;
      LAYER met2 ;
        RECT 208.565 2895.465 210.965 2895.745 ;
      LAYER met2 ;
        RECT 0.000 2893.265 208.565 2895.185 ;
        RECT 0.000 2892.425 208.285 2893.265 ;
        RECT 0.000 2890.045 208.565 2892.425 ;
        RECT 0.000 2889.205 208.285 2890.045 ;
        RECT 0.000 2886.825 208.565 2889.205 ;
        RECT 0.000 2885.985 208.285 2886.825 ;
        RECT 0.000 2884.065 208.565 2885.985 ;
        RECT 0.000 2883.225 208.285 2884.065 ;
        RECT 0.000 2880.845 208.565 2883.225 ;
      LAYER met2 ;
        RECT 208.940 2882.190 209.200 2882.510 ;
      LAYER met2 ;
        RECT 0.000 2880.005 208.285 2880.845 ;
      LAYER met2 ;
        RECT 209.000 2880.565 209.140 2882.190 ;
        RECT 211.300 2881.490 211.440 3074.550 ;
        RECT 212.220 3052.930 212.360 3092.310 ;
        RECT 213.140 3054.290 213.280 3125.290 ;
        RECT 213.600 3074.950 213.740 3293.250 ;
        RECT 213.540 3074.630 213.800 3074.950 ;
        RECT 213.140 3054.150 213.740 3054.290 ;
        RECT 212.220 3052.790 213.280 3052.930 ;
        RECT 212.620 3029.070 212.880 3029.390 ;
        RECT 212.160 2917.550 212.420 2917.870 ;
        RECT 212.220 2882.510 212.360 2917.550 ;
        RECT 212.680 2909.370 212.820 3029.070 ;
        RECT 212.620 2909.050 212.880 2909.370 ;
        RECT 212.160 2882.190 212.420 2882.510 ;
        RECT 211.240 2881.170 211.500 2881.490 ;
        RECT 208.565 2880.285 210.965 2880.565 ;
      LAYER met2 ;
        RECT 0.000 2877.625 208.565 2880.005 ;
        RECT 0.000 2876.785 208.285 2877.625 ;
        RECT 0.000 2874.405 208.565 2876.785 ;
        RECT 0.000 2873.565 208.285 2874.405 ;
      LAYER met2 ;
        RECT 208.565 2873.845 210.965 2874.125 ;
      LAYER met2 ;
        RECT 0.000 2871.645 208.565 2873.565 ;
      LAYER met2 ;
        RECT 209.000 2871.970 209.140 2873.845 ;
        RECT 208.940 2871.650 209.200 2871.970 ;
        RECT 212.160 2871.650 212.420 2871.970 ;
      LAYER met2 ;
        RECT 0.000 2870.805 208.285 2871.645 ;
        RECT 0.000 2868.425 208.565 2870.805 ;
        RECT 0.000 2867.585 208.285 2868.425 ;
        RECT 0.000 2865.205 208.565 2867.585 ;
        RECT 0.000 2864.365 208.285 2865.205 ;
        RECT 0.000 2862.445 208.565 2864.365 ;
        RECT 0.000 2861.605 208.285 2862.445 ;
        RECT 0.000 2859.225 208.565 2861.605 ;
        RECT 0.000 2858.385 208.285 2859.225 ;
      LAYER met2 ;
        RECT 208.565 2858.665 210.965 2858.945 ;
      LAYER met2 ;
        RECT 0.000 2856.005 208.565 2858.385 ;
      LAYER met2 ;
        RECT 209.000 2858.370 209.140 2858.665 ;
        RECT 208.940 2858.050 209.200 2858.370 ;
      LAYER met2 ;
        RECT 0.000 2855.165 208.285 2856.005 ;
        RECT 0.000 2853.245 208.565 2855.165 ;
        RECT 0.000 2852.405 208.285 2853.245 ;
        RECT 0.000 2850.025 208.565 2852.405 ;
        RECT 0.000 2849.185 208.285 2850.025 ;
        RECT 0.000 2846.805 208.565 2849.185 ;
        RECT 0.000 2845.965 208.285 2846.805 ;
        RECT 0.000 2844.045 208.565 2845.965 ;
        RECT 0.000 2843.205 208.285 2844.045 ;
      LAYER met2 ;
        RECT 208.565 2843.485 210.965 2843.765 ;
      LAYER met2 ;
        RECT 0.000 2842.210 208.565 2843.205 ;
        RECT 0.000 2704.865 208.565 2705.915 ;
        RECT 0.000 2704.025 208.285 2704.865 ;
      LAYER met2 ;
        RECT 208.565 2704.515 210.965 2704.585 ;
        RECT 208.565 2704.375 211.440 2704.515 ;
        RECT 208.565 2704.305 210.965 2704.375 ;
      LAYER met2 ;
        RECT 0.000 2701.645 208.565 2704.025 ;
        RECT 0.000 2700.805 208.285 2701.645 ;
        RECT 0.000 2698.425 208.565 2700.805 ;
        RECT 0.000 2697.585 208.285 2698.425 ;
      LAYER met2 ;
        RECT 208.565 2697.865 210.965 2698.145 ;
      LAYER met2 ;
        RECT 0.000 2695.665 208.565 2697.585 ;
        RECT 0.000 2694.825 208.285 2695.665 ;
      LAYER met2 ;
        RECT 208.940 2695.530 209.200 2695.850 ;
        RECT 209.000 2695.385 209.140 2695.530 ;
        RECT 208.565 2695.105 210.965 2695.385 ;
      LAYER met2 ;
        RECT 0.000 2692.445 208.565 2694.825 ;
        RECT 0.000 2691.605 208.285 2692.445 ;
        RECT 0.000 2689.225 208.565 2691.605 ;
        RECT 0.000 2688.385 208.285 2689.225 ;
        RECT 0.000 2686.465 208.565 2688.385 ;
        RECT 0.000 2685.625 208.285 2686.465 ;
      LAYER met2 ;
        RECT 208.565 2685.905 210.965 2686.185 ;
      LAYER met2 ;
        RECT 0.000 2683.245 208.565 2685.625 ;
        RECT 0.000 2682.405 208.285 2683.245 ;
        RECT 0.000 2680.025 208.565 2682.405 ;
        RECT 0.000 2679.185 208.285 2680.025 ;
      LAYER met2 ;
        RECT 208.565 2679.465 210.965 2679.745 ;
      LAYER met2 ;
        RECT 0.000 2677.265 208.565 2679.185 ;
        RECT 0.000 2676.425 208.285 2677.265 ;
        RECT 0.000 2674.045 208.565 2676.425 ;
        RECT 0.000 2673.205 208.285 2674.045 ;
        RECT 0.000 2670.825 208.565 2673.205 ;
        RECT 0.000 2669.985 208.285 2670.825 ;
        RECT 0.000 2668.065 208.565 2669.985 ;
        RECT 0.000 2667.225 208.285 2668.065 ;
        RECT 0.000 2664.845 208.565 2667.225 ;
      LAYER met2 ;
        RECT 211.300 2666.690 211.440 2704.375 ;
        RECT 209.000 2666.550 211.440 2666.690 ;
      LAYER met2 ;
        RECT 0.000 2664.005 208.285 2664.845 ;
      LAYER met2 ;
        RECT 209.000 2664.565 209.140 2666.550 ;
        RECT 208.565 2664.285 210.965 2664.565 ;
      LAYER met2 ;
        RECT 0.000 2661.625 208.565 2664.005 ;
        RECT 0.000 2660.785 208.285 2661.625 ;
      LAYER met2 ;
        RECT 212.220 2660.830 212.360 2871.650 ;
        RECT 212.680 2695.850 212.820 2909.050 ;
        RECT 213.140 2871.970 213.280 3052.790 ;
        RECT 213.600 3029.390 213.740 3054.150 ;
        RECT 213.540 3029.070 213.800 3029.390 ;
        RECT 213.540 2881.170 213.800 2881.490 ;
        RECT 213.080 2871.650 213.340 2871.970 ;
        RECT 213.600 2871.370 213.740 2881.170 ;
        RECT 213.140 2871.230 213.740 2871.370 ;
        RECT 213.140 2858.370 213.280 2871.230 ;
        RECT 213.080 2858.050 213.340 2858.370 ;
        RECT 212.620 2695.530 212.880 2695.850 ;
      LAYER met2 ;
        RECT 0.000 2658.405 208.565 2660.785 ;
      LAYER met2 ;
        RECT 208.940 2660.510 209.200 2660.830 ;
        RECT 212.160 2660.510 212.420 2660.830 ;
      LAYER met2 ;
        RECT 0.000 2657.565 208.285 2658.405 ;
      LAYER met2 ;
        RECT 209.000 2658.125 209.140 2660.510 ;
        RECT 208.565 2657.845 210.965 2658.125 ;
      LAYER met2 ;
        RECT 0.000 2655.645 208.565 2657.565 ;
        RECT 0.000 2654.805 208.285 2655.645 ;
        RECT 0.000 2652.425 208.565 2654.805 ;
        RECT 0.000 2651.585 208.285 2652.425 ;
        RECT 0.000 2649.205 208.565 2651.585 ;
        RECT 0.000 2648.365 208.285 2649.205 ;
        RECT 0.000 2646.445 208.565 2648.365 ;
        RECT 0.000 2645.605 208.285 2646.445 ;
        RECT 0.000 2643.225 208.565 2645.605 ;
        RECT 0.000 2642.385 208.285 2643.225 ;
      LAYER met2 ;
        RECT 208.565 2642.820 210.965 2642.945 ;
        RECT 208.540 2642.665 210.965 2642.820 ;
        RECT 208.540 2642.630 210.060 2642.665 ;
        RECT 209.920 2642.470 210.060 2642.630 ;
      LAYER met2 ;
        RECT 0.000 2640.005 208.565 2642.385 ;
      LAYER met2 ;
        RECT 209.860 2642.150 210.120 2642.470 ;
      LAYER met2 ;
        RECT 0.000 2639.165 208.285 2640.005 ;
        RECT 0.000 2637.245 208.565 2639.165 ;
        RECT 0.000 2636.405 208.285 2637.245 ;
        RECT 0.000 2634.025 208.565 2636.405 ;
        RECT 0.000 2633.185 208.285 2634.025 ;
        RECT 0.000 2630.805 208.565 2633.185 ;
        RECT 0.000 2629.965 208.285 2630.805 ;
        RECT 0.000 2628.045 208.565 2629.965 ;
        RECT 0.000 2627.205 208.285 2628.045 ;
      LAYER met2 ;
        RECT 208.565 2627.485 210.965 2627.765 ;
      LAYER met2 ;
        RECT 0.000 2626.210 208.565 2627.205 ;
        RECT 4.925 2465.390 200.000 2489.290 ;
        RECT 4.925 2439.395 197.965 2465.390 ;
        RECT 198.080 2440.895 200.000 2442.895 ;
        RECT 4.925 2415.495 200.000 2439.395 ;
        RECT 4.925 2415.265 197.965 2415.495 ;
        RECT 0.035 2280.200 151.405 2289.935 ;
        RECT 153.765 2279.000 158.415 2290.140 ;
        RECT 160.165 2280.200 174.575 2289.935 ;
        RECT 0.035 2278.700 197.965 2279.000 ;
        RECT 0.035 2258.095 198.000 2278.700 ;
        RECT 0.035 2257.535 197.965 2258.095 ;
        RECT 0.035 2224.925 198.000 2257.535 ;
        RECT 0.035 2224.495 197.965 2224.925 ;
        RECT 0.035 2204.500 198.000 2224.495 ;
        RECT 0.035 2204.000 197.965 2204.500 ;
        RECT 153.800 2193.025 158.450 2204.000 ;
        RECT 0.000 2066.865 208.565 2067.915 ;
        RECT 0.000 2066.025 208.285 2066.865 ;
      LAYER met2 ;
        RECT 208.565 2066.305 210.965 2066.585 ;
      LAYER met2 ;
        RECT 0.000 2063.645 208.565 2066.025 ;
      LAYER met2 ;
        RECT 209.000 2064.810 209.140 2066.305 ;
        RECT 208.940 2064.490 209.200 2064.810 ;
        RECT 211.700 2064.490 211.960 2064.810 ;
      LAYER met2 ;
        RECT 0.000 2062.805 208.285 2063.645 ;
        RECT 0.000 2060.425 208.565 2062.805 ;
        RECT 0.000 2059.585 208.285 2060.425 ;
      LAYER met2 ;
        RECT 208.565 2059.865 210.965 2060.145 ;
      LAYER met2 ;
        RECT 0.000 2057.665 208.565 2059.585 ;
        RECT 0.000 2056.825 208.285 2057.665 ;
      LAYER met2 ;
        RECT 208.610 2057.385 209.140 2057.410 ;
        RECT 208.565 2057.105 210.965 2057.385 ;
      LAYER met2 ;
        RECT 0.000 2054.445 208.565 2056.825 ;
      LAYER met2 ;
        RECT 209.000 2054.950 209.140 2057.105 ;
        RECT 208.940 2054.630 209.200 2054.950 ;
      LAYER met2 ;
        RECT 0.000 2053.605 208.285 2054.445 ;
        RECT 0.000 2051.225 208.565 2053.605 ;
        RECT 0.000 2050.385 208.285 2051.225 ;
        RECT 0.000 2048.465 208.565 2050.385 ;
        RECT 0.000 2047.625 208.285 2048.465 ;
      LAYER met2 ;
        RECT 208.565 2047.905 210.965 2048.185 ;
      LAYER met2 ;
        RECT 0.000 2045.245 208.565 2047.625 ;
        RECT 0.000 2044.405 208.285 2045.245 ;
        RECT 0.000 2042.025 208.565 2044.405 ;
        RECT 0.000 2041.185 208.285 2042.025 ;
      LAYER met2 ;
        RECT 208.565 2041.465 210.965 2041.745 ;
      LAYER met2 ;
        RECT 0.000 2039.265 208.565 2041.185 ;
        RECT 0.000 2038.425 208.285 2039.265 ;
        RECT 0.000 2036.045 208.565 2038.425 ;
        RECT 0.000 2035.205 208.285 2036.045 ;
        RECT 0.000 2032.825 208.565 2035.205 ;
        RECT 0.000 2031.985 208.285 2032.825 ;
        RECT 0.000 2030.065 208.565 2031.985 ;
        RECT 0.000 2029.225 208.285 2030.065 ;
        RECT 0.000 2026.845 208.565 2029.225 ;
      LAYER met2 ;
        RECT 211.760 2029.110 211.900 2064.490 ;
        RECT 208.940 2028.790 209.200 2029.110 ;
        RECT 211.700 2028.790 211.960 2029.110 ;
      LAYER met2 ;
        RECT 0.000 2026.005 208.285 2026.845 ;
      LAYER met2 ;
        RECT 209.000 2026.565 209.140 2028.790 ;
        RECT 208.565 2026.285 210.965 2026.565 ;
      LAYER met2 ;
        RECT 0.000 2023.625 208.565 2026.005 ;
        RECT 0.000 2022.785 208.285 2023.625 ;
        RECT 0.000 2020.405 208.565 2022.785 ;
      LAYER met2 ;
        RECT 212.220 2022.650 212.360 2660.510 ;
        RECT 212.680 2111.470 212.820 2695.530 ;
        RECT 213.140 2691.070 213.280 2858.050 ;
        RECT 213.140 2690.930 213.740 2691.070 ;
        RECT 213.600 2642.470 213.740 2690.930 ;
        RECT 213.540 2642.150 213.800 2642.470 ;
        RECT 212.680 2111.330 213.280 2111.470 ;
        RECT 213.140 2054.950 213.280 2111.330 ;
        RECT 213.080 2054.630 213.340 2054.950 ;
        RECT 208.940 2022.330 209.200 2022.650 ;
        RECT 212.160 2022.330 212.420 2022.650 ;
      LAYER met2 ;
        RECT 0.000 2019.565 208.285 2020.405 ;
      LAYER met2 ;
        RECT 209.000 2020.125 209.140 2022.330 ;
        RECT 208.565 2019.845 210.965 2020.125 ;
      LAYER met2 ;
        RECT 0.000 2017.645 208.565 2019.565 ;
        RECT 0.000 2016.805 208.285 2017.645 ;
        RECT 0.000 2014.425 208.565 2016.805 ;
      LAYER met2 ;
        RECT 212.220 2014.870 212.360 2022.330 ;
        RECT 212.220 2014.730 212.820 2014.870 ;
      LAYER met2 ;
        RECT 0.000 2013.585 208.285 2014.425 ;
        RECT 0.000 2011.205 208.565 2013.585 ;
        RECT 0.000 2010.365 208.285 2011.205 ;
        RECT 0.000 2008.445 208.565 2010.365 ;
        RECT 0.000 2007.605 208.285 2008.445 ;
        RECT 0.000 2005.225 208.565 2007.605 ;
        RECT 0.000 2004.385 208.285 2005.225 ;
      LAYER met2 ;
        RECT 208.565 2004.665 210.965 2004.945 ;
      LAYER met2 ;
        RECT 0.000 2002.005 208.565 2004.385 ;
      LAYER met2 ;
        RECT 209.000 2002.250 209.140 2004.665 ;
      LAYER met2 ;
        RECT 0.000 2001.165 208.285 2002.005 ;
      LAYER met2 ;
        RECT 208.940 2001.930 209.200 2002.250 ;
        RECT 212.160 2001.930 212.420 2002.250 ;
      LAYER met2 ;
        RECT 0.000 1999.245 208.565 2001.165 ;
        RECT 0.000 1998.405 208.285 1999.245 ;
        RECT 0.000 1996.025 208.565 1998.405 ;
        RECT 0.000 1995.185 208.285 1996.025 ;
        RECT 0.000 1992.805 208.565 1995.185 ;
        RECT 0.000 1991.965 208.285 1992.805 ;
        RECT 0.000 1990.045 208.565 1991.965 ;
        RECT 0.000 1989.205 208.285 1990.045 ;
      LAYER met2 ;
        RECT 208.565 1989.485 210.965 1989.765 ;
      LAYER met2 ;
        RECT 0.000 1988.210 208.565 1989.205 ;
        RECT 0.000 1850.865 208.565 1851.915 ;
        RECT 0.000 1850.025 208.285 1850.865 ;
      LAYER met2 ;
        RECT 208.565 1850.305 210.965 1850.585 ;
      LAYER met2 ;
        RECT 0.000 1847.645 208.565 1850.025 ;
      LAYER met2 ;
        RECT 209.000 1847.890 209.140 1850.305 ;
      LAYER met2 ;
        RECT 0.000 1846.805 208.285 1847.645 ;
      LAYER met2 ;
        RECT 208.940 1847.570 209.200 1847.890 ;
        RECT 211.700 1847.570 211.960 1847.890 ;
      LAYER met2 ;
        RECT 0.000 1844.425 208.565 1846.805 ;
        RECT 0.000 1843.585 208.285 1844.425 ;
      LAYER met2 ;
        RECT 208.565 1843.865 210.965 1844.145 ;
      LAYER met2 ;
        RECT 0.000 1841.665 208.565 1843.585 ;
      LAYER met2 ;
        RECT 208.940 1843.150 209.200 1843.470 ;
      LAYER met2 ;
        RECT 0.000 1840.825 208.285 1841.665 ;
      LAYER met2 ;
        RECT 209.000 1841.385 209.140 1843.150 ;
        RECT 208.565 1841.105 210.965 1841.385 ;
      LAYER met2 ;
        RECT 0.000 1838.445 208.565 1840.825 ;
        RECT 0.000 1837.605 208.285 1838.445 ;
        RECT 0.000 1835.225 208.565 1837.605 ;
        RECT 0.000 1834.385 208.285 1835.225 ;
        RECT 0.000 1832.465 208.565 1834.385 ;
        RECT 0.000 1831.625 208.285 1832.465 ;
      LAYER met2 ;
        RECT 208.565 1831.905 210.965 1832.185 ;
      LAYER met2 ;
        RECT 0.000 1829.245 208.565 1831.625 ;
        RECT 0.000 1828.405 208.285 1829.245 ;
        RECT 0.000 1826.025 208.565 1828.405 ;
        RECT 0.000 1825.185 208.285 1826.025 ;
      LAYER met2 ;
        RECT 208.565 1825.465 210.965 1825.745 ;
      LAYER met2 ;
        RECT 0.000 1823.265 208.565 1825.185 ;
        RECT 0.000 1822.425 208.285 1823.265 ;
        RECT 0.000 1820.045 208.565 1822.425 ;
        RECT 0.000 1819.205 208.285 1820.045 ;
        RECT 0.000 1816.825 208.565 1819.205 ;
        RECT 0.000 1815.985 208.285 1816.825 ;
        RECT 0.000 1814.065 208.565 1815.985 ;
        RECT 0.000 1813.225 208.285 1814.065 ;
        RECT 0.000 1810.845 208.565 1813.225 ;
      LAYER met2 ;
        RECT 211.760 1813.210 211.900 1847.570 ;
        RECT 208.940 1812.890 209.200 1813.210 ;
        RECT 211.700 1812.890 211.960 1813.210 ;
      LAYER met2 ;
        RECT 0.000 1810.005 208.285 1810.845 ;
      LAYER met2 ;
        RECT 209.000 1810.570 209.140 1812.890 ;
        RECT 208.610 1810.565 209.140 1810.570 ;
        RECT 208.565 1810.285 210.965 1810.565 ;
      LAYER met2 ;
        RECT 0.000 1807.625 208.565 1810.005 ;
        RECT 0.000 1806.785 208.285 1807.625 ;
        RECT 0.000 1804.405 208.565 1806.785 ;
        RECT 0.000 1803.565 208.285 1804.405 ;
      LAYER met2 ;
        RECT 208.565 1803.845 210.965 1804.125 ;
      LAYER met2 ;
        RECT 0.000 1801.645 208.565 1803.565 ;
      LAYER met2 ;
        RECT 209.000 1801.990 209.140 1803.845 ;
        RECT 208.940 1801.670 209.200 1801.990 ;
      LAYER met2 ;
        RECT 0.000 1800.805 208.285 1801.645 ;
        RECT 0.000 1798.425 208.565 1800.805 ;
        RECT 0.000 1797.585 208.285 1798.425 ;
        RECT 0.000 1795.205 208.565 1797.585 ;
        RECT 0.000 1794.365 208.285 1795.205 ;
        RECT 0.000 1792.445 208.565 1794.365 ;
        RECT 0.000 1791.605 208.285 1792.445 ;
        RECT 0.000 1789.225 208.565 1791.605 ;
        RECT 0.000 1788.385 208.285 1789.225 ;
      LAYER met2 ;
        RECT 208.565 1788.665 210.965 1788.945 ;
      LAYER met2 ;
        RECT 0.000 1786.005 208.565 1788.385 ;
      LAYER met2 ;
        RECT 209.000 1786.350 209.140 1788.665 ;
        RECT 212.220 1786.350 212.360 2001.930 ;
        RECT 212.680 1801.990 212.820 2014.730 ;
        RECT 213.140 1843.470 213.280 2054.630 ;
        RECT 213.600 2002.250 213.740 2642.150 ;
        RECT 3370.580 2139.270 3370.720 4950.410 ;
        RECT 3371.040 4766.790 3371.180 4965.370 ;
        RECT 3371.440 4965.030 3371.700 4965.350 ;
        RECT 3371.500 4820.850 3371.640 4965.030 ;
        RECT 3375.580 4964.350 3375.840 4964.670 ;
        RECT 3375.640 4912.870 3375.780 4964.350 ;
        RECT 3375.640 4912.730 3376.700 4912.870 ;
        RECT 3376.560 4821.265 3376.700 4912.730 ;
      LAYER met2 ;
        RECT 3379.435 4836.795 3588.000 4837.790 ;
      LAYER met2 ;
        RECT 3377.035 4836.235 3379.435 4836.515 ;
      LAYER met2 ;
        RECT 3379.715 4835.955 3588.000 4836.795 ;
        RECT 3379.435 4834.035 3588.000 4835.955 ;
        RECT 3379.715 4833.195 3588.000 4834.035 ;
        RECT 3379.435 4830.815 3588.000 4833.195 ;
        RECT 3379.715 4829.975 3588.000 4830.815 ;
        RECT 3379.435 4827.595 3588.000 4829.975 ;
        RECT 3379.715 4826.755 3588.000 4827.595 ;
        RECT 3379.435 4824.835 3588.000 4826.755 ;
        RECT 3379.715 4823.995 3588.000 4824.835 ;
        RECT 3379.435 4821.615 3588.000 4823.995 ;
      LAYER met2 ;
        RECT 3377.035 4821.265 3379.435 4821.335 ;
        RECT 3376.100 4821.125 3379.435 4821.265 ;
        RECT 3371.440 4820.530 3371.700 4820.850 ;
        RECT 3374.660 4803.190 3374.920 4803.510 ;
        RECT 3370.980 4766.470 3371.240 4766.790 ;
        RECT 3374.200 4372.410 3374.460 4372.730 ;
        RECT 3374.260 3926.650 3374.400 4372.410 ;
        RECT 3374.720 4358.530 3374.860 4803.190 ;
        RECT 3376.100 4801.130 3376.240 4821.125 ;
        RECT 3377.035 4821.055 3379.435 4821.125 ;
        RECT 3376.500 4820.530 3376.760 4820.850 ;
      LAYER met2 ;
        RECT 3379.715 4820.775 3588.000 4821.615 ;
      LAYER met2 ;
        RECT 3376.560 4805.970 3376.700 4820.530 ;
      LAYER met2 ;
        RECT 3379.435 4818.395 3588.000 4820.775 ;
        RECT 3379.715 4817.555 3588.000 4818.395 ;
        RECT 3379.435 4815.635 3588.000 4817.555 ;
        RECT 3379.715 4814.795 3588.000 4815.635 ;
        RECT 3379.435 4812.415 3588.000 4814.795 ;
        RECT 3379.715 4811.575 3588.000 4812.415 ;
        RECT 3379.435 4809.195 3588.000 4811.575 ;
        RECT 3379.715 4808.355 3588.000 4809.195 ;
        RECT 3379.435 4806.435 3588.000 4808.355 ;
      LAYER met2 ;
        RECT 3377.035 4805.970 3379.435 4806.155 ;
        RECT 3376.560 4805.875 3379.435 4805.970 ;
        RECT 3376.560 4805.830 3377.160 4805.875 ;
        RECT 3377.020 4803.510 3377.160 4805.830 ;
      LAYER met2 ;
        RECT 3379.715 4805.595 3588.000 4806.435 ;
      LAYER met2 ;
        RECT 3376.960 4803.190 3377.220 4803.510 ;
      LAYER met2 ;
        RECT 3379.435 4803.215 3588.000 4805.595 ;
        RECT 3379.715 4802.375 3588.000 4803.215 ;
      LAYER met2 ;
        RECT 3376.040 4800.810 3376.300 4801.130 ;
        RECT 3376.040 4799.790 3376.300 4800.110 ;
      LAYER met2 ;
        RECT 3379.435 4799.995 3588.000 4802.375 ;
      LAYER met2 ;
        RECT 3375.580 4766.470 3375.840 4766.790 ;
        RECT 3374.720 4358.450 3375.320 4358.530 ;
        RECT 3374.720 4358.390 3375.380 4358.450 ;
        RECT 3375.120 4358.130 3375.380 4358.390 ;
        RECT 3374.660 4320.390 3374.920 4320.710 ;
        RECT 3374.200 3926.330 3374.460 3926.650 ;
        RECT 3374.260 3701.910 3374.400 3926.330 ;
        RECT 3374.720 3875.310 3374.860 4320.390 ;
        RECT 3375.180 3916.450 3375.320 4358.130 ;
        RECT 3375.640 4320.710 3375.780 4766.470 ;
        RECT 3376.100 4372.730 3376.240 4799.790 ;
        RECT 3377.035 4799.645 3379.435 4799.715 ;
        RECT 3376.560 4799.505 3379.435 4799.645 ;
        RECT 3376.560 4759.050 3376.700 4799.505 ;
        RECT 3377.035 4799.435 3379.435 4799.505 ;
      LAYER met2 ;
        RECT 3379.715 4799.155 3588.000 4799.995 ;
        RECT 3379.435 4796.775 3588.000 4799.155 ;
        RECT 3379.715 4795.935 3588.000 4796.775 ;
        RECT 3379.435 4794.015 3588.000 4795.935 ;
        RECT 3379.715 4793.175 3588.000 4794.015 ;
        RECT 3379.435 4790.795 3588.000 4793.175 ;
        RECT 3379.715 4789.955 3588.000 4790.795 ;
        RECT 3379.435 4787.575 3588.000 4789.955 ;
        RECT 3379.715 4786.735 3588.000 4787.575 ;
        RECT 3379.435 4784.815 3588.000 4786.735 ;
      LAYER met2 ;
        RECT 3377.035 4784.255 3379.435 4784.535 ;
      LAYER met2 ;
        RECT 3379.715 4783.975 3588.000 4784.815 ;
        RECT 3379.435 4781.595 3588.000 4783.975 ;
        RECT 3379.715 4780.755 3588.000 4781.595 ;
        RECT 3379.435 4778.375 3588.000 4780.755 ;
      LAYER met2 ;
        RECT 3377.035 4777.815 3379.435 4778.095 ;
      LAYER met2 ;
        RECT 3379.715 4777.535 3588.000 4778.375 ;
        RECT 3379.435 4775.615 3588.000 4777.535 ;
        RECT 3379.715 4774.775 3588.000 4775.615 ;
        RECT 3379.435 4772.395 3588.000 4774.775 ;
        RECT 3379.715 4771.555 3588.000 4772.395 ;
        RECT 3379.435 4769.175 3588.000 4771.555 ;
      LAYER met2 ;
        RECT 3377.035 4768.755 3379.435 4768.895 ;
        RECT 3377.020 4768.615 3379.435 4768.755 ;
        RECT 3377.020 4767.970 3377.160 4768.615 ;
      LAYER met2 ;
        RECT 3379.715 4768.335 3588.000 4769.175 ;
      LAYER met2 ;
        RECT 3377.020 4767.830 3378.080 4767.970 ;
        RECT 3377.940 4766.790 3378.080 4767.830 ;
        RECT 3377.880 4766.470 3378.140 4766.790 ;
      LAYER met2 ;
        RECT 3379.435 4766.415 3588.000 4768.335 ;
      LAYER met2 ;
        RECT 3377.035 4765.855 3379.435 4766.135 ;
      LAYER met2 ;
        RECT 3379.715 4765.575 3588.000 4766.415 ;
        RECT 3379.435 4763.195 3588.000 4765.575 ;
        RECT 3379.715 4762.355 3588.000 4763.195 ;
        RECT 3379.435 4759.975 3588.000 4762.355 ;
      LAYER met2 ;
        RECT 3377.035 4759.660 3379.435 4759.695 ;
        RECT 3377.020 4759.415 3379.435 4759.660 ;
        RECT 3377.020 4759.050 3377.160 4759.415 ;
      LAYER met2 ;
        RECT 3379.715 4759.135 3588.000 4759.975 ;
      LAYER met2 ;
        RECT 3376.560 4758.910 3377.160 4759.050 ;
      LAYER met2 ;
        RECT 3379.435 4758.085 3588.000 4759.135 ;
        RECT 3429.550 4613.000 3434.200 4623.975 ;
        RECT 3390.035 4612.500 3587.965 4613.000 ;
        RECT 3390.000 4592.505 3587.965 4612.500 ;
        RECT 3390.035 4592.075 3587.965 4592.505 ;
        RECT 3390.000 4559.465 3587.965 4592.075 ;
        RECT 3390.035 4558.905 3587.965 4559.465 ;
        RECT 3390.000 4538.300 3587.965 4558.905 ;
        RECT 3390.035 4538.000 3587.965 4538.300 ;
        RECT 3413.425 4527.065 3427.835 4536.800 ;
        RECT 3429.585 4526.860 3434.235 4538.000 ;
        RECT 3436.595 4527.065 3587.965 4536.800 ;
        RECT 3379.435 4390.795 3588.000 4391.790 ;
      LAYER met2 ;
        RECT 3377.035 4390.235 3379.435 4390.515 ;
      LAYER met2 ;
        RECT 3379.715 4389.955 3588.000 4390.795 ;
        RECT 3379.435 4388.035 3588.000 4389.955 ;
        RECT 3379.715 4387.195 3588.000 4388.035 ;
        RECT 3379.435 4384.815 3588.000 4387.195 ;
        RECT 3379.715 4383.975 3588.000 4384.815 ;
        RECT 3379.435 4381.595 3588.000 4383.975 ;
        RECT 3379.715 4380.755 3588.000 4381.595 ;
        RECT 3379.435 4378.835 3588.000 4380.755 ;
        RECT 3379.715 4377.995 3588.000 4378.835 ;
        RECT 3379.435 4375.615 3588.000 4377.995 ;
      LAYER met2 ;
        RECT 3377.035 4375.195 3379.435 4375.335 ;
        RECT 3377.020 4375.055 3379.435 4375.195 ;
        RECT 3377.020 4372.730 3377.160 4375.055 ;
      LAYER met2 ;
        RECT 3379.715 4374.775 3588.000 4375.615 ;
      LAYER met2 ;
        RECT 3376.040 4372.410 3376.300 4372.730 ;
        RECT 3376.960 4372.410 3377.220 4372.730 ;
      LAYER met2 ;
        RECT 3379.435 4372.395 3588.000 4374.775 ;
        RECT 3379.715 4371.555 3588.000 4372.395 ;
        RECT 3379.435 4369.635 3588.000 4371.555 ;
        RECT 3379.715 4368.795 3588.000 4369.635 ;
        RECT 3379.435 4366.415 3588.000 4368.795 ;
        RECT 3379.715 4365.575 3588.000 4366.415 ;
        RECT 3379.435 4363.195 3588.000 4365.575 ;
        RECT 3379.715 4362.355 3588.000 4363.195 ;
        RECT 3379.435 4360.435 3588.000 4362.355 ;
      LAYER met2 ;
        RECT 3377.035 4360.015 3379.435 4360.155 ;
        RECT 3377.020 4359.875 3379.435 4360.015 ;
        RECT 3377.020 4358.450 3377.160 4359.875 ;
      LAYER met2 ;
        RECT 3379.715 4359.595 3588.000 4360.435 ;
      LAYER met2 ;
        RECT 3376.960 4358.130 3377.220 4358.450 ;
      LAYER met2 ;
        RECT 3379.435 4357.215 3588.000 4359.595 ;
        RECT 3379.715 4356.375 3588.000 4357.215 ;
        RECT 3379.435 4353.995 3588.000 4356.375 ;
      LAYER met2 ;
        RECT 3377.035 4353.700 3379.435 4353.715 ;
        RECT 3377.020 4353.435 3379.435 4353.700 ;
        RECT 3377.020 4351.050 3377.160 4353.435 ;
      LAYER met2 ;
        RECT 3379.715 4353.155 3588.000 4353.995 ;
      LAYER met2 ;
        RECT 3376.560 4350.910 3377.160 4351.050 ;
        RECT 3375.580 4320.390 3375.840 4320.710 ;
        RECT 3376.560 4313.650 3376.700 4350.910 ;
      LAYER met2 ;
        RECT 3379.435 4350.775 3588.000 4353.155 ;
        RECT 3379.715 4349.935 3588.000 4350.775 ;
        RECT 3379.435 4348.015 3588.000 4349.935 ;
        RECT 3379.715 4347.175 3588.000 4348.015 ;
        RECT 3379.435 4344.795 3588.000 4347.175 ;
        RECT 3379.715 4343.955 3588.000 4344.795 ;
        RECT 3379.435 4341.575 3588.000 4343.955 ;
        RECT 3379.715 4340.735 3588.000 4341.575 ;
        RECT 3379.435 4338.815 3588.000 4340.735 ;
      LAYER met2 ;
        RECT 3377.035 4338.255 3379.435 4338.535 ;
      LAYER met2 ;
        RECT 3379.715 4337.975 3588.000 4338.815 ;
        RECT 3379.435 4335.595 3588.000 4337.975 ;
        RECT 3379.715 4334.755 3588.000 4335.595 ;
        RECT 3379.435 4332.375 3588.000 4334.755 ;
      LAYER met2 ;
        RECT 3377.035 4331.815 3379.435 4332.095 ;
      LAYER met2 ;
        RECT 3379.715 4331.535 3588.000 4332.375 ;
        RECT 3379.435 4329.615 3588.000 4331.535 ;
        RECT 3379.715 4328.775 3588.000 4329.615 ;
        RECT 3379.435 4326.395 3588.000 4328.775 ;
        RECT 3379.715 4325.555 3588.000 4326.395 ;
        RECT 3379.435 4323.175 3588.000 4325.555 ;
      LAYER met2 ;
        RECT 3377.035 4322.755 3379.435 4322.895 ;
        RECT 3377.020 4322.615 3379.435 4322.755 ;
        RECT 3377.020 4320.710 3377.160 4322.615 ;
      LAYER met2 ;
        RECT 3379.715 4322.335 3588.000 4323.175 ;
      LAYER met2 ;
        RECT 3376.960 4320.390 3377.220 4320.710 ;
      LAYER met2 ;
        RECT 3379.435 4320.415 3588.000 4322.335 ;
      LAYER met2 ;
        RECT 3377.035 4319.855 3379.435 4320.135 ;
      LAYER met2 ;
        RECT 3379.715 4319.575 3588.000 4320.415 ;
        RECT 3379.435 4317.195 3588.000 4319.575 ;
        RECT 3379.715 4316.355 3588.000 4317.195 ;
        RECT 3379.435 4313.975 3588.000 4316.355 ;
      LAYER met2 ;
        RECT 3377.035 4313.650 3379.435 4313.695 ;
        RECT 3376.560 4313.510 3379.435 4313.650 ;
        RECT 3377.035 4313.415 3379.435 4313.510 ;
      LAYER met2 ;
        RECT 3379.715 4313.135 3588.000 4313.975 ;
        RECT 3379.435 4312.085 3588.000 4313.135 ;
        RECT 3390.035 4166.505 3583.075 4166.735 ;
        RECT 3388.000 4142.605 3583.075 4166.505 ;
        RECT 3388.000 4139.105 3389.920 4141.105 ;
        RECT 3390.035 4116.610 3583.075 4142.605 ;
        RECT 3388.000 4092.710 3583.075 4116.610 ;
      LAYER met2 ;
        RECT 3376.500 4091.570 3376.760 4091.890 ;
        RECT 3387.530 4091.715 3387.810 4092.085 ;
        RECT 3387.540 4091.570 3387.800 4091.715 ;
        RECT 3375.120 3916.130 3375.380 3916.450 ;
        RECT 3374.660 3874.990 3374.920 3875.310 ;
        RECT 3374.200 3701.590 3374.460 3701.910 ;
        RECT 3374.200 3679.830 3374.460 3680.150 ;
        RECT 3374.260 3645.470 3374.400 3679.830 ;
        RECT 3374.720 3649.890 3374.860 3874.990 ;
        RECT 3375.180 3686.610 3375.320 3916.130 ;
        RECT 3376.040 3904.910 3376.300 3905.230 ;
        RECT 3376.100 3870.210 3376.240 3904.910 ;
        RECT 3376.040 3869.890 3376.300 3870.210 ;
        RECT 3376.040 3701.590 3376.300 3701.910 ;
        RECT 3375.120 3686.290 3375.380 3686.610 ;
        RECT 3374.660 3649.570 3374.920 3649.890 ;
        RECT 3374.200 3645.150 3374.460 3645.470 ;
        RECT 3374.720 3632.550 3374.860 3649.570 ;
        RECT 3374.660 3632.230 3374.920 3632.550 ;
        RECT 3374.660 3494.870 3374.920 3495.190 ;
        RECT 3374.720 3481.250 3374.860 3494.870 ;
        RECT 3374.660 3480.930 3374.920 3481.250 ;
        RECT 3375.180 3480.650 3375.320 3686.290 ;
        RECT 3376.100 3632.970 3376.240 3701.590 ;
        RECT 3376.560 3633.570 3376.700 4091.570 ;
      LAYER met2 ;
        RECT 3379.435 3944.795 3588.000 3945.790 ;
      LAYER met2 ;
        RECT 3377.035 3944.235 3379.435 3944.515 ;
      LAYER met2 ;
        RECT 3379.715 3943.955 3588.000 3944.795 ;
        RECT 3379.435 3942.035 3588.000 3943.955 ;
        RECT 3379.715 3941.195 3588.000 3942.035 ;
        RECT 3379.435 3938.815 3588.000 3941.195 ;
        RECT 3379.715 3937.975 3588.000 3938.815 ;
        RECT 3379.435 3935.595 3588.000 3937.975 ;
        RECT 3379.715 3934.755 3588.000 3935.595 ;
        RECT 3379.435 3932.835 3588.000 3934.755 ;
        RECT 3379.715 3931.995 3588.000 3932.835 ;
        RECT 3379.435 3929.615 3588.000 3931.995 ;
      LAYER met2 ;
        RECT 3377.035 3929.195 3379.435 3929.335 ;
        RECT 3377.020 3929.055 3379.435 3929.195 ;
        RECT 3377.020 3926.650 3377.160 3929.055 ;
      LAYER met2 ;
        RECT 3379.715 3928.775 3588.000 3929.615 ;
      LAYER met2 ;
        RECT 3376.960 3926.330 3377.220 3926.650 ;
      LAYER met2 ;
        RECT 3379.435 3926.395 3588.000 3928.775 ;
        RECT 3379.715 3925.555 3588.000 3926.395 ;
        RECT 3379.435 3923.635 3588.000 3925.555 ;
        RECT 3379.715 3922.795 3588.000 3923.635 ;
        RECT 3379.435 3920.415 3588.000 3922.795 ;
        RECT 3379.715 3919.575 3588.000 3920.415 ;
        RECT 3379.435 3917.195 3588.000 3919.575 ;
      LAYER met2 ;
        RECT 3376.960 3916.130 3377.220 3916.450 ;
      LAYER met2 ;
        RECT 3379.715 3916.355 3588.000 3917.195 ;
      LAYER met2 ;
        RECT 3377.020 3914.155 3377.160 3916.130 ;
      LAYER met2 ;
        RECT 3379.435 3914.435 3588.000 3916.355 ;
      LAYER met2 ;
        RECT 3377.020 3914.015 3379.435 3914.155 ;
        RECT 3377.035 3913.875 3379.435 3914.015 ;
      LAYER met2 ;
        RECT 3379.715 3913.595 3588.000 3914.435 ;
        RECT 3379.435 3911.215 3588.000 3913.595 ;
        RECT 3379.715 3910.375 3588.000 3911.215 ;
        RECT 3379.435 3907.995 3588.000 3910.375 ;
      LAYER met2 ;
        RECT 3377.035 3907.620 3379.435 3907.715 ;
        RECT 3377.020 3907.435 3379.435 3907.620 ;
        RECT 3377.020 3905.230 3377.160 3907.435 ;
      LAYER met2 ;
        RECT 3379.715 3907.155 3588.000 3907.995 ;
      LAYER met2 ;
        RECT 3376.960 3904.910 3377.220 3905.230 ;
      LAYER met2 ;
        RECT 3379.435 3904.775 3588.000 3907.155 ;
        RECT 3379.715 3903.935 3588.000 3904.775 ;
        RECT 3379.435 3902.015 3588.000 3903.935 ;
        RECT 3379.715 3901.175 3588.000 3902.015 ;
        RECT 3379.435 3898.795 3588.000 3901.175 ;
        RECT 3379.715 3897.955 3588.000 3898.795 ;
        RECT 3379.435 3895.575 3588.000 3897.955 ;
        RECT 3379.715 3894.735 3588.000 3895.575 ;
        RECT 3379.435 3892.815 3588.000 3894.735 ;
      LAYER met2 ;
        RECT 3377.035 3892.255 3379.435 3892.535 ;
      LAYER met2 ;
        RECT 3379.715 3891.975 3588.000 3892.815 ;
        RECT 3379.435 3889.595 3588.000 3891.975 ;
        RECT 3379.715 3888.755 3588.000 3889.595 ;
        RECT 3379.435 3886.375 3588.000 3888.755 ;
      LAYER met2 ;
        RECT 3377.035 3885.815 3379.435 3886.095 ;
      LAYER met2 ;
        RECT 3379.715 3885.535 3588.000 3886.375 ;
        RECT 3379.435 3883.615 3588.000 3885.535 ;
        RECT 3379.715 3882.775 3588.000 3883.615 ;
        RECT 3379.435 3880.395 3588.000 3882.775 ;
        RECT 3379.715 3879.555 3588.000 3880.395 ;
        RECT 3379.435 3877.175 3588.000 3879.555 ;
      LAYER met2 ;
        RECT 3377.035 3876.755 3379.435 3876.895 ;
        RECT 3377.020 3876.615 3379.435 3876.755 ;
        RECT 3377.020 3875.310 3377.160 3876.615 ;
      LAYER met2 ;
        RECT 3379.715 3876.335 3588.000 3877.175 ;
      LAYER met2 ;
        RECT 3376.960 3874.990 3377.220 3875.310 ;
      LAYER met2 ;
        RECT 3379.435 3874.415 3588.000 3876.335 ;
      LAYER met2 ;
        RECT 3377.035 3873.855 3379.435 3874.135 ;
      LAYER met2 ;
        RECT 3379.715 3873.575 3588.000 3874.415 ;
        RECT 3379.435 3871.195 3588.000 3873.575 ;
        RECT 3379.715 3870.355 3588.000 3871.195 ;
      LAYER met2 ;
        RECT 3376.960 3869.890 3377.220 3870.210 ;
        RECT 3377.020 3867.695 3377.160 3869.890 ;
      LAYER met2 ;
        RECT 3379.435 3867.975 3588.000 3870.355 ;
      LAYER met2 ;
        RECT 3377.020 3867.500 3379.435 3867.695 ;
        RECT 3377.035 3867.415 3379.435 3867.500 ;
      LAYER met2 ;
        RECT 3379.715 3867.135 3588.000 3867.975 ;
        RECT 3379.435 3866.085 3588.000 3867.135 ;
        RECT 3379.435 3719.795 3588.000 3720.790 ;
      LAYER met2 ;
        RECT 3377.035 3719.235 3379.435 3719.515 ;
      LAYER met2 ;
        RECT 3379.715 3718.955 3588.000 3719.795 ;
        RECT 3379.435 3717.035 3588.000 3718.955 ;
        RECT 3379.715 3716.195 3588.000 3717.035 ;
        RECT 3379.435 3713.815 3588.000 3716.195 ;
        RECT 3379.715 3712.975 3588.000 3713.815 ;
        RECT 3379.435 3710.595 3588.000 3712.975 ;
        RECT 3379.715 3709.755 3588.000 3710.595 ;
        RECT 3379.435 3707.835 3588.000 3709.755 ;
        RECT 3379.715 3706.995 3588.000 3707.835 ;
        RECT 3379.435 3704.615 3588.000 3706.995 ;
      LAYER met2 ;
        RECT 3377.035 3704.300 3379.435 3704.335 ;
        RECT 3377.020 3704.055 3379.435 3704.300 ;
        RECT 3377.020 3701.910 3377.160 3704.055 ;
      LAYER met2 ;
        RECT 3379.715 3703.775 3588.000 3704.615 ;
      LAYER met2 ;
        RECT 3376.960 3701.590 3377.220 3701.910 ;
      LAYER met2 ;
        RECT 3379.435 3701.395 3588.000 3703.775 ;
        RECT 3379.715 3700.555 3588.000 3701.395 ;
        RECT 3379.435 3698.635 3588.000 3700.555 ;
        RECT 3379.715 3697.795 3588.000 3698.635 ;
        RECT 3379.435 3695.415 3588.000 3697.795 ;
        RECT 3379.715 3694.575 3588.000 3695.415 ;
        RECT 3379.435 3692.195 3588.000 3694.575 ;
        RECT 3379.715 3691.355 3588.000 3692.195 ;
        RECT 3379.435 3689.435 3588.000 3691.355 ;
      LAYER met2 ;
        RECT 3377.035 3689.015 3379.435 3689.155 ;
        RECT 3377.020 3688.875 3379.435 3689.015 ;
        RECT 3377.020 3686.610 3377.160 3688.875 ;
      LAYER met2 ;
        RECT 3379.715 3688.595 3588.000 3689.435 ;
      LAYER met2 ;
        RECT 3376.960 3686.290 3377.220 3686.610 ;
      LAYER met2 ;
        RECT 3379.435 3686.215 3588.000 3688.595 ;
        RECT 3379.715 3685.375 3588.000 3686.215 ;
        RECT 3379.435 3682.995 3588.000 3685.375 ;
      LAYER met2 ;
        RECT 3377.035 3682.540 3379.435 3682.715 ;
        RECT 3377.020 3682.435 3379.435 3682.540 ;
        RECT 3377.020 3680.150 3377.160 3682.435 ;
      LAYER met2 ;
        RECT 3379.715 3682.155 3588.000 3682.995 ;
      LAYER met2 ;
        RECT 3376.960 3679.830 3377.220 3680.150 ;
      LAYER met2 ;
        RECT 3379.435 3679.775 3588.000 3682.155 ;
        RECT 3379.715 3678.935 3588.000 3679.775 ;
        RECT 3379.435 3677.015 3588.000 3678.935 ;
        RECT 3379.715 3676.175 3588.000 3677.015 ;
        RECT 3379.435 3673.795 3588.000 3676.175 ;
        RECT 3379.715 3672.955 3588.000 3673.795 ;
        RECT 3379.435 3670.575 3588.000 3672.955 ;
        RECT 3379.715 3669.735 3588.000 3670.575 ;
        RECT 3379.435 3667.815 3588.000 3669.735 ;
      LAYER met2 ;
        RECT 3377.035 3667.255 3379.435 3667.535 ;
      LAYER met2 ;
        RECT 3379.715 3666.975 3588.000 3667.815 ;
        RECT 3379.435 3664.595 3588.000 3666.975 ;
        RECT 3379.715 3663.755 3588.000 3664.595 ;
        RECT 3379.435 3661.375 3588.000 3663.755 ;
      LAYER met2 ;
        RECT 3377.035 3660.815 3379.435 3661.095 ;
      LAYER met2 ;
        RECT 3379.715 3660.535 3588.000 3661.375 ;
        RECT 3379.435 3658.615 3588.000 3660.535 ;
        RECT 3379.715 3657.775 3588.000 3658.615 ;
        RECT 3379.435 3655.395 3588.000 3657.775 ;
        RECT 3379.715 3654.555 3588.000 3655.395 ;
        RECT 3379.435 3652.175 3588.000 3654.555 ;
      LAYER met2 ;
        RECT 3377.035 3651.755 3379.435 3651.895 ;
        RECT 3377.020 3651.615 3379.435 3651.755 ;
        RECT 3377.020 3649.890 3377.160 3651.615 ;
      LAYER met2 ;
        RECT 3379.715 3651.335 3588.000 3652.175 ;
      LAYER met2 ;
        RECT 3376.960 3649.570 3377.220 3649.890 ;
      LAYER met2 ;
        RECT 3379.435 3649.415 3588.000 3651.335 ;
      LAYER met2 ;
        RECT 3377.035 3648.855 3379.435 3649.135 ;
      LAYER met2 ;
        RECT 3379.715 3648.575 3588.000 3649.415 ;
        RECT 3379.435 3646.195 3588.000 3648.575 ;
      LAYER met2 ;
        RECT 3376.960 3645.150 3377.220 3645.470 ;
      LAYER met2 ;
        RECT 3379.715 3645.355 3588.000 3646.195 ;
      LAYER met2 ;
        RECT 3377.020 3642.695 3377.160 3645.150 ;
      LAYER met2 ;
        RECT 3379.435 3642.975 3588.000 3645.355 ;
      LAYER met2 ;
        RECT 3377.020 3642.420 3379.435 3642.695 ;
        RECT 3377.035 3642.415 3379.435 3642.420 ;
      LAYER met2 ;
        RECT 3379.715 3642.135 3588.000 3642.975 ;
        RECT 3379.435 3641.085 3588.000 3642.135 ;
      LAYER met2 ;
        RECT 3376.500 3633.250 3376.760 3633.570 ;
        RECT 3376.100 3632.830 3377.160 3632.970 ;
        RECT 3376.040 3632.230 3376.300 3632.550 ;
        RECT 3376.500 3632.230 3376.760 3632.550 ;
        RECT 3374.260 3480.510 3375.320 3480.650 ;
        RECT 3374.260 3466.290 3374.400 3480.510 ;
        RECT 3374.660 3479.910 3374.920 3480.230 ;
        RECT 3374.720 3476.830 3374.860 3479.910 ;
        RECT 3374.660 3476.510 3374.920 3476.830 ;
        RECT 3374.200 3465.970 3374.460 3466.290 ;
        RECT 3374.260 3240.190 3374.400 3465.970 ;
        RECT 3374.720 3250.730 3374.860 3476.510 ;
        RECT 3376.100 3467.050 3376.240 3632.230 ;
        RECT 3375.640 3466.910 3376.240 3467.050 ;
        RECT 3375.640 3426.170 3375.780 3466.910 ;
        RECT 3376.040 3458.150 3376.300 3458.470 ;
        RECT 3375.580 3425.850 3375.840 3426.170 ;
        RECT 3375.640 3419.450 3375.780 3425.850 ;
        RECT 3376.100 3420.390 3376.240 3458.150 ;
        RECT 3376.560 3458.130 3376.700 3632.230 ;
        RECT 3377.020 3495.190 3377.160 3632.830 ;
        RECT 3376.960 3494.870 3377.220 3495.190 ;
      LAYER met2 ;
        RECT 3379.435 3494.795 3588.000 3495.790 ;
      LAYER met2 ;
        RECT 3377.035 3494.235 3379.435 3494.515 ;
      LAYER met2 ;
        RECT 3379.715 3493.955 3588.000 3494.795 ;
        RECT 3379.435 3492.035 3588.000 3493.955 ;
        RECT 3379.715 3491.195 3588.000 3492.035 ;
        RECT 3379.435 3488.815 3588.000 3491.195 ;
        RECT 3379.715 3487.975 3588.000 3488.815 ;
        RECT 3379.435 3485.595 3588.000 3487.975 ;
        RECT 3379.715 3484.755 3588.000 3485.595 ;
        RECT 3379.435 3482.835 3588.000 3484.755 ;
        RECT 3379.715 3481.995 3588.000 3482.835 ;
        RECT 3379.435 3479.615 3588.000 3481.995 ;
      LAYER met2 ;
        RECT 3377.035 3479.220 3379.435 3479.335 ;
        RECT 3377.020 3479.055 3379.435 3479.220 ;
        RECT 3377.020 3476.830 3377.160 3479.055 ;
      LAYER met2 ;
        RECT 3379.715 3478.775 3588.000 3479.615 ;
      LAYER met2 ;
        RECT 3376.960 3476.510 3377.220 3476.830 ;
      LAYER met2 ;
        RECT 3379.435 3476.395 3588.000 3478.775 ;
        RECT 3379.715 3475.555 3588.000 3476.395 ;
        RECT 3379.435 3473.635 3588.000 3475.555 ;
        RECT 3379.715 3472.795 3588.000 3473.635 ;
        RECT 3379.435 3470.415 3588.000 3472.795 ;
        RECT 3379.715 3469.575 3588.000 3470.415 ;
        RECT 3379.435 3467.195 3588.000 3469.575 ;
        RECT 3379.715 3466.355 3588.000 3467.195 ;
      LAYER met2 ;
        RECT 3376.960 3465.970 3377.220 3466.290 ;
        RECT 3377.020 3464.155 3377.160 3465.970 ;
      LAYER met2 ;
        RECT 3379.435 3464.435 3588.000 3466.355 ;
      LAYER met2 ;
        RECT 3377.020 3464.015 3379.435 3464.155 ;
        RECT 3377.035 3463.875 3379.435 3464.015 ;
      LAYER met2 ;
        RECT 3379.715 3463.595 3588.000 3464.435 ;
        RECT 3379.435 3461.215 3588.000 3463.595 ;
        RECT 3379.715 3460.375 3588.000 3461.215 ;
      LAYER met2 ;
        RECT 3376.960 3458.150 3377.220 3458.470 ;
        RECT 3376.500 3457.810 3376.760 3458.130 ;
        RECT 3377.020 3457.715 3377.160 3458.150 ;
      LAYER met2 ;
        RECT 3379.435 3457.995 3588.000 3460.375 ;
      LAYER met2 ;
        RECT 3377.020 3457.460 3379.435 3457.715 ;
        RECT 3377.035 3457.435 3379.435 3457.460 ;
      LAYER met2 ;
        RECT 3379.715 3457.155 3588.000 3457.995 ;
      LAYER met2 ;
        RECT 3376.500 3456.790 3376.760 3457.110 ;
        RECT 3376.040 3420.070 3376.300 3420.390 ;
        RECT 3375.640 3419.310 3376.240 3419.450 ;
        RECT 3376.100 3357.150 3376.240 3419.310 ;
        RECT 3375.120 3356.830 3375.380 3357.150 ;
        RECT 3376.040 3356.830 3376.300 3357.150 ;
        RECT 3374.660 3250.410 3374.920 3250.730 ;
        RECT 3374.200 3239.870 3374.460 3240.190 ;
        RECT 3374.260 3012.050 3374.400 3239.870 ;
        RECT 3374.720 3027.690 3374.860 3250.410 ;
        RECT 3375.180 3199.050 3375.320 3356.830 ;
        RECT 3376.040 3228.650 3376.300 3228.970 ;
        RECT 3375.120 3198.730 3375.380 3199.050 ;
        RECT 3374.660 3027.370 3374.920 3027.690 ;
        RECT 3374.200 3011.730 3374.460 3012.050 ;
        RECT 3374.720 3011.450 3374.860 3027.370 ;
        RECT 3373.800 3011.310 3374.860 3011.450 ;
        RECT 3373.800 3010.090 3373.940 3011.310 ;
        RECT 3374.660 3010.370 3374.920 3010.690 ;
        RECT 3373.800 3009.950 3374.400 3010.090 ;
        RECT 3374.260 2804.990 3374.400 3009.950 ;
        RECT 3374.200 2804.670 3374.460 2804.990 ;
        RECT 3370.520 2138.950 3370.780 2139.270 ;
        RECT 213.540 2001.930 213.800 2002.250 ;
        RECT 3374.260 1918.950 3374.400 2804.670 ;
        RECT 3374.720 2789.350 3374.860 3010.370 ;
        RECT 3375.180 2973.630 3375.320 3198.730 ;
        RECT 3376.100 3194.290 3376.240 3228.650 ;
        RECT 3376.040 3193.970 3376.300 3194.290 ;
        RECT 3376.040 3003.910 3376.300 3004.230 ;
        RECT 3375.120 2973.310 3375.380 2973.630 ;
        RECT 3374.660 2789.030 3374.920 2789.350 ;
        RECT 3375.180 2752.630 3375.320 2973.310 ;
        RECT 3376.100 2969.210 3376.240 3003.910 ;
        RECT 3376.040 2968.890 3376.300 2969.210 ;
        RECT 3376.560 2787.670 3376.700 3456.790 ;
      LAYER met2 ;
        RECT 3379.435 3454.775 3588.000 3457.155 ;
        RECT 3379.715 3453.935 3588.000 3454.775 ;
        RECT 3379.435 3452.015 3588.000 3453.935 ;
        RECT 3379.715 3451.175 3588.000 3452.015 ;
        RECT 3379.435 3448.795 3588.000 3451.175 ;
        RECT 3379.715 3447.955 3588.000 3448.795 ;
        RECT 3379.435 3445.575 3588.000 3447.955 ;
        RECT 3379.715 3444.735 3588.000 3445.575 ;
        RECT 3379.435 3442.815 3588.000 3444.735 ;
      LAYER met2 ;
        RECT 3377.035 3442.255 3379.435 3442.535 ;
      LAYER met2 ;
        RECT 3379.715 3441.975 3588.000 3442.815 ;
        RECT 3379.435 3439.595 3588.000 3441.975 ;
        RECT 3379.715 3438.755 3588.000 3439.595 ;
        RECT 3379.435 3436.375 3588.000 3438.755 ;
      LAYER met2 ;
        RECT 3377.035 3435.815 3379.435 3436.095 ;
      LAYER met2 ;
        RECT 3379.715 3435.535 3588.000 3436.375 ;
        RECT 3379.435 3433.615 3588.000 3435.535 ;
        RECT 3379.715 3432.775 3588.000 3433.615 ;
        RECT 3379.435 3430.395 3588.000 3432.775 ;
        RECT 3379.715 3429.555 3588.000 3430.395 ;
        RECT 3379.435 3427.175 3588.000 3429.555 ;
      LAYER met2 ;
        RECT 3377.035 3426.860 3379.435 3426.895 ;
        RECT 3377.020 3426.615 3379.435 3426.860 ;
        RECT 3377.020 3426.170 3377.160 3426.615 ;
      LAYER met2 ;
        RECT 3379.715 3426.335 3588.000 3427.175 ;
      LAYER met2 ;
        RECT 3376.960 3425.850 3377.220 3426.170 ;
      LAYER met2 ;
        RECT 3379.435 3424.415 3588.000 3426.335 ;
      LAYER met2 ;
        RECT 3377.035 3423.855 3379.435 3424.135 ;
      LAYER met2 ;
        RECT 3379.715 3423.575 3588.000 3424.415 ;
        RECT 3379.435 3421.195 3588.000 3423.575 ;
      LAYER met2 ;
        RECT 3376.960 3420.070 3377.220 3420.390 ;
      LAYER met2 ;
        RECT 3379.715 3420.355 3588.000 3421.195 ;
      LAYER met2 ;
        RECT 3377.020 3417.695 3377.160 3420.070 ;
      LAYER met2 ;
        RECT 3379.435 3417.975 3588.000 3420.355 ;
      LAYER met2 ;
        RECT 3377.020 3417.555 3379.435 3417.695 ;
        RECT 3377.035 3417.415 3379.435 3417.555 ;
      LAYER met2 ;
        RECT 3379.715 3417.135 3588.000 3417.975 ;
        RECT 3379.435 3416.085 3588.000 3417.135 ;
        RECT 3379.435 3268.795 3588.000 3269.790 ;
      LAYER met2 ;
        RECT 3377.035 3268.235 3379.435 3268.515 ;
      LAYER met2 ;
        RECT 3379.715 3267.955 3588.000 3268.795 ;
        RECT 3379.435 3266.035 3588.000 3267.955 ;
        RECT 3379.715 3265.195 3588.000 3266.035 ;
        RECT 3379.435 3262.815 3588.000 3265.195 ;
        RECT 3379.715 3261.975 3588.000 3262.815 ;
        RECT 3379.435 3259.595 3588.000 3261.975 ;
        RECT 3379.715 3258.755 3588.000 3259.595 ;
        RECT 3379.435 3256.835 3588.000 3258.755 ;
        RECT 3379.715 3255.995 3588.000 3256.835 ;
        RECT 3379.435 3253.615 3588.000 3255.995 ;
      LAYER met2 ;
        RECT 3377.035 3253.195 3379.435 3253.335 ;
        RECT 3377.020 3253.055 3379.435 3253.195 ;
        RECT 3377.020 3250.730 3377.160 3253.055 ;
      LAYER met2 ;
        RECT 3379.715 3252.775 3588.000 3253.615 ;
      LAYER met2 ;
        RECT 3376.960 3250.410 3377.220 3250.730 ;
      LAYER met2 ;
        RECT 3379.435 3250.395 3588.000 3252.775 ;
        RECT 3379.715 3249.555 3588.000 3250.395 ;
        RECT 3379.435 3247.635 3588.000 3249.555 ;
        RECT 3379.715 3246.795 3588.000 3247.635 ;
        RECT 3379.435 3244.415 3588.000 3246.795 ;
        RECT 3379.715 3243.575 3588.000 3244.415 ;
        RECT 3379.435 3241.195 3588.000 3243.575 ;
        RECT 3379.715 3240.355 3588.000 3241.195 ;
      LAYER met2 ;
        RECT 3376.960 3239.870 3377.220 3240.190 ;
        RECT 3377.020 3238.155 3377.160 3239.870 ;
      LAYER met2 ;
        RECT 3379.435 3238.435 3588.000 3240.355 ;
      LAYER met2 ;
        RECT 3377.020 3238.015 3379.435 3238.155 ;
        RECT 3377.035 3237.875 3379.435 3238.015 ;
      LAYER met2 ;
        RECT 3379.715 3237.595 3588.000 3238.435 ;
        RECT 3379.435 3235.215 3588.000 3237.595 ;
        RECT 3379.715 3234.375 3588.000 3235.215 ;
        RECT 3379.435 3231.995 3588.000 3234.375 ;
      LAYER met2 ;
        RECT 3377.035 3231.700 3379.435 3231.715 ;
        RECT 3377.020 3231.435 3379.435 3231.700 ;
        RECT 3377.020 3228.970 3377.160 3231.435 ;
      LAYER met2 ;
        RECT 3379.715 3231.155 3588.000 3231.995 ;
      LAYER met2 ;
        RECT 3376.960 3228.650 3377.220 3228.970 ;
      LAYER met2 ;
        RECT 3379.435 3228.775 3588.000 3231.155 ;
        RECT 3379.715 3227.935 3588.000 3228.775 ;
        RECT 3379.435 3226.015 3588.000 3227.935 ;
        RECT 3379.715 3225.175 3588.000 3226.015 ;
        RECT 3379.435 3222.795 3588.000 3225.175 ;
        RECT 3379.715 3221.955 3588.000 3222.795 ;
        RECT 3379.435 3219.575 3588.000 3221.955 ;
        RECT 3379.715 3218.735 3588.000 3219.575 ;
        RECT 3379.435 3216.815 3588.000 3218.735 ;
      LAYER met2 ;
        RECT 3377.035 3216.255 3379.435 3216.535 ;
      LAYER met2 ;
        RECT 3379.715 3215.975 3588.000 3216.815 ;
        RECT 3379.435 3213.595 3588.000 3215.975 ;
        RECT 3379.715 3212.755 3588.000 3213.595 ;
        RECT 3379.435 3210.375 3588.000 3212.755 ;
      LAYER met2 ;
        RECT 3377.035 3209.815 3379.435 3210.095 ;
      LAYER met2 ;
        RECT 3379.715 3209.535 3588.000 3210.375 ;
        RECT 3379.435 3207.615 3588.000 3209.535 ;
        RECT 3379.715 3206.775 3588.000 3207.615 ;
        RECT 3379.435 3204.395 3588.000 3206.775 ;
        RECT 3379.715 3203.555 3588.000 3204.395 ;
        RECT 3379.435 3201.175 3588.000 3203.555 ;
      LAYER met2 ;
        RECT 3377.035 3200.755 3379.435 3200.895 ;
        RECT 3377.020 3200.615 3379.435 3200.755 ;
        RECT 3377.020 3199.050 3377.160 3200.615 ;
      LAYER met2 ;
        RECT 3379.715 3200.335 3588.000 3201.175 ;
      LAYER met2 ;
        RECT 3376.960 3198.730 3377.220 3199.050 ;
      LAYER met2 ;
        RECT 3379.435 3198.415 3588.000 3200.335 ;
      LAYER met2 ;
        RECT 3377.035 3197.855 3379.435 3198.135 ;
      LAYER met2 ;
        RECT 3379.715 3197.575 3588.000 3198.415 ;
        RECT 3379.435 3195.195 3588.000 3197.575 ;
        RECT 3379.715 3194.355 3588.000 3195.195 ;
      LAYER met2 ;
        RECT 3376.960 3193.970 3377.220 3194.290 ;
        RECT 3377.020 3191.695 3377.160 3193.970 ;
      LAYER met2 ;
        RECT 3379.435 3191.975 3588.000 3194.355 ;
      LAYER met2 ;
        RECT 3377.020 3191.580 3379.435 3191.695 ;
        RECT 3377.035 3191.415 3379.435 3191.580 ;
      LAYER met2 ;
        RECT 3379.715 3191.135 3588.000 3191.975 ;
        RECT 3379.435 3190.085 3588.000 3191.135 ;
        RECT 3379.435 3043.795 3588.000 3044.790 ;
      LAYER met2 ;
        RECT 3377.035 3043.235 3379.435 3043.515 ;
      LAYER met2 ;
        RECT 3379.715 3042.955 3588.000 3043.795 ;
        RECT 3379.435 3041.035 3588.000 3042.955 ;
        RECT 3379.715 3040.195 3588.000 3041.035 ;
        RECT 3379.435 3037.815 3588.000 3040.195 ;
        RECT 3379.715 3036.975 3588.000 3037.815 ;
        RECT 3379.435 3034.595 3588.000 3036.975 ;
        RECT 3379.715 3033.755 3588.000 3034.595 ;
        RECT 3379.435 3031.835 3588.000 3033.755 ;
        RECT 3379.715 3030.995 3588.000 3031.835 ;
        RECT 3379.435 3028.615 3588.000 3030.995 ;
      LAYER met2 ;
        RECT 3377.035 3028.195 3379.435 3028.335 ;
        RECT 3377.020 3028.055 3379.435 3028.195 ;
        RECT 3377.020 3027.690 3377.160 3028.055 ;
      LAYER met2 ;
        RECT 3379.715 3027.775 3588.000 3028.615 ;
      LAYER met2 ;
        RECT 3376.960 3027.370 3377.220 3027.690 ;
      LAYER met2 ;
        RECT 3379.435 3025.395 3588.000 3027.775 ;
        RECT 3379.715 3024.555 3588.000 3025.395 ;
        RECT 3379.435 3022.635 3588.000 3024.555 ;
        RECT 3379.715 3021.795 3588.000 3022.635 ;
        RECT 3379.435 3019.415 3588.000 3021.795 ;
        RECT 3379.715 3018.575 3588.000 3019.415 ;
        RECT 3379.435 3016.195 3588.000 3018.575 ;
        RECT 3379.715 3015.355 3588.000 3016.195 ;
        RECT 3379.435 3013.435 3588.000 3015.355 ;
      LAYER met2 ;
        RECT 3377.035 3013.015 3379.435 3013.155 ;
        RECT 3377.020 3012.875 3379.435 3013.015 ;
        RECT 3377.020 3010.690 3377.160 3012.875 ;
      LAYER met2 ;
        RECT 3379.715 3012.595 3588.000 3013.435 ;
      LAYER met2 ;
        RECT 3376.960 3010.370 3377.220 3010.690 ;
      LAYER met2 ;
        RECT 3379.435 3010.215 3588.000 3012.595 ;
        RECT 3379.715 3009.375 3588.000 3010.215 ;
        RECT 3379.435 3006.995 3588.000 3009.375 ;
      LAYER met2 ;
        RECT 3377.035 3006.620 3379.435 3006.715 ;
        RECT 3377.020 3006.435 3379.435 3006.620 ;
        RECT 3377.020 3004.230 3377.160 3006.435 ;
      LAYER met2 ;
        RECT 3379.715 3006.155 3588.000 3006.995 ;
      LAYER met2 ;
        RECT 3376.960 3003.910 3377.220 3004.230 ;
      LAYER met2 ;
        RECT 3379.435 3003.775 3588.000 3006.155 ;
        RECT 3379.715 3002.935 3588.000 3003.775 ;
        RECT 3379.435 3001.015 3588.000 3002.935 ;
        RECT 3379.715 3000.175 3588.000 3001.015 ;
        RECT 3379.435 2997.795 3588.000 3000.175 ;
        RECT 3379.715 2996.955 3588.000 2997.795 ;
        RECT 3379.435 2994.575 3588.000 2996.955 ;
        RECT 3379.715 2993.735 3588.000 2994.575 ;
        RECT 3379.435 2991.815 3588.000 2993.735 ;
      LAYER met2 ;
        RECT 3377.035 2991.255 3379.435 2991.535 ;
      LAYER met2 ;
        RECT 3379.715 2990.975 3588.000 2991.815 ;
        RECT 3379.435 2988.595 3588.000 2990.975 ;
        RECT 3379.715 2987.755 3588.000 2988.595 ;
        RECT 3379.435 2985.375 3588.000 2987.755 ;
      LAYER met2 ;
        RECT 3377.035 2984.815 3379.435 2985.095 ;
      LAYER met2 ;
        RECT 3379.715 2984.535 3588.000 2985.375 ;
        RECT 3379.435 2982.615 3588.000 2984.535 ;
        RECT 3379.715 2981.775 3588.000 2982.615 ;
        RECT 3379.435 2979.395 3588.000 2981.775 ;
        RECT 3379.715 2978.555 3588.000 2979.395 ;
        RECT 3379.435 2976.175 3588.000 2978.555 ;
      LAYER met2 ;
        RECT 3377.035 2975.755 3379.435 2975.895 ;
        RECT 3377.020 2975.615 3379.435 2975.755 ;
        RECT 3377.020 2973.630 3377.160 2975.615 ;
      LAYER met2 ;
        RECT 3379.715 2975.335 3588.000 2976.175 ;
      LAYER met2 ;
        RECT 3376.960 2973.310 3377.220 2973.630 ;
      LAYER met2 ;
        RECT 3379.435 2973.415 3588.000 2975.335 ;
      LAYER met2 ;
        RECT 3377.035 2972.855 3379.435 2973.135 ;
      LAYER met2 ;
        RECT 3379.715 2972.575 3588.000 2973.415 ;
        RECT 3379.435 2970.195 3588.000 2972.575 ;
        RECT 3379.715 2969.355 3588.000 2970.195 ;
      LAYER met2 ;
        RECT 3376.960 2968.890 3377.220 2969.210 ;
        RECT 3377.020 2966.695 3377.160 2968.890 ;
      LAYER met2 ;
        RECT 3379.435 2966.975 3588.000 2969.355 ;
      LAYER met2 ;
        RECT 3377.020 2966.500 3379.435 2966.695 ;
        RECT 3377.035 2966.415 3379.435 2966.500 ;
      LAYER met2 ;
        RECT 3379.715 2966.135 3588.000 2966.975 ;
        RECT 3379.435 2965.085 3588.000 2966.135 ;
        RECT 3379.435 2817.795 3588.000 2818.790 ;
      LAYER met2 ;
        RECT 3377.035 2817.235 3379.435 2817.515 ;
      LAYER met2 ;
        RECT 3379.715 2816.955 3588.000 2817.795 ;
        RECT 3379.435 2815.035 3588.000 2816.955 ;
        RECT 3379.715 2814.195 3588.000 2815.035 ;
        RECT 3379.435 2811.815 3588.000 2814.195 ;
        RECT 3379.715 2810.975 3588.000 2811.815 ;
        RECT 3379.435 2808.595 3588.000 2810.975 ;
        RECT 3379.715 2807.755 3588.000 2808.595 ;
        RECT 3379.435 2805.835 3588.000 2807.755 ;
        RECT 3379.715 2804.995 3588.000 2805.835 ;
      LAYER met2 ;
        RECT 3376.960 2804.670 3377.220 2804.990 ;
        RECT 3377.020 2802.335 3377.160 2804.670 ;
      LAYER met2 ;
        RECT 3379.435 2802.615 3588.000 2804.995 ;
      LAYER met2 ;
        RECT 3377.020 2802.195 3379.435 2802.335 ;
        RECT 3377.035 2802.055 3379.435 2802.195 ;
      LAYER met2 ;
        RECT 3379.715 2801.775 3588.000 2802.615 ;
        RECT 3379.435 2799.395 3588.000 2801.775 ;
        RECT 3379.715 2798.555 3588.000 2799.395 ;
        RECT 3379.435 2796.635 3588.000 2798.555 ;
        RECT 3379.715 2795.795 3588.000 2796.635 ;
        RECT 3379.435 2793.415 3588.000 2795.795 ;
        RECT 3379.715 2792.575 3588.000 2793.415 ;
        RECT 3379.435 2790.195 3588.000 2792.575 ;
        RECT 3379.715 2789.355 3588.000 2790.195 ;
      LAYER met2 ;
        RECT 3376.960 2789.030 3377.220 2789.350 ;
        RECT 3376.100 2787.530 3376.700 2787.670 ;
        RECT 3376.100 2778.890 3376.240 2787.530 ;
        RECT 3377.020 2787.155 3377.160 2789.030 ;
      LAYER met2 ;
        RECT 3379.435 2787.435 3588.000 2789.355 ;
      LAYER met2 ;
        RECT 3377.020 2786.980 3379.435 2787.155 ;
        RECT 3377.035 2786.875 3379.435 2786.980 ;
      LAYER met2 ;
        RECT 3379.715 2786.595 3588.000 2787.435 ;
        RECT 3379.435 2784.215 3588.000 2786.595 ;
        RECT 3379.715 2783.375 3588.000 2784.215 ;
        RECT 3379.435 2780.995 3588.000 2783.375 ;
      LAYER met2 ;
        RECT 3377.035 2780.575 3379.435 2780.715 ;
        RECT 3375.640 2778.750 3376.240 2778.890 ;
        RECT 3377.020 2780.435 3379.435 2780.575 ;
        RECT 3375.120 2752.310 3375.380 2752.630 ;
        RECT 3375.640 2739.370 3375.780 2778.750 ;
        RECT 3377.020 2778.130 3377.160 2780.435 ;
      LAYER met2 ;
        RECT 3379.715 2780.155 3588.000 2780.995 ;
      LAYER met2 ;
        RECT 3376.040 2777.810 3376.300 2778.130 ;
        RECT 3376.960 2777.810 3377.220 2778.130 ;
        RECT 3376.100 2740.625 3376.240 2777.810 ;
      LAYER met2 ;
        RECT 3379.435 2777.775 3588.000 2780.155 ;
        RECT 3379.715 2776.935 3588.000 2777.775 ;
        RECT 3379.435 2775.015 3588.000 2776.935 ;
        RECT 3379.715 2774.175 3588.000 2775.015 ;
        RECT 3379.435 2771.795 3588.000 2774.175 ;
        RECT 3379.715 2770.955 3588.000 2771.795 ;
        RECT 3379.435 2768.575 3588.000 2770.955 ;
        RECT 3379.715 2767.735 3588.000 2768.575 ;
        RECT 3379.435 2765.815 3588.000 2767.735 ;
      LAYER met2 ;
        RECT 3377.035 2765.255 3379.435 2765.535 ;
      LAYER met2 ;
        RECT 3379.715 2764.975 3588.000 2765.815 ;
        RECT 3379.435 2762.595 3588.000 2764.975 ;
        RECT 3379.715 2761.755 3588.000 2762.595 ;
        RECT 3379.435 2759.375 3588.000 2761.755 ;
      LAYER met2 ;
        RECT 3377.035 2758.815 3379.435 2759.095 ;
      LAYER met2 ;
        RECT 3379.715 2758.535 3588.000 2759.375 ;
        RECT 3379.435 2756.615 3588.000 2758.535 ;
        RECT 3379.715 2755.775 3588.000 2756.615 ;
        RECT 3379.435 2753.395 3588.000 2755.775 ;
      LAYER met2 ;
        RECT 3376.960 2752.310 3377.220 2752.630 ;
      LAYER met2 ;
        RECT 3379.715 2752.555 3588.000 2753.395 ;
      LAYER met2 ;
        RECT 3377.020 2749.895 3377.160 2752.310 ;
      LAYER met2 ;
        RECT 3379.435 2750.175 3588.000 2752.555 ;
      LAYER met2 ;
        RECT 3377.020 2749.755 3379.435 2749.895 ;
        RECT 3377.035 2749.615 3379.435 2749.755 ;
      LAYER met2 ;
        RECT 3379.715 2749.335 3588.000 2750.175 ;
        RECT 3379.435 2747.415 3588.000 2749.335 ;
      LAYER met2 ;
        RECT 3377.035 2746.855 3379.435 2747.135 ;
      LAYER met2 ;
        RECT 3379.715 2746.575 3588.000 2747.415 ;
        RECT 3379.435 2744.195 3588.000 2746.575 ;
        RECT 3379.715 2743.355 3588.000 2744.195 ;
        RECT 3379.435 2740.975 3588.000 2743.355 ;
      LAYER met2 ;
        RECT 3377.035 2740.625 3379.435 2740.695 ;
        RECT 3376.100 2740.485 3379.435 2740.625 ;
        RECT 3377.035 2740.415 3379.435 2740.485 ;
      LAYER met2 ;
        RECT 3379.715 2740.135 3588.000 2740.975 ;
      LAYER met2 ;
        RECT 3375.640 2739.230 3376.700 2739.370 ;
        RECT 3376.560 2519.730 3376.700 2739.230 ;
      LAYER met2 ;
        RECT 3379.435 2739.085 3588.000 2740.135 ;
        RECT 3390.035 2593.505 3583.075 2593.735 ;
        RECT 3388.000 2569.605 3583.075 2593.505 ;
        RECT 3388.000 2566.105 3389.920 2568.105 ;
        RECT 3390.035 2543.610 3583.075 2569.605 ;
      LAYER met2 ;
        RECT 3376.500 2519.410 3376.760 2519.730 ;
        RECT 3387.540 2519.410 3387.800 2519.730 ;
      LAYER met2 ;
        RECT 3388.000 2519.710 3583.075 2543.610 ;
      LAYER met2 ;
        RECT 3387.600 2519.245 3387.740 2519.410 ;
        RECT 3387.530 2518.875 3387.810 2519.245 ;
      LAYER met2 ;
        RECT 3429.550 2374.000 3434.200 2384.975 ;
        RECT 3390.035 2373.500 3587.965 2374.000 ;
        RECT 3390.000 2353.505 3587.965 2373.500 ;
        RECT 3390.035 2353.075 3587.965 2353.505 ;
        RECT 3390.000 2320.465 3587.965 2353.075 ;
        RECT 3390.035 2319.905 3587.965 2320.465 ;
        RECT 3390.000 2299.300 3587.965 2319.905 ;
        RECT 3390.035 2299.000 3587.965 2299.300 ;
        RECT 3413.425 2288.065 3427.835 2297.800 ;
        RECT 3429.585 2287.860 3434.235 2299.000 ;
        RECT 3436.595 2288.065 3587.965 2297.800 ;
        RECT 3390.035 2152.505 3583.075 2152.735 ;
      LAYER met2 ;
        RECT 3387.540 2138.950 3387.800 2139.270 ;
        RECT 3387.600 2128.245 3387.740 2138.950 ;
      LAYER met2 ;
        RECT 3388.000 2128.605 3583.075 2152.505 ;
      LAYER met2 ;
        RECT 3387.530 2127.875 3387.810 2128.245 ;
      LAYER met2 ;
        RECT 3388.000 2125.105 3389.920 2127.105 ;
        RECT 3390.035 2102.610 3583.075 2128.605 ;
        RECT 3388.000 2078.710 3583.075 2102.610 ;
        RECT 3379.435 1931.795 3588.000 1932.790 ;
      LAYER met2 ;
        RECT 3377.035 1931.235 3379.435 1931.515 ;
      LAYER met2 ;
        RECT 3379.715 1930.955 3588.000 1931.795 ;
        RECT 3379.435 1929.035 3588.000 1930.955 ;
        RECT 3379.715 1928.195 3588.000 1929.035 ;
        RECT 3379.435 1925.815 3588.000 1928.195 ;
        RECT 3379.715 1924.975 3588.000 1925.815 ;
        RECT 3379.435 1922.595 3588.000 1924.975 ;
        RECT 3379.715 1921.755 3588.000 1922.595 ;
        RECT 3379.435 1919.835 3588.000 1921.755 ;
        RECT 3379.715 1918.995 3588.000 1919.835 ;
      LAYER met2 ;
        RECT 3374.200 1918.630 3374.460 1918.950 ;
        RECT 3376.960 1918.630 3377.220 1918.950 ;
        RECT 3374.260 1897.570 3374.400 1918.630 ;
        RECT 3377.020 1916.335 3377.160 1918.630 ;
      LAYER met2 ;
        RECT 3379.435 1916.615 3588.000 1918.995 ;
      LAYER met2 ;
        RECT 3377.020 1916.195 3379.435 1916.335 ;
        RECT 3377.035 1916.055 3379.435 1916.195 ;
      LAYER met2 ;
        RECT 3379.715 1915.775 3588.000 1916.615 ;
        RECT 3379.435 1913.395 3588.000 1915.775 ;
        RECT 3379.715 1912.555 3588.000 1913.395 ;
        RECT 3379.435 1910.635 3588.000 1912.555 ;
        RECT 3379.715 1909.795 3588.000 1910.635 ;
        RECT 3379.435 1907.415 3588.000 1909.795 ;
        RECT 3379.715 1906.575 3588.000 1907.415 ;
        RECT 3379.435 1904.195 3588.000 1906.575 ;
        RECT 3379.715 1903.355 3588.000 1904.195 ;
        RECT 3379.435 1901.435 3588.000 1903.355 ;
      LAYER met2 ;
        RECT 3377.035 1900.940 3379.435 1901.155 ;
        RECT 3377.020 1900.875 3379.435 1900.940 ;
        RECT 3377.020 1899.230 3377.160 1900.875 ;
      LAYER met2 ;
        RECT 3379.715 1900.595 3588.000 1901.435 ;
      LAYER met2 ;
        RECT 3375.120 1898.910 3375.380 1899.230 ;
        RECT 3376.960 1898.910 3377.220 1899.230 ;
        RECT 3374.260 1897.430 3374.860 1897.570 ;
        RECT 3374.200 1891.770 3374.460 1892.090 ;
        RECT 3374.260 1857.410 3374.400 1891.770 ;
        RECT 3374.200 1857.090 3374.460 1857.410 ;
        RECT 213.080 1843.150 213.340 1843.470 ;
        RECT 212.620 1801.670 212.880 1801.990 ;
        RECT 208.940 1786.030 209.200 1786.350 ;
        RECT 212.160 1786.030 212.420 1786.350 ;
      LAYER met2 ;
        RECT 0.000 1785.165 208.285 1786.005 ;
        RECT 0.000 1783.245 208.565 1785.165 ;
      LAYER met2 ;
        RECT 211.240 1785.010 211.500 1785.330 ;
      LAYER met2 ;
        RECT 0.000 1782.405 208.285 1783.245 ;
        RECT 0.000 1780.025 208.565 1782.405 ;
        RECT 0.000 1779.185 208.285 1780.025 ;
        RECT 0.000 1776.805 208.565 1779.185 ;
        RECT 0.000 1775.965 208.285 1776.805 ;
        RECT 0.000 1774.045 208.565 1775.965 ;
        RECT 0.000 1773.205 208.285 1774.045 ;
      LAYER met2 ;
        RECT 208.565 1773.485 210.965 1773.765 ;
      LAYER met2 ;
        RECT 0.000 1772.210 208.565 1773.205 ;
        RECT 0.000 1634.865 208.565 1635.915 ;
        RECT 0.000 1634.025 208.285 1634.865 ;
      LAYER met2 ;
        RECT 208.565 1634.305 210.965 1634.585 ;
      LAYER met2 ;
        RECT 0.000 1631.645 208.565 1634.025 ;
      LAYER met2 ;
        RECT 209.000 1631.990 209.140 1634.305 ;
        RECT 208.940 1631.670 209.200 1631.990 ;
      LAYER met2 ;
        RECT 0.000 1630.805 208.285 1631.645 ;
        RECT 0.000 1628.425 208.565 1630.805 ;
        RECT 0.000 1627.585 208.285 1628.425 ;
      LAYER met2 ;
        RECT 208.565 1627.865 210.965 1628.145 ;
      LAYER met2 ;
        RECT 0.000 1625.665 208.565 1627.585 ;
        RECT 0.000 1624.825 208.285 1625.665 ;
      LAYER met2 ;
        RECT 208.940 1625.550 209.200 1625.870 ;
        RECT 209.000 1625.385 209.140 1625.550 ;
        RECT 208.565 1625.105 210.965 1625.385 ;
      LAYER met2 ;
        RECT 0.000 1622.445 208.565 1624.825 ;
        RECT 0.000 1621.605 208.285 1622.445 ;
        RECT 0.000 1619.225 208.565 1621.605 ;
        RECT 0.000 1618.385 208.285 1619.225 ;
        RECT 0.000 1616.465 208.565 1618.385 ;
        RECT 0.000 1615.625 208.285 1616.465 ;
      LAYER met2 ;
        RECT 208.565 1615.905 210.965 1616.185 ;
      LAYER met2 ;
        RECT 0.000 1613.245 208.565 1615.625 ;
        RECT 0.000 1612.405 208.285 1613.245 ;
        RECT 0.000 1610.025 208.565 1612.405 ;
        RECT 0.000 1609.185 208.285 1610.025 ;
      LAYER met2 ;
        RECT 208.565 1609.465 210.965 1609.745 ;
      LAYER met2 ;
        RECT 0.000 1607.265 208.565 1609.185 ;
        RECT 0.000 1606.425 208.285 1607.265 ;
        RECT 0.000 1604.045 208.565 1606.425 ;
        RECT 0.000 1603.205 208.285 1604.045 ;
        RECT 0.000 1600.825 208.565 1603.205 ;
        RECT 0.000 1599.985 208.285 1600.825 ;
        RECT 0.000 1598.065 208.565 1599.985 ;
        RECT 0.000 1597.225 208.285 1598.065 ;
        RECT 0.000 1594.845 208.565 1597.225 ;
      LAYER met2 ;
        RECT 208.940 1596.990 209.200 1597.310 ;
      LAYER met2 ;
        RECT 0.000 1594.005 208.285 1594.845 ;
      LAYER met2 ;
        RECT 209.000 1594.565 209.140 1596.990 ;
        RECT 208.565 1594.285 210.965 1594.565 ;
      LAYER met2 ;
        RECT 0.000 1591.625 208.565 1594.005 ;
        RECT 0.000 1590.785 208.285 1591.625 ;
        RECT 0.000 1588.405 208.565 1590.785 ;
      LAYER met2 ;
        RECT 208.940 1590.530 209.200 1590.850 ;
      LAYER met2 ;
        RECT 0.000 1587.565 208.285 1588.405 ;
      LAYER met2 ;
        RECT 209.000 1588.125 209.140 1590.530 ;
        RECT 208.565 1587.845 210.965 1588.125 ;
      LAYER met2 ;
        RECT 0.000 1585.645 208.565 1587.565 ;
        RECT 0.000 1584.805 208.285 1585.645 ;
        RECT 0.000 1582.425 208.565 1584.805 ;
        RECT 0.000 1581.585 208.285 1582.425 ;
        RECT 0.000 1579.205 208.565 1581.585 ;
        RECT 0.000 1578.365 208.285 1579.205 ;
        RECT 0.000 1576.445 208.565 1578.365 ;
        RECT 0.000 1575.605 208.285 1576.445 ;
        RECT 0.000 1573.225 208.565 1575.605 ;
        RECT 0.000 1572.385 208.285 1573.225 ;
      LAYER met2 ;
        RECT 208.565 1572.665 210.965 1572.945 ;
      LAYER met2 ;
        RECT 0.000 1570.005 208.565 1572.385 ;
      LAYER met2 ;
        RECT 209.000 1570.530 209.140 1572.665 ;
        RECT 211.300 1570.530 211.440 1785.010 ;
        RECT 212.160 1631.670 212.420 1631.990 ;
        RECT 212.220 1597.310 212.360 1631.670 ;
        RECT 213.140 1628.470 213.280 1843.150 ;
        RECT 213.540 1801.670 213.800 1801.990 ;
        RECT 212.680 1628.330 213.280 1628.470 ;
        RECT 212.680 1625.870 212.820 1628.330 ;
        RECT 212.620 1625.550 212.880 1625.870 ;
        RECT 212.160 1596.990 212.420 1597.310 ;
        RECT 209.000 1570.390 211.440 1570.530 ;
      LAYER met2 ;
        RECT 0.000 1569.165 208.285 1570.005 ;
        RECT 0.000 1567.245 208.565 1569.165 ;
        RECT 0.000 1566.405 208.285 1567.245 ;
        RECT 0.000 1564.025 208.565 1566.405 ;
        RECT 0.000 1563.185 208.285 1564.025 ;
        RECT 0.000 1560.805 208.565 1563.185 ;
        RECT 0.000 1559.965 208.285 1560.805 ;
        RECT 0.000 1558.045 208.565 1559.965 ;
        RECT 0.000 1557.205 208.285 1558.045 ;
      LAYER met2 ;
        RECT 208.565 1557.485 210.965 1557.765 ;
      LAYER met2 ;
        RECT 0.000 1556.210 208.565 1557.205 ;
        RECT 0.000 1418.865 208.565 1419.915 ;
        RECT 0.000 1418.025 208.285 1418.865 ;
      LAYER met2 ;
        RECT 208.565 1418.305 210.965 1418.585 ;
      LAYER met2 ;
        RECT 0.000 1415.645 208.565 1418.025 ;
      LAYER met2 ;
        RECT 209.000 1416.090 209.140 1418.305 ;
        RECT 208.940 1415.770 209.200 1416.090 ;
      LAYER met2 ;
        RECT 0.000 1414.805 208.285 1415.645 ;
        RECT 0.000 1412.425 208.565 1414.805 ;
        RECT 0.000 1411.585 208.285 1412.425 ;
      LAYER met2 ;
        RECT 208.565 1411.865 210.965 1412.145 ;
      LAYER met2 ;
        RECT 0.000 1409.665 208.565 1411.585 ;
      LAYER met2 ;
        RECT 208.940 1410.330 209.200 1410.650 ;
      LAYER met2 ;
        RECT 0.000 1408.825 208.285 1409.665 ;
      LAYER met2 ;
        RECT 209.000 1409.385 209.140 1410.330 ;
        RECT 208.565 1409.105 210.965 1409.385 ;
      LAYER met2 ;
        RECT 0.000 1406.445 208.565 1408.825 ;
        RECT 0.000 1405.605 208.285 1406.445 ;
        RECT 0.000 1403.225 208.565 1405.605 ;
        RECT 0.000 1402.385 208.285 1403.225 ;
        RECT 0.000 1400.465 208.565 1402.385 ;
        RECT 0.000 1399.625 208.285 1400.465 ;
      LAYER met2 ;
        RECT 208.565 1399.905 210.965 1400.185 ;
      LAYER met2 ;
        RECT 0.000 1397.245 208.565 1399.625 ;
        RECT 0.000 1396.405 208.285 1397.245 ;
        RECT 0.000 1394.025 208.565 1396.405 ;
        RECT 0.000 1393.185 208.285 1394.025 ;
      LAYER met2 ;
        RECT 208.565 1393.465 210.965 1393.745 ;
      LAYER met2 ;
        RECT 0.000 1391.265 208.565 1393.185 ;
        RECT 0.000 1390.425 208.285 1391.265 ;
        RECT 0.000 1388.045 208.565 1390.425 ;
        RECT 0.000 1387.205 208.285 1388.045 ;
        RECT 0.000 1384.825 208.565 1387.205 ;
        RECT 0.000 1383.985 208.285 1384.825 ;
        RECT 0.000 1382.065 208.565 1383.985 ;
        RECT 0.000 1381.225 208.285 1382.065 ;
        RECT 0.000 1378.845 208.565 1381.225 ;
      LAYER met2 ;
        RECT 208.940 1380.750 209.200 1381.070 ;
      LAYER met2 ;
        RECT 0.000 1378.005 208.285 1378.845 ;
      LAYER met2 ;
        RECT 209.000 1378.565 209.140 1380.750 ;
        RECT 208.565 1378.285 210.965 1378.565 ;
      LAYER met2 ;
        RECT 0.000 1375.625 208.565 1378.005 ;
        RECT 0.000 1374.785 208.285 1375.625 ;
        RECT 0.000 1372.405 208.565 1374.785 ;
        RECT 0.000 1371.565 208.285 1372.405 ;
      LAYER met2 ;
        RECT 208.565 1371.845 210.965 1372.125 ;
        RECT 208.610 1371.830 209.140 1371.845 ;
      LAYER met2 ;
        RECT 0.000 1369.645 208.565 1371.565 ;
      LAYER met2 ;
        RECT 209.000 1369.850 209.140 1371.830 ;
      LAYER met2 ;
        RECT 0.000 1368.805 208.285 1369.645 ;
      LAYER met2 ;
        RECT 208.940 1369.530 209.200 1369.850 ;
      LAYER met2 ;
        RECT 0.000 1366.425 208.565 1368.805 ;
        RECT 0.000 1365.585 208.285 1366.425 ;
        RECT 0.000 1363.205 208.565 1365.585 ;
        RECT 0.000 1362.365 208.285 1363.205 ;
        RECT 0.000 1360.445 208.565 1362.365 ;
        RECT 0.000 1359.605 208.285 1360.445 ;
        RECT 0.000 1357.225 208.565 1359.605 ;
      LAYER met2 ;
        RECT 211.300 1357.690 211.440 1570.390 ;
        RECT 212.160 1415.770 212.420 1416.090 ;
        RECT 212.220 1381.070 212.360 1415.770 ;
        RECT 212.680 1410.650 212.820 1625.550 ;
        RECT 213.600 1590.850 213.740 1801.670 ;
        RECT 3374.720 1687.750 3374.860 1897.430 ;
        RECT 3374.660 1687.430 3374.920 1687.750 ;
        RECT 3374.200 1640.170 3374.460 1640.490 ;
        RECT 213.540 1590.530 213.800 1590.850 ;
        RECT 213.600 1580.170 213.740 1590.530 ;
        RECT 213.140 1580.030 213.740 1580.170 ;
        RECT 212.620 1410.330 212.880 1410.650 ;
        RECT 212.160 1380.750 212.420 1381.070 ;
        RECT 209.000 1357.550 211.440 1357.690 ;
      LAYER met2 ;
        RECT 0.000 1356.385 208.285 1357.225 ;
      LAYER met2 ;
        RECT 209.000 1357.010 209.140 1357.550 ;
        RECT 208.610 1356.945 209.140 1357.010 ;
        RECT 208.565 1356.665 210.965 1356.945 ;
      LAYER met2 ;
        RECT 0.000 1354.005 208.565 1356.385 ;
        RECT 0.000 1353.165 208.285 1354.005 ;
        RECT 0.000 1351.245 208.565 1353.165 ;
        RECT 0.000 1350.405 208.285 1351.245 ;
        RECT 0.000 1348.025 208.565 1350.405 ;
        RECT 0.000 1347.185 208.285 1348.025 ;
        RECT 0.000 1344.805 208.565 1347.185 ;
        RECT 0.000 1343.965 208.285 1344.805 ;
        RECT 0.000 1342.045 208.565 1343.965 ;
        RECT 0.000 1341.205 208.285 1342.045 ;
      LAYER met2 ;
        RECT 208.565 1341.485 210.965 1341.765 ;
      LAYER met2 ;
        RECT 0.000 1340.210 208.565 1341.205 ;
        RECT 0.000 1202.865 208.565 1203.915 ;
        RECT 0.000 1202.025 208.285 1202.865 ;
      LAYER met2 ;
        RECT 208.610 1202.585 209.140 1202.650 ;
        RECT 208.565 1202.305 210.965 1202.585 ;
      LAYER met2 ;
        RECT 0.000 1199.645 208.565 1202.025 ;
      LAYER met2 ;
        RECT 209.000 1199.850 209.140 1202.305 ;
      LAYER met2 ;
        RECT 0.000 1198.805 208.285 1199.645 ;
      LAYER met2 ;
        RECT 208.940 1199.530 209.200 1199.850 ;
      LAYER met2 ;
        RECT 0.000 1196.425 208.565 1198.805 ;
        RECT 0.000 1195.585 208.285 1196.425 ;
      LAYER met2 ;
        RECT 208.565 1195.865 210.965 1196.145 ;
      LAYER met2 ;
        RECT 0.000 1193.665 208.565 1195.585 ;
        RECT 0.000 1192.825 208.285 1193.665 ;
      LAYER met2 ;
        RECT 208.565 1193.105 210.965 1193.385 ;
      LAYER met2 ;
        RECT 0.000 1190.445 208.565 1192.825 ;
      LAYER met2 ;
        RECT 209.000 1192.710 209.140 1193.105 ;
        RECT 208.940 1192.390 209.200 1192.710 ;
      LAYER met2 ;
        RECT 0.000 1189.605 208.285 1190.445 ;
        RECT 0.000 1187.225 208.565 1189.605 ;
        RECT 0.000 1186.385 208.285 1187.225 ;
      LAYER met2 ;
        RECT 208.565 1186.665 210.965 1186.945 ;
      LAYER met2 ;
        RECT 0.000 1184.465 208.565 1186.385 ;
        RECT 0.000 1183.625 208.285 1184.465 ;
      LAYER met2 ;
        RECT 208.565 1183.905 210.965 1184.185 ;
      LAYER met2 ;
        RECT 0.000 1181.245 208.565 1183.625 ;
        RECT 0.000 1180.405 208.285 1181.245 ;
        RECT 0.000 1178.025 208.565 1180.405 ;
        RECT 0.000 1177.185 208.285 1178.025 ;
      LAYER met2 ;
        RECT 208.565 1177.465 210.965 1177.745 ;
      LAYER met2 ;
        RECT 0.000 1175.265 208.565 1177.185 ;
        RECT 0.000 1174.425 208.285 1175.265 ;
        RECT 0.000 1172.045 208.565 1174.425 ;
        RECT 0.000 1171.205 208.285 1172.045 ;
        RECT 0.000 1168.825 208.565 1171.205 ;
        RECT 0.000 1167.985 208.285 1168.825 ;
        RECT 0.000 1166.065 208.565 1167.985 ;
        RECT 0.000 1165.225 208.285 1166.065 ;
        RECT 0.000 1162.845 208.565 1165.225 ;
      LAYER met2 ;
        RECT 208.940 1164.850 209.200 1165.170 ;
      LAYER met2 ;
        RECT 0.000 1162.005 208.285 1162.845 ;
      LAYER met2 ;
        RECT 209.000 1162.565 209.140 1164.850 ;
        RECT 208.565 1162.285 210.965 1162.565 ;
      LAYER met2 ;
        RECT 0.000 1159.625 208.565 1162.005 ;
        RECT 0.000 1158.785 208.285 1159.625 ;
        RECT 0.000 1156.405 208.565 1158.785 ;
      LAYER met2 ;
        RECT 208.940 1158.390 209.200 1158.710 ;
      LAYER met2 ;
        RECT 0.000 1155.565 208.285 1156.405 ;
      LAYER met2 ;
        RECT 209.000 1156.125 209.140 1158.390 ;
        RECT 208.565 1155.845 210.965 1156.125 ;
      LAYER met2 ;
        RECT 0.000 1153.645 208.565 1155.565 ;
        RECT 0.000 1152.805 208.285 1153.645 ;
        RECT 0.000 1150.425 208.565 1152.805 ;
        RECT 0.000 1149.585 208.285 1150.425 ;
        RECT 0.000 1147.205 208.565 1149.585 ;
        RECT 0.000 1146.365 208.285 1147.205 ;
        RECT 0.000 1144.445 208.565 1146.365 ;
        RECT 0.000 1143.605 208.285 1144.445 ;
        RECT 0.000 1141.225 208.565 1143.605 ;
        RECT 0.000 1140.385 208.285 1141.225 ;
      LAYER met2 ;
        RECT 208.565 1140.665 210.965 1140.945 ;
        RECT 208.610 1140.630 209.140 1140.665 ;
      LAYER met2 ;
        RECT 0.000 1138.005 208.565 1140.385 ;
      LAYER met2 ;
        RECT 209.000 1138.050 209.140 1140.630 ;
        RECT 211.300 1138.050 211.440 1357.550 ;
        RECT 212.160 1199.530 212.420 1199.850 ;
        RECT 212.220 1165.170 212.360 1199.530 ;
        RECT 212.680 1192.710 212.820 1410.330 ;
        RECT 213.140 1369.850 213.280 1580.030 ;
        RECT 3374.260 1411.670 3374.400 1640.170 ;
        RECT 3374.720 1466.410 3374.860 1687.430 ;
        RECT 3375.180 1677.210 3375.320 1898.910 ;
      LAYER met2 ;
        RECT 3379.435 1898.215 3588.000 1900.595 ;
        RECT 3379.715 1897.375 3588.000 1898.215 ;
        RECT 3379.435 1894.995 3588.000 1897.375 ;
      LAYER met2 ;
        RECT 3377.035 1894.575 3379.435 1894.715 ;
        RECT 3377.020 1894.435 3379.435 1894.575 ;
        RECT 3377.020 1892.090 3377.160 1894.435 ;
      LAYER met2 ;
        RECT 3379.715 1894.155 3588.000 1894.995 ;
      LAYER met2 ;
        RECT 3376.960 1891.770 3377.220 1892.090 ;
      LAYER met2 ;
        RECT 3379.435 1891.775 3588.000 1894.155 ;
        RECT 3379.715 1890.935 3588.000 1891.775 ;
        RECT 3379.435 1889.015 3588.000 1890.935 ;
        RECT 3379.715 1888.175 3588.000 1889.015 ;
        RECT 3379.435 1885.795 3588.000 1888.175 ;
        RECT 3379.715 1884.955 3588.000 1885.795 ;
        RECT 3379.435 1882.575 3588.000 1884.955 ;
        RECT 3379.715 1881.735 3588.000 1882.575 ;
        RECT 3379.435 1879.815 3588.000 1881.735 ;
      LAYER met2 ;
        RECT 3377.035 1879.255 3379.435 1879.535 ;
      LAYER met2 ;
        RECT 3379.715 1878.975 3588.000 1879.815 ;
        RECT 3379.435 1876.595 3588.000 1878.975 ;
        RECT 3379.715 1875.755 3588.000 1876.595 ;
        RECT 3379.435 1873.375 3588.000 1875.755 ;
      LAYER met2 ;
        RECT 3377.035 1872.815 3379.435 1873.095 ;
      LAYER met2 ;
        RECT 3379.715 1872.535 3588.000 1873.375 ;
        RECT 3379.435 1870.615 3588.000 1872.535 ;
      LAYER met2 ;
        RECT 3377.035 1870.055 3379.435 1870.335 ;
      LAYER met2 ;
        RECT 3379.715 1869.775 3588.000 1870.615 ;
        RECT 3379.435 1867.395 3588.000 1869.775 ;
        RECT 3379.715 1866.555 3588.000 1867.395 ;
        RECT 3379.435 1864.175 3588.000 1866.555 ;
      LAYER met2 ;
        RECT 3377.035 1863.825 3379.435 1863.895 ;
        RECT 3376.100 1863.685 3379.435 1863.825 ;
        RECT 3376.100 1680.010 3376.240 1863.685 ;
        RECT 3377.035 1863.615 3379.435 1863.685 ;
      LAYER met2 ;
        RECT 3379.715 1863.335 3588.000 1864.175 ;
        RECT 3379.435 1861.415 3588.000 1863.335 ;
      LAYER met2 ;
        RECT 3377.035 1860.855 3379.435 1861.135 ;
      LAYER met2 ;
        RECT 3379.715 1860.575 3588.000 1861.415 ;
        RECT 3379.435 1858.195 3588.000 1860.575 ;
      LAYER met2 ;
        RECT 3376.960 1857.090 3377.220 1857.410 ;
      LAYER met2 ;
        RECT 3379.715 1857.355 3588.000 1858.195 ;
      LAYER met2 ;
        RECT 3377.020 1854.695 3377.160 1857.090 ;
      LAYER met2 ;
        RECT 3379.435 1854.975 3588.000 1857.355 ;
      LAYER met2 ;
        RECT 3377.020 1854.555 3379.435 1854.695 ;
        RECT 3377.035 1854.415 3379.435 1854.555 ;
      LAYER met2 ;
        RECT 3379.715 1854.135 3588.000 1854.975 ;
        RECT 3379.435 1853.085 3588.000 1854.135 ;
        RECT 3379.435 1705.795 3588.000 1706.790 ;
      LAYER met2 ;
        RECT 3377.035 1705.235 3379.435 1705.515 ;
      LAYER met2 ;
        RECT 3379.715 1704.955 3588.000 1705.795 ;
        RECT 3379.435 1703.035 3588.000 1704.955 ;
        RECT 3379.715 1702.195 3588.000 1703.035 ;
        RECT 3379.435 1699.815 3588.000 1702.195 ;
        RECT 3379.715 1698.975 3588.000 1699.815 ;
        RECT 3379.435 1696.595 3588.000 1698.975 ;
        RECT 3379.715 1695.755 3588.000 1696.595 ;
        RECT 3379.435 1693.835 3588.000 1695.755 ;
        RECT 3379.715 1692.995 3588.000 1693.835 ;
        RECT 3379.435 1690.615 3588.000 1692.995 ;
      LAYER met2 ;
        RECT 3377.035 1690.140 3379.435 1690.335 ;
        RECT 3377.020 1690.055 3379.435 1690.140 ;
        RECT 3377.020 1687.750 3377.160 1690.055 ;
      LAYER met2 ;
        RECT 3379.715 1689.775 3588.000 1690.615 ;
      LAYER met2 ;
        RECT 3376.960 1687.430 3377.220 1687.750 ;
      LAYER met2 ;
        RECT 3379.435 1687.395 3588.000 1689.775 ;
        RECT 3379.715 1686.555 3588.000 1687.395 ;
        RECT 3379.435 1684.635 3588.000 1686.555 ;
        RECT 3379.715 1683.795 3588.000 1684.635 ;
        RECT 3379.435 1681.415 3588.000 1683.795 ;
        RECT 3379.715 1680.575 3588.000 1681.415 ;
      LAYER met2 ;
        RECT 3375.640 1679.870 3376.240 1680.010 ;
        RECT 3375.120 1676.890 3375.380 1677.210 ;
        RECT 3375.640 1640.490 3375.780 1679.870 ;
      LAYER met2 ;
        RECT 3379.435 1678.195 3588.000 1680.575 ;
        RECT 3379.715 1677.355 3588.000 1678.195 ;
      LAYER met2 ;
        RECT 3376.040 1676.890 3376.300 1677.210 ;
        RECT 3376.960 1676.890 3377.220 1677.210 ;
        RECT 3375.580 1640.170 3375.840 1640.490 ;
        RECT 3376.100 1580.170 3376.240 1676.890 ;
        RECT 3377.020 1675.155 3377.160 1676.890 ;
      LAYER met2 ;
        RECT 3379.435 1675.435 3588.000 1677.355 ;
      LAYER met2 ;
        RECT 3377.020 1675.015 3379.435 1675.155 ;
        RECT 3377.035 1674.875 3379.435 1675.015 ;
      LAYER met2 ;
        RECT 3379.715 1674.595 3588.000 1675.435 ;
        RECT 3379.435 1672.215 3588.000 1674.595 ;
        RECT 3379.715 1671.375 3588.000 1672.215 ;
        RECT 3379.435 1668.995 3588.000 1671.375 ;
      LAYER met2 ;
        RECT 3377.035 1668.645 3379.435 1668.715 ;
        RECT 3376.560 1668.505 3379.435 1668.645 ;
        RECT 3376.560 1628.625 3376.700 1668.505 ;
        RECT 3377.035 1668.435 3379.435 1668.505 ;
      LAYER met2 ;
        RECT 3379.715 1668.155 3588.000 1668.995 ;
        RECT 3379.435 1665.775 3588.000 1668.155 ;
        RECT 3379.715 1664.935 3588.000 1665.775 ;
        RECT 3379.435 1663.015 3588.000 1664.935 ;
        RECT 3379.715 1662.175 3588.000 1663.015 ;
        RECT 3379.435 1659.795 3588.000 1662.175 ;
        RECT 3379.715 1658.955 3588.000 1659.795 ;
        RECT 3379.435 1656.575 3588.000 1658.955 ;
        RECT 3379.715 1655.735 3588.000 1656.575 ;
        RECT 3379.435 1653.815 3588.000 1655.735 ;
      LAYER met2 ;
        RECT 3377.035 1653.255 3379.435 1653.535 ;
      LAYER met2 ;
        RECT 3379.715 1652.975 3588.000 1653.815 ;
        RECT 3379.435 1650.595 3588.000 1652.975 ;
        RECT 3379.715 1649.755 3588.000 1650.595 ;
        RECT 3379.435 1647.375 3588.000 1649.755 ;
      LAYER met2 ;
        RECT 3377.035 1646.815 3379.435 1647.095 ;
      LAYER met2 ;
        RECT 3379.715 1646.535 3588.000 1647.375 ;
        RECT 3379.435 1644.615 3588.000 1646.535 ;
      LAYER met2 ;
        RECT 3377.035 1644.055 3379.435 1644.335 ;
      LAYER met2 ;
        RECT 3379.715 1643.775 3588.000 1644.615 ;
        RECT 3379.435 1641.395 3588.000 1643.775 ;
        RECT 3379.715 1640.555 3588.000 1641.395 ;
      LAYER met2 ;
        RECT 3376.960 1640.170 3377.220 1640.490 ;
        RECT 3377.020 1637.895 3377.160 1640.170 ;
      LAYER met2 ;
        RECT 3379.435 1638.175 3588.000 1640.555 ;
      LAYER met2 ;
        RECT 3377.020 1637.780 3379.435 1637.895 ;
        RECT 3377.035 1637.615 3379.435 1637.780 ;
      LAYER met2 ;
        RECT 3379.715 1637.335 3588.000 1638.175 ;
        RECT 3379.435 1635.415 3588.000 1637.335 ;
      LAYER met2 ;
        RECT 3377.035 1634.855 3379.435 1635.135 ;
      LAYER met2 ;
        RECT 3379.715 1634.575 3588.000 1635.415 ;
        RECT 3379.435 1632.195 3588.000 1634.575 ;
        RECT 3379.715 1631.355 3588.000 1632.195 ;
        RECT 3379.435 1628.975 3588.000 1631.355 ;
      LAYER met2 ;
        RECT 3377.035 1628.625 3379.435 1628.695 ;
        RECT 3376.560 1628.485 3379.435 1628.625 ;
        RECT 3377.035 1628.415 3379.435 1628.485 ;
      LAYER met2 ;
        RECT 3379.715 1628.135 3588.000 1628.975 ;
        RECT 3379.435 1627.085 3588.000 1628.135 ;
      LAYER met2 ;
        RECT 3375.640 1580.030 3376.240 1580.170 ;
        RECT 3375.640 1531.870 3375.780 1580.030 ;
        RECT 3375.640 1531.730 3376.240 1531.870 ;
        RECT 3376.100 1511.170 3376.240 1531.730 ;
        RECT 3376.100 1511.030 3376.700 1511.170 ;
        RECT 3376.560 1469.890 3376.700 1511.030 ;
      LAYER met2 ;
        RECT 3379.435 1480.795 3588.000 1481.790 ;
      LAYER met2 ;
        RECT 3377.035 1480.235 3379.435 1480.515 ;
      LAYER met2 ;
        RECT 3379.715 1479.955 3588.000 1480.795 ;
        RECT 3379.435 1478.035 3588.000 1479.955 ;
        RECT 3379.715 1477.195 3588.000 1478.035 ;
        RECT 3379.435 1474.815 3588.000 1477.195 ;
        RECT 3379.715 1473.975 3588.000 1474.815 ;
        RECT 3379.435 1471.595 3588.000 1473.975 ;
        RECT 3379.715 1470.755 3588.000 1471.595 ;
      LAYER met2 ;
        RECT 3375.640 1469.750 3376.700 1469.890 ;
        RECT 3374.660 1466.090 3374.920 1466.410 ;
        RECT 3374.720 1449.070 3374.860 1466.090 ;
        RECT 3374.720 1448.930 3375.320 1449.070 ;
        RECT 3374.660 1447.390 3374.920 1447.710 ;
        RECT 3374.200 1411.350 3374.460 1411.670 ;
        RECT 213.080 1369.530 213.340 1369.850 ;
        RECT 212.620 1192.390 212.880 1192.710 ;
        RECT 212.160 1164.850 212.420 1165.170 ;
      LAYER met2 ;
        RECT 0.000 1137.165 208.285 1138.005 ;
      LAYER met2 ;
        RECT 209.000 1137.910 211.440 1138.050 ;
      LAYER met2 ;
        RECT 0.000 1135.245 208.565 1137.165 ;
        RECT 0.000 1134.405 208.285 1135.245 ;
        RECT 0.000 1132.025 208.565 1134.405 ;
        RECT 0.000 1131.185 208.285 1132.025 ;
        RECT 0.000 1128.805 208.565 1131.185 ;
        RECT 0.000 1127.965 208.285 1128.805 ;
        RECT 0.000 1126.045 208.565 1127.965 ;
        RECT 0.000 1125.205 208.285 1126.045 ;
      LAYER met2 ;
        RECT 208.565 1125.485 210.965 1125.765 ;
      LAYER met2 ;
        RECT 0.000 1124.210 208.565 1125.205 ;
        RECT 0.000 986.865 208.565 987.915 ;
        RECT 0.000 986.025 208.285 986.865 ;
      LAYER met2 ;
        RECT 208.565 986.305 210.965 986.585 ;
        RECT 208.610 986.270 209.140 986.305 ;
      LAYER met2 ;
        RECT 0.000 983.645 208.565 986.025 ;
      LAYER met2 ;
        RECT 209.000 983.950 209.140 986.270 ;
      LAYER met2 ;
        RECT 0.000 982.805 208.285 983.645 ;
      LAYER met2 ;
        RECT 208.940 983.630 209.200 983.950 ;
      LAYER met2 ;
        RECT 0.000 980.425 208.565 982.805 ;
        RECT 0.000 979.585 208.285 980.425 ;
      LAYER met2 ;
        RECT 208.565 979.865 210.965 980.145 ;
      LAYER met2 ;
        RECT 0.000 977.665 208.565 979.585 ;
        RECT 0.000 976.825 208.285 977.665 ;
      LAYER met2 ;
        RECT 208.565 977.105 210.965 977.385 ;
      LAYER met2 ;
        RECT 0.000 974.445 208.565 976.825 ;
      LAYER met2 ;
        RECT 209.000 976.810 209.140 977.105 ;
        RECT 208.940 976.490 209.200 976.810 ;
      LAYER met2 ;
        RECT 0.000 973.605 208.285 974.445 ;
        RECT 0.000 971.225 208.565 973.605 ;
        RECT 0.000 970.385 208.285 971.225 ;
      LAYER met2 ;
        RECT 208.565 970.665 210.965 970.945 ;
      LAYER met2 ;
        RECT 0.000 968.465 208.565 970.385 ;
        RECT 0.000 967.625 208.285 968.465 ;
      LAYER met2 ;
        RECT 208.565 967.905 210.965 968.185 ;
      LAYER met2 ;
        RECT 0.000 965.245 208.565 967.625 ;
        RECT 0.000 964.405 208.285 965.245 ;
        RECT 0.000 962.025 208.565 964.405 ;
        RECT 0.000 961.185 208.285 962.025 ;
      LAYER met2 ;
        RECT 208.565 961.465 210.965 961.745 ;
      LAYER met2 ;
        RECT 0.000 959.265 208.565 961.185 ;
        RECT 0.000 958.425 208.285 959.265 ;
        RECT 0.000 956.045 208.565 958.425 ;
        RECT 0.000 955.205 208.285 956.045 ;
        RECT 0.000 952.825 208.565 955.205 ;
        RECT 0.000 951.985 208.285 952.825 ;
        RECT 0.000 950.065 208.565 951.985 ;
        RECT 0.000 949.225 208.285 950.065 ;
        RECT 0.000 946.845 208.565 949.225 ;
      LAYER met2 ;
        RECT 208.940 948.950 209.200 949.270 ;
      LAYER met2 ;
        RECT 0.000 946.005 208.285 946.845 ;
      LAYER met2 ;
        RECT 209.000 946.565 209.140 948.950 ;
        RECT 208.565 946.285 210.965 946.565 ;
      LAYER met2 ;
        RECT 0.000 943.625 208.565 946.005 ;
        RECT 0.000 942.785 208.285 943.625 ;
        RECT 0.000 940.405 208.565 942.785 ;
        RECT 0.000 939.565 208.285 940.405 ;
      LAYER met2 ;
        RECT 208.610 940.125 209.140 940.170 ;
        RECT 208.565 939.845 210.965 940.125 ;
      LAYER met2 ;
        RECT 0.000 937.645 208.565 939.565 ;
      LAYER met2 ;
        RECT 209.000 938.050 209.140 939.845 ;
        RECT 208.940 937.730 209.200 938.050 ;
      LAYER met2 ;
        RECT 0.000 936.805 208.285 937.645 ;
        RECT 0.000 934.425 208.565 936.805 ;
        RECT 0.000 933.585 208.285 934.425 ;
        RECT 0.000 931.205 208.565 933.585 ;
        RECT 0.000 930.365 208.285 931.205 ;
        RECT 0.000 928.445 208.565 930.365 ;
        RECT 0.000 927.605 208.285 928.445 ;
        RECT 0.000 925.225 208.565 927.605 ;
        RECT 0.000 924.385 208.285 925.225 ;
      LAYER met2 ;
        RECT 208.565 924.875 210.965 924.945 ;
        RECT 211.300 924.875 211.440 1137.910 ;
        RECT 212.680 1000.570 212.820 1192.390 ;
        RECT 213.140 1158.710 213.280 1369.530 ;
        RECT 3374.260 1188.630 3374.400 1411.350 ;
        RECT 3374.720 1222.630 3374.860 1447.390 ;
        RECT 3375.180 1443.290 3375.320 1448.930 ;
        RECT 3375.640 1447.710 3375.780 1469.750 ;
      LAYER met2 ;
        RECT 3379.435 1468.835 3588.000 1470.755 ;
        RECT 3379.715 1467.995 3588.000 1468.835 ;
      LAYER met2 ;
        RECT 3376.960 1466.090 3377.220 1466.410 ;
        RECT 3377.020 1465.335 3377.160 1466.090 ;
      LAYER met2 ;
        RECT 3379.435 1465.615 3588.000 1467.995 ;
      LAYER met2 ;
        RECT 3377.020 1465.060 3379.435 1465.335 ;
        RECT 3377.035 1465.055 3379.435 1465.060 ;
      LAYER met2 ;
        RECT 3379.715 1464.775 3588.000 1465.615 ;
        RECT 3379.435 1462.395 3588.000 1464.775 ;
        RECT 3379.715 1461.555 3588.000 1462.395 ;
        RECT 3379.435 1459.635 3588.000 1461.555 ;
        RECT 3379.715 1458.795 3588.000 1459.635 ;
        RECT 3379.435 1456.415 3588.000 1458.795 ;
        RECT 3379.715 1455.575 3588.000 1456.415 ;
        RECT 3379.435 1453.195 3588.000 1455.575 ;
        RECT 3379.715 1452.355 3588.000 1453.195 ;
        RECT 3379.435 1450.435 3588.000 1452.355 ;
      LAYER met2 ;
        RECT 3377.035 1450.100 3379.435 1450.155 ;
        RECT 3377.020 1449.875 3379.435 1450.100 ;
        RECT 3377.020 1447.710 3377.160 1449.875 ;
      LAYER met2 ;
        RECT 3379.715 1449.595 3588.000 1450.435 ;
      LAYER met2 ;
        RECT 3375.580 1447.390 3375.840 1447.710 ;
        RECT 3376.960 1447.390 3377.220 1447.710 ;
      LAYER met2 ;
        RECT 3379.435 1447.215 3588.000 1449.595 ;
        RECT 3379.715 1446.375 3588.000 1447.215 ;
        RECT 3379.435 1443.995 3588.000 1446.375 ;
      LAYER met2 ;
        RECT 3377.035 1443.645 3379.435 1443.715 ;
        RECT 3376.100 1443.505 3379.435 1443.645 ;
        RECT 3375.120 1442.970 3375.380 1443.290 ;
        RECT 3376.100 1406.230 3376.240 1443.505 ;
        RECT 3377.035 1443.435 3379.435 1443.505 ;
        RECT 3376.500 1442.970 3376.760 1443.290 ;
      LAYER met2 ;
        RECT 3379.715 1443.155 3588.000 1443.995 ;
      LAYER met2 ;
        RECT 3376.040 1405.910 3376.300 1406.230 ;
        RECT 3376.560 1242.770 3376.700 1442.970 ;
      LAYER met2 ;
        RECT 3379.435 1440.775 3588.000 1443.155 ;
        RECT 3379.715 1439.935 3588.000 1440.775 ;
        RECT 3379.435 1438.015 3588.000 1439.935 ;
        RECT 3379.715 1437.175 3588.000 1438.015 ;
        RECT 3379.435 1434.795 3588.000 1437.175 ;
        RECT 3379.715 1433.955 3588.000 1434.795 ;
        RECT 3379.435 1431.575 3588.000 1433.955 ;
        RECT 3379.715 1430.735 3588.000 1431.575 ;
        RECT 3379.435 1428.815 3588.000 1430.735 ;
      LAYER met2 ;
        RECT 3377.035 1428.255 3379.435 1428.535 ;
      LAYER met2 ;
        RECT 3379.715 1427.975 3588.000 1428.815 ;
        RECT 3379.435 1425.595 3588.000 1427.975 ;
        RECT 3379.715 1424.755 3588.000 1425.595 ;
        RECT 3379.435 1422.375 3588.000 1424.755 ;
      LAYER met2 ;
        RECT 3377.035 1421.815 3379.435 1422.095 ;
      LAYER met2 ;
        RECT 3379.715 1421.535 3588.000 1422.375 ;
        RECT 3379.435 1419.615 3588.000 1421.535 ;
      LAYER met2 ;
        RECT 3377.035 1419.055 3379.435 1419.335 ;
      LAYER met2 ;
        RECT 3379.715 1418.775 3588.000 1419.615 ;
        RECT 3379.435 1416.395 3588.000 1418.775 ;
        RECT 3379.715 1415.555 3588.000 1416.395 ;
        RECT 3379.435 1413.175 3588.000 1415.555 ;
      LAYER met2 ;
        RECT 3377.035 1412.700 3379.435 1412.895 ;
        RECT 3377.020 1412.615 3379.435 1412.700 ;
        RECT 3377.020 1411.670 3377.160 1412.615 ;
      LAYER met2 ;
        RECT 3379.715 1412.335 3588.000 1413.175 ;
      LAYER met2 ;
        RECT 3376.960 1411.350 3377.220 1411.670 ;
      LAYER met2 ;
        RECT 3379.435 1410.415 3588.000 1412.335 ;
      LAYER met2 ;
        RECT 3377.035 1409.855 3379.435 1410.135 ;
      LAYER met2 ;
        RECT 3379.715 1409.575 3588.000 1410.415 ;
        RECT 3379.435 1407.195 3588.000 1409.575 ;
        RECT 3379.715 1406.355 3588.000 1407.195 ;
      LAYER met2 ;
        RECT 3376.960 1405.910 3377.220 1406.230 ;
        RECT 3377.020 1403.695 3377.160 1405.910 ;
      LAYER met2 ;
        RECT 3379.435 1403.975 3588.000 1406.355 ;
      LAYER met2 ;
        RECT 3377.020 1403.555 3379.435 1403.695 ;
        RECT 3377.035 1403.415 3379.435 1403.555 ;
      LAYER met2 ;
        RECT 3379.715 1403.135 3588.000 1403.975 ;
        RECT 3379.435 1402.085 3588.000 1403.135 ;
        RECT 3379.435 1255.795 3588.000 1256.790 ;
      LAYER met2 ;
        RECT 3377.035 1255.235 3379.435 1255.515 ;
      LAYER met2 ;
        RECT 3379.715 1254.955 3588.000 1255.795 ;
        RECT 3379.435 1253.035 3588.000 1254.955 ;
        RECT 3379.715 1252.195 3588.000 1253.035 ;
        RECT 3379.435 1249.815 3588.000 1252.195 ;
        RECT 3379.715 1248.975 3588.000 1249.815 ;
        RECT 3379.435 1246.595 3588.000 1248.975 ;
        RECT 3379.715 1245.755 3588.000 1246.595 ;
        RECT 3379.435 1243.835 3588.000 1245.755 ;
        RECT 3379.715 1242.995 3588.000 1243.835 ;
      LAYER met2 ;
        RECT 3376.560 1242.630 3377.160 1242.770 ;
        RECT 3377.020 1240.335 3377.160 1242.630 ;
      LAYER met2 ;
        RECT 3379.435 1240.615 3588.000 1242.995 ;
      LAYER met2 ;
        RECT 3377.020 1240.055 3379.435 1240.335 ;
        RECT 3377.020 1237.590 3377.160 1240.055 ;
      LAYER met2 ;
        RECT 3379.715 1239.775 3588.000 1240.615 ;
      LAYER met2 ;
        RECT 3375.120 1237.270 3375.380 1237.590 ;
        RECT 3376.960 1237.270 3377.220 1237.590 ;
      LAYER met2 ;
        RECT 3379.435 1237.395 3588.000 1239.775 ;
      LAYER met2 ;
        RECT 3374.660 1222.310 3374.920 1222.630 ;
        RECT 3374.200 1188.310 3374.460 1188.630 ;
        RECT 213.080 1158.390 213.340 1158.710 ;
        RECT 212.220 1000.430 212.820 1000.570 ;
        RECT 212.220 976.810 212.360 1000.430 ;
        RECT 212.160 976.490 212.420 976.810 ;
        RECT 208.565 924.735 211.440 924.875 ;
        RECT 208.565 924.665 210.965 924.735 ;
      LAYER met2 ;
        RECT 0.000 922.005 208.565 924.385 ;
        RECT 0.000 921.165 208.285 922.005 ;
        RECT 0.000 919.245 208.565 921.165 ;
        RECT 0.000 918.405 208.285 919.245 ;
        RECT 0.000 916.025 208.565 918.405 ;
        RECT 0.000 915.185 208.285 916.025 ;
        RECT 0.000 912.805 208.565 915.185 ;
        RECT 0.000 911.965 208.285 912.805 ;
        RECT 0.000 910.045 208.565 911.965 ;
        RECT 0.000 909.205 208.285 910.045 ;
      LAYER met2 ;
        RECT 208.565 909.485 210.965 909.765 ;
      LAYER met2 ;
        RECT 0.000 908.210 208.565 909.205 ;
        RECT 4.925 601.390 200.000 625.290 ;
        RECT 4.925 575.395 197.965 601.390 ;
        RECT 198.080 576.895 200.000 578.895 ;
        RECT 4.925 551.495 200.000 575.395 ;
      LAYER met2 ;
        RECT 210.310 565.915 210.590 566.285 ;
      LAYER met2 ;
        RECT 4.925 551.265 197.965 551.495 ;
        RECT 153.765 415.000 158.415 426.140 ;
        RECT 159.640 415.245 163.510 426.195 ;
        RECT 3.570 414.700 197.965 415.000 ;
        RECT 3.570 394.095 198.000 414.700 ;
        RECT 3.570 393.535 197.965 394.095 ;
        RECT 3.570 360.925 198.000 393.535 ;
        RECT 3.570 360.495 197.965 360.925 ;
        RECT 3.570 340.500 198.000 360.495 ;
        RECT 3.570 340.490 197.965 340.500 ;
      LAYER met2 ;
        RECT 210.380 224.390 210.520 565.915 ;
        RECT 210.770 391.155 211.050 391.525 ;
        RECT 210.840 224.730 210.980 391.155 ;
        RECT 210.780 224.410 211.040 224.730 ;
        RECT 210.320 224.070 210.580 224.390 ;
        RECT 211.300 210.790 211.440 924.735 ;
        RECT 212.220 391.525 212.360 976.490 ;
        RECT 213.140 952.270 213.280 1158.390 ;
        RECT 3374.720 1001.290 3374.860 1222.310 ;
        RECT 3375.180 1011.830 3375.320 1237.270 ;
      LAYER met2 ;
        RECT 3379.715 1236.555 3588.000 1237.395 ;
        RECT 3379.435 1234.635 3588.000 1236.555 ;
        RECT 3379.715 1233.795 3588.000 1234.635 ;
        RECT 3379.435 1231.415 3588.000 1233.795 ;
        RECT 3379.715 1230.575 3588.000 1231.415 ;
        RECT 3379.435 1228.195 3588.000 1230.575 ;
        RECT 3379.715 1227.355 3588.000 1228.195 ;
        RECT 3379.435 1225.435 3588.000 1227.355 ;
      LAYER met2 ;
        RECT 3377.035 1225.020 3379.435 1225.155 ;
        RECT 3377.020 1224.875 3379.435 1225.020 ;
        RECT 3377.020 1222.630 3377.160 1224.875 ;
      LAYER met2 ;
        RECT 3379.715 1224.595 3588.000 1225.435 ;
      LAYER met2 ;
        RECT 3376.960 1222.310 3377.220 1222.630 ;
      LAYER met2 ;
        RECT 3379.435 1222.215 3588.000 1224.595 ;
        RECT 3379.715 1221.375 3588.000 1222.215 ;
        RECT 3379.435 1218.995 3588.000 1221.375 ;
      LAYER met2 ;
        RECT 3377.035 1218.645 3379.435 1218.715 ;
        RECT 3376.100 1218.505 3379.435 1218.645 ;
        RECT 3376.100 1181.490 3376.240 1218.505 ;
        RECT 3377.035 1218.435 3379.435 1218.505 ;
      LAYER met2 ;
        RECT 3379.715 1218.155 3588.000 1218.995 ;
        RECT 3379.435 1215.775 3588.000 1218.155 ;
        RECT 3379.715 1214.935 3588.000 1215.775 ;
        RECT 3379.435 1213.015 3588.000 1214.935 ;
        RECT 3379.715 1212.175 3588.000 1213.015 ;
        RECT 3379.435 1209.795 3588.000 1212.175 ;
        RECT 3379.715 1208.955 3588.000 1209.795 ;
        RECT 3379.435 1206.575 3588.000 1208.955 ;
        RECT 3379.715 1205.735 3588.000 1206.575 ;
        RECT 3379.435 1203.815 3588.000 1205.735 ;
      LAYER met2 ;
        RECT 3377.035 1203.255 3379.435 1203.535 ;
      LAYER met2 ;
        RECT 3379.715 1202.975 3588.000 1203.815 ;
        RECT 3379.435 1200.595 3588.000 1202.975 ;
        RECT 3379.715 1199.755 3588.000 1200.595 ;
        RECT 3379.435 1197.375 3588.000 1199.755 ;
      LAYER met2 ;
        RECT 3377.035 1196.815 3379.435 1197.095 ;
      LAYER met2 ;
        RECT 3379.715 1196.535 3588.000 1197.375 ;
        RECT 3379.435 1194.615 3588.000 1196.535 ;
      LAYER met2 ;
        RECT 3377.035 1194.055 3379.435 1194.335 ;
      LAYER met2 ;
        RECT 3379.715 1193.775 3588.000 1194.615 ;
        RECT 3379.435 1191.395 3588.000 1193.775 ;
        RECT 3379.715 1190.555 3588.000 1191.395 ;
      LAYER met2 ;
        RECT 3376.960 1188.310 3377.220 1188.630 ;
        RECT 3377.020 1187.895 3377.160 1188.310 ;
      LAYER met2 ;
        RECT 3379.435 1188.175 3588.000 1190.555 ;
      LAYER met2 ;
        RECT 3377.020 1187.615 3379.435 1187.895 ;
        RECT 3377.020 1185.650 3377.160 1187.615 ;
      LAYER met2 ;
        RECT 3379.715 1187.335 3588.000 1188.175 ;
      LAYER met2 ;
        RECT 3376.560 1185.510 3377.160 1185.650 ;
        RECT 3376.040 1181.170 3376.300 1181.490 ;
        RECT 3376.560 1028.170 3376.700 1185.510 ;
      LAYER met2 ;
        RECT 3379.435 1185.415 3588.000 1187.335 ;
      LAYER met2 ;
        RECT 3377.035 1184.855 3379.435 1185.135 ;
      LAYER met2 ;
        RECT 3379.715 1184.575 3588.000 1185.415 ;
        RECT 3379.435 1182.195 3588.000 1184.575 ;
      LAYER met2 ;
        RECT 3376.960 1181.170 3377.220 1181.490 ;
      LAYER met2 ;
        RECT 3379.715 1181.355 3588.000 1182.195 ;
      LAYER met2 ;
        RECT 3377.020 1178.695 3377.160 1181.170 ;
      LAYER met2 ;
        RECT 3379.435 1178.975 3588.000 1181.355 ;
      LAYER met2 ;
        RECT 3377.020 1178.555 3379.435 1178.695 ;
        RECT 3377.035 1178.415 3379.435 1178.555 ;
      LAYER met2 ;
        RECT 3379.715 1178.135 3588.000 1178.975 ;
        RECT 3379.435 1177.085 3588.000 1178.135 ;
        RECT 3379.435 1029.795 3588.000 1030.790 ;
      LAYER met2 ;
        RECT 3377.035 1029.235 3379.435 1029.515 ;
      LAYER met2 ;
        RECT 3379.715 1028.955 3588.000 1029.795 ;
      LAYER met2 ;
        RECT 3376.100 1028.030 3376.700 1028.170 ;
        RECT 3375.120 1011.510 3375.380 1011.830 ;
        RECT 3374.660 1000.970 3374.920 1001.290 ;
        RECT 213.540 983.630 213.800 983.950 ;
        RECT 212.680 952.130 213.280 952.270 ;
        RECT 212.680 938.050 212.820 952.130 ;
        RECT 213.600 949.270 213.740 983.630 ;
        RECT 213.540 948.950 213.800 949.270 ;
        RECT 212.620 937.730 212.880 938.050 ;
        RECT 212.680 566.285 212.820 937.730 ;
        RECT 3374.200 786.430 3374.460 786.750 ;
        RECT 212.610 565.915 212.890 566.285 ;
        RECT 3374.260 562.690 3374.400 786.430 ;
        RECT 3374.720 776.210 3374.860 1000.970 ;
        RECT 3375.180 786.750 3375.320 1011.510 ;
        RECT 3376.100 996.530 3376.240 1028.030 ;
      LAYER met2 ;
        RECT 3379.435 1027.035 3588.000 1028.955 ;
        RECT 3379.715 1026.195 3588.000 1027.035 ;
        RECT 3379.435 1023.815 3588.000 1026.195 ;
        RECT 3379.715 1022.975 3588.000 1023.815 ;
        RECT 3379.435 1020.595 3588.000 1022.975 ;
        RECT 3379.715 1019.755 3588.000 1020.595 ;
        RECT 3379.435 1017.835 3588.000 1019.755 ;
        RECT 3379.715 1016.995 3588.000 1017.835 ;
        RECT 3379.435 1014.615 3588.000 1016.995 ;
      LAYER met2 ;
        RECT 3377.035 1014.220 3379.435 1014.335 ;
        RECT 3377.020 1014.055 3379.435 1014.220 ;
        RECT 3377.020 1011.830 3377.160 1014.055 ;
      LAYER met2 ;
        RECT 3379.715 1013.775 3588.000 1014.615 ;
      LAYER met2 ;
        RECT 3376.960 1011.510 3377.220 1011.830 ;
      LAYER met2 ;
        RECT 3379.435 1011.395 3588.000 1013.775 ;
        RECT 3379.715 1010.555 3588.000 1011.395 ;
        RECT 3379.435 1008.635 3588.000 1010.555 ;
        RECT 3379.715 1007.795 3588.000 1008.635 ;
        RECT 3379.435 1005.415 3588.000 1007.795 ;
        RECT 3379.715 1004.575 3588.000 1005.415 ;
        RECT 3379.435 1002.195 3588.000 1004.575 ;
        RECT 3379.715 1001.355 3588.000 1002.195 ;
      LAYER met2 ;
        RECT 3376.960 1000.970 3377.220 1001.290 ;
        RECT 3377.020 999.155 3377.160 1000.970 ;
      LAYER met2 ;
        RECT 3379.435 999.435 3588.000 1001.355 ;
      LAYER met2 ;
        RECT 3377.020 999.015 3379.435 999.155 ;
        RECT 3377.035 998.875 3379.435 999.015 ;
      LAYER met2 ;
        RECT 3379.715 998.595 3588.000 999.435 ;
      LAYER met2 ;
        RECT 3376.040 996.210 3376.300 996.530 ;
      LAYER met2 ;
        RECT 3379.435 996.215 3588.000 998.595 ;
      LAYER met2 ;
        RECT 3376.040 995.190 3376.300 995.510 ;
      LAYER met2 ;
        RECT 3379.715 995.375 3588.000 996.215 ;
      LAYER met2 ;
        RECT 3376.100 959.810 3376.240 995.190 ;
        RECT 3376.560 993.070 3377.160 993.210 ;
        RECT 3376.040 959.490 3376.300 959.810 ;
        RECT 3376.100 855.670 3376.240 959.490 ;
        RECT 3376.560 952.625 3376.700 993.070 ;
        RECT 3377.020 992.715 3377.160 993.070 ;
      LAYER met2 ;
        RECT 3379.435 992.995 3588.000 995.375 ;
      LAYER met2 ;
        RECT 3377.020 992.460 3379.435 992.715 ;
        RECT 3377.035 992.435 3379.435 992.460 ;
      LAYER met2 ;
        RECT 3379.715 992.155 3588.000 992.995 ;
        RECT 3379.435 989.775 3588.000 992.155 ;
        RECT 3379.715 988.935 3588.000 989.775 ;
        RECT 3379.435 987.015 3588.000 988.935 ;
        RECT 3379.715 986.175 3588.000 987.015 ;
        RECT 3379.435 983.795 3588.000 986.175 ;
        RECT 3379.715 982.955 3588.000 983.795 ;
        RECT 3379.435 980.575 3588.000 982.955 ;
        RECT 3379.715 979.735 3588.000 980.575 ;
        RECT 3379.435 977.815 3588.000 979.735 ;
      LAYER met2 ;
        RECT 3377.035 977.255 3379.435 977.535 ;
      LAYER met2 ;
        RECT 3379.715 976.975 3588.000 977.815 ;
        RECT 3379.435 974.595 3588.000 976.975 ;
        RECT 3379.715 973.755 3588.000 974.595 ;
        RECT 3379.435 971.375 3588.000 973.755 ;
      LAYER met2 ;
        RECT 3377.035 970.815 3379.435 971.095 ;
      LAYER met2 ;
        RECT 3379.715 970.535 3588.000 971.375 ;
        RECT 3379.435 968.615 3588.000 970.535 ;
      LAYER met2 ;
        RECT 3377.035 968.055 3379.435 968.335 ;
      LAYER met2 ;
        RECT 3379.715 967.775 3588.000 968.615 ;
        RECT 3379.435 965.395 3588.000 967.775 ;
        RECT 3379.715 964.555 3588.000 965.395 ;
        RECT 3379.435 962.175 3588.000 964.555 ;
      LAYER met2 ;
        RECT 3377.035 961.860 3379.435 961.895 ;
        RECT 3377.020 961.615 3379.435 961.860 ;
        RECT 3377.020 959.810 3377.160 961.615 ;
      LAYER met2 ;
        RECT 3379.715 961.335 3588.000 962.175 ;
      LAYER met2 ;
        RECT 3376.960 959.490 3377.220 959.810 ;
      LAYER met2 ;
        RECT 3379.435 959.415 3588.000 961.335 ;
      LAYER met2 ;
        RECT 3377.035 958.855 3379.435 959.135 ;
      LAYER met2 ;
        RECT 3379.715 958.575 3588.000 959.415 ;
        RECT 3379.435 956.195 3588.000 958.575 ;
        RECT 3379.715 955.355 3588.000 956.195 ;
        RECT 3379.435 952.975 3588.000 955.355 ;
      LAYER met2 ;
        RECT 3377.035 952.625 3379.435 952.695 ;
        RECT 3376.560 952.485 3379.435 952.625 ;
        RECT 3377.035 952.415 3379.435 952.485 ;
      LAYER met2 ;
        RECT 3379.715 952.135 3588.000 952.975 ;
        RECT 3379.435 951.085 3588.000 952.135 ;
      LAYER met2 ;
        RECT 3376.100 855.530 3376.700 855.670 ;
        RECT 3376.560 793.890 3376.700 855.530 ;
      LAYER met2 ;
        RECT 3379.435 804.795 3588.000 805.790 ;
      LAYER met2 ;
        RECT 3377.035 804.235 3379.435 804.515 ;
      LAYER met2 ;
        RECT 3379.715 803.955 3588.000 804.795 ;
        RECT 3379.435 802.035 3588.000 803.955 ;
        RECT 3379.715 801.195 3588.000 802.035 ;
        RECT 3379.435 798.815 3588.000 801.195 ;
        RECT 3379.715 797.975 3588.000 798.815 ;
        RECT 3379.435 795.595 3588.000 797.975 ;
        RECT 3379.715 794.755 3588.000 795.595 ;
      LAYER met2 ;
        RECT 3376.500 793.570 3376.760 793.890 ;
        RECT 3375.580 792.550 3375.840 792.870 ;
      LAYER met2 ;
        RECT 3379.435 792.835 3588.000 794.755 ;
      LAYER met2 ;
        RECT 3375.120 786.430 3375.380 786.750 ;
        RECT 3375.640 783.090 3375.780 792.550 ;
      LAYER met2 ;
        RECT 3379.715 791.995 3588.000 792.835 ;
        RECT 3379.435 789.615 3588.000 791.995 ;
      LAYER met2 ;
        RECT 3377.035 789.140 3379.435 789.335 ;
        RECT 3377.020 789.055 3379.435 789.140 ;
        RECT 3377.020 786.750 3377.160 789.055 ;
      LAYER met2 ;
        RECT 3379.715 788.775 3588.000 789.615 ;
      LAYER met2 ;
        RECT 3376.960 786.430 3377.220 786.750 ;
      LAYER met2 ;
        RECT 3379.435 786.395 3588.000 788.775 ;
        RECT 3379.715 785.555 3588.000 786.395 ;
        RECT 3379.435 783.635 3588.000 785.555 ;
      LAYER met2 ;
        RECT 3375.180 782.950 3375.780 783.090 ;
        RECT 3374.660 775.890 3374.920 776.210 ;
        RECT 3374.200 562.370 3374.460 562.690 ;
        RECT 212.150 391.155 212.430 391.525 ;
        RECT 738.400 224.410 738.660 224.730 ;
        RECT 2618.880 224.410 2619.140 224.730 ;
        RECT 444.000 222.030 444.260 222.350 ;
        RECT 211.240 210.470 211.500 210.790 ;
      LAYER met2 ;
        RECT 394.710 197.965 418.610 200.000 ;
        RECT 441.105 198.080 443.105 200.000 ;
      LAYER met2 ;
        RECT 444.060 199.765 444.200 222.030 ;
        RECT 738.460 221.330 738.600 224.410 ;
        RECT 979.900 224.070 980.160 224.390 ;
        RECT 2580.700 224.070 2580.960 224.390 ;
        RECT 942.640 221.690 942.900 222.010 ;
        RECT 964.260 221.690 964.520 222.010 ;
        RECT 942.700 221.330 942.840 221.690 ;
        RECT 738.400 221.010 738.660 221.330 ;
        RECT 942.640 221.010 942.900 221.330 ;
        RECT 704.820 210.470 705.080 210.790 ;
        RECT 704.880 201.010 705.020 210.470 ;
        RECT 715.400 207.070 715.660 207.390 ;
        RECT 715.460 201.805 715.600 207.070 ;
        RECT 723.220 206.730 723.480 207.050 ;
        RECT 715.390 201.435 715.670 201.805 ;
        RECT 704.880 200.870 705.180 201.010 ;
        RECT 705.040 200.590 705.180 200.870 ;
        RECT 715.460 200.590 715.600 201.435 ;
        RECT 704.980 200.270 705.240 200.590 ;
        RECT 715.400 200.270 715.660 200.590 ;
        RECT 705.040 200.000 705.180 200.270 ;
        RECT 715.460 200.000 715.600 200.270 ;
        RECT 723.280 200.000 723.420 206.730 ;
        RECT 443.990 199.395 444.270 199.765 ;
      LAYER met2 ;
        RECT 444.605 197.965 468.505 200.000 ;
        RECT 663.085 199.390 664.485 200.000 ;
      LAYER met2 ;
        RECT 664.765 199.670 665.785 200.000 ;
      LAYER met2 ;
        RECT 666.065 199.390 704.700 200.000 ;
        RECT 663.085 199.080 704.700 199.390 ;
      LAYER met2 ;
        RECT 704.980 199.360 705.240 200.000 ;
      LAYER met2 ;
        RECT 705.520 199.390 706.565 200.000 ;
      LAYER met2 ;
        RECT 706.845 199.670 707.495 200.000 ;
      LAYER met2 ;
        RECT 707.775 199.390 708.055 200.000 ;
      LAYER met2 ;
        RECT 708.335 199.670 709.065 200.000 ;
      LAYER met2 ;
        RECT 709.345 199.390 709.490 200.000 ;
      LAYER met2 ;
        RECT 709.770 199.670 710.420 200.000 ;
      LAYER met2 ;
        RECT 710.700 199.390 715.060 200.000 ;
        RECT 705.520 199.080 715.060 199.390 ;
        RECT 394.710 4.925 468.735 197.965 ;
        RECT 663.085 196.020 715.060 199.080 ;
        RECT 663.085 195.735 714.775 196.020 ;
      LAYER met2 ;
        RECT 715.340 195.755 715.640 200.000 ;
      LAYER met2 ;
        RECT 715.920 198.310 716.495 200.000 ;
      LAYER met2 ;
        RECT 716.775 198.590 717.925 200.000 ;
      LAYER met2 ;
        RECT 718.205 199.155 718.810 200.000 ;
      LAYER met2 ;
        RECT 719.090 199.435 720.755 200.000 ;
      LAYER met2 ;
        RECT 721.035 199.155 722.585 200.000 ;
        RECT 718.205 198.735 722.585 199.155 ;
      LAYER met2 ;
        RECT 722.865 199.015 723.445 200.000 ;
      LAYER met2 ;
        RECT 723.725 198.735 725.175 200.000 ;
        RECT 718.205 198.310 725.175 198.735 ;
        RECT 715.920 198.250 725.175 198.310 ;
        RECT 725.995 199.390 728.825 200.000 ;
      LAYER met2 ;
        RECT 729.105 199.670 729.575 200.000 ;
      LAYER met2 ;
        RECT 729.855 199.390 737.660 200.000 ;
      LAYER met2 ;
        RECT 738.460 199.765 738.600 221.010 ;
        RECT 933.440 220.670 933.700 220.990 ;
        RECT 933.500 210.965 933.640 220.670 ;
        RECT 942.700 210.965 942.840 221.010 ;
        RECT 964.320 210.965 964.460 221.690 ;
        RECT 979.960 221.330 980.100 224.070 ;
        RECT 2298.260 223.730 2298.520 224.050 ;
        RECT 2338.280 223.730 2338.540 224.050 ;
        RECT 2076.540 223.390 2076.800 223.710 ;
        RECT 1476.240 222.710 1476.500 223.030 ;
        RECT 1516.260 222.710 1516.520 223.030 ;
        RECT 1750.400 222.710 1750.660 223.030 ;
        RECT 1790.420 222.710 1790.680 223.030 ;
        RECT 1802.840 222.710 1803.100 223.030 ;
        RECT 2033.760 222.710 2034.020 223.030 ;
        RECT 995.080 222.030 995.340 222.350 ;
        RECT 1004.280 222.030 1004.540 222.350 ;
        RECT 1206.680 222.030 1206.940 222.350 ;
        RECT 979.900 221.010 980.160 221.330 ;
        RECT 973.460 220.670 973.720 220.990 ;
        RECT 973.520 210.965 973.660 220.670 ;
        RECT 979.960 210.965 980.100 221.010 ;
        RECT 995.140 210.965 995.280 222.030 ;
        RECT 1004.340 210.965 1004.480 222.030 ;
        RECT 1007.500 221.690 1007.760 222.010 ;
        RECT 1007.560 210.965 1007.700 221.690 ;
        RECT 933.415 208.565 933.695 210.965 ;
        RECT 939.855 208.565 940.135 210.965 ;
        RECT 942.615 208.565 942.895 210.965 ;
        RECT 945.835 209.170 946.115 210.965 ;
        RECT 945.835 209.090 946.520 209.170 ;
        RECT 945.835 209.030 946.580 209.090 ;
        RECT 945.835 208.565 946.115 209.030 ;
        RECT 946.320 208.770 946.580 209.030 ;
        RECT 949.055 208.565 949.335 210.965 ;
        RECT 951.815 208.565 952.095 210.965 ;
        RECT 955.035 209.170 955.315 210.965 ;
        RECT 955.035 209.090 955.720 209.170 ;
        RECT 955.035 209.030 955.780 209.090 ;
        RECT 955.035 208.565 955.315 209.030 ;
        RECT 955.520 208.770 955.780 209.030 ;
        RECT 958.255 208.565 958.535 210.965 ;
        RECT 961.015 209.170 961.295 210.965 ;
        RECT 961.015 209.090 961.700 209.170 ;
        RECT 961.015 209.030 961.760 209.090 ;
        RECT 961.015 208.565 961.295 209.030 ;
        RECT 961.500 208.770 961.760 209.030 ;
        RECT 964.235 208.565 964.515 210.965 ;
        RECT 967.455 209.170 967.735 210.965 ;
        RECT 967.455 209.090 968.140 209.170 ;
        RECT 967.455 209.030 968.200 209.090 ;
        RECT 967.455 208.565 967.735 209.030 ;
        RECT 967.940 208.770 968.200 209.030 ;
        RECT 973.435 208.565 973.715 210.965 ;
        RECT 979.875 208.565 980.155 210.965 ;
        RECT 982.635 209.170 982.915 210.965 ;
        RECT 985.855 209.170 986.135 210.965 ;
        RECT 989.075 209.170 989.355 210.965 ;
        RECT 991.835 209.170 992.115 210.965 ;
        RECT 992.320 209.450 992.580 209.770 ;
        RECT 992.380 209.170 992.520 209.450 ;
        RECT 982.260 209.090 992.520 209.170 ;
        RECT 982.200 209.030 992.520 209.090 ;
        RECT 982.200 208.770 982.460 209.030 ;
        RECT 982.635 208.565 982.915 209.030 ;
        RECT 985.855 208.565 986.135 209.030 ;
        RECT 989.075 208.565 989.355 209.030 ;
        RECT 991.835 208.565 992.115 209.030 ;
        RECT 995.055 208.565 995.335 210.965 ;
        RECT 1000.600 209.450 1000.860 209.770 ;
        RECT 1000.660 209.170 1000.800 209.450 ;
        RECT 1001.035 209.170 1001.315 210.965 ;
        RECT 1004.255 209.170 1004.535 210.965 ;
        RECT 1000.660 209.030 1004.535 209.170 ;
        RECT 1001.035 208.565 1001.315 209.030 ;
        RECT 1004.255 208.565 1004.535 209.030 ;
        RECT 1007.475 208.565 1007.755 210.965 ;
        RECT 1010.235 208.565 1010.515 210.965 ;
      LAYER met2 ;
        RECT 932.085 208.285 933.135 208.565 ;
        RECT 933.975 208.285 936.355 208.565 ;
        RECT 937.195 208.285 939.575 208.565 ;
        RECT 940.415 208.285 942.335 208.565 ;
        RECT 943.175 208.285 945.555 208.565 ;
        RECT 946.395 208.285 948.775 208.565 ;
        RECT 949.615 208.285 951.535 208.565 ;
        RECT 952.375 208.285 954.755 208.565 ;
        RECT 955.595 208.285 957.975 208.565 ;
        RECT 958.815 208.285 960.735 208.565 ;
        RECT 961.575 208.285 963.955 208.565 ;
        RECT 964.795 208.285 967.175 208.565 ;
        RECT 968.015 208.285 969.935 208.565 ;
        RECT 970.775 208.285 973.155 208.565 ;
        RECT 973.995 208.285 976.375 208.565 ;
        RECT 977.215 208.285 979.595 208.565 ;
        RECT 980.435 208.285 982.355 208.565 ;
        RECT 983.195 208.285 985.575 208.565 ;
        RECT 986.415 208.285 988.795 208.565 ;
        RECT 989.635 208.285 991.555 208.565 ;
        RECT 992.395 208.285 994.775 208.565 ;
        RECT 995.615 208.285 997.995 208.565 ;
        RECT 998.835 208.285 1000.755 208.565 ;
        RECT 1001.595 208.285 1003.975 208.565 ;
        RECT 1004.815 208.285 1007.195 208.565 ;
        RECT 1008.035 208.285 1009.955 208.565 ;
        RECT 1010.795 208.285 1011.790 208.565 ;
      LAYER met2 ;
        RECT 738.390 199.395 738.670 199.765 ;
      LAYER met2 ;
        RECT 725.995 198.250 737.660 199.390 ;
        RECT 715.920 196.845 737.660 198.250 ;
        RECT 715.920 196.485 722.475 196.845 ;
        RECT 727.600 196.705 737.660 196.845 ;
        RECT 715.920 196.215 722.205 196.485 ;
      LAYER met2 ;
        RECT 722.755 196.425 727.320 196.565 ;
        RECT 722.755 196.355 727.650 196.425 ;
      LAYER met2 ;
        RECT 727.930 196.375 737.660 196.705 ;
      LAYER met2 ;
        RECT 722.755 196.305 727.180 196.355 ;
      LAYER met2 ;
        RECT 715.920 196.035 721.835 196.215 ;
      LAYER met2 ;
        RECT 722.755 196.205 723.115 196.305 ;
        RECT 723.125 196.205 723.225 196.305 ;
        RECT 727.070 196.235 727.305 196.305 ;
        RECT 727.320 196.235 727.650 196.355 ;
      LAYER met2 ;
        RECT 716.220 195.845 721.835 196.035 ;
      LAYER met2 ;
        RECT 722.485 196.165 722.755 196.205 ;
        RECT 722.855 196.165 723.125 196.205 ;
        RECT 722.485 196.025 723.125 196.165 ;
        RECT 727.070 196.095 727.650 196.235 ;
        RECT 727.070 196.070 727.305 196.095 ;
        RECT 722.485 195.935 722.755 196.025 ;
        RECT 722.855 195.935 723.125 196.025 ;
        RECT 715.340 195.740 715.940 195.755 ;
      LAYER met2 ;
        RECT 663.085 195.380 708.600 195.735 ;
      LAYER met2 ;
        RECT 715.055 195.455 715.940 195.740 ;
      LAYER met2 ;
        RECT 716.220 195.735 721.725 195.845 ;
      LAYER met2 ;
        RECT 722.115 195.565 722.855 195.935 ;
      LAYER met2 ;
        RECT 723.505 195.925 726.790 196.025 ;
        RECT 723.405 195.790 726.790 195.925 ;
      LAYER met2 ;
        RECT 727.305 195.955 727.625 196.070 ;
        RECT 727.650 195.955 727.995 196.095 ;
      LAYER met2 ;
        RECT 728.275 196.030 737.660 196.375 ;
      LAYER met2 ;
        RECT 727.305 195.815 727.995 195.955 ;
      LAYER met2 ;
        RECT 723.405 195.655 727.025 195.790 ;
      LAYER met2 ;
        RECT 727.305 195.750 727.625 195.815 ;
        RECT 727.650 195.750 727.995 195.815 ;
        RECT 722.005 195.455 722.485 195.565 ;
      LAYER met2 ;
        RECT 663.085 195.050 708.270 195.380 ;
      LAYER met2 ;
        RECT 708.880 195.315 722.485 195.455 ;
        RECT 708.880 195.245 709.235 195.315 ;
        RECT 715.340 195.245 715.640 195.315 ;
        RECT 722.115 195.245 722.485 195.315 ;
      LAYER met2 ;
        RECT 723.135 195.470 727.025 195.655 ;
      LAYER met2 ;
        RECT 727.625 195.675 727.955 195.750 ;
        RECT 727.995 195.675 728.265 195.750 ;
      LAYER met2 ;
        RECT 723.135 195.285 727.345 195.470 ;
      LAYER met2 ;
        RECT 727.625 195.425 728.265 195.675 ;
        RECT 727.625 195.420 727.955 195.425 ;
        RECT 708.880 195.195 722.485 195.245 ;
        RECT 708.880 195.100 709.235 195.195 ;
        RECT 709.250 195.100 709.345 195.195 ;
      LAYER met2 ;
        RECT 722.765 195.140 727.345 195.285 ;
      LAYER met2 ;
        RECT 708.550 195.055 708.880 195.100 ;
        RECT 708.920 195.055 709.250 195.100 ;
      LAYER met2 ;
        RECT 663.085 189.305 708.140 195.050 ;
      LAYER met2 ;
        RECT 708.550 194.845 709.250 195.055 ;
      LAYER met2 ;
        RECT 722.765 194.915 727.725 195.140 ;
      LAYER met2 ;
        RECT 708.550 194.770 708.880 194.845 ;
        RECT 708.920 194.770 709.250 194.845 ;
      LAYER met2 ;
        RECT 709.625 194.820 727.725 194.915 ;
      LAYER met2 ;
        RECT 708.420 194.640 708.550 194.770 ;
        RECT 708.680 194.640 708.920 194.770 ;
        RECT 708.420 194.530 708.920 194.640 ;
      LAYER met2 ;
        RECT 663.085 189.115 707.950 189.305 ;
        RECT 663.085 184.635 707.690 189.115 ;
      LAYER met2 ;
        RECT 708.420 189.025 708.680 194.530 ;
      LAYER met2 ;
        RECT 709.530 194.490 727.725 194.820 ;
        RECT 709.200 194.250 727.725 194.490 ;
      LAYER met2 ;
        RECT 708.230 188.915 708.680 189.025 ;
        RECT 708.230 188.835 708.420 188.915 ;
        RECT 708.600 188.835 708.680 188.915 ;
      LAYER met2 ;
        RECT 708.960 191.420 727.725 194.250 ;
        RECT 708.960 191.080 727.385 191.420 ;
      LAYER met2 ;
        RECT 728.005 191.140 728.265 195.425 ;
      LAYER met2 ;
        RECT 708.960 190.880 727.185 191.080 ;
      LAYER met2 ;
        RECT 727.665 190.890 728.265 191.140 ;
      LAYER met2 ;
        RECT 708.960 190.550 726.855 190.880 ;
      LAYER met2 ;
        RECT 727.665 190.800 728.005 190.890 ;
        RECT 728.035 190.800 728.265 190.890 ;
        RECT 727.465 190.750 727.665 190.800 ;
        RECT 727.835 190.750 728.035 190.800 ;
        RECT 727.465 190.680 728.035 190.750 ;
        RECT 727.465 190.600 727.665 190.680 ;
        RECT 727.835 190.600 728.035 190.680 ;
        RECT 707.970 188.465 708.600 188.835 ;
      LAYER met2 ;
        RECT 708.960 188.555 726.595 190.550 ;
      LAYER met2 ;
        RECT 727.135 190.540 727.465 190.600 ;
        RECT 727.505 190.540 727.835 190.600 ;
        RECT 727.135 190.400 727.835 190.540 ;
      LAYER met2 ;
        RECT 728.545 190.520 737.660 196.030 ;
      LAYER met2 ;
        RECT 727.135 190.270 727.465 190.400 ;
        RECT 727.505 190.270 727.835 190.400 ;
      LAYER met2 ;
        RECT 728.315 190.320 737.660 190.520 ;
        RECT 663.085 184.300 707.355 184.635 ;
      LAYER met2 ;
        RECT 707.970 184.355 708.230 188.465 ;
      LAYER met2 ;
        RECT 708.880 188.185 726.595 188.555 ;
        RECT 663.085 179.225 707.095 184.300 ;
      LAYER met2 ;
        RECT 707.635 184.105 708.230 184.355 ;
        RECT 707.635 184.020 707.970 184.105 ;
        RECT 708.005 184.020 708.230 184.105 ;
        RECT 707.375 183.650 708.005 184.020 ;
      LAYER met2 ;
        RECT 708.510 183.740 726.595 188.185 ;
      LAYER met2 ;
        RECT 707.375 179.505 707.635 183.650 ;
      LAYER met2 ;
        RECT 708.285 183.370 726.595 183.740 ;
        RECT 707.915 179.225 726.595 183.370 ;
        RECT 663.085 172.420 726.595 179.225 ;
      LAYER met2 ;
        RECT 726.875 189.900 727.505 190.270 ;
      LAYER met2 ;
        RECT 728.115 189.990 737.660 190.320 ;
      LAYER met2 ;
        RECT 726.875 173.390 727.135 189.900 ;
      LAYER met2 ;
        RECT 727.785 189.620 737.660 189.990 ;
        RECT 727.415 173.670 737.660 189.620 ;
      LAYER met2 ;
        RECT 726.875 172.700 727.350 173.390 ;
      LAYER met2 ;
        RECT 663.085 172.345 726.810 172.420 ;
        RECT 663.085 169.195 726.595 172.345 ;
      LAYER met2 ;
        RECT 727.090 172.065 727.350 172.700 ;
        RECT 726.875 171.855 727.350 172.065 ;
        RECT 726.875 171.850 727.090 171.855 ;
        RECT 726.875 171.375 727.350 171.850 ;
      LAYER met2 ;
        RECT 663.085 169.050 726.450 169.195 ;
        RECT 663.085 168.825 726.225 169.050 ;
      LAYER met2 ;
        RECT 726.875 168.915 727.135 171.375 ;
      LAYER met2 ;
        RECT 727.630 171.095 737.660 173.670 ;
        RECT 663.085 164.260 726.200 168.825 ;
      LAYER met2 ;
        RECT 726.730 168.770 727.135 168.915 ;
        RECT 726.505 168.735 726.730 168.770 ;
        RECT 726.875 168.735 727.135 168.770 ;
        RECT 726.505 168.665 727.135 168.735 ;
        RECT 726.505 168.545 726.730 168.665 ;
        RECT 726.875 168.545 727.135 168.665 ;
        RECT 726.480 168.520 726.505 168.545 ;
        RECT 726.740 168.520 726.875 168.545 ;
        RECT 726.480 168.410 726.875 168.520 ;
      LAYER met2 ;
        RECT 663.085 163.440 725.570 164.260 ;
      LAYER met2 ;
        RECT 726.480 163.980 726.740 168.410 ;
      LAYER met2 ;
        RECT 727.415 168.265 737.660 171.095 ;
        RECT 727.155 168.130 737.660 168.265 ;
      LAYER met2 ;
        RECT 725.850 163.720 726.740 163.980 ;
      LAYER met2 ;
        RECT 727.020 163.440 737.660 168.130 ;
        RECT 663.085 0.790 737.660 163.440 ;
        RECT 932.085 0.000 1011.790 208.285 ;
      LAYER met2 ;
        RECT 1198.390 206.875 1198.670 207.245 ;
        RECT 1198.400 206.730 1198.660 206.875 ;
        RECT 1206.740 199.085 1206.880 222.030 ;
        RECT 1476.300 210.965 1476.440 222.710 ;
        RECT 1488.660 222.030 1488.920 222.350 ;
        RECT 1503.840 222.030 1504.100 222.350 ;
        RECT 1485.440 221.690 1485.700 222.010 ;
        RECT 1485.500 210.965 1485.640 221.690 ;
        RECT 1488.720 210.965 1488.860 222.030 ;
        RECT 1497.860 221.690 1498.120 222.010 ;
        RECT 1497.920 210.965 1498.060 221.690 ;
        RECT 1503.900 210.965 1504.040 222.030 ;
        RECT 1516.320 210.965 1516.460 222.710 ;
        RECT 1537.880 222.370 1538.140 222.690 ;
        RECT 1525.460 222.030 1525.720 222.350 ;
        RECT 1522.700 221.010 1522.960 221.330 ;
        RECT 1522.760 210.965 1522.900 221.010 ;
        RECT 1525.520 210.965 1525.660 222.030 ;
        RECT 1528.680 221.690 1528.940 222.010 ;
        RECT 1528.740 210.965 1528.880 221.690 ;
        RECT 1537.940 210.965 1538.080 222.370 ;
        RECT 1547.080 222.030 1547.340 222.350 ;
        RECT 1547.140 210.965 1547.280 222.030 ;
        RECT 1750.460 210.965 1750.600 222.710 ;
        RECT 1762.820 222.030 1763.080 222.350 ;
        RECT 1778.000 222.030 1778.260 222.350 ;
        RECT 1759.600 221.690 1759.860 222.010 ;
        RECT 1759.660 210.965 1759.800 221.690 ;
        RECT 1762.880 210.965 1763.020 222.030 ;
        RECT 1772.020 221.690 1772.280 222.010 ;
        RECT 1772.080 210.965 1772.220 221.690 ;
        RECT 1778.060 210.965 1778.200 222.030 ;
        RECT 1790.480 210.965 1790.620 222.710 ;
        RECT 1799.620 222.030 1799.880 222.350 ;
        RECT 1796.860 221.010 1797.120 221.330 ;
        RECT 1796.920 210.965 1797.060 221.010 ;
        RECT 1799.680 210.965 1799.820 222.030 ;
        RECT 1802.900 222.010 1803.040 222.710 ;
        RECT 1812.040 222.370 1812.300 222.690 ;
        RECT 1802.840 221.690 1803.100 222.010 ;
        RECT 1802.900 210.965 1803.040 221.690 ;
        RECT 1812.100 210.965 1812.240 222.370 ;
        RECT 1821.240 222.030 1821.500 222.350 ;
        RECT 1821.300 210.965 1821.440 222.030 ;
        RECT 2024.560 221.690 2024.820 222.010 ;
        RECT 2024.620 210.965 2024.760 221.690 ;
        RECT 2033.820 210.965 2033.960 222.710 ;
        RECT 2036.980 222.030 2037.240 222.350 ;
        RECT 2052.160 222.030 2052.420 222.350 ;
        RECT 2037.040 210.965 2037.180 222.030 ;
        RECT 2052.220 210.965 2052.360 222.030 ;
        RECT 2064.580 221.690 2064.840 222.010 ;
        RECT 2064.640 210.965 2064.780 221.690 ;
        RECT 2076.600 221.330 2076.740 223.390 ;
        RECT 2086.200 222.370 2086.460 222.690 ;
        RECT 2080.220 222.030 2080.480 222.350 ;
        RECT 2071.020 221.010 2071.280 221.330 ;
        RECT 2076.540 221.010 2076.800 221.330 ;
        RECT 2071.080 210.965 2071.220 221.010 ;
        RECT 2080.280 210.965 2080.420 222.030 ;
        RECT 2086.260 210.965 2086.400 222.370 ;
        RECT 2095.400 222.030 2095.660 222.350 ;
        RECT 2095.460 210.965 2095.600 222.030 ;
        RECT 2298.320 210.965 2298.460 223.730 ;
        RECT 2307.460 223.050 2307.720 223.370 ;
        RECT 2307.520 210.965 2307.660 223.050 ;
        RECT 2310.680 222.030 2310.940 222.350 ;
        RECT 2325.860 222.030 2326.120 222.350 ;
        RECT 2310.740 210.965 2310.880 222.030 ;
        RECT 2325.920 210.965 2326.060 222.030 ;
        RECT 2338.340 210.965 2338.480 223.730 ;
        RECT 2339.200 223.390 2339.460 223.710 ;
        RECT 2366.340 223.390 2366.600 223.710 ;
        RECT 2339.260 223.030 2339.400 223.390 ;
        RECT 2339.200 222.710 2339.460 223.030 ;
        RECT 2344.720 222.710 2344.980 223.030 ;
        RECT 2344.780 210.965 2344.920 222.710 ;
        RECT 2366.400 222.690 2366.540 223.390 ;
        RECT 2580.760 223.370 2580.900 224.070 ;
        RECT 2580.700 223.050 2580.960 223.370 ;
        RECT 2359.900 222.370 2360.160 222.690 ;
        RECT 2366.340 222.370 2366.600 222.690 ;
        RECT 2572.420 222.370 2572.680 222.690 ;
        RECT 2353.920 222.030 2354.180 222.350 ;
        RECT 2353.980 210.965 2354.120 222.030 ;
        RECT 2359.960 210.965 2360.100 222.370 ;
        RECT 2369.100 222.030 2369.360 222.350 ;
        RECT 2369.160 210.965 2369.300 222.030 ;
        RECT 2572.480 210.965 2572.620 222.370 ;
        RECT 1476.300 209.030 1476.695 210.965 ;
        RECT 1476.415 208.565 1476.695 209.030 ;
        RECT 1479.635 208.565 1479.915 210.965 ;
        RECT 1482.855 208.565 1483.135 210.965 ;
        RECT 1485.500 209.030 1485.895 210.965 ;
        RECT 1488.720 209.030 1489.115 210.965 ;
        RECT 1485.615 208.565 1485.895 209.030 ;
        RECT 1488.835 208.565 1489.115 209.030 ;
        RECT 1492.055 208.565 1492.335 210.965 ;
        RECT 1494.815 208.565 1495.095 210.965 ;
        RECT 1497.920 209.030 1498.315 210.965 ;
        RECT 1498.035 208.565 1498.315 209.030 ;
        RECT 1501.255 208.565 1501.535 210.965 ;
        RECT 1503.900 209.170 1504.295 210.965 ;
        RECT 1507.235 209.170 1507.515 210.965 ;
        RECT 1510.455 209.170 1510.735 210.965 ;
        RECT 1503.900 209.030 1510.735 209.170 ;
        RECT 1516.320 209.030 1516.715 210.965 ;
        RECT 1522.760 209.030 1523.155 210.965 ;
        RECT 1525.520 209.170 1525.915 210.965 ;
        RECT 1526.380 209.450 1526.640 209.770 ;
        RECT 1526.440 209.170 1526.580 209.450 ;
        RECT 1525.520 209.030 1526.580 209.170 ;
        RECT 1528.740 209.030 1529.135 210.965 ;
        RECT 1532.075 209.835 1532.355 210.965 ;
        RECT 1531.500 209.770 1532.355 209.835 ;
        RECT 1531.440 209.695 1532.355 209.770 ;
        RECT 1531.440 209.450 1531.700 209.695 ;
        RECT 1531.960 209.030 1532.355 209.695 ;
        RECT 1537.940 209.030 1538.335 210.965 ;
        RECT 1543.400 209.450 1543.660 209.770 ;
        RECT 1543.460 209.170 1543.600 209.450 ;
        RECT 1544.035 209.170 1544.315 210.965 ;
        RECT 1547.140 209.170 1547.535 210.965 ;
        RECT 1543.460 209.030 1547.535 209.170 ;
        RECT 1504.015 208.565 1504.295 209.030 ;
        RECT 1507.235 208.565 1507.515 209.030 ;
        RECT 1510.455 208.565 1510.735 209.030 ;
        RECT 1516.435 208.565 1516.715 209.030 ;
        RECT 1522.875 208.565 1523.155 209.030 ;
        RECT 1525.635 208.565 1525.915 209.030 ;
        RECT 1528.855 208.565 1529.135 209.030 ;
        RECT 1532.075 208.565 1532.355 209.030 ;
        RECT 1538.055 208.565 1538.335 209.030 ;
        RECT 1544.035 208.565 1544.315 209.030 ;
        RECT 1547.255 208.565 1547.535 209.030 ;
        RECT 1553.235 208.565 1553.515 210.965 ;
        RECT 1750.415 208.565 1750.695 210.965 ;
        RECT 1753.635 208.565 1753.915 210.965 ;
        RECT 1756.855 208.565 1757.135 210.965 ;
        RECT 1759.615 208.565 1759.895 210.965 ;
        RECT 1762.835 208.565 1763.115 210.965 ;
        RECT 1766.055 208.565 1766.335 210.965 ;
        RECT 1768.815 208.565 1769.095 210.965 ;
        RECT 1772.035 208.565 1772.315 210.965 ;
        RECT 1775.255 208.565 1775.535 210.965 ;
        RECT 1778.015 209.170 1778.295 210.965 ;
        RECT 1781.235 209.170 1781.515 210.965 ;
        RECT 1784.455 209.170 1784.735 210.965 ;
        RECT 1778.015 209.030 1784.735 209.170 ;
        RECT 1778.015 208.565 1778.295 209.030 ;
        RECT 1781.235 208.565 1781.515 209.030 ;
        RECT 1784.455 208.565 1784.735 209.030 ;
        RECT 1790.435 208.565 1790.715 210.965 ;
        RECT 1796.875 208.565 1797.155 210.965 ;
        RECT 1799.635 209.170 1799.915 210.965 ;
        RECT 1799.635 209.090 1800.280 209.170 ;
        RECT 1799.635 209.030 1800.340 209.090 ;
        RECT 1799.635 208.565 1799.915 209.030 ;
        RECT 1800.080 208.770 1800.340 209.030 ;
        RECT 1802.855 208.565 1803.135 210.965 ;
        RECT 1806.075 209.170 1806.355 210.965 ;
        RECT 1805.660 209.090 1806.355 209.170 ;
        RECT 1805.600 209.030 1806.355 209.090 ;
        RECT 1805.600 208.770 1805.860 209.030 ;
        RECT 1806.075 208.565 1806.355 209.030 ;
        RECT 1812.055 208.565 1812.335 210.965 ;
        RECT 1818.035 209.170 1818.315 210.965 ;
        RECT 1821.255 209.170 1821.535 210.965 ;
        RECT 1817.620 209.090 1821.535 209.170 ;
        RECT 1817.560 209.030 1821.535 209.090 ;
        RECT 1817.560 208.770 1817.820 209.030 ;
        RECT 1818.035 208.565 1818.315 209.030 ;
        RECT 1821.255 208.565 1821.535 209.030 ;
        RECT 1827.235 208.565 1827.515 210.965 ;
        RECT 2024.415 209.100 2024.760 210.965 ;
        RECT 2024.415 208.565 2024.695 209.100 ;
        RECT 2030.855 208.565 2031.135 210.965 ;
        RECT 2033.615 209.100 2033.960 210.965 ;
        RECT 2036.835 209.100 2037.180 210.965 ;
        RECT 2033.615 208.565 2033.895 209.100 ;
        RECT 2036.835 208.565 2037.115 209.100 ;
        RECT 2040.055 208.565 2040.335 210.965 ;
        RECT 2042.815 208.565 2043.095 210.965 ;
        RECT 2049.255 208.565 2049.535 210.965 ;
        RECT 2052.015 209.170 2052.360 210.965 ;
        RECT 2058.455 209.170 2058.735 210.965 ;
        RECT 2052.015 209.090 2052.820 209.170 ;
        RECT 2057.740 209.090 2058.735 209.170 ;
        RECT 2052.015 209.030 2052.880 209.090 ;
        RECT 2052.015 208.565 2052.295 209.030 ;
        RECT 2052.620 208.770 2052.880 209.030 ;
        RECT 2057.680 209.030 2058.735 209.090 ;
        RECT 2057.680 208.770 2057.940 209.030 ;
        RECT 2058.455 208.565 2058.735 209.030 ;
        RECT 2064.435 209.100 2064.780 210.965 ;
        RECT 2070.875 209.100 2071.220 210.965 ;
        RECT 2073.635 209.170 2073.915 210.965 ;
        RECT 2080.075 209.170 2080.420 210.965 ;
        RECT 2064.435 208.565 2064.715 209.100 ;
        RECT 2070.875 208.565 2071.155 209.100 ;
        RECT 2073.635 209.090 2074.440 209.170 ;
        RECT 2079.360 209.100 2080.420 209.170 ;
        RECT 2086.055 209.100 2086.400 210.965 ;
        RECT 2092.035 209.170 2092.315 210.965 ;
        RECT 2095.255 209.170 2095.600 210.965 ;
        RECT 2092.035 209.100 2095.600 209.170 ;
        RECT 2079.360 209.090 2080.355 209.100 ;
        RECT 2073.635 209.030 2074.500 209.090 ;
        RECT 2073.635 208.565 2073.915 209.030 ;
        RECT 2074.240 208.770 2074.500 209.030 ;
        RECT 2079.300 209.030 2080.355 209.090 ;
        RECT 2079.300 208.770 2079.560 209.030 ;
        RECT 2080.075 208.565 2080.355 209.030 ;
        RECT 2086.055 208.565 2086.335 209.100 ;
        RECT 2092.035 209.030 2095.535 209.100 ;
        RECT 2092.035 208.565 2092.315 209.030 ;
        RECT 2095.255 208.565 2095.535 209.030 ;
        RECT 2101.235 208.565 2101.515 210.965 ;
        RECT 2298.320 209.030 2298.695 210.965 ;
        RECT 2298.415 208.565 2298.695 209.030 ;
        RECT 2304.855 208.565 2305.135 210.965 ;
        RECT 2307.520 209.030 2307.895 210.965 ;
        RECT 2310.740 209.030 2311.115 210.965 ;
        RECT 2307.615 208.565 2307.895 209.030 ;
        RECT 2310.835 208.565 2311.115 209.030 ;
        RECT 2314.055 208.565 2314.335 210.965 ;
        RECT 2316.815 208.565 2317.095 210.965 ;
        RECT 2323.255 208.565 2323.535 210.965 ;
        RECT 2325.920 209.170 2326.295 210.965 ;
        RECT 2332.455 209.170 2332.735 210.965 ;
        RECT 2325.920 209.090 2326.980 209.170 ;
        RECT 2331.900 209.090 2332.735 209.170 ;
        RECT 2325.920 209.030 2327.040 209.090 ;
        RECT 2326.015 208.565 2326.295 209.030 ;
        RECT 2326.780 208.770 2327.040 209.030 ;
        RECT 2331.840 209.030 2332.735 209.090 ;
        RECT 2338.340 209.030 2338.715 210.965 ;
        RECT 2344.780 209.030 2345.155 210.965 ;
        RECT 2347.635 209.170 2347.915 210.965 ;
        RECT 2348.400 209.790 2348.660 210.110 ;
        RECT 2353.460 209.850 2353.720 210.110 ;
        RECT 2353.980 209.850 2354.355 210.965 ;
        RECT 2353.460 209.790 2354.355 209.850 ;
        RECT 2348.460 209.170 2348.600 209.790 ;
        RECT 2353.520 209.710 2354.355 209.790 ;
        RECT 2347.080 209.090 2348.600 209.170 ;
        RECT 2331.840 208.770 2332.100 209.030 ;
        RECT 2332.455 208.565 2332.735 209.030 ;
        RECT 2338.435 208.565 2338.715 209.030 ;
        RECT 2344.875 208.565 2345.155 209.030 ;
        RECT 2347.020 209.030 2348.600 209.090 ;
        RECT 2353.980 209.030 2354.355 209.710 ;
        RECT 2359.960 209.030 2360.335 210.965 ;
        RECT 2347.020 208.770 2347.280 209.030 ;
        RECT 2347.635 208.565 2347.915 209.030 ;
        RECT 2354.075 208.565 2354.355 209.030 ;
        RECT 2360.055 208.565 2360.335 209.030 ;
        RECT 2366.035 209.170 2366.315 210.965 ;
        RECT 2369.160 209.170 2369.535 210.965 ;
        RECT 2366.035 209.030 2369.535 209.170 ;
        RECT 2366.035 208.565 2366.315 209.030 ;
        RECT 2369.255 208.565 2369.535 209.030 ;
        RECT 2375.235 208.565 2375.515 210.965 ;
        RECT 2572.415 208.565 2572.695 210.965 ;
        RECT 2578.855 208.565 2579.135 210.965 ;
        RECT 2580.760 209.170 2580.900 223.050 ;
        RECT 2618.940 223.030 2619.080 224.410 ;
        RECT 2634.060 223.390 2634.320 223.710 ;
        RECT 2618.880 222.710 2619.140 223.030 ;
        RECT 2612.440 222.370 2612.700 222.690 ;
        RECT 2584.840 222.030 2585.100 222.350 ;
        RECT 2600.020 222.030 2600.280 222.350 ;
        RECT 2584.900 210.965 2585.040 222.030 ;
        RECT 2600.080 210.965 2600.220 222.030 ;
        RECT 2612.500 210.965 2612.640 222.370 ;
        RECT 2618.940 210.965 2619.080 222.710 ;
        RECT 2634.120 210.965 2634.260 223.390 ;
        RECT 2581.615 209.170 2581.895 210.965 ;
        RECT 2580.760 209.030 2581.895 209.170 ;
        RECT 2581.615 208.565 2581.895 209.030 ;
        RECT 2584.835 208.565 2585.115 210.965 ;
        RECT 2588.055 208.565 2588.335 210.965 ;
        RECT 2590.815 208.565 2591.095 210.965 ;
        RECT 2597.255 208.565 2597.535 210.965 ;
        RECT 2600.015 209.170 2600.295 210.965 ;
        RECT 2606.455 209.170 2606.735 210.965 ;
        RECT 2600.015 209.090 2600.680 209.170 ;
        RECT 2606.060 209.090 2606.735 209.170 ;
        RECT 2600.015 209.030 2600.740 209.090 ;
        RECT 2600.015 208.565 2600.295 209.030 ;
        RECT 2600.480 208.770 2600.740 209.030 ;
        RECT 2606.000 209.030 2606.735 209.090 ;
        RECT 2606.000 208.770 2606.260 209.030 ;
        RECT 2606.455 208.565 2606.735 209.030 ;
        RECT 2612.435 208.565 2612.715 210.965 ;
        RECT 2618.875 208.565 2619.155 210.965 ;
        RECT 2621.635 209.170 2621.915 210.965 ;
        RECT 2628.075 209.170 2628.355 210.965 ;
        RECT 2621.240 209.090 2621.915 209.170 ;
        RECT 2627.680 209.090 2628.355 209.170 ;
        RECT 2621.180 209.030 2621.915 209.090 ;
        RECT 2621.180 208.770 2621.440 209.030 ;
        RECT 2621.635 208.565 2621.915 209.030 ;
        RECT 2627.620 209.030 2628.355 209.090 ;
        RECT 2627.620 208.770 2627.880 209.030 ;
        RECT 2628.075 208.565 2628.355 209.030 ;
        RECT 2634.055 208.565 2634.335 210.965 ;
        RECT 2640.035 209.170 2640.315 210.965 ;
        RECT 2643.255 209.835 2643.535 210.965 ;
        RECT 2642.400 209.695 2643.535 209.835 ;
        RECT 2642.400 209.170 2642.540 209.695 ;
        RECT 2639.640 209.090 2642.540 209.170 ;
        RECT 2639.580 209.030 2642.540 209.090 ;
        RECT 2639.580 208.770 2639.840 209.030 ;
        RECT 2640.035 208.565 2640.315 209.030 ;
        RECT 2643.255 208.565 2643.535 209.695 ;
        RECT 2649.235 208.565 2649.515 210.965 ;
      LAYER met2 ;
        RECT 1475.085 208.285 1476.135 208.565 ;
        RECT 1476.975 208.285 1479.355 208.565 ;
        RECT 1480.195 208.285 1482.575 208.565 ;
        RECT 1483.415 208.285 1485.335 208.565 ;
        RECT 1486.175 208.285 1488.555 208.565 ;
        RECT 1489.395 208.285 1491.775 208.565 ;
        RECT 1492.615 208.285 1494.535 208.565 ;
        RECT 1495.375 208.285 1497.755 208.565 ;
        RECT 1498.595 208.285 1500.975 208.565 ;
        RECT 1501.815 208.285 1503.735 208.565 ;
        RECT 1504.575 208.285 1506.955 208.565 ;
        RECT 1507.795 208.285 1510.175 208.565 ;
        RECT 1511.015 208.285 1512.935 208.565 ;
        RECT 1513.775 208.285 1516.155 208.565 ;
        RECT 1516.995 208.285 1519.375 208.565 ;
        RECT 1520.215 208.285 1522.595 208.565 ;
        RECT 1523.435 208.285 1525.355 208.565 ;
        RECT 1526.195 208.285 1528.575 208.565 ;
        RECT 1529.415 208.285 1531.795 208.565 ;
        RECT 1532.635 208.285 1534.555 208.565 ;
        RECT 1535.395 208.285 1537.775 208.565 ;
        RECT 1538.615 208.285 1540.995 208.565 ;
        RECT 1541.835 208.285 1543.755 208.565 ;
        RECT 1544.595 208.285 1546.975 208.565 ;
        RECT 1547.815 208.285 1550.195 208.565 ;
        RECT 1551.035 208.285 1552.955 208.565 ;
        RECT 1553.795 208.285 1554.790 208.565 ;
      LAYER met2 ;
        RECT 1262.790 206.875 1263.070 207.245 ;
        RECT 1262.800 206.730 1263.060 206.875 ;
        RECT 1206.670 198.715 1206.950 199.085 ;
      LAYER met2 ;
        RECT 1206.300 197.965 1226.905 198.000 ;
        RECT 1227.465 197.965 1260.075 198.000 ;
        RECT 1260.505 197.965 1280.500 198.000 ;
        RECT 1194.805 159.640 1205.755 163.510 ;
        RECT 1206.000 158.415 1280.500 197.965 ;
        RECT 1194.860 153.765 1280.500 158.415 ;
        RECT 1206.000 3.570 1280.500 153.765 ;
        RECT 1475.085 0.000 1554.790 208.285 ;
        RECT 1749.085 208.285 1750.135 208.565 ;
        RECT 1750.975 208.285 1753.355 208.565 ;
        RECT 1754.195 208.285 1756.575 208.565 ;
        RECT 1757.415 208.285 1759.335 208.565 ;
        RECT 1760.175 208.285 1762.555 208.565 ;
        RECT 1763.395 208.285 1765.775 208.565 ;
        RECT 1766.615 208.285 1768.535 208.565 ;
        RECT 1769.375 208.285 1771.755 208.565 ;
        RECT 1772.595 208.285 1774.975 208.565 ;
        RECT 1775.815 208.285 1777.735 208.565 ;
        RECT 1778.575 208.285 1780.955 208.565 ;
        RECT 1781.795 208.285 1784.175 208.565 ;
        RECT 1785.015 208.285 1786.935 208.565 ;
        RECT 1787.775 208.285 1790.155 208.565 ;
        RECT 1790.995 208.285 1793.375 208.565 ;
        RECT 1794.215 208.285 1796.595 208.565 ;
        RECT 1797.435 208.285 1799.355 208.565 ;
        RECT 1800.195 208.285 1802.575 208.565 ;
        RECT 1803.415 208.285 1805.795 208.565 ;
        RECT 1806.635 208.285 1808.555 208.565 ;
        RECT 1809.395 208.285 1811.775 208.565 ;
        RECT 1812.615 208.285 1814.995 208.565 ;
        RECT 1815.835 208.285 1817.755 208.565 ;
        RECT 1818.595 208.285 1820.975 208.565 ;
        RECT 1821.815 208.285 1824.195 208.565 ;
        RECT 1825.035 208.285 1826.955 208.565 ;
        RECT 1827.795 208.285 1828.790 208.565 ;
        RECT 1749.085 0.000 1828.790 208.285 ;
        RECT 2023.085 208.285 2024.135 208.565 ;
        RECT 2024.975 208.285 2027.355 208.565 ;
        RECT 2028.195 208.285 2030.575 208.565 ;
        RECT 2031.415 208.285 2033.335 208.565 ;
        RECT 2034.175 208.285 2036.555 208.565 ;
        RECT 2037.395 208.285 2039.775 208.565 ;
        RECT 2040.615 208.285 2042.535 208.565 ;
        RECT 2043.375 208.285 2045.755 208.565 ;
        RECT 2046.595 208.285 2048.975 208.565 ;
        RECT 2049.815 208.285 2051.735 208.565 ;
        RECT 2052.575 208.285 2054.955 208.565 ;
        RECT 2055.795 208.285 2058.175 208.565 ;
        RECT 2059.015 208.285 2060.935 208.565 ;
        RECT 2061.775 208.285 2064.155 208.565 ;
        RECT 2064.995 208.285 2067.375 208.565 ;
        RECT 2068.215 208.285 2070.595 208.565 ;
        RECT 2071.435 208.285 2073.355 208.565 ;
        RECT 2074.195 208.285 2076.575 208.565 ;
        RECT 2077.415 208.285 2079.795 208.565 ;
        RECT 2080.635 208.285 2082.555 208.565 ;
        RECT 2083.395 208.285 2085.775 208.565 ;
        RECT 2086.615 208.285 2088.995 208.565 ;
        RECT 2089.835 208.285 2091.755 208.565 ;
        RECT 2092.595 208.285 2094.975 208.565 ;
        RECT 2095.815 208.285 2098.195 208.565 ;
        RECT 2099.035 208.285 2100.955 208.565 ;
        RECT 2101.795 208.285 2102.790 208.565 ;
        RECT 2023.085 0.000 2102.790 208.285 ;
        RECT 2297.085 208.285 2298.135 208.565 ;
        RECT 2298.975 208.285 2301.355 208.565 ;
        RECT 2302.195 208.285 2304.575 208.565 ;
        RECT 2305.415 208.285 2307.335 208.565 ;
        RECT 2308.175 208.285 2310.555 208.565 ;
        RECT 2311.395 208.285 2313.775 208.565 ;
        RECT 2314.615 208.285 2316.535 208.565 ;
        RECT 2317.375 208.285 2319.755 208.565 ;
        RECT 2320.595 208.285 2322.975 208.565 ;
        RECT 2323.815 208.285 2325.735 208.565 ;
        RECT 2326.575 208.285 2328.955 208.565 ;
        RECT 2329.795 208.285 2332.175 208.565 ;
        RECT 2333.015 208.285 2334.935 208.565 ;
        RECT 2335.775 208.285 2338.155 208.565 ;
        RECT 2338.995 208.285 2341.375 208.565 ;
        RECT 2342.215 208.285 2344.595 208.565 ;
        RECT 2345.435 208.285 2347.355 208.565 ;
        RECT 2348.195 208.285 2350.575 208.565 ;
        RECT 2351.415 208.285 2353.795 208.565 ;
        RECT 2354.635 208.285 2356.555 208.565 ;
        RECT 2357.395 208.285 2359.775 208.565 ;
        RECT 2360.615 208.285 2362.995 208.565 ;
        RECT 2363.835 208.285 2365.755 208.565 ;
        RECT 2366.595 208.285 2368.975 208.565 ;
        RECT 2369.815 208.285 2372.195 208.565 ;
        RECT 2373.035 208.285 2374.955 208.565 ;
        RECT 2375.795 208.285 2376.790 208.565 ;
        RECT 2297.085 0.000 2376.790 208.285 ;
        RECT 2571.085 208.285 2572.135 208.565 ;
        RECT 2572.975 208.285 2575.355 208.565 ;
        RECT 2576.195 208.285 2578.575 208.565 ;
        RECT 2579.415 208.285 2581.335 208.565 ;
        RECT 2582.175 208.285 2584.555 208.565 ;
        RECT 2585.395 208.285 2587.775 208.565 ;
        RECT 2588.615 208.285 2590.535 208.565 ;
        RECT 2591.375 208.285 2593.755 208.565 ;
        RECT 2594.595 208.285 2596.975 208.565 ;
        RECT 2597.815 208.285 2599.735 208.565 ;
        RECT 2600.575 208.285 2602.955 208.565 ;
        RECT 2603.795 208.285 2606.175 208.565 ;
        RECT 2607.015 208.285 2608.935 208.565 ;
        RECT 2609.775 208.285 2612.155 208.565 ;
        RECT 2612.995 208.285 2615.375 208.565 ;
        RECT 2616.215 208.285 2618.595 208.565 ;
        RECT 2619.435 208.285 2621.355 208.565 ;
        RECT 2622.195 208.285 2624.575 208.565 ;
        RECT 2625.415 208.285 2627.795 208.565 ;
        RECT 2628.635 208.285 2630.555 208.565 ;
        RECT 2631.395 208.285 2633.775 208.565 ;
        RECT 2634.615 208.285 2636.995 208.565 ;
        RECT 2637.835 208.285 2639.755 208.565 ;
        RECT 2640.595 208.285 2642.975 208.565 ;
        RECT 2643.815 208.285 2646.195 208.565 ;
        RECT 2647.035 208.285 2648.955 208.565 ;
        RECT 2649.795 208.285 2650.790 208.565 ;
        RECT 2571.085 0.000 2650.790 208.285 ;
      LAYER met2 ;
        RECT 2863.600 206.730 2863.860 207.050 ;
        RECT 2863.660 203.650 2863.800 206.730 ;
        RECT 3374.260 203.650 3374.400 562.370 ;
        RECT 3374.720 545.690 3374.860 775.890 ;
        RECT 3375.180 735.750 3375.320 782.950 ;
      LAYER met2 ;
        RECT 3379.715 782.795 3588.000 783.635 ;
        RECT 3379.435 780.415 3588.000 782.795 ;
        RECT 3379.715 779.575 3588.000 780.415 ;
        RECT 3379.435 777.195 3588.000 779.575 ;
        RECT 3379.715 776.355 3588.000 777.195 ;
      LAYER met2 ;
        RECT 3376.960 775.890 3377.220 776.210 ;
        RECT 3377.020 774.155 3377.160 775.890 ;
      LAYER met2 ;
        RECT 3379.435 774.435 3588.000 776.355 ;
      LAYER met2 ;
        RECT 3377.020 774.015 3379.435 774.155 ;
        RECT 3377.035 773.875 3379.435 774.015 ;
      LAYER met2 ;
        RECT 3379.715 773.595 3588.000 774.435 ;
        RECT 3379.435 771.215 3588.000 773.595 ;
        RECT 3379.715 770.375 3588.000 771.215 ;
        RECT 3379.435 767.995 3588.000 770.375 ;
      LAYER met2 ;
        RECT 3377.035 767.645 3379.435 767.715 ;
        RECT 3376.560 767.505 3379.435 767.645 ;
        RECT 3375.120 735.430 3375.380 735.750 ;
        RECT 3376.040 735.430 3376.300 735.750 ;
        RECT 3376.100 710.770 3376.240 735.430 ;
        RECT 3376.560 727.625 3376.700 767.505 ;
        RECT 3377.035 767.435 3379.435 767.505 ;
      LAYER met2 ;
        RECT 3379.715 767.155 3588.000 767.995 ;
        RECT 3379.435 764.775 3588.000 767.155 ;
        RECT 3379.715 763.935 3588.000 764.775 ;
        RECT 3379.435 762.015 3588.000 763.935 ;
        RECT 3379.715 761.175 3588.000 762.015 ;
        RECT 3379.435 758.795 3588.000 761.175 ;
        RECT 3379.715 757.955 3588.000 758.795 ;
        RECT 3379.435 755.575 3588.000 757.955 ;
        RECT 3379.715 754.735 3588.000 755.575 ;
        RECT 3379.435 752.815 3588.000 754.735 ;
      LAYER met2 ;
        RECT 3377.035 752.255 3379.435 752.535 ;
      LAYER met2 ;
        RECT 3379.715 751.975 3588.000 752.815 ;
        RECT 3379.435 749.595 3588.000 751.975 ;
        RECT 3379.715 748.755 3588.000 749.595 ;
        RECT 3379.435 746.375 3588.000 748.755 ;
      LAYER met2 ;
        RECT 3377.035 745.815 3379.435 746.095 ;
      LAYER met2 ;
        RECT 3379.715 745.535 3588.000 746.375 ;
        RECT 3379.435 743.615 3588.000 745.535 ;
      LAYER met2 ;
        RECT 3377.035 743.055 3379.435 743.335 ;
      LAYER met2 ;
        RECT 3379.715 742.775 3588.000 743.615 ;
        RECT 3379.435 740.395 3588.000 742.775 ;
        RECT 3379.715 739.555 3588.000 740.395 ;
        RECT 3379.435 737.175 3588.000 739.555 ;
      LAYER met2 ;
        RECT 3377.035 736.780 3379.435 736.895 ;
        RECT 3377.020 736.615 3379.435 736.780 ;
        RECT 3377.020 735.750 3377.160 736.615 ;
      LAYER met2 ;
        RECT 3379.715 736.335 3588.000 737.175 ;
      LAYER met2 ;
        RECT 3376.960 735.430 3377.220 735.750 ;
      LAYER met2 ;
        RECT 3379.435 734.415 3588.000 736.335 ;
      LAYER met2 ;
        RECT 3377.035 733.855 3379.435 734.135 ;
      LAYER met2 ;
        RECT 3379.715 733.575 3588.000 734.415 ;
        RECT 3379.435 731.195 3588.000 733.575 ;
        RECT 3379.715 730.355 3588.000 731.195 ;
        RECT 3379.435 727.975 3588.000 730.355 ;
      LAYER met2 ;
        RECT 3377.035 727.625 3379.435 727.695 ;
        RECT 3376.560 727.485 3379.435 727.625 ;
        RECT 3377.035 727.415 3379.435 727.485 ;
      LAYER met2 ;
        RECT 3379.715 727.135 3588.000 727.975 ;
        RECT 3379.435 726.085 3588.000 727.135 ;
      LAYER met2 ;
        RECT 3376.100 710.630 3376.700 710.770 ;
        RECT 3374.660 545.370 3374.920 545.690 ;
        RECT 3374.720 224.730 3374.860 545.370 ;
        RECT 3376.040 538.910 3376.300 539.230 ;
        RECT 3376.100 510.330 3376.240 538.910 ;
        RECT 3376.040 510.010 3376.300 510.330 ;
        RECT 3376.560 509.730 3376.700 710.630 ;
      LAYER met2 ;
        RECT 3379.435 578.795 3588.000 579.790 ;
      LAYER met2 ;
        RECT 3377.035 578.235 3379.435 578.515 ;
      LAYER met2 ;
        RECT 3379.715 577.955 3588.000 578.795 ;
        RECT 3379.435 576.035 3588.000 577.955 ;
        RECT 3379.715 575.195 3588.000 576.035 ;
        RECT 3379.435 572.815 3588.000 575.195 ;
        RECT 3379.715 571.975 3588.000 572.815 ;
        RECT 3379.435 569.595 3588.000 571.975 ;
        RECT 3379.715 568.755 3588.000 569.595 ;
        RECT 3379.435 566.835 3588.000 568.755 ;
        RECT 3379.715 565.995 3588.000 566.835 ;
        RECT 3379.435 563.615 3588.000 565.995 ;
      LAYER met2 ;
        RECT 3377.035 563.195 3379.435 563.335 ;
        RECT 3377.020 563.055 3379.435 563.195 ;
        RECT 3377.020 562.690 3377.160 563.055 ;
      LAYER met2 ;
        RECT 3379.715 562.775 3588.000 563.615 ;
      LAYER met2 ;
        RECT 3376.960 562.370 3377.220 562.690 ;
      LAYER met2 ;
        RECT 3379.435 560.395 3588.000 562.775 ;
        RECT 3379.715 559.555 3588.000 560.395 ;
        RECT 3379.435 557.635 3588.000 559.555 ;
        RECT 3379.715 556.795 3588.000 557.635 ;
        RECT 3379.435 554.415 3588.000 556.795 ;
        RECT 3379.715 553.575 3588.000 554.415 ;
        RECT 3379.435 551.195 3588.000 553.575 ;
        RECT 3379.715 550.355 3588.000 551.195 ;
        RECT 3379.435 548.435 3588.000 550.355 ;
      LAYER met2 ;
        RECT 3377.035 548.015 3379.435 548.155 ;
        RECT 3377.020 547.875 3379.435 548.015 ;
        RECT 3377.020 545.690 3377.160 547.875 ;
      LAYER met2 ;
        RECT 3379.715 547.595 3588.000 548.435 ;
      LAYER met2 ;
        RECT 3376.960 545.370 3377.220 545.690 ;
      LAYER met2 ;
        RECT 3379.435 545.215 3588.000 547.595 ;
        RECT 3379.715 544.375 3588.000 545.215 ;
        RECT 3379.435 541.995 3588.000 544.375 ;
      LAYER met2 ;
        RECT 3377.035 541.620 3379.435 541.715 ;
        RECT 3377.020 541.435 3379.435 541.620 ;
        RECT 3377.020 539.230 3377.160 541.435 ;
      LAYER met2 ;
        RECT 3379.715 541.155 3588.000 541.995 ;
      LAYER met2 ;
        RECT 3376.960 538.910 3377.220 539.230 ;
      LAYER met2 ;
        RECT 3379.435 538.775 3588.000 541.155 ;
        RECT 3379.715 537.935 3588.000 538.775 ;
        RECT 3379.435 536.015 3588.000 537.935 ;
        RECT 3379.715 535.175 3588.000 536.015 ;
        RECT 3379.435 532.795 3588.000 535.175 ;
        RECT 3379.715 531.955 3588.000 532.795 ;
        RECT 3379.435 529.575 3588.000 531.955 ;
        RECT 3379.715 528.735 3588.000 529.575 ;
        RECT 3379.435 526.815 3588.000 528.735 ;
      LAYER met2 ;
        RECT 3377.035 526.255 3379.435 526.535 ;
      LAYER met2 ;
        RECT 3379.715 525.975 3588.000 526.815 ;
        RECT 3379.435 523.595 3588.000 525.975 ;
        RECT 3379.715 522.755 3588.000 523.595 ;
        RECT 3379.435 520.375 3588.000 522.755 ;
      LAYER met2 ;
        RECT 3377.035 519.815 3379.435 520.095 ;
      LAYER met2 ;
        RECT 3379.715 519.535 3588.000 520.375 ;
        RECT 3379.435 517.615 3588.000 519.535 ;
      LAYER met2 ;
        RECT 3377.035 517.055 3379.435 517.335 ;
      LAYER met2 ;
        RECT 3379.715 516.775 3588.000 517.615 ;
        RECT 3379.435 514.395 3588.000 516.775 ;
        RECT 3379.715 513.555 3588.000 514.395 ;
        RECT 3379.435 511.175 3588.000 513.555 ;
      LAYER met2 ;
        RECT 3377.035 510.755 3379.435 510.895 ;
        RECT 3377.020 510.615 3379.435 510.755 ;
        RECT 3377.020 509.730 3377.160 510.615 ;
      LAYER met2 ;
        RECT 3379.715 510.335 3588.000 511.175 ;
      LAYER met2 ;
        RECT 3375.640 509.590 3377.160 509.730 ;
        RECT 3374.660 224.410 3374.920 224.730 ;
        RECT 3375.640 224.390 3375.780 509.590 ;
        RECT 3376.500 508.990 3376.760 509.310 ;
        RECT 3376.560 501.570 3376.700 508.990 ;
      LAYER met2 ;
        RECT 3379.435 508.415 3588.000 510.335 ;
      LAYER met2 ;
        RECT 3377.035 507.855 3379.435 508.135 ;
      LAYER met2 ;
        RECT 3379.715 507.575 3588.000 508.415 ;
        RECT 3379.435 505.195 3588.000 507.575 ;
        RECT 3379.715 504.355 3588.000 505.195 ;
        RECT 3379.435 501.975 3588.000 504.355 ;
      LAYER met2 ;
        RECT 3377.035 501.570 3379.435 501.695 ;
        RECT 3376.560 501.430 3379.435 501.570 ;
        RECT 3377.035 501.415 3379.435 501.430 ;
      LAYER met2 ;
        RECT 3379.715 501.135 3588.000 501.975 ;
        RECT 3379.435 500.085 3588.000 501.135 ;
      LAYER met2 ;
        RECT 3375.580 224.070 3375.840 224.390 ;
        RECT 2863.600 203.330 2863.860 203.650 ;
        RECT 3374.200 203.330 3374.460 203.650 ;
        RECT 2863.660 201.125 2863.800 203.330 ;
        RECT 2863.590 200.755 2863.870 201.125 ;
      LAYER met2 ;
        RECT 2845.710 197.965 2869.610 200.000 ;
        RECT 2892.105 198.080 2894.105 200.000 ;
        RECT 2895.605 197.965 2919.505 200.000 ;
        RECT 3114.710 197.965 3138.610 200.000 ;
        RECT 3161.105 198.080 3163.105 200.000 ;
        RECT 3164.605 197.965 3188.505 200.000 ;
        RECT 2845.710 4.925 2919.735 197.965 ;
        RECT 3114.710 4.925 3188.735 197.965 ;
      LAYER via2 ;
        RECT 1666.210 4989.360 1666.490 4989.640 ;
        RECT 207.090 4409.320 207.370 4409.600 ;
        RECT 207.090 4399.800 207.370 4400.080 ;
        RECT 211.230 4399.800 211.510 4400.080 ;
        RECT 2903.150 4989.360 2903.430 4989.640 ;
        RECT 213.070 4409.320 213.350 4409.600 ;
        RECT 3387.530 4091.760 3387.810 4092.040 ;
        RECT 3387.530 2518.920 3387.810 2519.200 ;
        RECT 3387.530 2127.920 3387.810 2128.200 ;
        RECT 210.310 565.960 210.590 566.240 ;
        RECT 210.770 391.200 211.050 391.480 ;
        RECT 212.610 565.960 212.890 566.240 ;
        RECT 212.150 391.200 212.430 391.480 ;
        RECT 715.390 201.480 715.670 201.760 ;
        RECT 443.990 199.440 444.270 199.720 ;
        RECT 738.390 199.440 738.670 199.720 ;
        RECT 1198.390 206.920 1198.670 207.200 ;
        RECT 1262.790 206.920 1263.070 207.200 ;
        RECT 1206.670 198.760 1206.950 199.040 ;
        RECT 2863.590 200.800 2863.870 201.080 ;
      LAYER met3 ;
        RECT 381.310 4986.690 460.570 5188.000 ;
        RECT 638.310 4986.690 717.570 5188.000 ;
        RECT 895.310 4986.690 974.570 5188.000 ;
        RECT 1152.310 4986.690 1231.570 5188.000 ;
        RECT 1410.310 4986.690 1489.570 5188.000 ;
        RECT 1667.240 5014.250 1741.290 5188.000 ;
      LAYER met3 ;
        RECT 1666.185 4989.650 1666.515 4989.665 ;
        RECT 1667.495 4989.650 1691.395 5013.850 ;
      LAYER met3 ;
        RECT 1691.795 4990.035 1716.990 5014.250 ;
      LAYER met3 ;
        RECT 1666.185 4989.350 1691.395 4989.650 ;
        RECT 1666.185 4989.335 1666.515 4989.350 ;
        RECT 1667.350 4988.140 1691.395 4989.350 ;
        RECT 1667.495 4988.000 1691.395 4988.140 ;
      LAYER met3 ;
        RECT 1692.895 4988.000 1703.895 4990.035 ;
        RECT 1704.890 4988.000 1715.890 4990.035 ;
      LAYER met3 ;
        RECT 1717.390 4988.000 1741.290 5013.850 ;
      LAYER met3 ;
        RECT 1919.310 4986.690 1998.570 5188.000 ;
        RECT 2364.310 4986.690 2443.570 5188.000 ;
        RECT 2621.310 4986.690 2700.570 5188.000 ;
        RECT 2878.240 5025.160 2952.290 5183.100 ;
        RECT 2878.240 5020.915 2927.990 5025.160 ;
      LAYER met3 ;
        RECT 2878.495 4989.650 2902.395 5020.515 ;
      LAYER met3 ;
        RECT 2902.795 4990.035 2927.990 5020.915 ;
      LAYER met3 ;
        RECT 2903.125 4989.650 2903.455 4989.665 ;
        RECT 2878.495 4989.350 2903.455 4989.650 ;
        RECT 2878.495 4988.000 2902.395 4989.350 ;
        RECT 2903.125 4989.335 2903.455 4989.350 ;
      LAYER met3 ;
        RECT 2903.895 4988.000 2914.895 4990.035 ;
        RECT 2915.890 4988.000 2926.890 4990.035 ;
      LAYER met3 ;
        RECT 2928.390 4988.000 2952.290 5024.760 ;
      LAYER met3 ;
        RECT 3130.310 4986.690 3209.570 5188.000 ;
        RECT 0.000 4771.310 201.310 4850.570 ;
        RECT 3386.690 4758.430 3588.000 4837.690 ;
        RECT 0.035 4636.200 24.250 4645.935 ;
        RECT 153.765 4635.605 158.415 4646.140 ;
        RECT 169.550 4636.200 174.200 4645.935 ;
        RECT 0.035 4610.355 190.700 4635.000 ;
      LAYER met3 ;
        RECT 191.100 4610.755 198.000 4634.700 ;
      LAYER met3 ;
        RECT 3429.550 4613.895 3434.200 4623.975 ;
        RECT 3390.035 4612.900 3587.965 4613.000 ;
        RECT 0.035 4609.255 197.965 4610.355 ;
        RECT 0.035 4598.380 198.000 4609.255 ;
        RECT 0.035 4596.880 197.965 4598.380 ;
        RECT 0.035 4586.000 198.000 4596.880 ;
      LAYER met3 ;
        RECT 3390.000 4588.500 3396.900 4612.500 ;
      LAYER met3 ;
        RECT 3397.300 4588.100 3587.965 4612.900 ;
        RECT 3390.035 4587.000 3587.965 4588.100 ;
        RECT 0.035 4584.900 197.965 4586.000 ;
        RECT 0.035 4560.100 190.700 4584.900 ;
      LAYER met3 ;
        RECT 191.100 4560.500 198.000 4584.500 ;
      LAYER met3 ;
        RECT 3390.000 4576.120 3587.965 4587.000 ;
        RECT 3390.035 4574.620 3587.965 4576.120 ;
        RECT 3390.000 4563.745 3587.965 4574.620 ;
        RECT 3390.035 4562.645 3587.965 4563.745 ;
        RECT 0.035 4560.000 197.965 4560.100 ;
        RECT 153.800 4549.025 158.450 4559.105 ;
      LAYER met3 ;
        RECT 3390.000 4538.300 3396.900 4562.245 ;
      LAYER met3 ;
        RECT 3397.300 4538.000 3587.965 4562.645 ;
        RECT 3413.800 4527.065 3418.450 4536.800 ;
        RECT 3429.585 4526.860 3434.235 4537.395 ;
        RECT 3563.750 4527.065 3587.965 4536.800 ;
        RECT 0.000 4398.990 179.800 4423.290 ;
      LAYER met3 ;
        RECT 180.200 4400.090 200.000 4423.290 ;
        RECT 207.065 4409.610 207.395 4409.625 ;
        RECT 213.045 4409.610 213.375 4409.625 ;
        RECT 207.065 4409.310 213.375 4409.610 ;
        RECT 207.065 4409.295 207.395 4409.310 ;
        RECT 213.045 4409.295 213.375 4409.310 ;
        RECT 207.065 4400.090 207.395 4400.105 ;
        RECT 211.205 4400.090 211.535 4400.105 ;
        RECT 180.200 4399.790 211.535 4400.090 ;
        RECT 180.200 4399.390 200.000 4399.790 ;
        RECT 207.065 4399.775 207.395 4399.790 ;
        RECT 211.205 4399.775 211.535 4399.790 ;
      LAYER met3 ;
        RECT 0.000 4397.890 197.965 4398.990 ;
        RECT 0.000 4386.890 200.000 4397.890 ;
        RECT 0.000 4385.895 197.965 4386.890 ;
        RECT 0.000 4374.895 200.000 4385.895 ;
        RECT 0.000 4373.795 197.965 4374.895 ;
        RECT 0.000 4349.240 179.800 4373.795 ;
      LAYER met3 ;
        RECT 180.200 4349.495 200.000 4373.395 ;
      LAYER met3 ;
        RECT 3386.690 4312.430 3588.000 4391.690 ;
        RECT 4.900 4187.990 162.840 4212.290 ;
      LAYER met3 ;
        RECT 163.240 4188.390 200.000 4212.290 ;
      LAYER met3 ;
        RECT 4.900 4186.890 197.965 4187.990 ;
        RECT 4.900 4175.890 200.000 4186.890 ;
        RECT 4.900 4174.895 197.965 4175.890 ;
        RECT 4.900 4163.895 200.000 4174.895 ;
        RECT 4.900 4162.795 197.965 4163.895 ;
        RECT 4.900 4138.240 167.085 4162.795 ;
      LAYER met3 ;
        RECT 167.485 4138.495 200.000 4162.395 ;
        RECT 3388.000 4142.605 3402.960 4166.505 ;
      LAYER met3 ;
        RECT 3403.360 4142.205 3588.000 4166.760 ;
        RECT 3390.035 4141.105 3588.000 4142.205 ;
        RECT 3388.000 4130.105 3588.000 4141.105 ;
        RECT 3390.035 4129.110 3588.000 4130.105 ;
        RECT 3388.000 4118.110 3588.000 4129.110 ;
        RECT 3390.035 4117.010 3588.000 4118.110 ;
      LAYER met3 ;
        RECT 3388.000 4092.710 3402.960 4116.610 ;
      LAYER met3 ;
        RECT 3403.360 4092.710 3588.000 4117.010 ;
      LAYER met3 ;
        RECT 3387.505 4092.050 3387.835 4092.065 ;
        RECT 3388.670 4092.050 3388.970 4092.710 ;
        RECT 3387.505 4091.750 3388.970 4092.050 ;
        RECT 3387.505 4091.735 3387.835 4091.750 ;
      LAYER met3 ;
        RECT 0.000 3922.310 201.310 4001.570 ;
        RECT 3386.690 3866.430 3588.000 3945.690 ;
        RECT 0.000 3706.310 201.310 3785.570 ;
        RECT 3386.690 3641.430 3588.000 3720.690 ;
        RECT 0.000 3490.310 201.310 3569.570 ;
        RECT 3386.690 3416.430 3588.000 3495.690 ;
        RECT 0.000 3274.310 201.310 3353.570 ;
        RECT 3386.690 3190.430 3588.000 3269.690 ;
        RECT 0.000 3058.310 201.310 3137.570 ;
        RECT 3386.690 2965.430 3588.000 3044.690 ;
        RECT 0.000 2842.310 201.310 2921.570 ;
        RECT 3386.690 2739.430 3588.000 2818.690 ;
        RECT 0.000 2626.310 201.310 2705.570 ;
      LAYER met3 ;
        RECT 3388.000 2569.605 3402.960 2593.505 ;
      LAYER met3 ;
        RECT 3403.360 2569.205 3588.000 2593.760 ;
        RECT 3390.035 2568.105 3588.000 2569.205 ;
        RECT 3388.000 2557.105 3588.000 2568.105 ;
        RECT 3390.035 2556.110 3588.000 2557.105 ;
        RECT 3388.000 2545.110 3588.000 2556.110 ;
        RECT 3390.035 2544.010 3588.000 2545.110 ;
      LAYER met3 ;
        RECT 3388.000 2519.710 3402.960 2543.610 ;
      LAYER met3 ;
        RECT 3403.360 2519.710 3588.000 2544.010 ;
      LAYER met3 ;
        RECT 3387.505 2519.210 3387.835 2519.225 ;
        RECT 3388.670 2519.210 3388.970 2519.710 ;
        RECT 3387.505 2518.910 3388.970 2519.210 ;
        RECT 3387.505 2518.895 3387.835 2518.910 ;
      LAYER met3 ;
        RECT 0.000 2464.990 184.640 2489.290 ;
      LAYER met3 ;
        RECT 185.040 2465.390 200.000 2489.290 ;
      LAYER met3 ;
        RECT 0.000 2463.890 197.965 2464.990 ;
        RECT 0.000 2452.890 200.000 2463.890 ;
        RECT 0.000 2451.895 197.965 2452.890 ;
        RECT 0.000 2440.895 200.000 2451.895 ;
        RECT 0.000 2439.795 197.965 2440.895 ;
        RECT 0.000 2415.240 184.640 2439.795 ;
      LAYER met3 ;
        RECT 185.040 2415.495 200.000 2439.395 ;
      LAYER met3 ;
        RECT 3429.550 2374.895 3434.200 2384.975 ;
        RECT 3390.035 2373.900 3587.965 2374.000 ;
        RECT 3430.000 2349.100 3587.965 2373.900 ;
        RECT 3390.035 2348.000 3587.965 2349.100 ;
        RECT 3390.000 2337.120 3587.965 2348.000 ;
        RECT 3390.035 2335.620 3587.965 2337.120 ;
        RECT 3390.000 2324.745 3587.965 2335.620 ;
        RECT 3390.035 2323.645 3587.965 2324.745 ;
      LAYER met3 ;
        RECT 3390.000 2299.300 3429.600 2323.245 ;
      LAYER met3 ;
        RECT 3430.000 2299.000 3587.965 2323.645 ;
        RECT 0.035 2280.200 24.250 2289.935 ;
        RECT 153.765 2279.605 158.415 2290.140 ;
        RECT 169.550 2280.200 174.200 2289.935 ;
        RECT 3413.800 2288.065 3418.450 2297.800 ;
        RECT 3429.585 2287.860 3434.235 2298.395 ;
        RECT 3563.750 2288.065 3587.965 2297.800 ;
        RECT 0.035 2254.355 158.000 2279.000 ;
      LAYER met3 ;
        RECT 158.400 2254.755 198.000 2278.700 ;
      LAYER met3 ;
        RECT 0.035 2253.255 197.965 2254.355 ;
        RECT 0.035 2242.380 198.000 2253.255 ;
        RECT 0.035 2240.880 197.965 2242.380 ;
        RECT 0.035 2230.000 198.000 2240.880 ;
        RECT 0.035 2228.900 197.965 2230.000 ;
        RECT 0.035 2204.100 158.000 2228.900 ;
        RECT 0.035 2204.000 197.965 2204.100 ;
        RECT 153.800 2193.025 158.450 2203.105 ;
      LAYER met3 ;
        RECT 3388.000 2128.605 3420.515 2152.505 ;
        RECT 3387.505 2128.210 3387.835 2128.225 ;
        RECT 3388.670 2128.210 3388.970 2128.605 ;
        RECT 3387.505 2127.910 3388.970 2128.210 ;
      LAYER met3 ;
        RECT 3420.915 2128.205 3583.100 2152.760 ;
      LAYER met3 ;
        RECT 3387.505 2127.895 3387.835 2127.910 ;
      LAYER met3 ;
        RECT 3390.035 2127.105 3583.100 2128.205 ;
        RECT 3388.000 2116.105 3583.100 2127.105 ;
        RECT 3390.035 2115.110 3583.100 2116.105 ;
        RECT 3388.000 2104.110 3583.100 2115.110 ;
        RECT 3390.035 2103.010 3583.100 2104.110 ;
      LAYER met3 ;
        RECT 3388.000 2078.710 3424.760 2102.610 ;
      LAYER met3 ;
        RECT 3425.160 2078.710 3583.100 2103.010 ;
        RECT 0.000 1988.310 201.310 2067.570 ;
        RECT 3386.690 1853.430 3588.000 1932.690 ;
        RECT 0.000 1772.310 201.310 1851.570 ;
        RECT 0.000 1556.310 201.310 1635.570 ;
        RECT 3386.690 1627.430 3588.000 1706.690 ;
        RECT 0.000 1340.310 201.310 1419.570 ;
        RECT 3386.690 1402.430 3588.000 1481.690 ;
        RECT 0.000 1124.310 201.310 1203.570 ;
        RECT 3386.690 1177.430 3588.000 1256.690 ;
        RECT 0.000 908.310 201.310 987.570 ;
        RECT 3386.690 951.430 3588.000 1030.690 ;
        RECT 3386.690 726.430 3588.000 805.690 ;
        RECT 0.000 600.990 179.800 625.290 ;
      LAYER met3 ;
        RECT 180.200 601.390 200.000 625.290 ;
      LAYER met3 ;
        RECT 0.000 599.890 197.965 600.990 ;
        RECT 0.000 588.890 200.000 599.890 ;
        RECT 0.000 587.895 197.965 588.890 ;
        RECT 0.000 576.895 200.000 587.895 ;
        RECT 0.000 575.795 197.965 576.895 ;
        RECT 0.000 551.240 179.800 575.795 ;
      LAYER met3 ;
        RECT 180.200 566.250 200.000 575.395 ;
        RECT 210.285 566.250 210.615 566.265 ;
        RECT 212.585 566.250 212.915 566.265 ;
        RECT 180.200 565.950 212.915 566.250 ;
        RECT 180.200 551.495 200.000 565.950 ;
        RECT 210.285 565.935 210.615 565.950 ;
        RECT 212.585 565.935 212.915 565.950 ;
      LAYER met3 ;
        RECT 3386.690 500.430 3588.000 579.690 ;
        RECT 153.765 415.605 158.415 426.140 ;
        RECT 159.805 415.440 163.270 426.140 ;
        RECT 4.395 390.355 190.700 415.000 ;
      LAYER met3 ;
        RECT 191.100 391.490 198.000 414.700 ;
        RECT 210.745 391.490 211.075 391.505 ;
        RECT 212.125 391.490 212.455 391.505 ;
        RECT 191.100 391.190 212.455 391.490 ;
        RECT 191.100 390.755 198.000 391.190 ;
        RECT 210.745 391.175 211.075 391.190 ;
        RECT 212.125 391.175 212.455 391.190 ;
      LAYER met3 ;
        RECT 4.395 389.255 197.965 390.355 ;
        RECT 4.395 378.380 198.000 389.255 ;
        RECT 4.395 376.880 197.965 378.380 ;
        RECT 4.395 366.000 198.000 376.880 ;
        RECT 4.395 364.900 197.965 366.000 ;
        RECT 4.395 340.490 190.700 364.900 ;
      LAYER met3 ;
        RECT 191.100 340.500 198.000 364.500 ;
        RECT 1198.365 207.210 1198.695 207.225 ;
        RECT 1262.765 207.210 1263.095 207.225 ;
        RECT 1198.365 206.910 1263.095 207.210 ;
        RECT 1198.365 206.895 1198.695 206.910 ;
        RECT 1262.765 206.895 1263.095 206.910 ;
        RECT 710.550 202.150 720.050 202.450 ;
        RECT 710.550 201.090 710.850 202.150 ;
        RECT 715.365 201.770 715.695 201.785 ;
        RECT 715.365 201.470 717.290 201.770 ;
        RECT 715.365 201.455 715.695 201.470 ;
        RECT 665.470 200.790 710.850 201.090 ;
        RECT 665.470 200.000 665.770 200.790 ;
        RECT 716.990 200.000 717.290 201.470 ;
        RECT 719.750 200.000 720.050 202.150 ;
        RECT 731.710 200.110 738.450 200.410 ;
        RECT 731.710 200.070 732.010 200.110 ;
        RECT 729.100 200.000 732.010 200.070 ;
        RECT 238.000 164.765 256.010 180.085 ;
        RECT 258.000 164.765 276.010 180.085 ;
        RECT 278.000 164.765 296.010 180.085 ;
        RECT 298.000 164.765 316.010 180.085 ;
        RECT 318.000 164.765 336.010 180.085 ;
        RECT 338.000 164.765 356.010 180.085 ;
        RECT 394.710 163.240 418.610 200.000 ;
      LAYER met3 ;
        RECT 420.110 197.965 431.110 200.000 ;
        RECT 432.105 197.965 443.105 200.000 ;
      LAYER met3 ;
        RECT 443.965 199.730 444.295 199.745 ;
        RECT 444.605 199.730 468.505 200.000 ;
        RECT 443.965 199.430 468.505 199.730 ;
        RECT 443.965 199.415 444.295 199.430 ;
      LAYER met3 ;
        RECT 419.010 167.085 444.205 197.965 ;
      LAYER met3 ;
        RECT 444.605 167.485 468.505 199.430 ;
      LAYER met3 ;
        RECT 419.010 162.840 468.760 167.085 ;
      LAYER met3 ;
        RECT 507.000 164.765 525.010 180.085 ;
        RECT 527.000 164.765 545.010 180.085 ;
        RECT 547.000 164.765 565.010 180.085 ;
        RECT 567.000 164.765 585.010 180.085 ;
        RECT 587.000 164.765 605.010 180.085 ;
        RECT 607.000 164.765 625.010 180.085 ;
      LAYER met3 ;
        RECT 394.710 4.900 468.760 162.840 ;
        RECT 663.300 151.080 664.340 199.375 ;
        RECT 663.300 133.400 663.675 151.080 ;
      LAYER met3 ;
        RECT 664.740 150.680 665.810 200.000 ;
        RECT 664.075 135.400 665.810 150.680 ;
      LAYER met3 ;
        RECT 666.210 188.690 707.935 199.375 ;
        RECT 709.465 193.730 716.375 199.375 ;
        RECT 709.465 192.265 714.910 193.730 ;
      LAYER met3 ;
        RECT 716.775 193.330 717.925 200.000 ;
      LAYER met3 ;
        RECT 709.465 191.985 714.630 192.265 ;
        RECT 709.465 190.555 713.550 191.985 ;
      LAYER met3 ;
        RECT 715.310 191.950 717.925 193.330 ;
        RECT 715.310 191.865 716.875 191.950 ;
        RECT 716.940 191.865 717.925 191.950 ;
      LAYER met3 ;
        RECT 718.325 196.465 718.690 199.375 ;
      LAYER met3 ;
        RECT 719.090 196.865 720.755 200.000 ;
        RECT 729.080 199.770 732.010 200.000 ;
      LAYER met3 ;
        RECT 721.155 196.465 728.680 199.375 ;
      LAYER met3 ;
        RECT 715.030 191.800 715.310 191.865 ;
        RECT 715.395 191.800 716.940 191.865 ;
        RECT 715.030 191.650 716.940 191.800 ;
        RECT 715.030 191.585 716.575 191.650 ;
        RECT 716.660 191.585 716.940 191.650 ;
      LAYER met3 ;
        RECT 709.765 190.255 713.550 190.555 ;
        RECT 666.210 184.830 708.700 188.690 ;
        RECT 710.230 187.335 713.550 190.255 ;
      LAYER met3 ;
        RECT 713.950 191.500 715.030 191.585 ;
        RECT 715.095 191.500 716.660 191.585 ;
        RECT 713.950 190.020 716.660 191.500 ;
      LAYER met3 ;
        RECT 718.325 191.465 728.680 196.465 ;
        RECT 717.340 191.185 728.680 191.465 ;
      LAYER met3 ;
        RECT 713.950 187.735 715.095 190.020 ;
      LAYER met3 ;
        RECT 717.060 189.620 728.680 191.185 ;
        RECT 715.495 187.335 728.680 189.620 ;
        RECT 710.230 184.830 728.680 187.335 ;
        RECT 666.210 183.015 728.680 184.830 ;
      LAYER met3 ;
        RECT 729.080 184.215 729.600 199.770 ;
        RECT 738.150 199.745 738.450 200.110 ;
        RECT 738.150 199.430 738.695 199.745 ;
        RECT 738.365 199.415 738.695 199.430 ;
      LAYER met3 ;
        RECT 730.000 184.615 737.035 199.375 ;
        RECT 730.210 184.405 737.035 184.615 ;
      LAYER met3 ;
        RECT 729.080 184.005 729.810 184.215 ;
        RECT 729.080 183.555 730.260 184.005 ;
      LAYER met3 ;
        RECT 730.660 183.955 737.035 184.405 ;
      LAYER met3 ;
        RECT 729.080 183.415 729.670 183.555 ;
        RECT 729.680 183.415 730.710 183.555 ;
      LAYER met3 ;
        RECT 731.110 183.505 737.035 183.955 ;
      LAYER met3 ;
        RECT 729.670 183.105 730.710 183.415 ;
      LAYER met3 ;
        RECT 666.210 182.555 729.270 183.015 ;
      LAYER met3 ;
        RECT 729.670 182.955 731.225 183.105 ;
      LAYER met3 ;
        RECT 666.210 181.980 729.730 182.555 ;
      LAYER met3 ;
        RECT 730.130 182.380 731.225 182.955 ;
      LAYER met3 ;
        RECT 666.210 169.105 730.305 181.980 ;
        RECT 666.210 168.520 729.720 169.105 ;
      LAYER met3 ;
        RECT 730.705 168.705 731.225 182.380 ;
      LAYER met3 ;
        RECT 666.210 167.805 729.005 168.520 ;
      LAYER met3 ;
        RECT 730.120 168.195 731.225 168.705 ;
        RECT 730.120 168.120 730.775 168.195 ;
        RECT 730.850 168.120 731.225 168.195 ;
        RECT 729.405 168.045 730.120 168.120 ;
        RECT 730.135 168.045 730.850 168.120 ;
      LAYER met3 ;
        RECT 666.210 167.220 728.420 167.805 ;
      LAYER met3 ;
        RECT 729.405 167.445 730.850 168.045 ;
      LAYER met3 ;
        RECT 731.625 167.720 737.035 183.505 ;
      LAYER met3 ;
        RECT 729.405 167.405 730.120 167.445 ;
        RECT 730.135 167.405 730.850 167.445 ;
        RECT 728.820 167.295 729.405 167.405 ;
        RECT 729.445 167.295 730.135 167.405 ;
      LAYER met3 ;
        RECT 666.210 167.005 728.205 167.220 ;
        RECT 666.210 165.475 715.325 167.005 ;
      LAYER met3 ;
        RECT 728.820 166.845 730.135 167.295 ;
      LAYER met3 ;
        RECT 731.250 167.005 737.035 167.720 ;
      LAYER met3 ;
        RECT 728.820 166.820 729.425 166.845 ;
        RECT 729.550 166.820 730.135 166.845 ;
        RECT 728.605 166.695 728.820 166.820 ;
        RECT 728.845 166.695 729.550 166.820 ;
        RECT 728.605 166.605 729.550 166.695 ;
        RECT 715.725 166.305 729.550 166.605 ;
      LAYER met3 ;
        RECT 730.535 166.420 737.035 167.005 ;
      LAYER met3 ;
        RECT 715.725 166.300 728.885 166.305 ;
        RECT 729.030 166.300 729.550 166.305 ;
        RECT 715.725 165.875 729.030 166.300 ;
      LAYER met3 ;
        RECT 729.950 165.900 737.035 166.420 ;
        RECT 729.430 165.475 737.035 165.900 ;
        RECT 666.210 135.800 737.035 165.475 ;
      LAYER met3 ;
        RECT 776.000 164.765 794.010 180.085 ;
        RECT 796.000 164.765 814.010 180.085 ;
        RECT 816.000 164.765 834.010 180.085 ;
        RECT 836.000 164.765 854.010 180.085 ;
        RECT 856.000 164.765 874.010 180.085 ;
        RECT 876.000 164.765 894.010 180.085 ;
        RECT 664.075 133.800 667.410 135.400 ;
      LAYER met3 ;
        RECT 667.810 134.200 737.035 135.800 ;
        RECT 663.300 131.800 665.410 133.400 ;
      LAYER met3 ;
        RECT 665.810 132.400 668.810 133.800 ;
      LAYER met3 ;
        RECT 669.210 132.800 737.035 134.200 ;
      LAYER met3 ;
        RECT 665.810 132.250 669.745 132.400 ;
        RECT 665.810 132.200 667.410 132.250 ;
        RECT 667.510 132.200 669.745 132.250 ;
      LAYER met3 ;
        RECT 663.300 130.515 667.010 131.800 ;
      LAYER met3 ;
        RECT 667.410 131.465 669.745 132.200 ;
      LAYER met3 ;
        RECT 670.145 131.865 737.035 132.800 ;
      LAYER met3 ;
        RECT 667.410 131.350 669.710 131.465 ;
        RECT 669.745 131.350 670.610 131.465 ;
        RECT 667.410 131.050 670.610 131.350 ;
        RECT 667.410 130.915 668.695 131.050 ;
        RECT 668.710 130.915 670.610 131.050 ;
      LAYER met3 ;
        RECT 671.010 131.000 737.035 131.865 ;
      LAYER met3 ;
        RECT 668.695 130.600 670.610 130.915 ;
      LAYER met3 ;
        RECT 663.300 129.565 668.295 130.515 ;
      LAYER met3 ;
        RECT 668.695 130.000 671.960 130.600 ;
        RECT 668.695 129.965 669.645 130.000 ;
        RECT 669.760 129.965 671.960 130.000 ;
      LAYER met3 ;
        RECT 663.300 128.600 669.245 129.565 ;
      LAYER met3 ;
        RECT 669.645 129.250 671.960 129.965 ;
      LAYER met3 ;
        RECT 672.360 129.650 737.035 131.000 ;
      LAYER met3 ;
        RECT 669.645 129.100 673.140 129.250 ;
        RECT 669.645 129.000 670.610 129.100 ;
        RECT 670.660 129.000 673.140 129.100 ;
      LAYER met3 ;
        RECT 663.300 127.390 670.210 128.600 ;
      LAYER met3 ;
        RECT 670.610 127.920 673.140 129.000 ;
        RECT 670.610 127.790 671.820 127.920 ;
        RECT 671.840 127.790 673.140 127.920 ;
        RECT 671.820 127.600 673.140 127.790 ;
      LAYER met3 ;
        RECT 663.300 127.200 671.420 127.390 ;
        RECT 663.300 104.955 671.610 127.200 ;
      LAYER met3 ;
        RECT 672.010 105.355 673.140 127.600 ;
      LAYER met3 ;
        RECT 673.540 104.955 737.035 129.650 ;
        RECT 663.300 0.000 737.035 104.955 ;
        RECT 932.430 0.000 1011.690 201.310 ;
      LAYER met3 ;
        RECT 1206.645 199.050 1206.975 199.065 ;
        RECT 1206.430 198.735 1206.975 199.050 ;
        RECT 1206.430 198.000 1206.730 198.735 ;
        RECT 1050.000 164.765 1068.010 180.085 ;
        RECT 1070.000 164.765 1088.010 180.085 ;
        RECT 1090.000 164.765 1108.010 180.085 ;
        RECT 1110.000 164.765 1128.010 180.085 ;
        RECT 1130.000 164.765 1148.010 180.085 ;
        RECT 1150.000 164.765 1168.010 180.085 ;
      LAYER met3 ;
        RECT 1194.860 159.805 1205.560 163.270 ;
        RECT 1194.860 153.765 1205.395 158.415 ;
      LAYER met3 ;
        RECT 1206.300 158.400 1230.245 198.000 ;
      LAYER met3 ;
        RECT 1231.745 197.965 1242.620 198.000 ;
        RECT 1244.120 197.965 1255.000 198.000 ;
        RECT 1230.645 158.000 1256.100 197.965 ;
      LAYER met3 ;
        RECT 1256.500 158.400 1280.500 198.000 ;
        RECT 1319.000 164.765 1337.010 180.085 ;
        RECT 1339.000 164.765 1357.010 180.085 ;
        RECT 1359.000 164.765 1377.010 180.085 ;
        RECT 1379.000 164.765 1397.010 180.085 ;
        RECT 1399.000 164.765 1417.010 180.085 ;
        RECT 1419.000 164.765 1437.010 180.085 ;
      LAYER met3 ;
        RECT 1206.000 4.395 1280.500 158.000 ;
        RECT 1475.430 0.000 1554.690 201.310 ;
      LAYER met3 ;
        RECT 1593.000 164.765 1611.010 180.085 ;
        RECT 1613.000 164.765 1631.010 180.085 ;
        RECT 1633.000 164.765 1651.010 180.085 ;
        RECT 1653.000 164.765 1671.010 180.085 ;
        RECT 1673.000 164.765 1691.010 180.085 ;
        RECT 1693.000 164.765 1711.010 180.085 ;
      LAYER met3 ;
        RECT 1749.430 0.000 1828.690 201.310 ;
      LAYER met3 ;
        RECT 1867.000 164.765 1885.010 180.085 ;
        RECT 1887.000 164.765 1905.010 180.085 ;
        RECT 1907.000 164.765 1925.010 180.085 ;
        RECT 1927.000 164.765 1945.010 180.085 ;
        RECT 1947.000 164.765 1965.010 180.085 ;
        RECT 1967.000 164.765 1985.010 180.085 ;
      LAYER met3 ;
        RECT 2023.430 0.000 2102.690 201.310 ;
      LAYER met3 ;
        RECT 2141.000 164.765 2159.010 180.085 ;
        RECT 2161.000 164.765 2179.010 180.085 ;
        RECT 2181.000 164.765 2199.010 180.085 ;
        RECT 2201.000 164.765 2219.010 180.085 ;
        RECT 2221.000 164.765 2239.010 180.085 ;
        RECT 2241.000 164.765 2259.010 180.085 ;
      LAYER met3 ;
        RECT 2297.430 0.000 2376.690 201.310 ;
      LAYER met3 ;
        RECT 2415.000 164.765 2433.010 180.085 ;
        RECT 2435.000 164.765 2453.010 180.085 ;
        RECT 2455.000 164.765 2473.010 180.085 ;
        RECT 2475.000 164.765 2493.010 180.085 ;
        RECT 2495.000 164.765 2513.010 180.085 ;
        RECT 2515.000 164.765 2533.010 180.085 ;
      LAYER met3 ;
        RECT 2571.430 0.000 2650.690 201.310 ;
      LAYER met3 ;
        RECT 2863.565 201.090 2863.895 201.105 ;
        RECT 2863.350 200.775 2863.895 201.090 ;
        RECT 2863.350 200.000 2863.650 200.775 ;
        RECT 2689.000 164.765 2707.010 180.085 ;
        RECT 2709.000 164.765 2727.010 180.085 ;
        RECT 2729.000 164.765 2747.010 180.085 ;
        RECT 2749.000 164.765 2767.010 180.085 ;
        RECT 2769.000 164.765 2787.010 180.085 ;
        RECT 2789.000 164.765 2807.010 180.085 ;
        RECT 2845.710 174.150 2869.610 200.000 ;
      LAYER met3 ;
        RECT 2871.110 197.965 2882.110 200.000 ;
        RECT 2883.105 197.965 2894.105 200.000 ;
        RECT 2870.010 173.750 2895.205 197.965 ;
      LAYER met3 ;
        RECT 2895.605 174.150 2919.505 200.000 ;
        RECT 3114.710 185.040 3138.610 200.000 ;
      LAYER met3 ;
        RECT 3140.110 197.965 3151.110 200.000 ;
        RECT 3152.105 197.965 3163.105 200.000 ;
        RECT 3139.010 184.640 3164.205 197.965 ;
      LAYER met3 ;
        RECT 3164.605 185.040 3188.505 200.000 ;
      LAYER met3 ;
        RECT 2845.710 0.000 2919.760 173.750 ;
      LAYER met3 ;
        RECT 2958.000 164.765 2976.010 180.085 ;
        RECT 2978.000 164.765 2996.010 180.085 ;
        RECT 2998.000 164.765 3016.010 180.085 ;
        RECT 3018.000 164.765 3036.010 180.085 ;
        RECT 3038.000 164.765 3056.010 180.085 ;
        RECT 3058.000 164.765 3076.010 180.085 ;
      LAYER met3 ;
        RECT 3114.710 0.000 3188.760 184.640 ;
      LAYER met3 ;
        RECT 3227.000 164.765 3245.010 180.085 ;
        RECT 3247.000 164.765 3265.010 180.085 ;
        RECT 3267.000 164.765 3285.010 180.085 ;
        RECT 3287.000 164.765 3305.010 180.085 ;
        RECT 3307.000 164.765 3325.010 180.085 ;
        RECT 3327.000 164.765 3345.010 180.085 ;
      LAYER via3 ;
        RECT 238.230 175.875 255.720 179.885 ;
        RECT 238.260 164.935 255.910 167.885 ;
        RECT 258.230 175.875 275.720 179.885 ;
        RECT 258.260 164.935 275.910 167.885 ;
        RECT 278.230 175.875 295.720 179.885 ;
        RECT 278.260 164.935 295.910 167.885 ;
        RECT 298.230 175.875 315.720 179.885 ;
        RECT 298.260 164.935 315.910 167.885 ;
        RECT 318.230 175.875 335.720 179.885 ;
        RECT 318.260 164.935 335.910 167.885 ;
        RECT 338.230 175.875 355.720 179.885 ;
        RECT 338.260 164.935 355.910 167.885 ;
        RECT 507.230 175.875 524.720 179.885 ;
        RECT 507.260 164.935 524.910 167.885 ;
        RECT 527.230 175.875 544.720 179.885 ;
        RECT 527.260 164.935 544.910 167.885 ;
        RECT 547.230 175.875 564.720 179.885 ;
        RECT 547.260 164.935 564.910 167.885 ;
        RECT 567.230 175.875 584.720 179.885 ;
        RECT 567.260 164.935 584.910 167.885 ;
        RECT 587.230 175.875 604.720 179.885 ;
        RECT 587.260 164.935 604.910 167.885 ;
        RECT 607.230 175.875 624.720 179.885 ;
        RECT 607.260 164.935 624.910 167.885 ;
        RECT 776.230 175.875 793.720 179.885 ;
        RECT 776.260 164.935 793.910 167.885 ;
        RECT 796.230 175.875 813.720 179.885 ;
        RECT 796.260 164.935 813.910 167.885 ;
        RECT 816.230 175.875 833.720 179.885 ;
        RECT 816.260 164.935 833.910 167.885 ;
        RECT 836.230 175.875 853.720 179.885 ;
        RECT 836.260 164.935 853.910 167.885 ;
        RECT 856.230 175.875 873.720 179.885 ;
        RECT 856.260 164.935 873.910 167.885 ;
        RECT 876.230 175.875 893.720 179.885 ;
        RECT 876.260 164.935 893.910 167.885 ;
        RECT 1050.230 175.875 1067.720 179.885 ;
        RECT 1050.260 164.935 1067.910 167.885 ;
        RECT 1070.230 175.875 1087.720 179.885 ;
        RECT 1070.260 164.935 1087.910 167.885 ;
        RECT 1090.230 175.875 1107.720 179.885 ;
        RECT 1090.260 164.935 1107.910 167.885 ;
        RECT 1110.230 175.875 1127.720 179.885 ;
        RECT 1110.260 164.935 1127.910 167.885 ;
        RECT 1130.230 175.875 1147.720 179.885 ;
        RECT 1130.260 164.935 1147.910 167.885 ;
        RECT 1150.230 175.875 1167.720 179.885 ;
        RECT 1150.260 164.935 1167.910 167.885 ;
        RECT 1319.230 175.875 1336.720 179.885 ;
        RECT 1319.260 164.935 1336.910 167.885 ;
        RECT 1339.230 175.875 1356.720 179.885 ;
        RECT 1339.260 164.935 1356.910 167.885 ;
        RECT 1359.230 175.875 1376.720 179.885 ;
        RECT 1359.260 164.935 1376.910 167.885 ;
        RECT 1379.230 175.875 1396.720 179.885 ;
        RECT 1379.260 164.935 1396.910 167.885 ;
        RECT 1399.230 175.875 1416.720 179.885 ;
        RECT 1399.260 164.935 1416.910 167.885 ;
        RECT 1419.230 175.875 1436.720 179.885 ;
        RECT 1419.260 164.935 1436.910 167.885 ;
        RECT 1593.230 175.875 1610.720 179.885 ;
        RECT 1593.260 164.935 1610.910 167.885 ;
        RECT 1613.230 175.875 1630.720 179.885 ;
        RECT 1613.260 164.935 1630.910 167.885 ;
        RECT 1633.230 175.875 1650.720 179.885 ;
        RECT 1633.260 164.935 1650.910 167.885 ;
        RECT 1653.230 175.875 1670.720 179.885 ;
        RECT 1653.260 164.935 1670.910 167.885 ;
        RECT 1673.230 175.875 1690.720 179.885 ;
        RECT 1673.260 164.935 1690.910 167.885 ;
        RECT 1693.230 175.875 1710.720 179.885 ;
        RECT 1693.260 164.935 1710.910 167.885 ;
        RECT 1867.230 175.875 1884.720 179.885 ;
        RECT 1867.260 164.935 1884.910 167.885 ;
        RECT 1887.230 175.875 1904.720 179.885 ;
        RECT 1887.260 164.935 1904.910 167.885 ;
        RECT 1907.230 175.875 1924.720 179.885 ;
        RECT 1907.260 164.935 1924.910 167.885 ;
        RECT 1927.230 175.875 1944.720 179.885 ;
        RECT 1927.260 164.935 1944.910 167.885 ;
        RECT 1947.230 175.875 1964.720 179.885 ;
        RECT 1947.260 164.935 1964.910 167.885 ;
        RECT 1967.230 175.875 1984.720 179.885 ;
        RECT 1967.260 164.935 1984.910 167.885 ;
        RECT 2141.230 175.875 2158.720 179.885 ;
        RECT 2141.260 164.935 2158.910 167.885 ;
        RECT 2161.230 175.875 2178.720 179.885 ;
        RECT 2161.260 164.935 2178.910 167.885 ;
        RECT 2181.230 175.875 2198.720 179.885 ;
        RECT 2181.260 164.935 2198.910 167.885 ;
        RECT 2201.230 175.875 2218.720 179.885 ;
        RECT 2201.260 164.935 2218.910 167.885 ;
        RECT 2221.230 175.875 2238.720 179.885 ;
        RECT 2221.260 164.935 2238.910 167.885 ;
        RECT 2241.230 175.875 2258.720 179.885 ;
        RECT 2241.260 164.935 2258.910 167.885 ;
        RECT 2415.230 175.875 2432.720 179.885 ;
        RECT 2415.260 164.935 2432.910 167.885 ;
        RECT 2435.230 175.875 2452.720 179.885 ;
        RECT 2435.260 164.935 2452.910 167.885 ;
        RECT 2455.230 175.875 2472.720 179.885 ;
        RECT 2455.260 164.935 2472.910 167.885 ;
        RECT 2475.230 175.875 2492.720 179.885 ;
        RECT 2475.260 164.935 2492.910 167.885 ;
        RECT 2495.230 175.875 2512.720 179.885 ;
        RECT 2495.260 164.935 2512.910 167.885 ;
        RECT 2515.230 175.875 2532.720 179.885 ;
        RECT 2515.260 164.935 2532.910 167.885 ;
        RECT 2689.230 175.875 2706.720 179.885 ;
        RECT 2689.260 164.935 2706.910 167.885 ;
        RECT 2709.230 175.875 2726.720 179.885 ;
        RECT 2709.260 164.935 2726.910 167.885 ;
        RECT 2729.230 175.875 2746.720 179.885 ;
        RECT 2729.260 164.935 2746.910 167.885 ;
        RECT 2749.230 175.875 2766.720 179.885 ;
        RECT 2749.260 164.935 2766.910 167.885 ;
        RECT 2769.230 175.875 2786.720 179.885 ;
        RECT 2769.260 164.935 2786.910 167.885 ;
        RECT 2789.230 175.875 2806.720 179.885 ;
        RECT 2958.230 175.875 2975.720 179.885 ;
        RECT 2789.260 164.935 2806.910 167.885 ;
        RECT 2958.260 164.935 2975.910 167.885 ;
        RECT 2978.230 175.875 2995.720 179.885 ;
        RECT 2978.260 164.935 2995.910 167.885 ;
        RECT 2998.230 175.875 3015.720 179.885 ;
        RECT 2998.260 164.935 3015.910 167.885 ;
        RECT 3018.230 175.875 3035.720 179.885 ;
        RECT 3018.260 164.935 3035.910 167.885 ;
        RECT 3038.230 175.875 3055.720 179.885 ;
        RECT 3038.260 164.935 3055.910 167.885 ;
        RECT 3058.230 175.875 3075.720 179.885 ;
        RECT 3058.260 164.935 3075.910 167.885 ;
        RECT 3227.230 175.875 3244.720 179.885 ;
        RECT 3227.260 164.935 3244.910 167.885 ;
        RECT 3247.230 175.875 3264.720 179.885 ;
        RECT 3247.260 164.935 3264.910 167.885 ;
        RECT 3267.230 175.875 3284.720 179.885 ;
        RECT 3267.260 164.935 3284.910 167.885 ;
        RECT 3287.230 175.875 3304.720 179.885 ;
        RECT 3287.260 164.935 3304.910 167.885 ;
        RECT 3307.230 175.875 3324.720 179.885 ;
        RECT 3307.260 164.935 3324.910 167.885 ;
        RECT 3327.230 175.875 3344.720 179.885 ;
        RECT 3327.260 164.935 3344.910 167.885 ;
      LAYER met4 ;
        RECT 0.000 5163.385 202.330 5188.000 ;
      LAYER met4 ;
        RECT 202.730 5163.785 204.000 5188.000 ;
      LAYER met4 ;
        RECT 0.000 5083.400 202.745 5163.385 ;
        RECT 204.000 5083.400 381.000 5188.000 ;
      LAYER met4 ;
        RECT 381.000 5163.785 382.270 5188.000 ;
      LAYER met4 ;
        RECT 382.670 5163.385 459.330 5188.000 ;
      LAYER met4 ;
        RECT 459.730 5163.785 461.000 5188.000 ;
      LAYER met4 ;
        RECT 381.965 5083.400 459.970 5163.385 ;
        RECT 461.000 5083.400 638.000 5188.000 ;
      LAYER met4 ;
        RECT 638.000 5163.785 639.270 5188.000 ;
      LAYER met4 ;
        RECT 639.670 5163.385 716.330 5188.000 ;
      LAYER met4 ;
        RECT 716.730 5163.785 718.000 5188.000 ;
      LAYER met4 ;
        RECT 638.965 5083.400 716.970 5163.385 ;
        RECT 718.000 5083.400 895.000 5188.000 ;
      LAYER met4 ;
        RECT 895.000 5163.785 896.270 5188.000 ;
      LAYER met4 ;
        RECT 896.670 5163.385 973.330 5188.000 ;
      LAYER met4 ;
        RECT 973.730 5163.785 975.000 5188.000 ;
      LAYER met4 ;
        RECT 895.965 5083.400 973.970 5163.385 ;
        RECT 975.000 5083.400 1152.000 5188.000 ;
      LAYER met4 ;
        RECT 1152.000 5163.785 1153.270 5188.000 ;
      LAYER met4 ;
        RECT 1153.670 5163.385 1230.330 5188.000 ;
      LAYER met4 ;
        RECT 1230.730 5163.785 1232.000 5188.000 ;
      LAYER met4 ;
        RECT 1152.965 5083.400 1230.970 5163.385 ;
        RECT 1232.000 5083.400 1410.000 5188.000 ;
      LAYER met4 ;
        RECT 1410.000 5163.785 1411.270 5188.000 ;
      LAYER met4 ;
        RECT 1411.670 5163.385 1488.330 5188.000 ;
      LAYER met4 ;
        RECT 1488.730 5163.785 1490.000 5188.000 ;
      LAYER met4 ;
        RECT 1410.965 5083.400 1488.970 5163.385 ;
        RECT 1490.000 5083.400 1667.000 5188.000 ;
      LAYER met4 ;
        RECT 1667.000 5163.785 1668.270 5188.000 ;
      LAYER met4 ;
        RECT 1668.670 5163.385 1740.330 5188.000 ;
      LAYER met4 ;
        RECT 1740.730 5163.785 1742.000 5188.000 ;
      LAYER met4 ;
        RECT 1742.000 5163.785 1919.000 5188.000 ;
      LAYER met4 ;
        RECT 1919.000 5163.785 1920.270 5188.000 ;
      LAYER met4 ;
        RECT 1667.965 5083.400 1741.035 5163.385 ;
        RECT 1747.000 5083.400 1919.000 5163.785 ;
        RECT 1920.670 5163.385 1997.330 5188.000 ;
      LAYER met4 ;
        RECT 1997.730 5163.785 1999.000 5188.000 ;
      LAYER met4 ;
        RECT 1919.965 5083.400 1997.970 5163.385 ;
        RECT 1999.000 5083.400 2364.000 5188.000 ;
      LAYER met4 ;
        RECT 2364.000 5163.785 2365.270 5188.000 ;
      LAYER met4 ;
        RECT 2365.670 5163.385 2442.330 5188.000 ;
      LAYER met4 ;
        RECT 2442.730 5163.785 2444.000 5188.000 ;
      LAYER met4 ;
        RECT 2364.965 5083.400 2442.970 5163.385 ;
        RECT 2444.000 5083.400 2621.000 5188.000 ;
      LAYER met4 ;
        RECT 2621.000 5163.785 2622.270 5188.000 ;
      LAYER met4 ;
        RECT 2622.670 5163.385 2699.330 5188.000 ;
      LAYER met4 ;
        RECT 2699.730 5163.785 2701.000 5188.000 ;
      LAYER met4 ;
        RECT 2621.965 5083.400 2699.970 5163.385 ;
        RECT 2701.000 5083.400 2878.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.000 5163.785 2879.270 5188.000 ;
      LAYER met4 ;
        RECT 2879.670 5163.385 2951.330 5188.000 ;
      LAYER met4 ;
        RECT 2951.730 5163.785 2953.000 5188.000 ;
      LAYER met4 ;
        RECT 2878.965 5083.400 2952.035 5163.385 ;
        RECT 2953.000 5083.400 3130.000 5188.000 ;
      LAYER met4 ;
        RECT 3130.000 5163.785 3131.270 5188.000 ;
      LAYER met4 ;
        RECT 3131.670 5163.385 3208.330 5188.000 ;
      LAYER met4 ;
        RECT 3208.730 5163.785 3210.000 5188.000 ;
      LAYER met4 ;
        RECT 3210.000 5163.385 3388.000 5188.000 ;
      LAYER met4 ;
        RECT 3388.000 5163.785 3389.435 5188.000 ;
      LAYER met4 ;
        RECT 3389.835 5163.385 3588.000 5188.000 ;
        RECT 3130.965 5083.400 3208.970 5163.385 ;
        RECT 3210.000 5083.400 3588.000 5163.385 ;
        RECT 0.000 5057.635 201.745 5083.400 ;
      LAYER met4 ;
        RECT 202.145 5058.035 382.270 5083.000 ;
      LAYER met4 ;
        RECT 382.670 5057.635 459.330 5083.400 ;
      LAYER met4 ;
        RECT 459.730 5058.035 639.270 5083.000 ;
      LAYER met4 ;
        RECT 639.670 5057.635 716.330 5083.400 ;
      LAYER met4 ;
        RECT 716.730 5058.035 896.270 5083.000 ;
      LAYER met4 ;
        RECT 896.670 5057.635 973.330 5083.400 ;
      LAYER met4 ;
        RECT 973.730 5058.035 1153.270 5083.000 ;
      LAYER met4 ;
        RECT 1153.670 5057.635 1230.330 5083.400 ;
      LAYER met4 ;
        RECT 1230.730 5058.035 1411.270 5083.000 ;
      LAYER met4 ;
        RECT 1411.670 5057.635 1488.330 5083.400 ;
      LAYER met4 ;
        RECT 1488.730 5058.035 1668.270 5083.000 ;
      LAYER met4 ;
        RECT 1668.670 5057.635 1740.330 5083.400 ;
      LAYER met4 ;
        RECT 1740.730 5058.035 1920.270 5083.000 ;
      LAYER met4 ;
        RECT 1920.670 5057.635 1997.330 5083.400 ;
      LAYER met4 ;
        RECT 1997.730 5058.035 2365.270 5083.000 ;
      LAYER met4 ;
        RECT 2365.670 5057.635 2442.330 5083.400 ;
      LAYER met4 ;
        RECT 2442.730 5058.035 2622.270 5083.000 ;
      LAYER met4 ;
        RECT 2622.670 5057.635 2699.330 5083.400 ;
      LAYER met4 ;
        RECT 2699.730 5058.035 2879.270 5083.000 ;
      LAYER met4 ;
        RECT 2879.670 5057.635 2951.330 5083.400 ;
      LAYER met4 ;
        RECT 2951.730 5058.035 3131.270 5083.000 ;
      LAYER met4 ;
        RECT 3131.670 5057.635 3208.330 5083.400 ;
      LAYER met4 ;
        RECT 3208.730 5058.035 3390.645 5083.000 ;
      LAYER met4 ;
        RECT 3391.045 5057.635 3588.000 5083.400 ;
        RECT 0.000 5056.935 202.745 5057.635 ;
        RECT 204.000 5056.935 381.000 5057.635 ;
        RECT 381.965 5056.935 459.970 5057.635 ;
        RECT 461.000 5056.935 638.000 5057.635 ;
        RECT 638.965 5056.935 716.970 5057.635 ;
        RECT 718.000 5056.935 895.000 5057.635 ;
        RECT 895.965 5056.935 973.970 5057.635 ;
        RECT 975.000 5056.935 1152.000 5057.635 ;
        RECT 1152.965 5056.935 1230.970 5057.635 ;
        RECT 1232.000 5056.935 1410.000 5057.635 ;
        RECT 1410.965 5056.935 1488.970 5057.635 ;
        RECT 1490.000 5056.935 1667.000 5057.635 ;
        RECT 1667.965 5056.935 1741.035 5057.635 ;
        RECT 1747.000 5056.935 1919.000 5057.635 ;
        RECT 1919.965 5056.935 1997.970 5057.635 ;
        RECT 1999.000 5056.935 2364.000 5057.635 ;
        RECT 2364.965 5056.935 2442.970 5057.635 ;
        RECT 2444.000 5056.935 2621.000 5057.635 ;
        RECT 2621.965 5056.935 2699.970 5057.635 ;
        RECT 2701.000 5056.935 2878.000 5057.635 ;
        RECT 2878.965 5056.935 2952.035 5057.635 ;
        RECT 2953.000 5056.935 3130.000 5057.635 ;
        RECT 3130.965 5056.935 3208.970 5057.635 ;
        RECT 3210.000 5056.935 3588.000 5057.635 ;
        RECT 0.000 5051.685 202.330 5056.935 ;
      LAYER met4 ;
        RECT 202.730 5052.085 382.270 5056.535 ;
      LAYER met4 ;
        RECT 382.670 5051.685 459.330 5056.935 ;
      LAYER met4 ;
        RECT 459.730 5052.085 639.270 5056.535 ;
      LAYER met4 ;
        RECT 639.670 5051.685 716.330 5056.935 ;
      LAYER met4 ;
        RECT 716.730 5052.085 896.270 5056.535 ;
      LAYER met4 ;
        RECT 896.670 5051.685 973.330 5056.935 ;
      LAYER met4 ;
        RECT 973.730 5052.085 1153.270 5056.535 ;
      LAYER met4 ;
        RECT 1153.670 5051.685 1230.330 5056.935 ;
      LAYER met4 ;
        RECT 1230.730 5052.085 1411.270 5056.535 ;
      LAYER met4 ;
        RECT 1411.670 5051.685 1488.330 5056.935 ;
      LAYER met4 ;
        RECT 1488.730 5052.085 1668.270 5056.535 ;
      LAYER met4 ;
        RECT 1668.670 5051.685 1740.330 5056.935 ;
      LAYER met4 ;
        RECT 1740.730 5052.085 1920.270 5056.535 ;
      LAYER met4 ;
        RECT 1920.670 5051.685 1997.330 5056.935 ;
      LAYER met4 ;
        RECT 1997.730 5052.085 2365.270 5056.535 ;
      LAYER met4 ;
        RECT 2365.670 5051.685 2442.330 5056.935 ;
      LAYER met4 ;
        RECT 2442.730 5052.085 2622.270 5056.535 ;
      LAYER met4 ;
        RECT 2622.670 5051.685 2699.330 5056.935 ;
      LAYER met4 ;
        RECT 2699.730 5052.085 2879.270 5056.535 ;
      LAYER met4 ;
        RECT 2879.670 5051.685 2951.330 5056.935 ;
      LAYER met4 ;
        RECT 2951.730 5052.085 3131.270 5056.535 ;
      LAYER met4 ;
        RECT 3131.670 5051.685 3208.330 5056.935 ;
      LAYER met4 ;
        RECT 3208.730 5052.085 3389.480 5056.535 ;
      LAYER met4 ;
        RECT 3389.880 5051.685 3588.000 5056.935 ;
        RECT 0.000 5051.085 202.745 5051.685 ;
        RECT 204.000 5051.085 381.000 5051.685 ;
        RECT 381.965 5051.085 459.970 5051.685 ;
        RECT 461.000 5051.085 638.000 5051.685 ;
        RECT 638.965 5051.085 716.970 5051.685 ;
        RECT 718.000 5051.085 895.000 5051.685 ;
        RECT 895.965 5051.085 973.970 5051.685 ;
        RECT 975.000 5051.085 1152.000 5051.685 ;
        RECT 1152.965 5051.085 1230.970 5051.685 ;
        RECT 1232.000 5051.085 1410.000 5051.685 ;
        RECT 1410.965 5051.085 1488.970 5051.685 ;
        RECT 1490.000 5051.085 1667.000 5051.685 ;
        RECT 1667.965 5051.085 1741.035 5051.685 ;
        RECT 1747.000 5051.085 1919.000 5051.685 ;
        RECT 1919.965 5051.085 1997.970 5051.685 ;
        RECT 1999.000 5051.085 2364.000 5051.685 ;
        RECT 2364.965 5051.085 2442.970 5051.685 ;
        RECT 2444.000 5051.085 2621.000 5051.685 ;
        RECT 2621.965 5051.085 2699.970 5051.685 ;
        RECT 2701.000 5051.085 2878.000 5051.685 ;
        RECT 2878.965 5051.085 2952.035 5051.685 ;
        RECT 2953.000 5051.085 3130.000 5051.685 ;
        RECT 3130.965 5051.085 3208.970 5051.685 ;
        RECT 3210.000 5051.085 3588.000 5051.685 ;
        RECT 0.000 5045.835 202.330 5051.085 ;
      LAYER met4 ;
        RECT 202.730 5046.235 382.270 5050.685 ;
      LAYER met4 ;
        RECT 382.670 5045.835 459.330 5051.085 ;
      LAYER met4 ;
        RECT 459.730 5046.235 639.270 5050.685 ;
      LAYER met4 ;
        RECT 639.670 5045.835 716.330 5051.085 ;
      LAYER met4 ;
        RECT 716.730 5046.235 896.270 5050.685 ;
      LAYER met4 ;
        RECT 896.670 5045.835 973.330 5051.085 ;
      LAYER met4 ;
        RECT 973.730 5046.235 1153.270 5050.685 ;
      LAYER met4 ;
        RECT 1153.670 5045.835 1230.330 5051.085 ;
      LAYER met4 ;
        RECT 1230.730 5046.235 1411.270 5050.685 ;
      LAYER met4 ;
        RECT 1411.670 5045.835 1488.330 5051.085 ;
      LAYER met4 ;
        RECT 1488.730 5046.235 1668.270 5050.685 ;
      LAYER met4 ;
        RECT 1668.670 5045.835 1740.330 5051.085 ;
      LAYER met4 ;
        RECT 1740.730 5046.235 1920.270 5050.685 ;
      LAYER met4 ;
        RECT 1920.670 5045.835 1997.330 5051.085 ;
      LAYER met4 ;
        RECT 1997.730 5046.235 2365.270 5050.685 ;
      LAYER met4 ;
        RECT 2365.670 5045.835 2442.330 5051.085 ;
      LAYER met4 ;
        RECT 2442.730 5046.235 2622.270 5050.685 ;
      LAYER met4 ;
        RECT 2622.670 5045.835 2699.330 5051.085 ;
      LAYER met4 ;
        RECT 2699.730 5046.235 2879.270 5050.685 ;
      LAYER met4 ;
        RECT 2879.670 5045.835 2951.330 5051.085 ;
      LAYER met4 ;
        RECT 2951.730 5046.235 3131.270 5050.685 ;
      LAYER met4 ;
        RECT 3131.670 5045.835 3208.330 5051.085 ;
      LAYER met4 ;
        RECT 3208.730 5046.235 3389.625 5050.685 ;
      LAYER met4 ;
        RECT 3390.025 5045.835 3588.000 5051.085 ;
        RECT 0.000 5045.135 202.745 5045.835 ;
        RECT 204.000 5045.135 381.000 5045.835 ;
        RECT 381.965 5045.135 459.970 5045.835 ;
        RECT 461.000 5045.135 638.000 5045.835 ;
        RECT 638.965 5045.135 716.970 5045.835 ;
        RECT 718.000 5045.135 895.000 5045.835 ;
        RECT 895.965 5045.135 973.970 5045.835 ;
        RECT 975.000 5045.135 1152.000 5045.835 ;
        RECT 1152.965 5045.135 1230.970 5045.835 ;
        RECT 1232.000 5045.135 1410.000 5045.835 ;
        RECT 1410.965 5045.135 1488.970 5045.835 ;
        RECT 1490.000 5045.135 1667.000 5045.835 ;
        RECT 1667.965 5045.135 1741.035 5045.835 ;
        RECT 1747.000 5045.135 1919.000 5045.835 ;
        RECT 1919.965 5045.135 1997.970 5045.835 ;
        RECT 1999.000 5045.135 2364.000 5045.835 ;
        RECT 2364.965 5045.135 2442.970 5045.835 ;
        RECT 2444.000 5045.135 2621.000 5045.835 ;
        RECT 2621.965 5045.135 2699.970 5045.835 ;
        RECT 2701.000 5045.135 2878.000 5045.835 ;
        RECT 2878.965 5045.135 2952.035 5045.835 ;
        RECT 2953.000 5045.135 3130.000 5045.835 ;
        RECT 3130.965 5045.135 3208.970 5045.835 ;
        RECT 3210.000 5045.135 3588.000 5045.835 ;
        RECT 0.000 5044.005 176.425 5045.135 ;
      LAYER met4 ;
        RECT 176.825 5044.405 383.610 5044.735 ;
      LAYER met4 ;
        RECT 384.010 5044.505 427.690 5045.135 ;
        RECT 0.000 5040.725 176.690 5044.005 ;
      LAYER met4 ;
        RECT 177.090 5041.125 417.440 5044.105 ;
      LAYER met4 ;
        RECT 0.000 5039.245 182.045 5040.725 ;
      LAYER met4 ;
        RECT 182.445 5039.645 204.000 5040.825 ;
      LAYER met4 ;
        RECT 204.000 5039.645 381.000 5040.825 ;
      LAYER met4 ;
        RECT 381.000 5039.645 382.270 5040.825 ;
      LAYER met4 ;
        RECT 417.840 5040.725 419.360 5044.505 ;
      LAYER met4 ;
        RECT 428.090 5044.405 640.610 5044.735 ;
      LAYER met4 ;
        RECT 641.010 5044.505 684.690 5045.135 ;
      LAYER met4 ;
        RECT 419.760 5041.125 674.440 5044.105 ;
      LAYER met4 ;
        RECT 382.670 5039.745 459.330 5040.725 ;
        RECT 0.000 5036.465 182.725 5039.245 ;
        RECT 0.000 5035.335 180.025 5036.465 ;
      LAYER met4 ;
        RECT 183.125 5036.365 433.145 5039.345 ;
      LAYER met4 ;
        RECT 433.545 5036.465 435.065 5039.745 ;
      LAYER met4 ;
        RECT 459.730 5039.645 461.000 5040.825 ;
      LAYER met4 ;
        RECT 461.000 5039.645 638.000 5040.825 ;
      LAYER met4 ;
        RECT 638.000 5039.645 639.270 5040.825 ;
      LAYER met4 ;
        RECT 674.840 5040.725 676.360 5044.505 ;
      LAYER met4 ;
        RECT 685.090 5044.405 897.610 5044.735 ;
      LAYER met4 ;
        RECT 898.010 5044.505 941.690 5045.135 ;
      LAYER met4 ;
        RECT 676.760 5041.125 931.440 5044.105 ;
      LAYER met4 ;
        RECT 639.670 5039.745 716.330 5040.725 ;
      LAYER met4 ;
        RECT 435.465 5036.365 690.145 5039.345 ;
      LAYER met4 ;
        RECT 690.545 5036.465 692.065 5039.745 ;
      LAYER met4 ;
        RECT 716.730 5039.645 718.000 5040.825 ;
      LAYER met4 ;
        RECT 718.000 5039.645 895.000 5040.825 ;
      LAYER met4 ;
        RECT 895.000 5039.645 896.270 5040.825 ;
      LAYER met4 ;
        RECT 931.840 5040.725 933.360 5044.505 ;
      LAYER met4 ;
        RECT 942.090 5044.405 1154.610 5044.735 ;
      LAYER met4 ;
        RECT 1155.010 5044.505 1198.690 5045.135 ;
      LAYER met4 ;
        RECT 933.760 5041.125 1188.440 5044.105 ;
      LAYER met4 ;
        RECT 896.670 5039.745 973.330 5040.725 ;
      LAYER met4 ;
        RECT 692.465 5036.365 947.145 5039.345 ;
      LAYER met4 ;
        RECT 947.545 5036.465 949.065 5039.745 ;
      LAYER met4 ;
        RECT 973.730 5039.645 975.000 5040.825 ;
      LAYER met4 ;
        RECT 975.000 5039.645 1152.000 5040.825 ;
      LAYER met4 ;
        RECT 1152.000 5039.645 1153.270 5040.825 ;
      LAYER met4 ;
        RECT 1188.840 5040.725 1190.360 5044.505 ;
      LAYER met4 ;
        RECT 1199.090 5044.405 1412.610 5044.735 ;
      LAYER met4 ;
        RECT 1413.010 5044.505 1456.690 5045.135 ;
      LAYER met4 ;
        RECT 1190.760 5041.125 1446.440 5044.105 ;
      LAYER met4 ;
        RECT 1153.670 5039.745 1230.330 5040.725 ;
      LAYER met4 ;
        RECT 949.465 5036.365 1204.145 5039.345 ;
      LAYER met4 ;
        RECT 1204.545 5036.465 1206.065 5039.745 ;
      LAYER met4 ;
        RECT 1230.730 5039.645 1232.000 5040.825 ;
      LAYER met4 ;
        RECT 1232.000 5039.645 1410.000 5040.825 ;
      LAYER met4 ;
        RECT 1410.000 5039.645 1411.270 5040.825 ;
      LAYER met4 ;
        RECT 1446.840 5040.725 1448.360 5044.505 ;
      LAYER met4 ;
        RECT 1457.090 5044.405 1742.000 5044.735 ;
        RECT 1747.000 5044.405 1921.610 5044.735 ;
      LAYER met4 ;
        RECT 1922.010 5044.505 1965.690 5045.135 ;
      LAYER met4 ;
        RECT 1448.760 5041.125 1955.440 5044.105 ;
      LAYER met4 ;
        RECT 1411.670 5039.745 1488.330 5040.725 ;
      LAYER met4 ;
        RECT 1206.465 5036.365 1462.145 5039.345 ;
      LAYER met4 ;
        RECT 1462.545 5036.465 1464.065 5039.745 ;
      LAYER met4 ;
        RECT 1488.730 5039.645 1490.000 5040.825 ;
      LAYER met4 ;
        RECT 1490.000 5039.645 1667.000 5040.825 ;
      LAYER met4 ;
        RECT 1667.000 5039.645 1668.270 5040.825 ;
      LAYER met4 ;
        RECT 1668.670 5039.745 1740.330 5040.725 ;
      LAYER met4 ;
        RECT 1740.730 5039.645 1742.000 5040.825 ;
      LAYER met4 ;
        RECT 1747.000 5039.645 1919.000 5040.825 ;
      LAYER met4 ;
        RECT 1919.000 5039.645 1920.270 5040.825 ;
      LAYER met4 ;
        RECT 1955.840 5040.725 1957.360 5044.505 ;
      LAYER met4 ;
        RECT 1966.090 5044.405 2366.610 5044.735 ;
      LAYER met4 ;
        RECT 2367.010 5044.505 2410.690 5045.135 ;
      LAYER met4 ;
        RECT 1957.760 5041.125 2400.440 5044.105 ;
      LAYER met4 ;
        RECT 1920.670 5039.745 1997.330 5040.725 ;
      LAYER met4 ;
        RECT 1464.465 5036.365 1971.145 5039.345 ;
      LAYER met4 ;
        RECT 1971.545 5036.465 1973.065 5039.745 ;
      LAYER met4 ;
        RECT 1997.730 5039.645 1999.000 5040.825 ;
      LAYER met4 ;
        RECT 1999.000 5039.645 2364.000 5040.825 ;
      LAYER met4 ;
        RECT 2364.000 5039.645 2365.270 5040.825 ;
      LAYER met4 ;
        RECT 2400.840 5040.725 2402.360 5044.505 ;
      LAYER met4 ;
        RECT 2411.090 5044.405 2623.610 5044.735 ;
      LAYER met4 ;
        RECT 2624.010 5044.505 2667.690 5045.135 ;
      LAYER met4 ;
        RECT 2402.760 5041.125 2657.440 5044.105 ;
      LAYER met4 ;
        RECT 2365.670 5039.745 2442.330 5040.725 ;
      LAYER met4 ;
        RECT 1973.465 5036.365 2416.145 5039.345 ;
      LAYER met4 ;
        RECT 2416.545 5036.465 2418.065 5039.745 ;
      LAYER met4 ;
        RECT 2442.730 5039.645 2444.000 5040.825 ;
      LAYER met4 ;
        RECT 2444.000 5039.645 2621.000 5040.825 ;
      LAYER met4 ;
        RECT 2621.000 5039.645 2622.270 5040.825 ;
      LAYER met4 ;
        RECT 2657.840 5040.725 2659.360 5044.505 ;
      LAYER met4 ;
        RECT 2668.090 5044.405 2879.270 5044.735 ;
      LAYER met4 ;
        RECT 2879.670 5044.505 2951.330 5045.135 ;
      LAYER met4 ;
        RECT 2951.730 5044.405 3132.610 5044.735 ;
      LAYER met4 ;
        RECT 3133.010 5044.505 3176.690 5045.135 ;
      LAYER met4 ;
        RECT 2659.760 5041.125 3166.440 5044.105 ;
      LAYER met4 ;
        RECT 2622.670 5039.745 2699.330 5040.725 ;
      LAYER met4 ;
        RECT 2418.465 5036.365 2673.145 5039.345 ;
      LAYER met4 ;
        RECT 2673.545 5036.465 2675.065 5039.745 ;
      LAYER met4 ;
        RECT 2699.730 5039.645 2701.000 5040.825 ;
      LAYER met4 ;
        RECT 2701.000 5039.645 2878.000 5040.825 ;
      LAYER met4 ;
        RECT 2878.000 5039.645 2879.270 5040.825 ;
      LAYER met4 ;
        RECT 2879.670 5039.745 2951.330 5040.725 ;
      LAYER met4 ;
        RECT 2951.730 5039.645 2953.000 5040.825 ;
      LAYER met4 ;
        RECT 2953.000 5039.645 3130.000 5040.825 ;
      LAYER met4 ;
        RECT 3130.000 5039.645 3131.270 5040.825 ;
      LAYER met4 ;
        RECT 3166.840 5040.725 3168.360 5044.505 ;
      LAYER met4 ;
        RECT 3177.090 5044.405 3411.175 5044.735 ;
        RECT 3168.760 5041.125 3410.910 5044.105 ;
      LAYER met4 ;
        RECT 3411.575 5044.005 3588.000 5045.135 ;
        RECT 3131.670 5039.745 3208.330 5040.725 ;
      LAYER met4 ;
        RECT 2675.465 5036.365 3182.145 5039.345 ;
      LAYER met4 ;
        RECT 3182.545 5036.465 3184.065 5039.745 ;
      LAYER met4 ;
        RECT 3208.730 5039.645 3210.000 5040.825 ;
      LAYER met4 ;
        RECT 3210.000 5039.645 3388.000 5040.825 ;
      LAYER met4 ;
        RECT 3388.000 5039.645 3409.550 5040.825 ;
      LAYER met4 ;
        RECT 3411.310 5040.725 3588.000 5044.005 ;
      LAYER met4 ;
        RECT 3184.465 5036.365 3408.935 5039.345 ;
      LAYER met4 ;
        RECT 3409.950 5039.245 3588.000 5040.725 ;
      LAYER met4 ;
        RECT 180.425 5035.735 383.610 5036.065 ;
      LAYER met4 ;
        RECT 384.010 5035.335 427.690 5035.965 ;
      LAYER met4 ;
        RECT 428.090 5035.735 640.610 5036.065 ;
      LAYER met4 ;
        RECT 641.010 5035.335 684.690 5035.965 ;
      LAYER met4 ;
        RECT 685.090 5035.735 897.610 5036.065 ;
      LAYER met4 ;
        RECT 898.010 5035.335 941.690 5035.965 ;
      LAYER met4 ;
        RECT 942.090 5035.735 1154.610 5036.065 ;
      LAYER met4 ;
        RECT 1155.010 5035.335 1198.690 5035.965 ;
      LAYER met4 ;
        RECT 1199.090 5035.735 1412.610 5036.065 ;
      LAYER met4 ;
        RECT 1413.010 5035.335 1456.690 5035.965 ;
      LAYER met4 ;
        RECT 1457.090 5035.735 1742.000 5036.065 ;
        RECT 1747.000 5035.735 1921.610 5036.065 ;
      LAYER met4 ;
        RECT 1922.010 5035.335 1965.690 5035.965 ;
      LAYER met4 ;
        RECT 1966.090 5035.735 2366.610 5036.065 ;
      LAYER met4 ;
        RECT 2367.010 5035.335 2410.690 5035.965 ;
      LAYER met4 ;
        RECT 2411.090 5035.735 2623.610 5036.065 ;
      LAYER met4 ;
        RECT 2624.010 5035.335 2667.690 5035.965 ;
      LAYER met4 ;
        RECT 2668.090 5035.735 2879.270 5036.065 ;
      LAYER met4 ;
        RECT 2879.670 5035.335 2951.330 5035.965 ;
      LAYER met4 ;
        RECT 2951.730 5035.735 3132.610 5036.065 ;
      LAYER met4 ;
        RECT 3133.010 5035.335 3176.690 5035.965 ;
      LAYER met4 ;
        RECT 3177.090 5035.735 3407.575 5036.065 ;
      LAYER met4 ;
        RECT 3409.335 5035.965 3588.000 5039.245 ;
        RECT 3407.975 5035.335 3588.000 5035.965 ;
        RECT 0.000 5034.635 202.745 5035.335 ;
        RECT 381.965 5034.635 459.970 5035.335 ;
        RECT 638.965 5034.635 716.970 5035.335 ;
        RECT 895.965 5034.635 973.970 5035.335 ;
        RECT 1152.965 5034.635 1230.970 5035.335 ;
        RECT 1410.965 5034.635 1488.970 5035.335 ;
        RECT 1667.965 5034.635 1741.035 5035.335 ;
        RECT 1919.965 5034.635 1997.970 5035.335 ;
        RECT 2364.965 5034.635 2442.970 5035.335 ;
        RECT 2621.965 5034.635 2699.970 5035.335 ;
        RECT 2878.965 5034.635 2952.035 5035.335 ;
        RECT 3130.965 5034.635 3208.970 5035.335 ;
        RECT 3388.000 5034.635 3588.000 5035.335 ;
        RECT 0.000 5029.185 202.330 5034.635 ;
      LAYER met4 ;
        RECT 202.730 5029.585 382.270 5034.235 ;
      LAYER met4 ;
        RECT 382.670 5029.185 459.330 5034.635 ;
      LAYER met4 ;
        RECT 459.730 5029.585 639.270 5034.235 ;
      LAYER met4 ;
        RECT 639.670 5029.185 716.330 5034.635 ;
      LAYER met4 ;
        RECT 716.730 5029.585 896.270 5034.235 ;
      LAYER met4 ;
        RECT 896.670 5029.185 973.330 5034.635 ;
      LAYER met4 ;
        RECT 973.730 5029.585 1153.270 5034.235 ;
      LAYER met4 ;
        RECT 1153.670 5029.185 1230.330 5034.635 ;
      LAYER met4 ;
        RECT 1230.730 5029.585 1411.270 5034.235 ;
      LAYER met4 ;
        RECT 1411.670 5029.185 1488.330 5034.635 ;
      LAYER met4 ;
        RECT 1488.730 5029.585 1668.270 5034.235 ;
      LAYER met4 ;
        RECT 1668.670 5029.185 1740.330 5034.635 ;
      LAYER met4 ;
        RECT 1740.730 5029.585 1747.000 5034.235 ;
        RECT 1752.000 5029.585 1920.270 5034.235 ;
      LAYER met4 ;
        RECT 1920.670 5029.185 1997.330 5034.635 ;
      LAYER met4 ;
        RECT 1997.730 5029.585 2365.270 5034.235 ;
      LAYER met4 ;
        RECT 2365.670 5029.185 2442.330 5034.635 ;
      LAYER met4 ;
        RECT 2442.730 5029.585 2622.270 5034.235 ;
      LAYER met4 ;
        RECT 2622.670 5029.185 2699.330 5034.635 ;
      LAYER met4 ;
        RECT 2699.730 5029.585 2879.270 5034.235 ;
      LAYER met4 ;
        RECT 2879.670 5029.185 2951.330 5034.635 ;
      LAYER met4 ;
        RECT 2951.730 5029.585 3131.270 5034.235 ;
      LAYER met4 ;
        RECT 3131.670 5029.185 3208.330 5034.635 ;
      LAYER met4 ;
        RECT 3208.730 5029.585 3389.475 5034.235 ;
      LAYER met4 ;
        RECT 3389.875 5029.185 3588.000 5034.635 ;
        RECT 0.000 5028.585 202.745 5029.185 ;
        RECT 381.965 5028.585 459.970 5029.185 ;
        RECT 638.965 5028.585 716.970 5029.185 ;
        RECT 895.965 5028.585 973.970 5029.185 ;
        RECT 1152.965 5028.585 1230.970 5029.185 ;
        RECT 1410.965 5028.585 1488.970 5029.185 ;
        RECT 1667.965 5028.585 1741.035 5029.185 ;
        RECT 1919.965 5028.585 1997.970 5029.185 ;
        RECT 2364.965 5028.585 2442.970 5029.185 ;
        RECT 2621.965 5028.585 2699.970 5029.185 ;
        RECT 2878.965 5028.585 2952.035 5029.185 ;
        RECT 3130.965 5028.585 3208.970 5029.185 ;
        RECT 3388.000 5028.585 3588.000 5029.185 ;
        RECT 0.000 5024.335 202.330 5028.585 ;
      LAYER met4 ;
        RECT 202.730 5024.735 382.270 5028.185 ;
      LAYER met4 ;
        RECT 382.670 5024.335 459.330 5028.585 ;
      LAYER met4 ;
        RECT 459.730 5024.735 639.270 5028.185 ;
      LAYER met4 ;
        RECT 639.670 5024.335 716.330 5028.585 ;
      LAYER met4 ;
        RECT 716.730 5024.735 896.270 5028.185 ;
      LAYER met4 ;
        RECT 896.670 5024.335 973.330 5028.585 ;
      LAYER met4 ;
        RECT 973.730 5024.735 1153.270 5028.185 ;
      LAYER met4 ;
        RECT 1153.670 5024.335 1230.330 5028.585 ;
      LAYER met4 ;
        RECT 1230.730 5024.735 1411.270 5028.185 ;
      LAYER met4 ;
        RECT 1411.670 5024.335 1488.330 5028.585 ;
      LAYER met4 ;
        RECT 1488.730 5024.735 1668.270 5028.185 ;
      LAYER met4 ;
        RECT 1668.670 5024.335 1740.330 5028.585 ;
      LAYER met4 ;
        RECT 1740.730 5024.735 1742.000 5028.185 ;
        RECT 1747.000 5024.735 1920.270 5028.185 ;
      LAYER met4 ;
        RECT 1920.670 5024.335 1997.330 5028.585 ;
      LAYER met4 ;
        RECT 1997.730 5024.735 2365.270 5028.185 ;
      LAYER met4 ;
        RECT 2365.670 5024.335 2442.330 5028.585 ;
      LAYER met4 ;
        RECT 2442.730 5024.735 2622.270 5028.185 ;
      LAYER met4 ;
        RECT 2622.670 5024.335 2699.330 5028.585 ;
      LAYER met4 ;
        RECT 2699.730 5024.735 2879.270 5028.185 ;
      LAYER met4 ;
        RECT 2879.670 5024.335 2951.330 5028.585 ;
      LAYER met4 ;
        RECT 2951.730 5024.735 3131.270 5028.185 ;
      LAYER met4 ;
        RECT 3131.670 5024.335 3208.330 5028.585 ;
      LAYER met4 ;
        RECT 3208.730 5024.735 3389.335 5028.185 ;
      LAYER met4 ;
        RECT 3389.735 5024.335 3588.000 5028.585 ;
        RECT 0.000 5023.735 202.745 5024.335 ;
        RECT 381.965 5023.735 459.970 5024.335 ;
        RECT 638.965 5023.735 716.970 5024.335 ;
        RECT 895.965 5023.735 973.970 5024.335 ;
        RECT 1152.965 5023.735 1230.970 5024.335 ;
        RECT 1410.965 5023.735 1488.970 5024.335 ;
        RECT 1667.965 5023.735 1741.035 5024.335 ;
        RECT 1919.965 5023.735 1997.970 5024.335 ;
        RECT 2364.965 5023.735 2442.970 5024.335 ;
        RECT 2621.965 5023.735 2699.970 5024.335 ;
        RECT 2878.965 5023.735 2952.035 5024.335 ;
        RECT 3130.965 5023.735 3208.970 5024.335 ;
        RECT 3388.000 5023.735 3588.000 5024.335 ;
        RECT 0.000 5019.485 202.330 5023.735 ;
      LAYER met4 ;
        RECT 202.730 5019.885 382.270 5023.335 ;
      LAYER met4 ;
        RECT 382.670 5019.485 459.330 5023.735 ;
      LAYER met4 ;
        RECT 459.730 5019.885 639.270 5023.335 ;
      LAYER met4 ;
        RECT 639.670 5019.485 716.330 5023.735 ;
      LAYER met4 ;
        RECT 716.730 5019.885 896.270 5023.335 ;
      LAYER met4 ;
        RECT 896.670 5019.485 973.330 5023.735 ;
      LAYER met4 ;
        RECT 973.730 5019.885 1153.270 5023.335 ;
      LAYER met4 ;
        RECT 1153.670 5019.485 1230.330 5023.735 ;
      LAYER met4 ;
        RECT 1230.730 5019.885 1411.270 5023.335 ;
      LAYER met4 ;
        RECT 1411.670 5019.485 1488.330 5023.735 ;
      LAYER met4 ;
        RECT 1488.730 5019.885 1668.270 5023.335 ;
      LAYER met4 ;
        RECT 1668.670 5019.485 1740.330 5023.735 ;
      LAYER met4 ;
        RECT 1740.730 5019.885 1920.270 5023.335 ;
      LAYER met4 ;
        RECT 1920.670 5019.485 1997.330 5023.735 ;
      LAYER met4 ;
        RECT 1997.730 5019.885 2365.270 5023.335 ;
      LAYER met4 ;
        RECT 2365.670 5019.485 2442.330 5023.735 ;
      LAYER met4 ;
        RECT 2442.730 5019.885 2622.270 5023.335 ;
      LAYER met4 ;
        RECT 2622.670 5019.485 2699.330 5023.735 ;
      LAYER met4 ;
        RECT 2699.730 5019.885 2879.270 5023.335 ;
      LAYER met4 ;
        RECT 2879.670 5019.485 2951.330 5023.735 ;
      LAYER met4 ;
        RECT 2951.730 5019.885 3131.270 5023.335 ;
      LAYER met4 ;
        RECT 3131.670 5019.485 3208.330 5023.735 ;
      LAYER met4 ;
        RECT 3208.730 5019.885 3389.385 5023.335 ;
      LAYER met4 ;
        RECT 3389.785 5019.485 3588.000 5023.735 ;
        RECT 0.000 5018.885 202.745 5019.485 ;
        RECT 381.965 5018.885 459.970 5019.485 ;
        RECT 638.965 5018.885 716.970 5019.485 ;
        RECT 895.965 5018.885 973.970 5019.485 ;
        RECT 1152.965 5018.885 1230.970 5019.485 ;
        RECT 1410.965 5018.885 1488.970 5019.485 ;
        RECT 1667.965 5018.885 1741.035 5019.485 ;
        RECT 1919.965 5018.885 1997.970 5019.485 ;
        RECT 2364.965 5018.885 2442.970 5019.485 ;
        RECT 2621.965 5018.885 2699.970 5019.485 ;
        RECT 2878.965 5018.885 2952.035 5019.485 ;
        RECT 3130.965 5018.885 3208.970 5019.485 ;
        RECT 3388.000 5018.885 3588.000 5019.485 ;
        RECT 0.000 5013.435 202.330 5018.885 ;
      LAYER met4 ;
        RECT 202.730 5013.835 382.270 5018.485 ;
      LAYER met4 ;
        RECT 382.670 5013.435 459.330 5018.885 ;
      LAYER met4 ;
        RECT 459.730 5013.835 639.270 5018.485 ;
      LAYER met4 ;
        RECT 639.670 5013.435 716.330 5018.885 ;
      LAYER met4 ;
        RECT 716.730 5013.835 896.270 5018.485 ;
      LAYER met4 ;
        RECT 896.670 5013.435 973.330 5018.885 ;
      LAYER met4 ;
        RECT 973.730 5013.835 1153.270 5018.485 ;
      LAYER met4 ;
        RECT 1153.670 5013.435 1230.330 5018.885 ;
      LAYER met4 ;
        RECT 1230.730 5013.835 1411.270 5018.485 ;
      LAYER met4 ;
        RECT 1411.670 5013.435 1488.330 5018.885 ;
      LAYER met4 ;
        RECT 1488.730 5013.835 1668.270 5018.485 ;
      LAYER met4 ;
        RECT 1668.670 5013.435 1740.330 5018.885 ;
      LAYER met4 ;
        RECT 1740.730 5013.835 1920.270 5018.485 ;
      LAYER met4 ;
        RECT 1920.670 5013.435 1997.330 5018.885 ;
      LAYER met4 ;
        RECT 1997.730 5013.835 2365.270 5018.485 ;
      LAYER met4 ;
        RECT 2365.670 5013.435 2442.330 5018.885 ;
      LAYER met4 ;
        RECT 2442.730 5013.835 2622.270 5018.485 ;
      LAYER met4 ;
        RECT 2622.670 5013.435 2699.330 5018.885 ;
      LAYER met4 ;
        RECT 2699.730 5013.835 2879.270 5018.485 ;
      LAYER met4 ;
        RECT 2879.670 5013.435 2951.330 5018.885 ;
      LAYER met4 ;
        RECT 2951.730 5013.835 3131.270 5018.485 ;
      LAYER met4 ;
        RECT 3131.670 5013.435 3208.330 5018.885 ;
      LAYER met4 ;
        RECT 3208.730 5013.835 3389.600 5018.485 ;
      LAYER met4 ;
        RECT 3390.000 5013.435 3588.000 5018.885 ;
        RECT 0.000 5012.835 202.745 5013.435 ;
        RECT 381.965 5012.835 459.970 5013.435 ;
        RECT 638.965 5012.835 716.970 5013.435 ;
        RECT 895.965 5012.835 973.970 5013.435 ;
        RECT 1152.965 5012.835 1230.970 5013.435 ;
        RECT 1410.965 5012.835 1488.970 5013.435 ;
        RECT 1667.965 5012.835 1741.035 5013.435 ;
        RECT 1919.965 5012.835 1997.970 5013.435 ;
        RECT 2364.965 5012.835 2442.970 5013.435 ;
        RECT 2621.965 5012.835 2699.970 5013.435 ;
        RECT 2878.965 5012.835 2952.035 5013.435 ;
        RECT 3130.965 5012.835 3208.970 5013.435 ;
        RECT 3388.000 5012.835 3588.000 5013.435 ;
        RECT 0.000 5011.575 202.330 5012.835 ;
        RECT 0.000 4991.045 142.865 5011.575 ;
        RECT 143.995 5011.310 202.330 5011.575 ;
        RECT 0.000 4989.835 104.600 4991.045 ;
      LAYER met4 ;
        RECT 0.000 4988.000 24.215 4989.435 ;
      LAYER met4 ;
        RECT 24.615 4988.000 104.600 4989.835 ;
        RECT 0.000 4851.000 104.600 4988.000 ;
      LAYER met4 ;
        RECT 0.000 4849.730 24.215 4851.000 ;
      LAYER met4 ;
        RECT 24.615 4849.330 104.600 4849.970 ;
      LAYER met4 ;
        RECT 105.000 4849.730 129.965 4990.645 ;
      LAYER met4 ;
        RECT 130.365 4990.025 142.865 4991.045 ;
        RECT 130.365 4989.880 136.915 4990.025 ;
        RECT 130.365 4851.000 131.065 4989.880 ;
        RECT 130.365 4849.330 131.065 4849.970 ;
      LAYER met4 ;
        RECT 131.465 4849.730 135.915 4989.480 ;
      LAYER met4 ;
        RECT 136.315 4851.000 136.915 4989.880 ;
        RECT 136.315 4849.330 136.915 4849.970 ;
      LAYER met4 ;
        RECT 137.315 4849.730 141.765 4989.625 ;
      LAYER met4 ;
        RECT 142.165 4851.000 142.865 4990.025 ;
        RECT 142.165 4849.330 142.865 4849.970 ;
        RECT 0.000 4817.690 142.865 4849.330 ;
      LAYER met4 ;
        RECT 143.265 4818.090 143.595 5011.175 ;
      LAYER met4 ;
        RECT 0.000 4809.360 143.495 4817.690 ;
      LAYER met4 ;
        RECT 143.895 4809.760 146.875 5010.910 ;
      LAYER met4 ;
        RECT 147.275 5009.950 202.330 5011.310 ;
      LAYER met4 ;
        RECT 147.175 4988.000 148.355 5009.550 ;
      LAYER met4 ;
        RECT 148.755 5009.335 202.330 5009.950 ;
        RECT 147.175 4851.000 148.355 4988.000 ;
      LAYER met4 ;
        RECT 147.175 4849.730 148.355 4851.000 ;
      LAYER met4 ;
        RECT 147.275 4825.065 148.255 4849.330 ;
      LAYER met4 ;
        RECT 148.655 4825.465 151.635 5008.935 ;
      LAYER met4 ;
        RECT 152.035 5007.975 202.330 5009.335 ;
        RECT 147.275 4823.545 151.535 4825.065 ;
        RECT 147.275 4809.360 148.255 4823.545 ;
        RECT 0.000 4807.840 148.255 4809.360 ;
        RECT 0.000 4774.010 143.495 4807.840 ;
        RECT 0.000 4772.670 142.865 4774.010 ;
      LAYER met4 ;
        RECT 0.000 4771.000 24.215 4772.270 ;
      LAYER met4 ;
        RECT 24.615 4771.965 104.600 4772.670 ;
        RECT 0.000 4635.000 104.600 4771.000 ;
      LAYER met4 ;
        RECT 0.000 4633.730 24.215 4635.000 ;
      LAYER met4 ;
        RECT 24.215 4634.785 24.250 4635.000 ;
        RECT 24.615 4633.330 104.600 4635.000 ;
      LAYER met4 ;
        RECT 105.000 4633.730 129.965 4772.270 ;
      LAYER met4 ;
        RECT 130.365 4771.965 131.065 4772.670 ;
        RECT 130.365 4633.330 131.065 4771.000 ;
      LAYER met4 ;
        RECT 131.465 4633.730 135.915 4772.270 ;
      LAYER met4 ;
        RECT 136.315 4771.965 136.915 4772.670 ;
        RECT 136.315 4633.330 136.915 4771.000 ;
      LAYER met4 ;
        RECT 137.315 4633.730 141.765 4772.270 ;
      LAYER met4 ;
        RECT 142.165 4771.965 142.865 4772.670 ;
        RECT 142.165 4633.330 142.865 4771.000 ;
        RECT 0.000 4561.670 142.865 4633.330 ;
      LAYER met4 ;
        RECT 0.000 4560.000 24.215 4561.270 ;
      LAYER met4 ;
        RECT 24.615 4560.000 104.600 4561.670 ;
        RECT 0.000 4424.000 104.600 4560.000 ;
      LAYER met4 ;
        RECT 0.000 4422.730 24.215 4424.000 ;
      LAYER met4 ;
        RECT 24.615 4422.330 104.600 4423.035 ;
      LAYER met4 ;
        RECT 105.000 4422.730 129.965 4561.270 ;
      LAYER met4 ;
        RECT 130.365 4424.000 131.065 4561.670 ;
        RECT 130.365 4422.330 131.065 4423.035 ;
      LAYER met4 ;
        RECT 131.465 4422.730 135.915 4561.270 ;
      LAYER met4 ;
        RECT 136.315 4424.000 136.915 4561.670 ;
        RECT 136.315 4422.330 136.915 4423.035 ;
      LAYER met4 ;
        RECT 137.315 4422.730 141.765 4561.270 ;
      LAYER met4 ;
        RECT 142.165 4424.000 142.865 4561.670 ;
        RECT 142.165 4422.330 142.865 4423.035 ;
        RECT 0.000 4350.670 142.865 4422.330 ;
      LAYER met4 ;
        RECT 0.000 4349.000 24.215 4350.270 ;
      LAYER met4 ;
        RECT 24.615 4349.965 104.600 4350.670 ;
        RECT 0.000 4213.000 104.600 4349.000 ;
      LAYER met4 ;
        RECT 0.000 4211.730 24.215 4213.000 ;
      LAYER met4 ;
        RECT 24.615 4211.330 104.600 4212.035 ;
      LAYER met4 ;
        RECT 105.000 4211.730 129.965 4350.270 ;
      LAYER met4 ;
        RECT 130.365 4349.965 131.065 4350.670 ;
        RECT 130.365 4213.000 131.065 4349.000 ;
        RECT 130.365 4211.330 131.065 4212.035 ;
      LAYER met4 ;
        RECT 131.465 4211.730 135.915 4350.270 ;
      LAYER met4 ;
        RECT 136.315 4349.965 136.915 4350.670 ;
        RECT 136.315 4213.000 136.915 4349.000 ;
        RECT 136.315 4211.330 136.915 4212.035 ;
      LAYER met4 ;
        RECT 137.315 4211.730 141.765 4350.270 ;
      LAYER met4 ;
        RECT 142.165 4349.965 142.865 4350.670 ;
        RECT 142.165 4213.000 142.865 4349.000 ;
        RECT 142.165 4211.330 142.865 4212.035 ;
      LAYER met4 ;
        RECT 143.265 4211.730 143.595 4773.610 ;
      LAYER met4 ;
        RECT 0.000 4139.670 143.495 4211.330 ;
      LAYER met4 ;
        RECT 0.000 4138.000 24.215 4139.270 ;
      LAYER met4 ;
        RECT 24.615 4138.965 104.600 4139.670 ;
        RECT 0.000 4002.000 104.600 4138.000 ;
      LAYER met4 ;
        RECT 0.000 4000.730 24.215 4002.000 ;
      LAYER met4 ;
        RECT 24.615 4000.330 104.600 4000.970 ;
      LAYER met4 ;
        RECT 105.000 4000.730 129.965 4139.270 ;
      LAYER met4 ;
        RECT 130.365 4138.965 131.065 4139.670 ;
        RECT 130.365 4002.000 131.065 4138.000 ;
        RECT 130.365 4000.330 131.065 4000.970 ;
      LAYER met4 ;
        RECT 131.465 4000.730 135.915 4139.270 ;
      LAYER met4 ;
        RECT 136.315 4138.965 136.915 4139.670 ;
        RECT 136.315 4002.000 136.915 4138.000 ;
        RECT 136.315 4000.330 136.915 4000.970 ;
      LAYER met4 ;
        RECT 137.315 4000.730 141.765 4139.270 ;
      LAYER met4 ;
        RECT 142.165 4138.965 142.865 4139.670 ;
        RECT 142.165 4002.000 142.865 4138.000 ;
        RECT 142.165 4000.330 142.865 4000.970 ;
        RECT 0.000 3968.690 142.865 4000.330 ;
      LAYER met4 ;
        RECT 143.265 3969.090 143.595 4139.270 ;
      LAYER met4 ;
        RECT 0.000 3960.360 143.495 3968.690 ;
      LAYER met4 ;
        RECT 143.895 3960.760 146.875 4807.440 ;
      LAYER met4 ;
        RECT 147.275 4772.670 148.255 4807.840 ;
      LAYER met4 ;
        RECT 147.175 4771.000 148.355 4772.270 ;
      LAYER met4 ;
        RECT 147.175 4635.000 148.355 4771.000 ;
      LAYER met4 ;
        RECT 147.175 4633.730 148.355 4635.000 ;
      LAYER met4 ;
        RECT 147.275 4561.670 148.255 4633.330 ;
      LAYER met4 ;
        RECT 147.175 4560.000 148.355 4561.270 ;
      LAYER met4 ;
        RECT 147.175 4424.000 148.355 4560.000 ;
      LAYER met4 ;
        RECT 147.175 4422.730 148.355 4424.000 ;
      LAYER met4 ;
        RECT 147.275 4350.670 148.255 4422.330 ;
      LAYER met4 ;
        RECT 147.175 4349.000 148.355 4350.270 ;
      LAYER met4 ;
        RECT 147.175 4213.000 148.355 4349.000 ;
      LAYER met4 ;
        RECT 147.175 4211.730 148.355 4213.000 ;
      LAYER met4 ;
        RECT 147.275 4139.670 148.255 4211.330 ;
      LAYER met4 ;
        RECT 147.175 4138.000 148.355 4139.270 ;
      LAYER met4 ;
        RECT 147.175 4002.000 148.355 4138.000 ;
      LAYER met4 ;
        RECT 147.175 4000.730 148.355 4002.000 ;
      LAYER met4 ;
        RECT 147.275 3976.065 148.255 4000.330 ;
      LAYER met4 ;
        RECT 148.655 3976.465 151.635 4823.145 ;
        RECT 151.935 4818.090 152.265 5007.575 ;
      LAYER met4 ;
        RECT 152.665 5007.385 202.330 5007.975 ;
      LAYER met4 ;
        RECT 202.730 5007.785 382.270 5012.435 ;
      LAYER met4 ;
        RECT 382.670 5007.385 459.330 5012.835 ;
      LAYER met4 ;
        RECT 459.730 5007.785 639.270 5012.435 ;
      LAYER met4 ;
        RECT 639.670 5007.385 716.330 5012.835 ;
      LAYER met4 ;
        RECT 716.730 5007.785 896.270 5012.435 ;
      LAYER met4 ;
        RECT 896.670 5007.385 973.330 5012.835 ;
      LAYER met4 ;
        RECT 973.730 5007.785 1153.270 5012.435 ;
      LAYER met4 ;
        RECT 1153.670 5007.385 1230.330 5012.835 ;
      LAYER met4 ;
        RECT 1230.730 5007.785 1411.270 5012.435 ;
      LAYER met4 ;
        RECT 1411.670 5007.385 1488.330 5012.835 ;
      LAYER met4 ;
        RECT 1488.730 5007.785 1668.270 5012.435 ;
      LAYER met4 ;
        RECT 1668.670 5007.385 1740.330 5012.835 ;
      LAYER met4 ;
        RECT 1740.730 5007.785 1920.270 5012.435 ;
      LAYER met4 ;
        RECT 1920.670 5007.385 1997.330 5012.835 ;
      LAYER met4 ;
        RECT 1997.730 5007.785 2365.270 5012.435 ;
      LAYER met4 ;
        RECT 2365.670 5007.385 2442.330 5012.835 ;
      LAYER met4 ;
        RECT 2442.730 5007.785 2622.270 5012.435 ;
      LAYER met4 ;
        RECT 2622.670 5007.385 2699.330 5012.835 ;
      LAYER met4 ;
        RECT 2699.730 5007.785 2879.270 5012.435 ;
      LAYER met4 ;
        RECT 2879.670 5007.385 2951.330 5012.835 ;
      LAYER met4 ;
        RECT 2951.730 5007.785 3131.270 5012.435 ;
      LAYER met4 ;
        RECT 3131.670 5007.385 3208.330 5012.835 ;
      LAYER met4 ;
        RECT 3208.730 5007.785 3389.525 5012.435 ;
      LAYER met4 ;
        RECT 3389.925 5011.575 3588.000 5012.835 ;
        RECT 3389.925 5011.310 3444.005 5011.575 ;
        RECT 3389.925 5007.975 3440.725 5011.310 ;
        RECT 3389.925 5007.385 3435.335 5007.975 ;
        RECT 152.665 5006.785 202.745 5007.385 ;
        RECT 381.965 5006.785 459.970 5007.385 ;
        RECT 638.965 5006.785 716.970 5007.385 ;
        RECT 895.965 5006.785 973.970 5007.385 ;
        RECT 1152.965 5006.785 1230.970 5007.385 ;
        RECT 1410.965 5006.785 1488.970 5007.385 ;
        RECT 1667.965 5006.785 1741.035 5007.385 ;
        RECT 1919.965 5006.785 1997.970 5007.385 ;
        RECT 2364.965 5006.785 2442.970 5007.385 ;
        RECT 2621.965 5006.785 2699.970 5007.385 ;
        RECT 2878.965 5006.785 2952.035 5007.385 ;
        RECT 3130.965 5006.785 3208.970 5007.385 ;
        RECT 3388.000 5006.785 3435.335 5007.385 ;
        RECT 152.665 5002.535 202.345 5006.785 ;
      LAYER met4 ;
        RECT 202.745 5002.935 381.965 5006.385 ;
      LAYER met4 ;
        RECT 382.365 5002.535 459.570 5006.785 ;
      LAYER met4 ;
        RECT 459.970 5002.935 638.965 5006.385 ;
      LAYER met4 ;
        RECT 639.365 5002.535 716.570 5006.785 ;
      LAYER met4 ;
        RECT 716.970 5002.935 895.965 5006.385 ;
      LAYER met4 ;
        RECT 896.365 5002.535 973.570 5006.785 ;
      LAYER met4 ;
        RECT 973.970 5002.935 1152.965 5006.385 ;
      LAYER met4 ;
        RECT 1153.365 5002.535 1230.570 5006.785 ;
      LAYER met4 ;
        RECT 1230.970 5002.935 1410.965 5006.385 ;
      LAYER met4 ;
        RECT 1411.365 5002.535 1488.570 5006.785 ;
      LAYER met4 ;
        RECT 1488.970 5002.935 1667.965 5006.385 ;
      LAYER met4 ;
        RECT 1668.365 5002.535 1740.635 5006.785 ;
      LAYER met4 ;
        RECT 1741.035 5002.935 1742.000 5006.385 ;
        RECT 1747.000 5002.935 1919.965 5006.385 ;
      LAYER met4 ;
        RECT 1920.365 5002.535 1997.570 5006.785 ;
      LAYER met4 ;
        RECT 1997.970 5002.935 2364.965 5006.385 ;
      LAYER met4 ;
        RECT 2365.365 5002.535 2442.570 5006.785 ;
      LAYER met4 ;
        RECT 2442.970 5002.935 2621.965 5006.385 ;
      LAYER met4 ;
        RECT 2622.365 5002.535 2699.570 5006.785 ;
      LAYER met4 ;
        RECT 2699.970 5002.935 2878.965 5006.385 ;
      LAYER met4 ;
        RECT 2879.365 5002.535 2951.635 5006.785 ;
      LAYER met4 ;
        RECT 2952.035 5002.935 3130.965 5006.385 ;
      LAYER met4 ;
        RECT 3131.365 5002.535 3208.570 5006.785 ;
      LAYER met4 ;
        RECT 3208.970 5002.935 3389.470 5006.385 ;
      LAYER met4 ;
        RECT 3389.870 5002.535 3435.335 5006.785 ;
        RECT 152.665 5001.935 202.745 5002.535 ;
        RECT 381.965 5001.935 459.970 5002.535 ;
        RECT 638.965 5001.935 716.970 5002.535 ;
        RECT 895.965 5001.935 973.970 5002.535 ;
        RECT 1152.965 5001.935 1230.970 5002.535 ;
        RECT 1410.965 5001.935 1488.970 5002.535 ;
        RECT 1667.965 5001.935 1741.035 5002.535 ;
        RECT 1919.965 5001.935 1997.970 5002.535 ;
        RECT 2364.965 5001.935 2442.970 5002.535 ;
        RECT 2621.965 5001.935 2699.970 5002.535 ;
        RECT 2878.965 5001.935 2952.035 5002.535 ;
        RECT 3130.965 5001.935 3208.970 5002.535 ;
        RECT 3388.000 5001.935 3435.335 5002.535 ;
        RECT 152.665 4996.485 202.330 5001.935 ;
      LAYER met4 ;
        RECT 202.730 4996.885 382.270 5001.535 ;
      LAYER met4 ;
        RECT 382.670 4996.485 459.330 5001.935 ;
      LAYER met4 ;
        RECT 459.730 4996.885 639.270 5001.535 ;
      LAYER met4 ;
        RECT 639.670 4996.485 716.330 5001.935 ;
      LAYER met4 ;
        RECT 716.730 4996.885 896.270 5001.535 ;
      LAYER met4 ;
        RECT 896.670 4996.485 973.330 5001.935 ;
      LAYER met4 ;
        RECT 973.730 4996.885 1153.270 5001.535 ;
      LAYER met4 ;
        RECT 1153.670 4996.485 1230.330 5001.935 ;
      LAYER met4 ;
        RECT 1230.730 4996.885 1411.270 5001.535 ;
      LAYER met4 ;
        RECT 1411.670 4996.485 1488.330 5001.935 ;
      LAYER met4 ;
        RECT 1488.730 4996.885 1668.270 5001.535 ;
      LAYER met4 ;
        RECT 1668.670 4996.485 1740.330 5001.935 ;
      LAYER met4 ;
        RECT 1740.730 4996.885 1747.000 5001.535 ;
        RECT 1752.000 4996.885 1920.270 5001.535 ;
      LAYER met4 ;
        RECT 1920.670 4996.485 1997.330 5001.935 ;
      LAYER met4 ;
        RECT 1997.730 4996.885 2365.270 5001.535 ;
      LAYER met4 ;
        RECT 2365.670 4996.485 2442.330 5001.935 ;
      LAYER met4 ;
        RECT 2442.730 4996.885 2622.270 5001.535 ;
      LAYER met4 ;
        RECT 2622.670 4996.485 2699.330 5001.935 ;
      LAYER met4 ;
        RECT 2699.730 4996.885 2879.270 5001.535 ;
      LAYER met4 ;
        RECT 2879.670 4996.485 2951.330 5001.935 ;
      LAYER met4 ;
        RECT 2951.730 4996.885 3131.270 5001.535 ;
      LAYER met4 ;
        RECT 3131.670 4996.485 3208.330 5001.935 ;
      LAYER met4 ;
        RECT 3208.730 4996.885 3391.785 5001.535 ;
      LAYER met4 ;
        RECT 3392.185 4996.485 3435.335 5001.935 ;
        RECT 152.665 4995.885 202.745 4996.485 ;
        RECT 381.965 4995.885 459.970 4996.485 ;
        RECT 638.965 4995.885 716.970 4996.485 ;
        RECT 895.965 4995.885 973.970 4996.485 ;
        RECT 1152.965 4995.885 1230.970 4996.485 ;
        RECT 1410.965 4995.885 1488.970 4996.485 ;
        RECT 1667.965 4995.885 1741.035 4996.485 ;
        RECT 1919.965 4995.885 1997.970 4996.485 ;
        RECT 2364.965 4995.885 2442.970 4996.485 ;
        RECT 2621.965 4995.885 2699.970 4996.485 ;
        RECT 2878.965 4995.885 2952.035 4996.485 ;
        RECT 3130.965 4995.885 3208.970 4996.485 ;
        RECT 3388.000 4995.885 3435.335 4996.485 ;
        RECT 152.665 4992.185 202.330 4995.885 ;
        RECT 152.665 4990.000 186.065 4992.185 ;
        RECT 152.665 4989.875 169.115 4990.000 ;
        RECT 152.665 4988.000 153.365 4989.875 ;
        RECT 158.815 4989.785 169.115 4989.875 ;
        RECT 158.815 4989.735 164.265 4989.785 ;
        RECT 152.665 4849.330 153.365 4849.970 ;
      LAYER met4 ;
        RECT 153.765 4849.730 158.415 4989.475 ;
      LAYER met4 ;
        RECT 158.815 4988.000 159.415 4989.735 ;
        RECT 158.815 4849.330 159.415 4849.970 ;
      LAYER met4 ;
        RECT 159.815 4849.730 163.265 4989.335 ;
      LAYER met4 ;
        RECT 163.665 4988.000 164.265 4989.735 ;
        RECT 163.665 4849.330 164.265 4849.970 ;
      LAYER met4 ;
        RECT 164.665 4849.730 168.115 4989.385 ;
      LAYER met4 ;
        RECT 168.515 4988.000 169.115 4989.785 ;
        RECT 174.565 4989.925 186.065 4990.000 ;
        RECT 168.515 4849.330 169.115 4849.970 ;
      LAYER met4 ;
        RECT 169.515 4849.730 174.165 4989.600 ;
      LAYER met4 ;
        RECT 174.565 4988.000 175.165 4989.925 ;
        RECT 180.615 4989.870 186.065 4989.925 ;
        RECT 174.565 4849.330 175.165 4849.970 ;
      LAYER met4 ;
        RECT 175.565 4849.730 180.215 4989.525 ;
      LAYER met4 ;
        RECT 180.615 4988.000 181.215 4989.870 ;
      LAYER met4 ;
        RECT 181.615 4849.970 185.065 4989.470 ;
      LAYER met4 ;
        RECT 185.465 4988.000 186.065 4989.870 ;
        RECT 180.615 4849.570 181.215 4849.970 ;
        RECT 185.465 4849.570 186.065 4849.970 ;
      LAYER met4 ;
        RECT 186.465 4849.730 191.115 4991.785 ;
      LAYER met4 ;
        RECT 191.515 4990.750 202.330 4992.185 ;
        RECT 191.515 4988.000 192.115 4990.750 ;
        RECT 180.615 4849.330 186.065 4849.570 ;
        RECT 191.515 4849.330 192.115 4849.970 ;
      LAYER met4 ;
        RECT 192.515 4849.730 197.965 4990.350 ;
      LAYER met4 ;
        RECT 198.365 4989.635 202.330 4990.750 ;
      LAYER met4 ;
        RECT 202.730 4990.035 382.270 4995.485 ;
      LAYER met4 ;
        RECT 382.670 4989.635 459.330 4995.885 ;
      LAYER met4 ;
        RECT 459.730 4990.035 639.270 4995.485 ;
      LAYER met4 ;
        RECT 639.670 4989.635 716.330 4995.885 ;
      LAYER met4 ;
        RECT 716.730 4990.035 896.270 4995.485 ;
      LAYER met4 ;
        RECT 896.670 4989.635 973.330 4995.885 ;
      LAYER met4 ;
        RECT 973.730 4990.035 1153.270 4995.485 ;
      LAYER met4 ;
        RECT 1153.670 4989.635 1230.330 4995.885 ;
      LAYER met4 ;
        RECT 1230.730 4990.035 1411.270 4995.485 ;
      LAYER met4 ;
        RECT 1411.670 4989.635 1488.330 4995.885 ;
      LAYER met4 ;
        RECT 1488.730 4990.035 1668.270 4995.485 ;
      LAYER met4 ;
        RECT 1668.670 4990.035 1740.330 4995.885 ;
      LAYER met4 ;
        RECT 1740.730 4990.035 1920.270 4995.485 ;
      LAYER met4 ;
        RECT 1920.670 4989.635 1997.330 4995.885 ;
      LAYER met4 ;
        RECT 1997.730 4990.035 2365.270 4995.485 ;
      LAYER met4 ;
        RECT 2365.670 4989.635 2442.330 4995.885 ;
      LAYER met4 ;
        RECT 2442.730 4990.035 2622.270 4995.485 ;
      LAYER met4 ;
        RECT 2622.670 4989.635 2699.330 4995.885 ;
      LAYER met4 ;
        RECT 2699.730 4990.035 2879.270 4995.485 ;
      LAYER met4 ;
        RECT 2879.670 4990.035 2951.330 4995.885 ;
      LAYER met4 ;
        RECT 2951.730 4990.035 3131.270 4995.485 ;
      LAYER met4 ;
        RECT 3131.670 4989.635 3208.330 4995.885 ;
      LAYER met4 ;
        RECT 3208.730 4990.035 3390.350 4995.485 ;
      LAYER met4 ;
        RECT 3390.750 4989.635 3435.335 4995.885 ;
        RECT 198.365 4988.000 202.745 4989.635 ;
        RECT 381.965 4988.535 459.970 4989.635 ;
        RECT 638.965 4988.535 716.970 4989.635 ;
        RECT 895.965 4988.535 973.970 4989.635 ;
        RECT 1152.965 4988.535 1230.970 4989.635 ;
        RECT 1410.965 4988.535 1488.970 4989.635 ;
        RECT 1919.965 4988.535 1997.970 4989.635 ;
        RECT 2364.965 4988.535 2442.970 4989.635 ;
        RECT 2621.965 4988.535 2699.970 4989.635 ;
        RECT 3130.965 4988.535 3208.970 4989.635 ;
        RECT 3388.000 4985.670 3435.335 4989.635 ;
        RECT 3388.000 4985.255 3389.635 4985.670 ;
        RECT 198.365 4849.330 199.465 4849.970 ;
        RECT 152.665 4817.690 199.465 4849.330 ;
        RECT 152.035 4774.010 199.465 4817.690 ;
      LAYER met4 ;
        RECT 151.935 4211.730 152.265 4773.610 ;
      LAYER met4 ;
        RECT 152.665 4772.670 199.465 4774.010 ;
        RECT 152.665 4771.965 153.365 4772.670 ;
        RECT 152.665 4633.330 153.365 4635.000 ;
      LAYER met4 ;
        RECT 153.765 4633.730 158.415 4772.270 ;
      LAYER met4 ;
        RECT 158.815 4771.965 159.415 4772.670 ;
        RECT 158.815 4633.330 159.415 4635.000 ;
      LAYER met4 ;
        RECT 159.815 4633.730 163.265 4772.270 ;
      LAYER met4 ;
        RECT 163.665 4771.965 164.265 4772.670 ;
        RECT 163.665 4633.330 164.265 4635.000 ;
      LAYER met4 ;
        RECT 164.665 4633.730 168.115 4772.270 ;
      LAYER met4 ;
        RECT 168.515 4771.965 169.115 4772.670 ;
        RECT 168.515 4633.330 169.115 4635.000 ;
      LAYER met4 ;
        RECT 169.515 4633.730 174.165 4772.270 ;
      LAYER met4 ;
        RECT 174.565 4771.965 175.165 4772.670 ;
        RECT 180.615 4772.365 186.065 4772.670 ;
        RECT 174.165 4634.935 174.200 4645.935 ;
        RECT 174.565 4633.330 175.165 4635.000 ;
      LAYER met4 ;
        RECT 175.565 4633.730 180.215 4772.270 ;
      LAYER met4 ;
        RECT 180.615 4771.965 181.215 4772.365 ;
        RECT 185.465 4771.965 186.065 4772.365 ;
        RECT 180.615 4633.635 181.215 4635.000 ;
      LAYER met4 ;
        RECT 181.615 4634.035 185.065 4771.965 ;
      LAYER met4 ;
        RECT 185.465 4633.635 186.065 4635.000 ;
      LAYER met4 ;
        RECT 186.465 4633.730 191.115 4772.270 ;
      LAYER met4 ;
        RECT 191.515 4771.965 192.115 4772.670 ;
        RECT 180.615 4633.330 186.065 4633.635 ;
        RECT 191.515 4633.330 192.115 4635.000 ;
      LAYER met4 ;
        RECT 192.515 4633.730 197.965 4772.270 ;
      LAYER met4 ;
        RECT 198.365 4771.965 199.465 4772.670 ;
        RECT 3388.535 4836.330 3389.635 4837.035 ;
      LAYER met4 ;
        RECT 3390.035 4836.730 3395.485 4985.270 ;
      LAYER met4 ;
        RECT 3395.885 4985.255 3396.485 4985.670 ;
        RECT 3401.935 4985.655 3407.385 4985.670 ;
        RECT 3395.885 4836.330 3396.485 4837.035 ;
      LAYER met4 ;
        RECT 3396.885 4836.730 3401.535 4985.270 ;
      LAYER met4 ;
        RECT 3401.935 4985.255 3402.535 4985.655 ;
        RECT 3406.785 4985.255 3407.385 4985.655 ;
      LAYER met4 ;
        RECT 3402.935 4837.035 3406.385 4985.255 ;
      LAYER met4 ;
        RECT 3401.935 4836.635 3402.535 4837.035 ;
        RECT 3406.785 4836.635 3407.385 4837.035 ;
      LAYER met4 ;
        RECT 3407.785 4836.730 3412.435 4985.270 ;
      LAYER met4 ;
        RECT 3412.835 4985.255 3413.435 4985.670 ;
        RECT 3401.935 4836.330 3407.385 4836.635 ;
        RECT 3412.835 4836.330 3413.435 4837.035 ;
      LAYER met4 ;
        RECT 3413.835 4836.730 3418.485 4985.270 ;
      LAYER met4 ;
        RECT 3418.885 4985.255 3419.485 4985.670 ;
        RECT 3418.885 4836.330 3419.485 4837.035 ;
      LAYER met4 ;
        RECT 3419.885 4836.730 3423.335 4985.270 ;
      LAYER met4 ;
        RECT 3423.735 4985.255 3424.335 4985.670 ;
        RECT 3423.735 4836.330 3424.335 4837.035 ;
      LAYER met4 ;
        RECT 3424.735 4836.730 3428.185 4985.270 ;
      LAYER met4 ;
        RECT 3428.585 4985.255 3429.185 4985.670 ;
        RECT 3428.585 4836.330 3429.185 4837.035 ;
      LAYER met4 ;
        RECT 3429.585 4836.730 3434.235 4985.270 ;
      LAYER met4 ;
        RECT 3434.635 4985.255 3435.335 4985.670 ;
        RECT 3434.635 4836.330 3435.335 4837.035 ;
        RECT 3388.535 4834.990 3435.335 4836.330 ;
      LAYER met4 ;
        RECT 3435.735 4835.390 3436.065 5007.575 ;
      LAYER met4 ;
        RECT 3436.465 5005.955 3440.725 5007.975 ;
        RECT 3436.465 5005.275 3439.245 5005.955 ;
        RECT 3388.535 4791.310 3435.965 4834.990 ;
        RECT 3388.535 4759.670 3435.335 4791.310 ;
        RECT 3388.535 4759.030 3389.635 4759.670 ;
        RECT 152.665 4561.670 197.965 4633.330 ;
      LAYER met4 ;
        RECT 3390.035 4611.730 3395.485 4759.270 ;
      LAYER met4 ;
        RECT 3395.885 4759.030 3396.485 4759.670 ;
        RECT 3401.935 4759.430 3407.385 4759.670 ;
        RECT 3395.885 4611.330 3396.485 4613.000 ;
      LAYER met4 ;
        RECT 3396.885 4611.730 3401.535 4759.270 ;
      LAYER met4 ;
        RECT 3401.935 4759.030 3402.535 4759.430 ;
        RECT 3406.785 4759.030 3407.385 4759.430 ;
        RECT 3401.935 4611.635 3402.535 4613.000 ;
      LAYER met4 ;
        RECT 3402.935 4612.035 3406.385 4759.030 ;
      LAYER met4 ;
        RECT 3406.785 4611.635 3407.385 4613.000 ;
      LAYER met4 ;
        RECT 3407.785 4611.730 3412.435 4759.270 ;
      LAYER met4 ;
        RECT 3412.835 4759.030 3413.435 4759.670 ;
        RECT 3401.935 4611.330 3407.385 4611.635 ;
        RECT 3412.835 4611.330 3413.435 4613.000 ;
      LAYER met4 ;
        RECT 3413.835 4611.730 3418.485 4759.270 ;
      LAYER met4 ;
        RECT 3418.885 4759.030 3419.485 4759.670 ;
        RECT 3418.885 4611.330 3419.485 4613.000 ;
      LAYER met4 ;
        RECT 3419.885 4611.730 3423.335 4759.270 ;
      LAYER met4 ;
        RECT 3423.735 4759.030 3424.335 4759.670 ;
        RECT 3423.735 4611.330 3424.335 4613.000 ;
      LAYER met4 ;
        RECT 3424.735 4611.730 3428.185 4759.270 ;
      LAYER met4 ;
        RECT 3428.585 4759.030 3429.185 4759.670 ;
        RECT 3428.585 4611.330 3429.185 4613.000 ;
        RECT 3429.550 4612.930 3429.585 4623.975 ;
      LAYER met4 ;
        RECT 3429.585 4611.730 3434.235 4759.270 ;
      LAYER met4 ;
        RECT 3434.635 4759.030 3435.335 4759.670 ;
        RECT 3434.635 4611.330 3435.335 4613.000 ;
        RECT 152.665 4560.000 153.365 4561.670 ;
        RECT 152.665 4422.330 153.365 4423.035 ;
      LAYER met4 ;
        RECT 153.765 4422.730 158.415 4561.270 ;
      LAYER met4 ;
        RECT 158.415 4549.025 158.450 4560.070 ;
        RECT 158.815 4560.000 159.415 4561.670 ;
        RECT 158.815 4422.330 159.415 4423.035 ;
      LAYER met4 ;
        RECT 159.815 4422.730 163.265 4561.270 ;
      LAYER met4 ;
        RECT 163.665 4560.000 164.265 4561.670 ;
        RECT 163.665 4422.330 164.265 4423.035 ;
      LAYER met4 ;
        RECT 164.665 4422.730 168.115 4561.270 ;
      LAYER met4 ;
        RECT 168.515 4560.000 169.115 4561.670 ;
        RECT 168.515 4422.330 169.115 4423.035 ;
      LAYER met4 ;
        RECT 169.515 4422.730 174.165 4561.270 ;
      LAYER met4 ;
        RECT 174.565 4560.000 175.165 4561.670 ;
        RECT 180.615 4561.365 186.065 4561.670 ;
        RECT 174.565 4422.330 175.165 4423.035 ;
      LAYER met4 ;
        RECT 175.565 4422.730 180.215 4561.270 ;
      LAYER met4 ;
        RECT 180.615 4560.000 181.215 4561.365 ;
      LAYER met4 ;
        RECT 181.615 4423.035 185.065 4560.965 ;
      LAYER met4 ;
        RECT 185.465 4560.000 186.065 4561.365 ;
        RECT 180.615 4422.635 181.215 4423.035 ;
        RECT 185.465 4422.635 186.065 4423.035 ;
      LAYER met4 ;
        RECT 186.465 4422.730 191.115 4561.270 ;
      LAYER met4 ;
        RECT 191.515 4560.000 192.115 4561.670 ;
        RECT 180.615 4422.330 186.065 4422.635 ;
        RECT 191.515 4422.330 192.115 4423.035 ;
      LAYER met4 ;
        RECT 192.515 4422.730 197.965 4561.270 ;
      LAYER met4 ;
        RECT 3390.035 4539.670 3435.335 4611.330 ;
        RECT 152.665 4350.670 197.965 4422.330 ;
        RECT 3388.535 4390.330 3389.635 4391.035 ;
      LAYER met4 ;
        RECT 3390.035 4390.730 3395.485 4539.270 ;
      LAYER met4 ;
        RECT 3395.885 4538.000 3396.485 4539.670 ;
        RECT 3401.935 4539.365 3407.385 4539.670 ;
        RECT 3395.885 4390.330 3396.485 4391.035 ;
      LAYER met4 ;
        RECT 3396.885 4390.730 3401.535 4539.270 ;
      LAYER met4 ;
        RECT 3401.935 4538.000 3402.535 4539.365 ;
      LAYER met4 ;
        RECT 3402.935 4391.035 3406.385 4538.965 ;
      LAYER met4 ;
        RECT 3406.785 4538.000 3407.385 4539.365 ;
        RECT 3401.935 4390.635 3402.535 4391.035 ;
        RECT 3406.785 4390.635 3407.385 4391.035 ;
      LAYER met4 ;
        RECT 3407.785 4390.730 3412.435 4539.270 ;
      LAYER met4 ;
        RECT 3412.835 4538.000 3413.435 4539.670 ;
        RECT 3413.800 4527.065 3413.835 4538.065 ;
        RECT 3401.935 4390.330 3407.385 4390.635 ;
        RECT 3412.835 4390.330 3413.435 4391.035 ;
      LAYER met4 ;
        RECT 3413.835 4390.730 3418.485 4539.270 ;
      LAYER met4 ;
        RECT 3418.885 4538.000 3419.485 4539.670 ;
        RECT 3418.885 4390.330 3419.485 4391.035 ;
      LAYER met4 ;
        RECT 3419.885 4390.730 3423.335 4539.270 ;
      LAYER met4 ;
        RECT 3423.735 4538.000 3424.335 4539.670 ;
        RECT 3423.735 4390.330 3424.335 4391.035 ;
      LAYER met4 ;
        RECT 3424.735 4390.730 3428.185 4539.270 ;
      LAYER met4 ;
        RECT 3428.585 4538.000 3429.185 4539.670 ;
        RECT 3428.585 4390.330 3429.185 4391.035 ;
      LAYER met4 ;
        RECT 3429.585 4390.730 3434.235 4539.270 ;
      LAYER met4 ;
        RECT 3434.635 4538.000 3435.335 4539.670 ;
        RECT 3434.635 4390.330 3435.335 4391.035 ;
        RECT 3388.535 4388.990 3435.335 4390.330 ;
      LAYER met4 ;
        RECT 3435.735 4389.390 3436.065 4790.910 ;
        RECT 3436.365 4785.855 3439.345 5004.875 ;
        RECT 3439.645 4984.000 3440.825 5005.555 ;
      LAYER met4 ;
        RECT 3439.645 4838.000 3440.825 4984.000 ;
      LAYER met4 ;
        RECT 3439.645 4836.730 3440.825 4838.000 ;
      LAYER met4 ;
        RECT 3439.745 4801.160 3440.725 4836.330 ;
      LAYER met4 ;
        RECT 3441.125 4801.560 3444.105 5010.910 ;
        RECT 3444.405 4835.390 3444.735 5011.175 ;
      LAYER met4 ;
        RECT 3445.135 4986.255 3588.000 5011.575 ;
        RECT 3445.135 4985.670 3457.635 4986.255 ;
        RECT 3445.135 4985.255 3445.835 4985.670 ;
        RECT 3445.135 4838.000 3445.835 4984.000 ;
        RECT 3445.135 4836.330 3445.835 4837.035 ;
      LAYER met4 ;
        RECT 3446.235 4836.730 3450.685 4985.270 ;
      LAYER met4 ;
        RECT 3451.085 4985.255 3451.685 4985.670 ;
        RECT 3451.085 4838.000 3451.685 4984.000 ;
        RECT 3451.085 4836.330 3451.685 4837.035 ;
      LAYER met4 ;
        RECT 3452.085 4836.730 3456.535 4985.270 ;
      LAYER met4 ;
        RECT 3456.935 4985.255 3457.635 4985.670 ;
        RECT 3456.935 4838.000 3457.635 4984.000 ;
        RECT 3456.935 4836.330 3457.635 4837.035 ;
      LAYER met4 ;
        RECT 3458.035 4836.730 3483.000 4985.855 ;
      LAYER met4 ;
        RECT 3483.400 4985.670 3588.000 4986.255 ;
        RECT 3483.400 4985.255 3563.385 4985.670 ;
      LAYER met4 ;
        RECT 3563.785 4984.000 3588.000 4985.270 ;
      LAYER met4 ;
        RECT 3483.400 4838.000 3588.000 4984.000 ;
        RECT 3483.400 4836.330 3563.385 4837.035 ;
      LAYER met4 ;
        RECT 3563.785 4836.730 3588.000 4838.000 ;
      LAYER met4 ;
        RECT 3445.135 4834.990 3588.000 4836.330 ;
        RECT 3444.505 4801.160 3588.000 4834.990 ;
        RECT 3439.745 4799.640 3588.000 4801.160 ;
        RECT 3439.745 4785.455 3440.725 4799.640 ;
        RECT 3436.465 4783.935 3440.725 4785.455 ;
        RECT 152.665 4349.965 153.365 4350.670 ;
        RECT 152.665 4211.330 153.365 4212.035 ;
      LAYER met4 ;
        RECT 153.765 4211.730 158.415 4350.270 ;
      LAYER met4 ;
        RECT 158.815 4349.965 159.415 4350.670 ;
        RECT 158.815 4211.330 159.415 4212.035 ;
      LAYER met4 ;
        RECT 159.815 4211.730 163.265 4350.270 ;
      LAYER met4 ;
        RECT 163.665 4349.965 164.265 4350.670 ;
        RECT 163.665 4211.330 164.265 4212.035 ;
      LAYER met4 ;
        RECT 164.665 4211.730 168.115 4350.270 ;
      LAYER met4 ;
        RECT 168.515 4349.965 169.115 4350.670 ;
        RECT 168.515 4211.330 169.115 4212.035 ;
      LAYER met4 ;
        RECT 169.515 4211.730 174.165 4350.270 ;
      LAYER met4 ;
        RECT 174.565 4349.965 175.165 4350.670 ;
        RECT 180.615 4350.365 186.065 4350.670 ;
        RECT 174.565 4211.330 175.165 4212.035 ;
      LAYER met4 ;
        RECT 175.565 4211.730 180.215 4350.270 ;
      LAYER met4 ;
        RECT 180.615 4349.965 181.215 4350.365 ;
        RECT 185.465 4349.965 186.065 4350.365 ;
      LAYER met4 ;
        RECT 181.615 4212.035 185.065 4349.965 ;
      LAYER met4 ;
        RECT 180.615 4211.635 181.215 4212.035 ;
        RECT 185.465 4211.635 186.065 4212.035 ;
      LAYER met4 ;
        RECT 186.465 4211.730 191.115 4350.270 ;
      LAYER met4 ;
        RECT 191.515 4349.965 192.115 4350.670 ;
        RECT 180.615 4211.330 186.065 4211.635 ;
        RECT 191.515 4211.330 192.115 4212.035 ;
      LAYER met4 ;
        RECT 192.515 4211.730 197.965 4350.270 ;
      LAYER met4 ;
        RECT 3388.535 4345.310 3435.965 4388.990 ;
        RECT 3388.535 4313.670 3435.335 4345.310 ;
        RECT 3388.535 4313.030 3389.635 4313.670 ;
        RECT 152.035 4139.670 197.965 4211.330 ;
      LAYER met4 ;
        RECT 3390.035 4165.730 3395.485 4313.270 ;
      LAYER met4 ;
        RECT 3395.885 4313.030 3396.485 4313.670 ;
        RECT 3401.935 4313.430 3407.385 4313.670 ;
        RECT 3395.885 4165.330 3396.485 4166.035 ;
      LAYER met4 ;
        RECT 3396.885 4165.730 3401.535 4313.270 ;
      LAYER met4 ;
        RECT 3401.935 4313.030 3402.535 4313.430 ;
        RECT 3406.785 4313.030 3407.385 4313.430 ;
      LAYER met4 ;
        RECT 3402.935 4166.035 3406.385 4313.030 ;
      LAYER met4 ;
        RECT 3401.935 4165.635 3402.535 4166.035 ;
        RECT 3406.785 4165.635 3407.385 4166.035 ;
      LAYER met4 ;
        RECT 3407.785 4165.730 3412.435 4313.270 ;
      LAYER met4 ;
        RECT 3412.835 4313.030 3413.435 4313.670 ;
        RECT 3401.935 4165.330 3407.385 4165.635 ;
        RECT 3412.835 4165.330 3413.435 4166.035 ;
      LAYER met4 ;
        RECT 3413.835 4165.730 3418.485 4313.270 ;
      LAYER met4 ;
        RECT 3418.885 4313.030 3419.485 4313.670 ;
        RECT 3418.885 4165.330 3419.485 4166.035 ;
      LAYER met4 ;
        RECT 3419.885 4165.730 3423.335 4313.270 ;
      LAYER met4 ;
        RECT 3423.735 4313.030 3424.335 4313.670 ;
        RECT 3423.735 4165.330 3424.335 4166.035 ;
      LAYER met4 ;
        RECT 3424.735 4165.730 3428.185 4313.270 ;
      LAYER met4 ;
        RECT 3428.585 4313.030 3429.185 4313.670 ;
        RECT 3428.585 4165.330 3429.185 4166.035 ;
      LAYER met4 ;
        RECT 3429.585 4165.730 3434.235 4313.270 ;
      LAYER met4 ;
        RECT 3434.635 4313.030 3435.335 4313.670 ;
        RECT 3434.635 4165.330 3435.335 4166.035 ;
        RECT 147.275 3974.545 151.535 3976.065 ;
        RECT 147.275 3960.360 148.255 3974.545 ;
        RECT 0.000 3958.840 148.255 3960.360 ;
        RECT 0.000 3925.010 143.495 3958.840 ;
        RECT 0.000 3923.670 142.865 3925.010 ;
      LAYER met4 ;
        RECT 0.000 3922.000 24.215 3923.270 ;
      LAYER met4 ;
        RECT 24.615 3922.965 104.600 3923.670 ;
        RECT 0.000 3786.000 104.600 3922.000 ;
      LAYER met4 ;
        RECT 0.000 3784.730 24.215 3786.000 ;
      LAYER met4 ;
        RECT 24.615 3784.330 104.600 3784.970 ;
      LAYER met4 ;
        RECT 105.000 3784.730 129.965 3923.270 ;
      LAYER met4 ;
        RECT 130.365 3922.965 131.065 3923.670 ;
        RECT 130.365 3786.000 131.065 3922.000 ;
        RECT 130.365 3784.330 131.065 3784.970 ;
      LAYER met4 ;
        RECT 131.465 3784.730 135.915 3923.270 ;
      LAYER met4 ;
        RECT 136.315 3922.965 136.915 3923.670 ;
        RECT 136.315 3786.000 136.915 3922.000 ;
        RECT 136.315 3784.330 136.915 3784.970 ;
      LAYER met4 ;
        RECT 137.315 3784.730 141.765 3923.270 ;
      LAYER met4 ;
        RECT 142.165 3922.965 142.865 3923.670 ;
        RECT 142.165 3786.000 142.865 3922.000 ;
        RECT 142.165 3784.330 142.865 3784.970 ;
        RECT 0.000 3752.690 142.865 3784.330 ;
      LAYER met4 ;
        RECT 143.265 3753.090 143.595 3924.610 ;
      LAYER met4 ;
        RECT 0.000 3744.360 143.495 3752.690 ;
      LAYER met4 ;
        RECT 143.895 3744.760 146.875 3958.440 ;
      LAYER met4 ;
        RECT 147.275 3923.670 148.255 3958.840 ;
      LAYER met4 ;
        RECT 147.175 3922.000 148.355 3923.270 ;
      LAYER met4 ;
        RECT 147.175 3786.000 148.355 3922.000 ;
      LAYER met4 ;
        RECT 147.175 3784.730 148.355 3786.000 ;
      LAYER met4 ;
        RECT 147.275 3760.065 148.255 3784.330 ;
      LAYER met4 ;
        RECT 148.655 3760.465 151.635 3974.145 ;
        RECT 151.935 3969.090 152.265 4139.270 ;
      LAYER met4 ;
        RECT 152.665 4138.965 153.365 4139.670 ;
        RECT 152.665 4000.330 153.365 4000.970 ;
      LAYER met4 ;
        RECT 153.765 4000.730 158.415 4139.270 ;
      LAYER met4 ;
        RECT 158.815 4138.965 159.415 4139.670 ;
        RECT 158.815 4000.330 159.415 4000.970 ;
      LAYER met4 ;
        RECT 159.815 4000.730 163.265 4139.270 ;
      LAYER met4 ;
        RECT 163.665 4138.965 164.265 4139.670 ;
        RECT 163.665 4000.330 164.265 4000.970 ;
      LAYER met4 ;
        RECT 164.665 4000.730 168.115 4139.270 ;
      LAYER met4 ;
        RECT 168.515 4138.965 169.115 4139.670 ;
        RECT 168.515 4000.330 169.115 4000.970 ;
      LAYER met4 ;
        RECT 169.515 4000.730 174.165 4139.270 ;
      LAYER met4 ;
        RECT 174.565 4138.965 175.165 4139.670 ;
        RECT 180.615 4139.365 186.065 4139.670 ;
        RECT 174.565 4000.330 175.165 4000.970 ;
      LAYER met4 ;
        RECT 175.565 4000.730 180.215 4139.270 ;
      LAYER met4 ;
        RECT 180.615 4138.965 181.215 4139.365 ;
        RECT 185.465 4138.965 186.065 4139.365 ;
      LAYER met4 ;
        RECT 181.615 4000.970 185.065 4138.965 ;
      LAYER met4 ;
        RECT 180.615 4000.570 181.215 4000.970 ;
        RECT 185.465 4000.570 186.065 4000.970 ;
      LAYER met4 ;
        RECT 186.465 4000.730 191.115 4139.270 ;
      LAYER met4 ;
        RECT 191.515 4138.965 192.115 4139.670 ;
        RECT 180.615 4000.330 186.065 4000.570 ;
        RECT 191.515 4000.330 192.115 4000.970 ;
      LAYER met4 ;
        RECT 192.515 4000.730 197.965 4139.270 ;
      LAYER met4 ;
        RECT 3390.035 4093.670 3435.335 4165.330 ;
        RECT 198.365 4000.330 199.465 4000.970 ;
        RECT 152.665 3968.690 199.465 4000.330 ;
        RECT 152.035 3925.010 199.465 3968.690 ;
        RECT 147.275 3758.545 151.535 3760.065 ;
        RECT 147.275 3744.360 148.255 3758.545 ;
        RECT 0.000 3742.840 148.255 3744.360 ;
        RECT 0.000 3709.010 143.495 3742.840 ;
        RECT 0.000 3707.670 142.865 3709.010 ;
      LAYER met4 ;
        RECT 0.000 3706.000 24.215 3707.270 ;
      LAYER met4 ;
        RECT 24.615 3706.965 104.600 3707.670 ;
        RECT 0.000 3570.000 104.600 3706.000 ;
      LAYER met4 ;
        RECT 0.000 3568.730 24.215 3570.000 ;
      LAYER met4 ;
        RECT 24.615 3568.330 104.600 3568.970 ;
      LAYER met4 ;
        RECT 105.000 3568.730 129.965 3707.270 ;
      LAYER met4 ;
        RECT 130.365 3706.965 131.065 3707.670 ;
        RECT 130.365 3570.000 131.065 3706.000 ;
        RECT 130.365 3568.330 131.065 3568.970 ;
      LAYER met4 ;
        RECT 131.465 3568.730 135.915 3707.270 ;
      LAYER met4 ;
        RECT 136.315 3706.965 136.915 3707.670 ;
        RECT 136.315 3570.000 136.915 3706.000 ;
        RECT 136.315 3568.330 136.915 3568.970 ;
      LAYER met4 ;
        RECT 137.315 3568.730 141.765 3707.270 ;
      LAYER met4 ;
        RECT 142.165 3706.965 142.865 3707.670 ;
        RECT 142.165 3570.000 142.865 3706.000 ;
        RECT 142.165 3568.330 142.865 3568.970 ;
        RECT 0.000 3536.690 142.865 3568.330 ;
      LAYER met4 ;
        RECT 143.265 3537.090 143.595 3708.610 ;
      LAYER met4 ;
        RECT 0.000 3528.360 143.495 3536.690 ;
      LAYER met4 ;
        RECT 143.895 3528.760 146.875 3742.440 ;
      LAYER met4 ;
        RECT 147.275 3707.670 148.255 3742.840 ;
      LAYER met4 ;
        RECT 147.175 3706.000 148.355 3707.270 ;
      LAYER met4 ;
        RECT 147.175 3570.000 148.355 3706.000 ;
      LAYER met4 ;
        RECT 147.175 3568.730 148.355 3570.000 ;
      LAYER met4 ;
        RECT 147.275 3544.065 148.255 3568.330 ;
      LAYER met4 ;
        RECT 148.655 3544.465 151.635 3758.145 ;
        RECT 151.935 3753.090 152.265 3924.610 ;
      LAYER met4 ;
        RECT 152.665 3923.670 199.465 3925.010 ;
        RECT 152.665 3922.965 153.365 3923.670 ;
        RECT 152.665 3784.330 153.365 3784.970 ;
      LAYER met4 ;
        RECT 153.765 3784.730 158.415 3923.270 ;
      LAYER met4 ;
        RECT 158.815 3922.965 159.415 3923.670 ;
        RECT 158.815 3784.330 159.415 3784.970 ;
      LAYER met4 ;
        RECT 159.815 3784.730 163.265 3923.270 ;
      LAYER met4 ;
        RECT 163.665 3922.965 164.265 3923.670 ;
        RECT 163.665 3784.330 164.265 3784.970 ;
      LAYER met4 ;
        RECT 164.665 3784.730 168.115 3923.270 ;
      LAYER met4 ;
        RECT 168.515 3922.965 169.115 3923.670 ;
        RECT 168.515 3784.330 169.115 3784.970 ;
      LAYER met4 ;
        RECT 169.515 3784.730 174.165 3923.270 ;
      LAYER met4 ;
        RECT 174.565 3922.965 175.165 3923.670 ;
        RECT 180.615 3923.365 186.065 3923.670 ;
        RECT 174.565 3784.330 175.165 3784.970 ;
      LAYER met4 ;
        RECT 175.565 3784.730 180.215 3923.270 ;
      LAYER met4 ;
        RECT 180.615 3922.965 181.215 3923.365 ;
        RECT 185.465 3922.965 186.065 3923.365 ;
      LAYER met4 ;
        RECT 181.615 3784.970 185.065 3922.965 ;
      LAYER met4 ;
        RECT 180.615 3784.570 181.215 3784.970 ;
        RECT 185.465 3784.570 186.065 3784.970 ;
      LAYER met4 ;
        RECT 186.465 3784.730 191.115 3923.270 ;
      LAYER met4 ;
        RECT 191.515 3922.965 192.115 3923.670 ;
        RECT 180.615 3784.330 186.065 3784.570 ;
        RECT 191.515 3784.330 192.115 3784.970 ;
      LAYER met4 ;
        RECT 192.515 3784.730 197.965 3923.270 ;
      LAYER met4 ;
        RECT 198.365 3922.965 199.465 3923.670 ;
        RECT 3388.535 3944.330 3389.635 3945.035 ;
      LAYER met4 ;
        RECT 3390.035 3944.730 3395.485 4093.270 ;
      LAYER met4 ;
        RECT 3395.885 4092.965 3396.485 4093.670 ;
        RECT 3401.935 4093.365 3407.385 4093.670 ;
        RECT 3395.885 3944.330 3396.485 3945.035 ;
      LAYER met4 ;
        RECT 3396.885 3944.730 3401.535 4093.270 ;
      LAYER met4 ;
        RECT 3401.935 4092.965 3402.535 4093.365 ;
        RECT 3406.785 4092.965 3407.385 4093.365 ;
      LAYER met4 ;
        RECT 3402.935 3945.035 3406.385 4092.965 ;
      LAYER met4 ;
        RECT 3401.935 3944.635 3402.535 3945.035 ;
        RECT 3406.785 3944.635 3407.385 3945.035 ;
      LAYER met4 ;
        RECT 3407.785 3944.730 3412.435 4093.270 ;
      LAYER met4 ;
        RECT 3412.835 4092.965 3413.435 4093.670 ;
        RECT 3401.935 3944.330 3407.385 3944.635 ;
        RECT 3412.835 3944.330 3413.435 3945.035 ;
      LAYER met4 ;
        RECT 3413.835 3944.730 3418.485 4093.270 ;
      LAYER met4 ;
        RECT 3418.885 4092.965 3419.485 4093.670 ;
        RECT 3418.885 3944.330 3419.485 3945.035 ;
      LAYER met4 ;
        RECT 3419.885 3944.730 3423.335 4093.270 ;
      LAYER met4 ;
        RECT 3423.735 4092.965 3424.335 4093.670 ;
        RECT 3423.735 3944.330 3424.335 3945.035 ;
      LAYER met4 ;
        RECT 3424.735 3944.730 3428.185 4093.270 ;
      LAYER met4 ;
        RECT 3428.585 4092.965 3429.185 4093.670 ;
        RECT 3428.585 3944.330 3429.185 3945.035 ;
      LAYER met4 ;
        RECT 3429.585 3944.730 3434.235 4093.270 ;
      LAYER met4 ;
        RECT 3434.635 4092.965 3435.335 4093.670 ;
        RECT 3434.635 3944.330 3435.335 3945.035 ;
        RECT 3388.535 3942.990 3435.335 3944.330 ;
      LAYER met4 ;
        RECT 3435.735 3943.390 3436.065 4344.910 ;
        RECT 3436.365 4339.855 3439.345 4783.535 ;
      LAYER met4 ;
        RECT 3439.745 4759.670 3440.725 4783.935 ;
      LAYER met4 ;
        RECT 3439.645 4758.000 3440.825 4759.270 ;
      LAYER met4 ;
        RECT 3439.645 4613.000 3440.825 4758.000 ;
      LAYER met4 ;
        RECT 3439.645 4611.730 3440.825 4613.000 ;
      LAYER met4 ;
        RECT 3439.745 4539.670 3440.725 4611.330 ;
      LAYER met4 ;
        RECT 3439.645 4538.000 3440.825 4539.270 ;
      LAYER met4 ;
        RECT 3439.645 4392.000 3440.825 4538.000 ;
      LAYER met4 ;
        RECT 3439.645 4390.730 3440.825 4392.000 ;
      LAYER met4 ;
        RECT 3439.745 4355.160 3440.725 4390.330 ;
      LAYER met4 ;
        RECT 3441.125 4355.560 3444.105 4799.240 ;
      LAYER met4 ;
        RECT 3444.505 4791.310 3588.000 4799.640 ;
      LAYER met4 ;
        RECT 3444.405 4389.390 3444.735 4790.910 ;
      LAYER met4 ;
        RECT 3445.135 4759.670 3588.000 4791.310 ;
        RECT 3445.135 4759.030 3445.835 4759.670 ;
        RECT 3445.135 4611.330 3445.835 4758.000 ;
      LAYER met4 ;
        RECT 3446.235 4611.730 3450.685 4759.270 ;
      LAYER met4 ;
        RECT 3451.085 4759.030 3451.685 4759.670 ;
        RECT 3451.085 4611.330 3451.685 4758.000 ;
      LAYER met4 ;
        RECT 3452.085 4611.730 3456.535 4759.270 ;
      LAYER met4 ;
        RECT 3456.935 4759.030 3457.635 4759.670 ;
        RECT 3456.935 4611.330 3457.635 4758.000 ;
      LAYER met4 ;
        RECT 3458.035 4611.730 3483.000 4759.270 ;
      LAYER met4 ;
        RECT 3483.400 4759.030 3563.385 4759.670 ;
      LAYER met4 ;
        RECT 3563.785 4758.000 3588.000 4759.270 ;
      LAYER met4 ;
        RECT 3483.400 4613.000 3588.000 4758.000 ;
        RECT 3483.400 4611.330 3563.385 4613.000 ;
      LAYER met4 ;
        RECT 3563.785 4611.730 3588.000 4613.000 ;
      LAYER met4 ;
        RECT 3445.135 4539.670 3588.000 4611.330 ;
        RECT 3445.135 4392.000 3445.835 4539.670 ;
        RECT 3445.135 4390.330 3445.835 4391.035 ;
      LAYER met4 ;
        RECT 3446.235 4390.730 3450.685 4539.270 ;
      LAYER met4 ;
        RECT 3451.085 4392.000 3451.685 4539.670 ;
        RECT 3451.085 4390.330 3451.685 4391.035 ;
      LAYER met4 ;
        RECT 3452.085 4390.730 3456.535 4539.270 ;
      LAYER met4 ;
        RECT 3456.935 4392.000 3457.635 4539.670 ;
        RECT 3456.935 4390.330 3457.635 4391.035 ;
      LAYER met4 ;
        RECT 3458.035 4390.730 3483.000 4539.270 ;
      LAYER met4 ;
        RECT 3483.400 4538.000 3563.385 4539.670 ;
        RECT 3563.750 4538.000 3563.785 4538.215 ;
      LAYER met4 ;
        RECT 3563.785 4538.000 3588.000 4539.270 ;
      LAYER met4 ;
        RECT 3483.400 4392.000 3588.000 4538.000 ;
        RECT 3483.400 4390.330 3563.385 4391.035 ;
      LAYER met4 ;
        RECT 3563.785 4390.730 3588.000 4392.000 ;
      LAYER met4 ;
        RECT 3445.135 4388.990 3588.000 4390.330 ;
        RECT 3444.505 4355.160 3588.000 4388.990 ;
        RECT 3439.745 4353.640 3588.000 4355.160 ;
        RECT 3439.745 4339.455 3440.725 4353.640 ;
        RECT 3436.465 4337.935 3440.725 4339.455 ;
        RECT 3388.535 3899.310 3435.965 3942.990 ;
        RECT 3388.535 3867.670 3435.335 3899.310 ;
        RECT 3388.535 3867.030 3389.635 3867.670 ;
        RECT 198.365 3784.330 199.465 3784.970 ;
        RECT 152.665 3752.690 199.465 3784.330 ;
        RECT 152.035 3709.010 199.465 3752.690 ;
        RECT 147.275 3542.545 151.535 3544.065 ;
        RECT 147.275 3528.360 148.255 3542.545 ;
        RECT 0.000 3526.840 148.255 3528.360 ;
        RECT 0.000 3493.010 143.495 3526.840 ;
        RECT 0.000 3491.670 142.865 3493.010 ;
      LAYER met4 ;
        RECT 0.000 3490.000 24.215 3491.270 ;
      LAYER met4 ;
        RECT 24.615 3490.965 104.600 3491.670 ;
        RECT 0.000 3354.000 104.600 3490.000 ;
      LAYER met4 ;
        RECT 0.000 3352.730 24.215 3354.000 ;
      LAYER met4 ;
        RECT 24.615 3352.330 104.600 3352.970 ;
      LAYER met4 ;
        RECT 105.000 3352.730 129.965 3491.270 ;
      LAYER met4 ;
        RECT 130.365 3490.965 131.065 3491.670 ;
        RECT 130.365 3354.000 131.065 3490.000 ;
        RECT 130.365 3352.330 131.065 3352.970 ;
      LAYER met4 ;
        RECT 131.465 3352.730 135.915 3491.270 ;
      LAYER met4 ;
        RECT 136.315 3490.965 136.915 3491.670 ;
        RECT 136.315 3354.000 136.915 3490.000 ;
        RECT 136.315 3352.330 136.915 3352.970 ;
      LAYER met4 ;
        RECT 137.315 3352.730 141.765 3491.270 ;
      LAYER met4 ;
        RECT 142.165 3490.965 142.865 3491.670 ;
        RECT 142.165 3354.000 142.865 3490.000 ;
        RECT 142.165 3352.330 142.865 3352.970 ;
        RECT 0.000 3320.690 142.865 3352.330 ;
      LAYER met4 ;
        RECT 143.265 3321.090 143.595 3492.610 ;
      LAYER met4 ;
        RECT 0.000 3312.360 143.495 3320.690 ;
      LAYER met4 ;
        RECT 143.895 3312.760 146.875 3526.440 ;
      LAYER met4 ;
        RECT 147.275 3491.670 148.255 3526.840 ;
      LAYER met4 ;
        RECT 147.175 3490.000 148.355 3491.270 ;
      LAYER met4 ;
        RECT 147.175 3354.000 148.355 3490.000 ;
      LAYER met4 ;
        RECT 147.175 3352.730 148.355 3354.000 ;
      LAYER met4 ;
        RECT 147.275 3328.065 148.255 3352.330 ;
      LAYER met4 ;
        RECT 148.655 3328.465 151.635 3542.145 ;
        RECT 151.935 3537.090 152.265 3708.610 ;
      LAYER met4 ;
        RECT 152.665 3707.670 199.465 3709.010 ;
        RECT 152.665 3706.965 153.365 3707.670 ;
        RECT 152.665 3568.330 153.365 3568.970 ;
      LAYER met4 ;
        RECT 153.765 3568.730 158.415 3707.270 ;
      LAYER met4 ;
        RECT 158.815 3706.965 159.415 3707.670 ;
        RECT 158.815 3568.330 159.415 3568.970 ;
      LAYER met4 ;
        RECT 159.815 3568.730 163.265 3707.270 ;
      LAYER met4 ;
        RECT 163.665 3706.965 164.265 3707.670 ;
        RECT 163.665 3568.330 164.265 3568.970 ;
      LAYER met4 ;
        RECT 164.665 3568.730 168.115 3707.270 ;
      LAYER met4 ;
        RECT 168.515 3706.965 169.115 3707.670 ;
        RECT 168.515 3568.330 169.115 3568.970 ;
      LAYER met4 ;
        RECT 169.515 3568.730 174.165 3707.270 ;
      LAYER met4 ;
        RECT 174.565 3706.965 175.165 3707.670 ;
        RECT 180.615 3707.365 186.065 3707.670 ;
        RECT 174.565 3568.330 175.165 3568.970 ;
      LAYER met4 ;
        RECT 175.565 3568.730 180.215 3707.270 ;
      LAYER met4 ;
        RECT 180.615 3706.965 181.215 3707.365 ;
        RECT 185.465 3706.965 186.065 3707.365 ;
      LAYER met4 ;
        RECT 181.615 3568.970 185.065 3706.965 ;
      LAYER met4 ;
        RECT 180.615 3568.570 181.215 3568.970 ;
        RECT 185.465 3568.570 186.065 3568.970 ;
      LAYER met4 ;
        RECT 186.465 3568.730 191.115 3707.270 ;
      LAYER met4 ;
        RECT 191.515 3706.965 192.115 3707.670 ;
        RECT 180.615 3568.330 186.065 3568.570 ;
        RECT 191.515 3568.330 192.115 3568.970 ;
      LAYER met4 ;
        RECT 192.515 3568.730 197.965 3707.270 ;
      LAYER met4 ;
        RECT 198.365 3706.965 199.465 3707.670 ;
        RECT 3388.535 3719.330 3389.635 3720.035 ;
      LAYER met4 ;
        RECT 3390.035 3719.730 3395.485 3867.270 ;
      LAYER met4 ;
        RECT 3395.885 3867.030 3396.485 3867.670 ;
        RECT 3401.935 3867.430 3407.385 3867.670 ;
        RECT 3395.885 3719.330 3396.485 3720.035 ;
      LAYER met4 ;
        RECT 3396.885 3719.730 3401.535 3867.270 ;
      LAYER met4 ;
        RECT 3401.935 3867.030 3402.535 3867.430 ;
        RECT 3406.785 3867.030 3407.385 3867.430 ;
      LAYER met4 ;
        RECT 3402.935 3720.035 3406.385 3867.030 ;
      LAYER met4 ;
        RECT 3401.935 3719.635 3402.535 3720.035 ;
        RECT 3406.785 3719.635 3407.385 3720.035 ;
      LAYER met4 ;
        RECT 3407.785 3719.730 3412.435 3867.270 ;
      LAYER met4 ;
        RECT 3412.835 3867.030 3413.435 3867.670 ;
        RECT 3401.935 3719.330 3407.385 3719.635 ;
        RECT 3412.835 3719.330 3413.435 3720.035 ;
      LAYER met4 ;
        RECT 3413.835 3719.730 3418.485 3867.270 ;
      LAYER met4 ;
        RECT 3418.885 3867.030 3419.485 3867.670 ;
        RECT 3418.885 3719.330 3419.485 3720.035 ;
      LAYER met4 ;
        RECT 3419.885 3719.730 3423.335 3867.270 ;
      LAYER met4 ;
        RECT 3423.735 3867.030 3424.335 3867.670 ;
        RECT 3423.735 3719.330 3424.335 3720.035 ;
      LAYER met4 ;
        RECT 3424.735 3719.730 3428.185 3867.270 ;
      LAYER met4 ;
        RECT 3428.585 3867.030 3429.185 3867.670 ;
        RECT 3428.585 3719.330 3429.185 3720.035 ;
      LAYER met4 ;
        RECT 3429.585 3719.730 3434.235 3867.270 ;
      LAYER met4 ;
        RECT 3434.635 3867.030 3435.335 3867.670 ;
        RECT 3434.635 3719.330 3435.335 3720.035 ;
        RECT 3388.535 3717.990 3435.335 3719.330 ;
      LAYER met4 ;
        RECT 3435.735 3718.390 3436.065 3898.910 ;
        RECT 3436.365 3893.855 3439.345 4337.535 ;
      LAYER met4 ;
        RECT 3439.745 4313.670 3440.725 4337.935 ;
      LAYER met4 ;
        RECT 3439.645 4312.000 3440.825 4313.270 ;
      LAYER met4 ;
        RECT 3439.645 4167.000 3440.825 4312.000 ;
      LAYER met4 ;
        RECT 3439.645 4165.730 3440.825 4167.000 ;
      LAYER met4 ;
        RECT 3439.745 4093.670 3440.725 4165.330 ;
      LAYER met4 ;
        RECT 3439.645 4092.000 3440.825 4093.270 ;
      LAYER met4 ;
        RECT 3439.645 3946.000 3440.825 4092.000 ;
      LAYER met4 ;
        RECT 3439.645 3944.730 3440.825 3946.000 ;
      LAYER met4 ;
        RECT 3439.745 3909.160 3440.725 3944.330 ;
      LAYER met4 ;
        RECT 3441.125 3909.560 3444.105 4353.240 ;
      LAYER met4 ;
        RECT 3444.505 4345.310 3588.000 4353.640 ;
      LAYER met4 ;
        RECT 3444.405 3943.390 3444.735 4344.910 ;
      LAYER met4 ;
        RECT 3445.135 4313.670 3588.000 4345.310 ;
        RECT 3445.135 4313.030 3445.835 4313.670 ;
        RECT 3445.135 4167.000 3445.835 4312.000 ;
        RECT 3445.135 4165.330 3445.835 4166.035 ;
      LAYER met4 ;
        RECT 3446.235 4165.730 3450.685 4313.270 ;
      LAYER met4 ;
        RECT 3451.085 4313.030 3451.685 4313.670 ;
        RECT 3451.085 4167.000 3451.685 4312.000 ;
        RECT 3451.085 4165.330 3451.685 4166.035 ;
      LAYER met4 ;
        RECT 3452.085 4165.730 3456.535 4313.270 ;
      LAYER met4 ;
        RECT 3456.935 4313.030 3457.635 4313.670 ;
        RECT 3456.935 4167.000 3457.635 4312.000 ;
        RECT 3456.935 4165.330 3457.635 4166.035 ;
      LAYER met4 ;
        RECT 3458.035 4165.730 3483.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4313.030 3563.385 4313.670 ;
      LAYER met4 ;
        RECT 3563.785 4312.000 3588.000 4313.270 ;
      LAYER met4 ;
        RECT 3483.400 4167.000 3588.000 4312.000 ;
        RECT 3483.400 4165.330 3563.385 4166.035 ;
      LAYER met4 ;
        RECT 3563.785 4165.730 3588.000 4167.000 ;
      LAYER met4 ;
        RECT 3445.135 4093.670 3588.000 4165.330 ;
        RECT 3445.135 4092.965 3445.835 4093.670 ;
        RECT 3445.135 3946.000 3445.835 4092.000 ;
        RECT 3445.135 3944.330 3445.835 3945.035 ;
      LAYER met4 ;
        RECT 3446.235 3944.730 3450.685 4093.270 ;
      LAYER met4 ;
        RECT 3451.085 4092.965 3451.685 4093.670 ;
        RECT 3451.085 3946.000 3451.685 4092.000 ;
        RECT 3451.085 3944.330 3451.685 3945.035 ;
      LAYER met4 ;
        RECT 3452.085 3944.730 3456.535 4093.270 ;
      LAYER met4 ;
        RECT 3456.935 4092.965 3457.635 4093.670 ;
        RECT 3456.935 3946.000 3457.635 4092.000 ;
        RECT 3456.935 3944.330 3457.635 3945.035 ;
      LAYER met4 ;
        RECT 3458.035 3944.730 3483.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 4092.965 3563.385 4093.670 ;
      LAYER met4 ;
        RECT 3563.785 4092.000 3588.000 4093.270 ;
      LAYER met4 ;
        RECT 3483.400 3946.000 3588.000 4092.000 ;
        RECT 3483.400 3944.330 3563.385 3945.035 ;
      LAYER met4 ;
        RECT 3563.785 3944.730 3588.000 3946.000 ;
      LAYER met4 ;
        RECT 3445.135 3942.990 3588.000 3944.330 ;
        RECT 3444.505 3909.160 3588.000 3942.990 ;
        RECT 3439.745 3907.640 3588.000 3909.160 ;
        RECT 3439.745 3893.455 3440.725 3907.640 ;
        RECT 3436.465 3891.935 3440.725 3893.455 ;
        RECT 3388.535 3674.310 3435.965 3717.990 ;
        RECT 3388.535 3642.670 3435.335 3674.310 ;
        RECT 3388.535 3642.030 3389.635 3642.670 ;
        RECT 198.365 3568.330 199.465 3568.970 ;
        RECT 152.665 3536.690 199.465 3568.330 ;
        RECT 152.035 3493.010 199.465 3536.690 ;
        RECT 147.275 3326.545 151.535 3328.065 ;
        RECT 147.275 3312.360 148.255 3326.545 ;
        RECT 0.000 3310.840 148.255 3312.360 ;
        RECT 0.000 3277.010 143.495 3310.840 ;
        RECT 0.000 3275.670 142.865 3277.010 ;
      LAYER met4 ;
        RECT 0.000 3274.000 24.215 3275.270 ;
      LAYER met4 ;
        RECT 24.615 3274.965 104.600 3275.670 ;
        RECT 0.000 3138.000 104.600 3274.000 ;
      LAYER met4 ;
        RECT 0.000 3136.730 24.215 3138.000 ;
      LAYER met4 ;
        RECT 24.615 3136.330 104.600 3136.970 ;
      LAYER met4 ;
        RECT 105.000 3136.730 129.965 3275.270 ;
      LAYER met4 ;
        RECT 130.365 3274.965 131.065 3275.670 ;
        RECT 130.365 3138.000 131.065 3274.000 ;
        RECT 130.365 3136.330 131.065 3136.970 ;
      LAYER met4 ;
        RECT 131.465 3136.730 135.915 3275.270 ;
      LAYER met4 ;
        RECT 136.315 3274.965 136.915 3275.670 ;
        RECT 136.315 3138.000 136.915 3274.000 ;
        RECT 136.315 3136.330 136.915 3136.970 ;
      LAYER met4 ;
        RECT 137.315 3136.730 141.765 3275.270 ;
      LAYER met4 ;
        RECT 142.165 3274.965 142.865 3275.670 ;
        RECT 142.165 3138.000 142.865 3274.000 ;
        RECT 142.165 3136.330 142.865 3136.970 ;
        RECT 0.000 3104.690 142.865 3136.330 ;
      LAYER met4 ;
        RECT 143.265 3105.090 143.595 3276.610 ;
      LAYER met4 ;
        RECT 0.000 3096.360 143.495 3104.690 ;
      LAYER met4 ;
        RECT 143.895 3096.760 146.875 3310.440 ;
      LAYER met4 ;
        RECT 147.275 3275.670 148.255 3310.840 ;
      LAYER met4 ;
        RECT 147.175 3274.000 148.355 3275.270 ;
      LAYER met4 ;
        RECT 147.175 3138.000 148.355 3274.000 ;
      LAYER met4 ;
        RECT 147.175 3136.730 148.355 3138.000 ;
      LAYER met4 ;
        RECT 147.275 3112.065 148.255 3136.330 ;
      LAYER met4 ;
        RECT 148.655 3112.465 151.635 3326.145 ;
        RECT 151.935 3321.090 152.265 3492.610 ;
      LAYER met4 ;
        RECT 152.665 3491.670 199.465 3493.010 ;
        RECT 152.665 3490.965 153.365 3491.670 ;
        RECT 152.665 3352.330 153.365 3352.970 ;
      LAYER met4 ;
        RECT 153.765 3352.730 158.415 3491.270 ;
      LAYER met4 ;
        RECT 158.815 3490.965 159.415 3491.670 ;
        RECT 158.815 3352.330 159.415 3352.970 ;
      LAYER met4 ;
        RECT 159.815 3352.730 163.265 3491.270 ;
      LAYER met4 ;
        RECT 163.665 3490.965 164.265 3491.670 ;
        RECT 163.665 3352.330 164.265 3352.970 ;
      LAYER met4 ;
        RECT 164.665 3352.730 168.115 3491.270 ;
      LAYER met4 ;
        RECT 168.515 3490.965 169.115 3491.670 ;
        RECT 168.515 3352.330 169.115 3352.970 ;
      LAYER met4 ;
        RECT 169.515 3352.730 174.165 3491.270 ;
      LAYER met4 ;
        RECT 174.565 3490.965 175.165 3491.670 ;
        RECT 180.615 3491.365 186.065 3491.670 ;
        RECT 174.565 3352.330 175.165 3352.970 ;
      LAYER met4 ;
        RECT 175.565 3352.730 180.215 3491.270 ;
      LAYER met4 ;
        RECT 180.615 3490.965 181.215 3491.365 ;
        RECT 185.465 3490.965 186.065 3491.365 ;
      LAYER met4 ;
        RECT 181.615 3352.970 185.065 3490.965 ;
      LAYER met4 ;
        RECT 180.615 3352.570 181.215 3352.970 ;
        RECT 185.465 3352.570 186.065 3352.970 ;
      LAYER met4 ;
        RECT 186.465 3352.730 191.115 3491.270 ;
      LAYER met4 ;
        RECT 191.515 3490.965 192.115 3491.670 ;
        RECT 180.615 3352.330 186.065 3352.570 ;
        RECT 191.515 3352.330 192.115 3352.970 ;
      LAYER met4 ;
        RECT 192.515 3352.730 197.965 3491.270 ;
      LAYER met4 ;
        RECT 198.365 3490.965 199.465 3491.670 ;
        RECT 3388.535 3494.330 3389.635 3495.035 ;
      LAYER met4 ;
        RECT 3390.035 3494.730 3395.485 3642.270 ;
      LAYER met4 ;
        RECT 3395.885 3642.030 3396.485 3642.670 ;
        RECT 3401.935 3642.430 3407.385 3642.670 ;
        RECT 3395.885 3494.330 3396.485 3495.035 ;
      LAYER met4 ;
        RECT 3396.885 3494.730 3401.535 3642.270 ;
      LAYER met4 ;
        RECT 3401.935 3642.030 3402.535 3642.430 ;
        RECT 3406.785 3642.030 3407.385 3642.430 ;
      LAYER met4 ;
        RECT 3402.935 3495.035 3406.385 3642.030 ;
      LAYER met4 ;
        RECT 3401.935 3494.635 3402.535 3495.035 ;
        RECT 3406.785 3494.635 3407.385 3495.035 ;
      LAYER met4 ;
        RECT 3407.785 3494.730 3412.435 3642.270 ;
      LAYER met4 ;
        RECT 3412.835 3642.030 3413.435 3642.670 ;
        RECT 3401.935 3494.330 3407.385 3494.635 ;
        RECT 3412.835 3494.330 3413.435 3495.035 ;
      LAYER met4 ;
        RECT 3413.835 3494.730 3418.485 3642.270 ;
      LAYER met4 ;
        RECT 3418.885 3642.030 3419.485 3642.670 ;
        RECT 3418.885 3494.330 3419.485 3495.035 ;
      LAYER met4 ;
        RECT 3419.885 3494.730 3423.335 3642.270 ;
      LAYER met4 ;
        RECT 3423.735 3642.030 3424.335 3642.670 ;
        RECT 3423.735 3494.330 3424.335 3495.035 ;
      LAYER met4 ;
        RECT 3424.735 3494.730 3428.185 3642.270 ;
      LAYER met4 ;
        RECT 3428.585 3642.030 3429.185 3642.670 ;
        RECT 3428.585 3494.330 3429.185 3495.035 ;
      LAYER met4 ;
        RECT 3429.585 3494.730 3434.235 3642.270 ;
      LAYER met4 ;
        RECT 3434.635 3642.030 3435.335 3642.670 ;
        RECT 3434.635 3494.330 3435.335 3495.035 ;
        RECT 3388.535 3492.990 3435.335 3494.330 ;
      LAYER met4 ;
        RECT 3435.735 3493.390 3436.065 3673.910 ;
        RECT 3436.365 3668.855 3439.345 3891.535 ;
      LAYER met4 ;
        RECT 3439.745 3867.670 3440.725 3891.935 ;
      LAYER met4 ;
        RECT 3439.645 3866.000 3440.825 3867.270 ;
      LAYER met4 ;
        RECT 3439.645 3721.000 3440.825 3866.000 ;
      LAYER met4 ;
        RECT 3439.645 3719.730 3440.825 3721.000 ;
      LAYER met4 ;
        RECT 3439.745 3684.160 3440.725 3719.330 ;
      LAYER met4 ;
        RECT 3441.125 3684.560 3444.105 3907.240 ;
      LAYER met4 ;
        RECT 3444.505 3899.310 3588.000 3907.640 ;
      LAYER met4 ;
        RECT 3444.405 3718.390 3444.735 3898.910 ;
      LAYER met4 ;
        RECT 3445.135 3867.670 3588.000 3899.310 ;
        RECT 3445.135 3867.030 3445.835 3867.670 ;
        RECT 3445.135 3721.000 3445.835 3866.000 ;
        RECT 3445.135 3719.330 3445.835 3720.035 ;
      LAYER met4 ;
        RECT 3446.235 3719.730 3450.685 3867.270 ;
      LAYER met4 ;
        RECT 3451.085 3867.030 3451.685 3867.670 ;
        RECT 3451.085 3721.000 3451.685 3866.000 ;
        RECT 3451.085 3719.330 3451.685 3720.035 ;
      LAYER met4 ;
        RECT 3452.085 3719.730 3456.535 3867.270 ;
      LAYER met4 ;
        RECT 3456.935 3867.030 3457.635 3867.670 ;
        RECT 3456.935 3721.000 3457.635 3866.000 ;
        RECT 3456.935 3719.330 3457.635 3720.035 ;
      LAYER met4 ;
        RECT 3458.035 3719.730 3483.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3867.030 3563.385 3867.670 ;
      LAYER met4 ;
        RECT 3563.785 3866.000 3588.000 3867.270 ;
      LAYER met4 ;
        RECT 3483.400 3721.000 3588.000 3866.000 ;
        RECT 3483.400 3719.330 3563.385 3720.035 ;
      LAYER met4 ;
        RECT 3563.785 3719.730 3588.000 3721.000 ;
      LAYER met4 ;
        RECT 3445.135 3717.990 3588.000 3719.330 ;
        RECT 3444.505 3684.160 3588.000 3717.990 ;
        RECT 3439.745 3682.640 3588.000 3684.160 ;
        RECT 3439.745 3668.455 3440.725 3682.640 ;
        RECT 3436.465 3666.935 3440.725 3668.455 ;
        RECT 3388.535 3449.310 3435.965 3492.990 ;
        RECT 3388.535 3417.670 3435.335 3449.310 ;
        RECT 3388.535 3417.030 3389.635 3417.670 ;
        RECT 198.365 3352.330 199.465 3352.970 ;
        RECT 152.665 3320.690 199.465 3352.330 ;
        RECT 152.035 3277.010 199.465 3320.690 ;
        RECT 147.275 3110.545 151.535 3112.065 ;
        RECT 147.275 3096.360 148.255 3110.545 ;
        RECT 0.000 3094.840 148.255 3096.360 ;
        RECT 0.000 3061.010 143.495 3094.840 ;
        RECT 0.000 3059.670 142.865 3061.010 ;
      LAYER met4 ;
        RECT 0.000 3058.000 24.215 3059.270 ;
      LAYER met4 ;
        RECT 24.615 3058.965 104.600 3059.670 ;
        RECT 0.000 2922.000 104.600 3058.000 ;
      LAYER met4 ;
        RECT 0.000 2920.730 24.215 2922.000 ;
      LAYER met4 ;
        RECT 24.615 2920.330 104.600 2920.970 ;
      LAYER met4 ;
        RECT 105.000 2920.730 129.965 3059.270 ;
      LAYER met4 ;
        RECT 130.365 3058.965 131.065 3059.670 ;
        RECT 130.365 2922.000 131.065 3058.000 ;
        RECT 130.365 2920.330 131.065 2920.970 ;
      LAYER met4 ;
        RECT 131.465 2920.730 135.915 3059.270 ;
      LAYER met4 ;
        RECT 136.315 3058.965 136.915 3059.670 ;
        RECT 136.315 2922.000 136.915 3058.000 ;
        RECT 136.315 2920.330 136.915 2920.970 ;
      LAYER met4 ;
        RECT 137.315 2920.730 141.765 3059.270 ;
      LAYER met4 ;
        RECT 142.165 3058.965 142.865 3059.670 ;
        RECT 142.165 2922.000 142.865 3058.000 ;
        RECT 142.165 2920.330 142.865 2920.970 ;
        RECT 0.000 2888.690 142.865 2920.330 ;
      LAYER met4 ;
        RECT 143.265 2889.090 143.595 3060.610 ;
      LAYER met4 ;
        RECT 0.000 2880.360 143.495 2888.690 ;
      LAYER met4 ;
        RECT 143.895 2880.760 146.875 3094.440 ;
      LAYER met4 ;
        RECT 147.275 3059.670 148.255 3094.840 ;
      LAYER met4 ;
        RECT 147.175 3058.000 148.355 3059.270 ;
      LAYER met4 ;
        RECT 147.175 2922.000 148.355 3058.000 ;
      LAYER met4 ;
        RECT 147.175 2920.730 148.355 2922.000 ;
      LAYER met4 ;
        RECT 147.275 2896.065 148.255 2920.330 ;
      LAYER met4 ;
        RECT 148.655 2896.465 151.635 3110.145 ;
        RECT 151.935 3105.090 152.265 3276.610 ;
      LAYER met4 ;
        RECT 152.665 3275.670 199.465 3277.010 ;
        RECT 152.665 3274.965 153.365 3275.670 ;
        RECT 152.665 3136.330 153.365 3136.970 ;
      LAYER met4 ;
        RECT 153.765 3136.730 158.415 3275.270 ;
      LAYER met4 ;
        RECT 158.815 3274.965 159.415 3275.670 ;
        RECT 158.815 3136.330 159.415 3136.970 ;
      LAYER met4 ;
        RECT 159.815 3136.730 163.265 3275.270 ;
      LAYER met4 ;
        RECT 163.665 3274.965 164.265 3275.670 ;
        RECT 163.665 3136.330 164.265 3136.970 ;
      LAYER met4 ;
        RECT 164.665 3136.730 168.115 3275.270 ;
      LAYER met4 ;
        RECT 168.515 3274.965 169.115 3275.670 ;
        RECT 168.515 3136.330 169.115 3136.970 ;
      LAYER met4 ;
        RECT 169.515 3136.730 174.165 3275.270 ;
      LAYER met4 ;
        RECT 174.565 3274.965 175.165 3275.670 ;
        RECT 180.615 3275.365 186.065 3275.670 ;
        RECT 174.565 3136.330 175.165 3136.970 ;
      LAYER met4 ;
        RECT 175.565 3136.730 180.215 3275.270 ;
      LAYER met4 ;
        RECT 180.615 3274.965 181.215 3275.365 ;
        RECT 185.465 3274.965 186.065 3275.365 ;
      LAYER met4 ;
        RECT 181.615 3136.970 185.065 3274.965 ;
      LAYER met4 ;
        RECT 180.615 3136.570 181.215 3136.970 ;
        RECT 185.465 3136.570 186.065 3136.970 ;
      LAYER met4 ;
        RECT 186.465 3136.730 191.115 3275.270 ;
      LAYER met4 ;
        RECT 191.515 3274.965 192.115 3275.670 ;
        RECT 180.615 3136.330 186.065 3136.570 ;
        RECT 191.515 3136.330 192.115 3136.970 ;
      LAYER met4 ;
        RECT 192.515 3136.730 197.965 3275.270 ;
      LAYER met4 ;
        RECT 198.365 3274.965 199.465 3275.670 ;
        RECT 3388.535 3268.330 3389.635 3269.035 ;
      LAYER met4 ;
        RECT 3390.035 3268.730 3395.485 3417.270 ;
      LAYER met4 ;
        RECT 3395.885 3417.030 3396.485 3417.670 ;
        RECT 3401.935 3417.430 3407.385 3417.670 ;
        RECT 3395.885 3268.330 3396.485 3269.035 ;
      LAYER met4 ;
        RECT 3396.885 3268.730 3401.535 3417.270 ;
      LAYER met4 ;
        RECT 3401.935 3417.030 3402.535 3417.430 ;
        RECT 3406.785 3417.030 3407.385 3417.430 ;
      LAYER met4 ;
        RECT 3402.935 3269.035 3406.385 3417.030 ;
      LAYER met4 ;
        RECT 3401.935 3268.635 3402.535 3269.035 ;
        RECT 3406.785 3268.635 3407.385 3269.035 ;
      LAYER met4 ;
        RECT 3407.785 3268.730 3412.435 3417.270 ;
      LAYER met4 ;
        RECT 3412.835 3417.030 3413.435 3417.670 ;
        RECT 3401.935 3268.330 3407.385 3268.635 ;
        RECT 3412.835 3268.330 3413.435 3269.035 ;
      LAYER met4 ;
        RECT 3413.835 3268.730 3418.485 3417.270 ;
      LAYER met4 ;
        RECT 3418.885 3417.030 3419.485 3417.670 ;
        RECT 3418.885 3268.330 3419.485 3269.035 ;
      LAYER met4 ;
        RECT 3419.885 3268.730 3423.335 3417.270 ;
      LAYER met4 ;
        RECT 3423.735 3417.030 3424.335 3417.670 ;
        RECT 3423.735 3268.330 3424.335 3269.035 ;
      LAYER met4 ;
        RECT 3424.735 3268.730 3428.185 3417.270 ;
      LAYER met4 ;
        RECT 3428.585 3417.030 3429.185 3417.670 ;
        RECT 3428.585 3268.330 3429.185 3269.035 ;
      LAYER met4 ;
        RECT 3429.585 3268.730 3434.235 3417.270 ;
      LAYER met4 ;
        RECT 3434.635 3417.030 3435.335 3417.670 ;
        RECT 3434.635 3268.330 3435.335 3269.035 ;
        RECT 3388.535 3266.990 3435.335 3268.330 ;
      LAYER met4 ;
        RECT 3435.735 3267.390 3436.065 3448.910 ;
        RECT 3436.365 3443.855 3439.345 3666.535 ;
      LAYER met4 ;
        RECT 3439.745 3642.670 3440.725 3666.935 ;
      LAYER met4 ;
        RECT 3439.645 3641.000 3440.825 3642.270 ;
      LAYER met4 ;
        RECT 3439.645 3496.000 3440.825 3641.000 ;
      LAYER met4 ;
        RECT 3439.645 3494.730 3440.825 3496.000 ;
      LAYER met4 ;
        RECT 3439.745 3459.160 3440.725 3494.330 ;
      LAYER met4 ;
        RECT 3441.125 3459.560 3444.105 3682.240 ;
      LAYER met4 ;
        RECT 3444.505 3674.310 3588.000 3682.640 ;
      LAYER met4 ;
        RECT 3444.405 3493.390 3444.735 3673.910 ;
      LAYER met4 ;
        RECT 3445.135 3642.670 3588.000 3674.310 ;
        RECT 3445.135 3642.030 3445.835 3642.670 ;
        RECT 3445.135 3496.000 3445.835 3641.000 ;
        RECT 3445.135 3494.330 3445.835 3495.035 ;
      LAYER met4 ;
        RECT 3446.235 3494.730 3450.685 3642.270 ;
      LAYER met4 ;
        RECT 3451.085 3642.030 3451.685 3642.670 ;
        RECT 3451.085 3496.000 3451.685 3641.000 ;
        RECT 3451.085 3494.330 3451.685 3495.035 ;
      LAYER met4 ;
        RECT 3452.085 3494.730 3456.535 3642.270 ;
      LAYER met4 ;
        RECT 3456.935 3642.030 3457.635 3642.670 ;
        RECT 3456.935 3496.000 3457.635 3641.000 ;
        RECT 3456.935 3494.330 3457.635 3495.035 ;
      LAYER met4 ;
        RECT 3458.035 3494.730 3483.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3642.030 3563.385 3642.670 ;
      LAYER met4 ;
        RECT 3563.785 3641.000 3588.000 3642.270 ;
      LAYER met4 ;
        RECT 3483.400 3496.000 3588.000 3641.000 ;
        RECT 3483.400 3494.330 3563.385 3495.035 ;
      LAYER met4 ;
        RECT 3563.785 3494.730 3588.000 3496.000 ;
      LAYER met4 ;
        RECT 3445.135 3492.990 3588.000 3494.330 ;
        RECT 3444.505 3459.160 3588.000 3492.990 ;
        RECT 3439.745 3457.640 3588.000 3459.160 ;
        RECT 3439.745 3443.455 3440.725 3457.640 ;
        RECT 3436.465 3441.935 3440.725 3443.455 ;
        RECT 3388.535 3223.310 3435.965 3266.990 ;
        RECT 3388.535 3191.670 3435.335 3223.310 ;
        RECT 3388.535 3191.030 3389.635 3191.670 ;
        RECT 198.365 3136.330 199.465 3136.970 ;
        RECT 152.665 3104.690 199.465 3136.330 ;
        RECT 152.035 3061.010 199.465 3104.690 ;
        RECT 147.275 2894.545 151.535 2896.065 ;
        RECT 147.275 2880.360 148.255 2894.545 ;
        RECT 0.000 2878.840 148.255 2880.360 ;
        RECT 0.000 2845.010 143.495 2878.840 ;
        RECT 0.000 2843.670 142.865 2845.010 ;
      LAYER met4 ;
        RECT 0.000 2842.000 24.215 2843.270 ;
      LAYER met4 ;
        RECT 24.615 2842.965 104.600 2843.670 ;
        RECT 0.000 2706.000 104.600 2842.000 ;
      LAYER met4 ;
        RECT 0.000 2704.730 24.215 2706.000 ;
      LAYER met4 ;
        RECT 24.615 2704.330 104.600 2704.970 ;
      LAYER met4 ;
        RECT 105.000 2704.730 129.965 2843.270 ;
      LAYER met4 ;
        RECT 130.365 2842.965 131.065 2843.670 ;
        RECT 130.365 2706.000 131.065 2842.000 ;
        RECT 130.365 2704.330 131.065 2704.970 ;
      LAYER met4 ;
        RECT 131.465 2704.730 135.915 2843.270 ;
      LAYER met4 ;
        RECT 136.315 2842.965 136.915 2843.670 ;
        RECT 136.315 2706.000 136.915 2842.000 ;
        RECT 136.315 2704.330 136.915 2704.970 ;
      LAYER met4 ;
        RECT 137.315 2704.730 141.765 2843.270 ;
      LAYER met4 ;
        RECT 142.165 2842.965 142.865 2843.670 ;
        RECT 142.165 2706.000 142.865 2842.000 ;
        RECT 142.165 2704.330 142.865 2704.970 ;
        RECT 0.000 2672.690 142.865 2704.330 ;
      LAYER met4 ;
        RECT 143.265 2673.090 143.595 2844.610 ;
      LAYER met4 ;
        RECT 0.000 2664.360 143.495 2672.690 ;
      LAYER met4 ;
        RECT 143.895 2664.760 146.875 2878.440 ;
      LAYER met4 ;
        RECT 147.275 2843.670 148.255 2878.840 ;
      LAYER met4 ;
        RECT 147.175 2842.000 148.355 2843.270 ;
      LAYER met4 ;
        RECT 147.175 2706.000 148.355 2842.000 ;
      LAYER met4 ;
        RECT 147.175 2704.730 148.355 2706.000 ;
      LAYER met4 ;
        RECT 147.275 2680.065 148.255 2704.330 ;
      LAYER met4 ;
        RECT 148.655 2680.465 151.635 2894.145 ;
        RECT 151.935 2889.090 152.265 3060.610 ;
      LAYER met4 ;
        RECT 152.665 3059.670 199.465 3061.010 ;
        RECT 152.665 3058.965 153.365 3059.670 ;
        RECT 152.665 2920.330 153.365 2920.970 ;
      LAYER met4 ;
        RECT 153.765 2920.730 158.415 3059.270 ;
      LAYER met4 ;
        RECT 158.815 3058.965 159.415 3059.670 ;
        RECT 158.815 2920.330 159.415 2920.970 ;
      LAYER met4 ;
        RECT 159.815 2920.730 163.265 3059.270 ;
      LAYER met4 ;
        RECT 163.665 3058.965 164.265 3059.670 ;
        RECT 163.665 2920.330 164.265 2920.970 ;
      LAYER met4 ;
        RECT 164.665 2920.730 168.115 3059.270 ;
      LAYER met4 ;
        RECT 168.515 3058.965 169.115 3059.670 ;
        RECT 168.515 2920.330 169.115 2920.970 ;
      LAYER met4 ;
        RECT 169.515 2920.730 174.165 3059.270 ;
      LAYER met4 ;
        RECT 174.565 3058.965 175.165 3059.670 ;
        RECT 180.615 3059.365 186.065 3059.670 ;
        RECT 174.565 2920.330 175.165 2920.970 ;
      LAYER met4 ;
        RECT 175.565 2920.730 180.215 3059.270 ;
      LAYER met4 ;
        RECT 180.615 3058.965 181.215 3059.365 ;
        RECT 185.465 3058.965 186.065 3059.365 ;
      LAYER met4 ;
        RECT 181.615 2920.970 185.065 3058.965 ;
      LAYER met4 ;
        RECT 180.615 2920.570 181.215 2920.970 ;
        RECT 185.465 2920.570 186.065 2920.970 ;
      LAYER met4 ;
        RECT 186.465 2920.730 191.115 3059.270 ;
      LAYER met4 ;
        RECT 191.515 3058.965 192.115 3059.670 ;
        RECT 180.615 2920.330 186.065 2920.570 ;
        RECT 191.515 2920.330 192.115 2920.970 ;
      LAYER met4 ;
        RECT 192.515 2920.730 197.965 3059.270 ;
      LAYER met4 ;
        RECT 198.365 3058.965 199.465 3059.670 ;
        RECT 3388.535 3043.330 3389.635 3044.035 ;
      LAYER met4 ;
        RECT 3390.035 3043.730 3395.485 3191.270 ;
      LAYER met4 ;
        RECT 3395.885 3191.030 3396.485 3191.670 ;
        RECT 3401.935 3191.430 3407.385 3191.670 ;
        RECT 3395.885 3043.330 3396.485 3044.035 ;
      LAYER met4 ;
        RECT 3396.885 3043.730 3401.535 3191.270 ;
      LAYER met4 ;
        RECT 3401.935 3191.030 3402.535 3191.430 ;
        RECT 3406.785 3191.030 3407.385 3191.430 ;
      LAYER met4 ;
        RECT 3402.935 3044.035 3406.385 3191.030 ;
      LAYER met4 ;
        RECT 3401.935 3043.635 3402.535 3044.035 ;
        RECT 3406.785 3043.635 3407.385 3044.035 ;
      LAYER met4 ;
        RECT 3407.785 3043.730 3412.435 3191.270 ;
      LAYER met4 ;
        RECT 3412.835 3191.030 3413.435 3191.670 ;
        RECT 3401.935 3043.330 3407.385 3043.635 ;
        RECT 3412.835 3043.330 3413.435 3044.035 ;
      LAYER met4 ;
        RECT 3413.835 3043.730 3418.485 3191.270 ;
      LAYER met4 ;
        RECT 3418.885 3191.030 3419.485 3191.670 ;
        RECT 3418.885 3043.330 3419.485 3044.035 ;
      LAYER met4 ;
        RECT 3419.885 3043.730 3423.335 3191.270 ;
      LAYER met4 ;
        RECT 3423.735 3191.030 3424.335 3191.670 ;
        RECT 3423.735 3043.330 3424.335 3044.035 ;
      LAYER met4 ;
        RECT 3424.735 3043.730 3428.185 3191.270 ;
      LAYER met4 ;
        RECT 3428.585 3191.030 3429.185 3191.670 ;
        RECT 3428.585 3043.330 3429.185 3044.035 ;
      LAYER met4 ;
        RECT 3429.585 3043.730 3434.235 3191.270 ;
      LAYER met4 ;
        RECT 3434.635 3191.030 3435.335 3191.670 ;
        RECT 3434.635 3043.330 3435.335 3044.035 ;
        RECT 3388.535 3041.990 3435.335 3043.330 ;
      LAYER met4 ;
        RECT 3435.735 3042.390 3436.065 3222.910 ;
        RECT 3436.365 3217.855 3439.345 3441.535 ;
      LAYER met4 ;
        RECT 3439.745 3417.670 3440.725 3441.935 ;
      LAYER met4 ;
        RECT 3439.645 3416.000 3440.825 3417.270 ;
      LAYER met4 ;
        RECT 3439.645 3270.000 3440.825 3416.000 ;
      LAYER met4 ;
        RECT 3439.645 3268.730 3440.825 3270.000 ;
      LAYER met4 ;
        RECT 3439.745 3233.160 3440.725 3268.330 ;
      LAYER met4 ;
        RECT 3441.125 3233.560 3444.105 3457.240 ;
      LAYER met4 ;
        RECT 3444.505 3449.310 3588.000 3457.640 ;
      LAYER met4 ;
        RECT 3444.405 3267.390 3444.735 3448.910 ;
      LAYER met4 ;
        RECT 3445.135 3417.670 3588.000 3449.310 ;
        RECT 3445.135 3417.030 3445.835 3417.670 ;
        RECT 3445.135 3270.000 3445.835 3416.000 ;
        RECT 3445.135 3268.330 3445.835 3269.035 ;
      LAYER met4 ;
        RECT 3446.235 3268.730 3450.685 3417.270 ;
      LAYER met4 ;
        RECT 3451.085 3417.030 3451.685 3417.670 ;
        RECT 3451.085 3270.000 3451.685 3416.000 ;
        RECT 3451.085 3268.330 3451.685 3269.035 ;
      LAYER met4 ;
        RECT 3452.085 3268.730 3456.535 3417.270 ;
      LAYER met4 ;
        RECT 3456.935 3417.030 3457.635 3417.670 ;
        RECT 3456.935 3270.000 3457.635 3416.000 ;
        RECT 3456.935 3268.330 3457.635 3269.035 ;
      LAYER met4 ;
        RECT 3458.035 3268.730 3483.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3417.030 3563.385 3417.670 ;
      LAYER met4 ;
        RECT 3563.785 3416.000 3588.000 3417.270 ;
      LAYER met4 ;
        RECT 3483.400 3270.000 3588.000 3416.000 ;
        RECT 3483.400 3268.330 3563.385 3269.035 ;
      LAYER met4 ;
        RECT 3563.785 3268.730 3588.000 3270.000 ;
      LAYER met4 ;
        RECT 3445.135 3266.990 3588.000 3268.330 ;
        RECT 3444.505 3233.160 3588.000 3266.990 ;
        RECT 3439.745 3231.640 3588.000 3233.160 ;
        RECT 3439.745 3217.455 3440.725 3231.640 ;
        RECT 3436.465 3215.935 3440.725 3217.455 ;
        RECT 3388.535 2998.310 3435.965 3041.990 ;
        RECT 3388.535 2966.670 3435.335 2998.310 ;
        RECT 3388.535 2966.030 3389.635 2966.670 ;
        RECT 198.365 2920.330 199.465 2920.970 ;
        RECT 152.665 2888.690 199.465 2920.330 ;
        RECT 152.035 2845.010 199.465 2888.690 ;
        RECT 147.275 2678.545 151.535 2680.065 ;
        RECT 147.275 2664.360 148.255 2678.545 ;
        RECT 0.000 2662.840 148.255 2664.360 ;
        RECT 0.000 2629.010 143.495 2662.840 ;
        RECT 0.000 2627.670 142.865 2629.010 ;
      LAYER met4 ;
        RECT 0.000 2626.000 24.215 2627.270 ;
      LAYER met4 ;
        RECT 24.615 2626.965 104.600 2627.670 ;
        RECT 0.000 2490.000 104.600 2626.000 ;
      LAYER met4 ;
        RECT 0.000 2488.730 24.215 2490.000 ;
      LAYER met4 ;
        RECT 24.615 2488.330 104.600 2489.035 ;
      LAYER met4 ;
        RECT 105.000 2488.730 129.965 2627.270 ;
      LAYER met4 ;
        RECT 130.365 2626.965 131.065 2627.670 ;
        RECT 130.365 2490.000 131.065 2626.000 ;
        RECT 130.365 2488.330 131.065 2489.035 ;
      LAYER met4 ;
        RECT 131.465 2488.730 135.915 2627.270 ;
      LAYER met4 ;
        RECT 136.315 2626.965 136.915 2627.670 ;
        RECT 136.315 2490.000 136.915 2626.000 ;
        RECT 136.315 2488.330 136.915 2489.035 ;
      LAYER met4 ;
        RECT 137.315 2488.730 141.765 2627.270 ;
      LAYER met4 ;
        RECT 142.165 2626.965 142.865 2627.670 ;
        RECT 142.165 2490.000 142.865 2626.000 ;
        RECT 142.165 2488.330 142.865 2489.035 ;
        RECT 0.000 2416.670 142.865 2488.330 ;
      LAYER met4 ;
        RECT 0.000 2415.000 24.215 2416.270 ;
      LAYER met4 ;
        RECT 24.615 2415.965 104.600 2416.670 ;
        RECT 0.000 2280.465 104.600 2415.000 ;
        RECT 0.000 2279.000 0.035 2280.465 ;
        RECT 24.215 2279.000 104.600 2280.465 ;
        RECT 24.215 2278.785 24.250 2279.000 ;
        RECT 24.615 2277.330 104.600 2279.000 ;
      LAYER met4 ;
        RECT 105.000 2277.730 129.965 2416.270 ;
      LAYER met4 ;
        RECT 130.365 2415.965 131.065 2416.670 ;
        RECT 130.365 2277.330 131.065 2415.000 ;
      LAYER met4 ;
        RECT 131.465 2277.730 135.915 2416.270 ;
      LAYER met4 ;
        RECT 136.315 2415.965 136.915 2416.670 ;
        RECT 136.315 2277.330 136.915 2415.000 ;
      LAYER met4 ;
        RECT 137.315 2277.730 141.765 2416.270 ;
      LAYER met4 ;
        RECT 142.165 2415.965 142.865 2416.670 ;
        RECT 142.165 2277.330 142.865 2415.000 ;
        RECT 0.000 2205.670 142.865 2277.330 ;
      LAYER met4 ;
        RECT 0.000 2204.000 24.215 2205.270 ;
      LAYER met4 ;
        RECT 24.615 2204.000 104.600 2205.670 ;
        RECT 0.000 2068.000 104.600 2204.000 ;
      LAYER met4 ;
        RECT 0.000 2066.730 24.215 2068.000 ;
      LAYER met4 ;
        RECT 24.615 2066.330 104.600 2066.970 ;
      LAYER met4 ;
        RECT 105.000 2066.730 129.965 2205.270 ;
      LAYER met4 ;
        RECT 130.365 2068.000 131.065 2205.670 ;
        RECT 130.365 2066.330 131.065 2066.970 ;
      LAYER met4 ;
        RECT 131.465 2066.730 135.915 2205.270 ;
      LAYER met4 ;
        RECT 136.315 2068.000 136.915 2205.670 ;
        RECT 136.315 2066.330 136.915 2066.970 ;
      LAYER met4 ;
        RECT 137.315 2066.730 141.765 2205.270 ;
      LAYER met4 ;
        RECT 142.165 2068.000 142.865 2205.670 ;
        RECT 142.165 2066.330 142.865 2066.970 ;
        RECT 0.000 2034.690 142.865 2066.330 ;
        RECT 0.000 2026.360 143.495 2034.690 ;
      LAYER met4 ;
        RECT 143.895 2026.760 146.875 2662.440 ;
      LAYER met4 ;
        RECT 147.275 2627.670 148.255 2662.840 ;
      LAYER met4 ;
        RECT 147.175 2626.000 148.355 2627.270 ;
      LAYER met4 ;
        RECT 147.175 2490.000 148.355 2626.000 ;
      LAYER met4 ;
        RECT 147.175 2488.730 148.355 2490.000 ;
      LAYER met4 ;
        RECT 147.275 2416.670 148.255 2488.330 ;
      LAYER met4 ;
        RECT 147.175 2415.000 148.355 2416.270 ;
      LAYER met4 ;
        RECT 147.175 2279.000 148.355 2415.000 ;
      LAYER met4 ;
        RECT 147.175 2277.730 148.355 2279.000 ;
      LAYER met4 ;
        RECT 147.275 2205.670 148.255 2277.330 ;
      LAYER met4 ;
        RECT 147.175 2204.000 148.355 2205.270 ;
      LAYER met4 ;
        RECT 147.175 2068.000 148.355 2204.000 ;
      LAYER met4 ;
        RECT 147.175 2066.730 148.355 2068.000 ;
      LAYER met4 ;
        RECT 147.275 2042.065 148.255 2066.330 ;
      LAYER met4 ;
        RECT 148.655 2042.465 151.635 2678.145 ;
        RECT 151.935 2673.090 152.265 2844.610 ;
      LAYER met4 ;
        RECT 152.665 2843.670 199.465 2845.010 ;
        RECT 152.665 2842.965 153.365 2843.670 ;
        RECT 152.665 2704.330 153.365 2704.970 ;
      LAYER met4 ;
        RECT 153.765 2704.730 158.415 2843.270 ;
      LAYER met4 ;
        RECT 158.815 2842.965 159.415 2843.670 ;
        RECT 158.815 2704.330 159.415 2704.970 ;
      LAYER met4 ;
        RECT 159.815 2704.730 163.265 2843.270 ;
      LAYER met4 ;
        RECT 163.665 2842.965 164.265 2843.670 ;
        RECT 163.665 2704.330 164.265 2704.970 ;
      LAYER met4 ;
        RECT 164.665 2704.730 168.115 2843.270 ;
      LAYER met4 ;
        RECT 168.515 2842.965 169.115 2843.670 ;
        RECT 168.515 2704.330 169.115 2704.970 ;
      LAYER met4 ;
        RECT 169.515 2704.730 174.165 2843.270 ;
      LAYER met4 ;
        RECT 174.565 2842.965 175.165 2843.670 ;
        RECT 180.615 2843.365 186.065 2843.670 ;
        RECT 174.565 2704.330 175.165 2704.970 ;
      LAYER met4 ;
        RECT 175.565 2704.730 180.215 2843.270 ;
      LAYER met4 ;
        RECT 180.615 2842.965 181.215 2843.365 ;
        RECT 185.465 2842.965 186.065 2843.365 ;
      LAYER met4 ;
        RECT 181.615 2704.970 185.065 2842.965 ;
      LAYER met4 ;
        RECT 180.615 2704.570 181.215 2704.970 ;
        RECT 185.465 2704.570 186.065 2704.970 ;
      LAYER met4 ;
        RECT 186.465 2704.730 191.115 2843.270 ;
      LAYER met4 ;
        RECT 191.515 2842.965 192.115 2843.670 ;
        RECT 180.615 2704.330 186.065 2704.570 ;
        RECT 191.515 2704.330 192.115 2704.970 ;
      LAYER met4 ;
        RECT 192.515 2704.730 197.965 2843.270 ;
      LAYER met4 ;
        RECT 198.365 2842.965 199.465 2843.670 ;
        RECT 3388.535 2817.330 3389.635 2818.035 ;
      LAYER met4 ;
        RECT 3390.035 2817.730 3395.485 2966.270 ;
      LAYER met4 ;
        RECT 3395.885 2966.030 3396.485 2966.670 ;
        RECT 3401.935 2966.430 3407.385 2966.670 ;
        RECT 3395.885 2817.330 3396.485 2818.035 ;
      LAYER met4 ;
        RECT 3396.885 2817.730 3401.535 2966.270 ;
      LAYER met4 ;
        RECT 3401.935 2966.030 3402.535 2966.430 ;
        RECT 3406.785 2966.030 3407.385 2966.430 ;
      LAYER met4 ;
        RECT 3402.935 2818.035 3406.385 2966.030 ;
      LAYER met4 ;
        RECT 3401.935 2817.635 3402.535 2818.035 ;
        RECT 3406.785 2817.635 3407.385 2818.035 ;
      LAYER met4 ;
        RECT 3407.785 2817.730 3412.435 2966.270 ;
      LAYER met4 ;
        RECT 3412.835 2966.030 3413.435 2966.670 ;
        RECT 3401.935 2817.330 3407.385 2817.635 ;
        RECT 3412.835 2817.330 3413.435 2818.035 ;
      LAYER met4 ;
        RECT 3413.835 2817.730 3418.485 2966.270 ;
      LAYER met4 ;
        RECT 3418.885 2966.030 3419.485 2966.670 ;
        RECT 3418.885 2817.330 3419.485 2818.035 ;
      LAYER met4 ;
        RECT 3419.885 2817.730 3423.335 2966.270 ;
      LAYER met4 ;
        RECT 3423.735 2966.030 3424.335 2966.670 ;
        RECT 3423.735 2817.330 3424.335 2818.035 ;
      LAYER met4 ;
        RECT 3424.735 2817.730 3428.185 2966.270 ;
      LAYER met4 ;
        RECT 3428.585 2966.030 3429.185 2966.670 ;
        RECT 3428.585 2817.330 3429.185 2818.035 ;
      LAYER met4 ;
        RECT 3429.585 2817.730 3434.235 2966.270 ;
      LAYER met4 ;
        RECT 3434.635 2966.030 3435.335 2966.670 ;
        RECT 3434.635 2817.330 3435.335 2818.035 ;
        RECT 3388.535 2815.990 3435.335 2817.330 ;
      LAYER met4 ;
        RECT 3435.735 2816.390 3436.065 2997.910 ;
        RECT 3436.365 2992.855 3439.345 3215.535 ;
      LAYER met4 ;
        RECT 3439.745 3191.670 3440.725 3215.935 ;
      LAYER met4 ;
        RECT 3439.645 3190.000 3440.825 3191.270 ;
      LAYER met4 ;
        RECT 3439.645 3045.000 3440.825 3190.000 ;
      LAYER met4 ;
        RECT 3439.645 3043.730 3440.825 3045.000 ;
      LAYER met4 ;
        RECT 3439.745 3008.160 3440.725 3043.330 ;
      LAYER met4 ;
        RECT 3441.125 3008.560 3444.105 3231.240 ;
      LAYER met4 ;
        RECT 3444.505 3223.310 3588.000 3231.640 ;
      LAYER met4 ;
        RECT 3444.405 3042.390 3444.735 3222.910 ;
      LAYER met4 ;
        RECT 3445.135 3191.670 3588.000 3223.310 ;
        RECT 3445.135 3191.030 3445.835 3191.670 ;
        RECT 3445.135 3045.000 3445.835 3190.000 ;
        RECT 3445.135 3043.330 3445.835 3044.035 ;
      LAYER met4 ;
        RECT 3446.235 3043.730 3450.685 3191.270 ;
      LAYER met4 ;
        RECT 3451.085 3191.030 3451.685 3191.670 ;
        RECT 3451.085 3045.000 3451.685 3190.000 ;
        RECT 3451.085 3043.330 3451.685 3044.035 ;
      LAYER met4 ;
        RECT 3452.085 3043.730 3456.535 3191.270 ;
      LAYER met4 ;
        RECT 3456.935 3191.030 3457.635 3191.670 ;
        RECT 3456.935 3045.000 3457.635 3190.000 ;
        RECT 3456.935 3043.330 3457.635 3044.035 ;
      LAYER met4 ;
        RECT 3458.035 3043.730 3483.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3191.030 3563.385 3191.670 ;
      LAYER met4 ;
        RECT 3563.785 3190.000 3588.000 3191.270 ;
      LAYER met4 ;
        RECT 3483.400 3045.000 3588.000 3190.000 ;
        RECT 3483.400 3043.330 3563.385 3044.035 ;
      LAYER met4 ;
        RECT 3563.785 3043.730 3588.000 3045.000 ;
      LAYER met4 ;
        RECT 3445.135 3041.990 3588.000 3043.330 ;
        RECT 3444.505 3008.160 3588.000 3041.990 ;
        RECT 3439.745 3006.640 3588.000 3008.160 ;
        RECT 3439.745 2992.455 3440.725 3006.640 ;
        RECT 3436.465 2990.935 3440.725 2992.455 ;
        RECT 3388.535 2772.310 3435.965 2815.990 ;
        RECT 3388.535 2740.670 3435.335 2772.310 ;
        RECT 3388.535 2740.030 3389.635 2740.670 ;
        RECT 198.365 2704.330 199.465 2704.970 ;
        RECT 152.665 2672.690 199.465 2704.330 ;
        RECT 152.035 2629.010 199.465 2672.690 ;
        RECT 147.275 2040.545 151.535 2042.065 ;
        RECT 147.275 2026.360 148.255 2040.545 ;
        RECT 0.000 2024.840 148.255 2026.360 ;
        RECT 0.000 1991.010 143.495 2024.840 ;
        RECT 0.000 1989.670 142.865 1991.010 ;
      LAYER met4 ;
        RECT 0.000 1988.000 24.215 1989.270 ;
      LAYER met4 ;
        RECT 24.615 1988.965 104.600 1989.670 ;
        RECT 0.000 1852.000 104.600 1988.000 ;
      LAYER met4 ;
        RECT 0.000 1850.730 24.215 1852.000 ;
      LAYER met4 ;
        RECT 24.615 1850.330 104.600 1850.970 ;
      LAYER met4 ;
        RECT 105.000 1850.730 129.965 1989.270 ;
      LAYER met4 ;
        RECT 130.365 1988.965 131.065 1989.670 ;
        RECT 130.365 1852.000 131.065 1988.000 ;
        RECT 130.365 1850.330 131.065 1850.970 ;
      LAYER met4 ;
        RECT 131.465 1850.730 135.915 1989.270 ;
      LAYER met4 ;
        RECT 136.315 1988.965 136.915 1989.670 ;
        RECT 136.315 1852.000 136.915 1988.000 ;
        RECT 136.315 1850.330 136.915 1850.970 ;
      LAYER met4 ;
        RECT 137.315 1850.730 141.765 1989.270 ;
      LAYER met4 ;
        RECT 142.165 1988.965 142.865 1989.670 ;
        RECT 142.165 1852.000 142.865 1988.000 ;
        RECT 142.165 1850.330 142.865 1850.970 ;
        RECT 0.000 1818.690 142.865 1850.330 ;
      LAYER met4 ;
        RECT 143.265 1819.090 143.595 1990.610 ;
      LAYER met4 ;
        RECT 0.000 1810.360 143.495 1818.690 ;
      LAYER met4 ;
        RECT 143.895 1810.760 146.875 2024.440 ;
      LAYER met4 ;
        RECT 147.275 1989.670 148.255 2024.840 ;
      LAYER met4 ;
        RECT 147.175 1988.000 148.355 1989.270 ;
      LAYER met4 ;
        RECT 147.175 1852.000 148.355 1988.000 ;
      LAYER met4 ;
        RECT 147.175 1850.730 148.355 1852.000 ;
      LAYER met4 ;
        RECT 147.275 1826.065 148.255 1850.330 ;
      LAYER met4 ;
        RECT 148.655 1826.465 151.635 2040.145 ;
        RECT 151.935 2035.090 152.265 2628.610 ;
      LAYER met4 ;
        RECT 152.665 2627.670 199.465 2629.010 ;
        RECT 152.665 2626.965 153.365 2627.670 ;
        RECT 152.665 2488.330 153.365 2489.035 ;
      LAYER met4 ;
        RECT 153.765 2488.730 158.415 2627.270 ;
      LAYER met4 ;
        RECT 158.815 2626.965 159.415 2627.670 ;
        RECT 158.815 2488.330 159.415 2489.035 ;
      LAYER met4 ;
        RECT 159.815 2488.730 163.265 2627.270 ;
      LAYER met4 ;
        RECT 163.665 2626.965 164.265 2627.670 ;
        RECT 163.665 2488.330 164.265 2489.035 ;
      LAYER met4 ;
        RECT 164.665 2488.730 168.115 2627.270 ;
      LAYER met4 ;
        RECT 168.515 2626.965 169.115 2627.670 ;
        RECT 168.515 2488.330 169.115 2489.035 ;
      LAYER met4 ;
        RECT 169.515 2488.730 174.165 2627.270 ;
      LAYER met4 ;
        RECT 174.565 2626.965 175.165 2627.670 ;
        RECT 180.615 2627.365 186.065 2627.670 ;
        RECT 174.565 2488.330 175.165 2489.035 ;
      LAYER met4 ;
        RECT 175.565 2488.730 180.215 2627.270 ;
      LAYER met4 ;
        RECT 180.615 2626.965 181.215 2627.365 ;
        RECT 185.465 2626.965 186.065 2627.365 ;
      LAYER met4 ;
        RECT 181.615 2489.035 185.065 2626.965 ;
      LAYER met4 ;
        RECT 180.615 2488.635 181.215 2489.035 ;
        RECT 185.465 2488.635 186.065 2489.035 ;
      LAYER met4 ;
        RECT 186.465 2488.730 191.115 2627.270 ;
      LAYER met4 ;
        RECT 191.515 2626.965 192.115 2627.670 ;
        RECT 180.615 2488.330 186.065 2488.635 ;
        RECT 191.515 2488.330 192.115 2489.035 ;
      LAYER met4 ;
        RECT 192.515 2488.730 197.965 2627.270 ;
      LAYER met4 ;
        RECT 198.365 2626.965 199.465 2627.670 ;
      LAYER met4 ;
        RECT 3390.035 2592.730 3395.485 2740.270 ;
      LAYER met4 ;
        RECT 3395.885 2740.030 3396.485 2740.670 ;
        RECT 3401.935 2740.430 3407.385 2740.670 ;
        RECT 3395.885 2592.330 3396.485 2593.035 ;
      LAYER met4 ;
        RECT 3396.885 2592.730 3401.535 2740.270 ;
      LAYER met4 ;
        RECT 3401.935 2740.030 3402.535 2740.430 ;
        RECT 3406.785 2740.030 3407.385 2740.430 ;
      LAYER met4 ;
        RECT 3402.935 2593.035 3406.385 2740.030 ;
      LAYER met4 ;
        RECT 3401.935 2592.635 3402.535 2593.035 ;
        RECT 3406.785 2592.635 3407.385 2593.035 ;
      LAYER met4 ;
        RECT 3407.785 2592.730 3412.435 2740.270 ;
      LAYER met4 ;
        RECT 3412.835 2740.030 3413.435 2740.670 ;
        RECT 3401.935 2592.330 3407.385 2592.635 ;
        RECT 3412.835 2592.330 3413.435 2593.035 ;
      LAYER met4 ;
        RECT 3413.835 2592.730 3418.485 2740.270 ;
      LAYER met4 ;
        RECT 3418.885 2740.030 3419.485 2740.670 ;
        RECT 3418.885 2592.330 3419.485 2593.035 ;
      LAYER met4 ;
        RECT 3419.885 2592.730 3423.335 2740.270 ;
      LAYER met4 ;
        RECT 3423.735 2740.030 3424.335 2740.670 ;
        RECT 3423.735 2592.330 3424.335 2593.035 ;
      LAYER met4 ;
        RECT 3424.735 2592.730 3428.185 2740.270 ;
      LAYER met4 ;
        RECT 3428.585 2740.030 3429.185 2740.670 ;
        RECT 3428.585 2592.330 3429.185 2593.035 ;
      LAYER met4 ;
        RECT 3429.585 2592.730 3434.235 2740.270 ;
      LAYER met4 ;
        RECT 3434.635 2740.030 3435.335 2740.670 ;
        RECT 3434.635 2592.330 3435.335 2593.035 ;
        RECT 3390.035 2520.670 3435.335 2592.330 ;
        RECT 152.665 2416.670 197.965 2488.330 ;
        RECT 152.665 2415.965 153.365 2416.670 ;
        RECT 152.665 2277.330 153.365 2279.000 ;
      LAYER met4 ;
        RECT 153.765 2277.730 158.415 2416.270 ;
      LAYER met4 ;
        RECT 158.815 2415.965 159.415 2416.670 ;
        RECT 158.815 2277.330 159.415 2279.000 ;
      LAYER met4 ;
        RECT 159.815 2277.730 163.265 2416.270 ;
      LAYER met4 ;
        RECT 163.665 2415.965 164.265 2416.670 ;
        RECT 168.515 2415.965 169.115 2416.670 ;
        RECT 163.665 2277.330 164.265 2279.000 ;
        RECT 168.515 2277.330 169.115 2279.000 ;
      LAYER met4 ;
        RECT 169.515 2277.730 174.165 2416.270 ;
      LAYER met4 ;
        RECT 174.565 2415.965 175.165 2416.670 ;
        RECT 180.615 2416.365 186.065 2416.670 ;
        RECT 174.165 2278.935 174.200 2289.935 ;
        RECT 174.565 2277.330 175.165 2279.000 ;
      LAYER met4 ;
        RECT 175.565 2277.730 180.215 2416.270 ;
      LAYER met4 ;
        RECT 180.615 2415.965 181.215 2416.365 ;
        RECT 185.465 2415.965 186.065 2416.365 ;
        RECT 191.515 2415.965 192.115 2416.670 ;
      LAYER met4 ;
        RECT 3390.035 2372.730 3395.485 2520.270 ;
      LAYER met4 ;
        RECT 3395.885 2519.965 3396.485 2520.670 ;
        RECT 3401.935 2520.365 3407.385 2520.670 ;
        RECT 3395.885 2372.330 3396.485 2374.000 ;
      LAYER met4 ;
        RECT 3396.885 2372.730 3401.535 2520.270 ;
      LAYER met4 ;
        RECT 3401.935 2519.965 3402.535 2520.365 ;
        RECT 3406.785 2519.965 3407.385 2520.365 ;
        RECT 3401.935 2372.635 3402.535 2374.000 ;
      LAYER met4 ;
        RECT 3402.935 2373.035 3406.385 2519.965 ;
      LAYER met4 ;
        RECT 3406.785 2372.635 3407.385 2374.000 ;
      LAYER met4 ;
        RECT 3407.785 2372.730 3412.435 2520.270 ;
      LAYER met4 ;
        RECT 3412.835 2519.965 3413.435 2520.670 ;
        RECT 3401.935 2372.330 3407.385 2372.635 ;
        RECT 3412.835 2372.330 3413.435 2374.000 ;
      LAYER met4 ;
        RECT 3413.835 2372.730 3418.485 2520.270 ;
      LAYER met4 ;
        RECT 3418.885 2519.965 3419.485 2520.670 ;
        RECT 3418.885 2372.330 3419.485 2374.000 ;
      LAYER met4 ;
        RECT 3419.885 2372.730 3423.335 2520.270 ;
      LAYER met4 ;
        RECT 3423.735 2519.965 3424.335 2520.670 ;
        RECT 3423.735 2372.330 3424.335 2374.000 ;
      LAYER met4 ;
        RECT 3424.735 2372.730 3428.185 2520.270 ;
      LAYER met4 ;
        RECT 3428.585 2519.965 3429.185 2520.670 ;
        RECT 3428.585 2372.330 3429.185 2374.000 ;
        RECT 3429.550 2373.930 3429.585 2384.975 ;
      LAYER met4 ;
        RECT 3429.585 2372.730 3434.235 2520.270 ;
      LAYER met4 ;
        RECT 3434.635 2519.965 3435.335 2520.670 ;
        RECT 3434.635 2372.330 3435.335 2374.000 ;
        RECT 3390.035 2300.670 3435.335 2372.330 ;
        RECT 180.615 2277.635 181.215 2279.000 ;
        RECT 185.465 2277.635 186.065 2279.000 ;
        RECT 180.615 2277.330 186.065 2277.635 ;
        RECT 191.515 2277.330 192.115 2279.000 ;
        RECT 152.665 2205.670 197.965 2277.330 ;
        RECT 152.665 2204.000 153.365 2205.670 ;
        RECT 152.665 2066.330 153.365 2066.970 ;
      LAYER met4 ;
        RECT 153.765 2066.730 158.415 2205.270 ;
      LAYER met4 ;
        RECT 158.415 2193.025 158.450 2204.070 ;
        RECT 158.815 2204.000 159.415 2205.670 ;
        RECT 158.815 2066.330 159.415 2066.970 ;
      LAYER met4 ;
        RECT 159.815 2066.730 163.265 2205.270 ;
      LAYER met4 ;
        RECT 163.665 2204.000 164.265 2205.670 ;
        RECT 163.665 2066.330 164.265 2066.970 ;
      LAYER met4 ;
        RECT 164.665 2066.730 168.115 2205.270 ;
      LAYER met4 ;
        RECT 168.515 2204.000 169.115 2205.670 ;
        RECT 168.515 2066.330 169.115 2066.970 ;
      LAYER met4 ;
        RECT 169.515 2066.730 174.165 2205.270 ;
      LAYER met4 ;
        RECT 174.565 2204.000 175.165 2205.670 ;
        RECT 180.615 2205.365 186.065 2205.670 ;
        RECT 174.565 2066.330 175.165 2066.970 ;
      LAYER met4 ;
        RECT 175.565 2066.730 180.215 2205.270 ;
      LAYER met4 ;
        RECT 180.615 2204.000 181.215 2205.365 ;
      LAYER met4 ;
        RECT 181.615 2066.970 185.065 2204.965 ;
      LAYER met4 ;
        RECT 185.465 2204.000 186.065 2205.365 ;
        RECT 180.615 2066.570 181.215 2066.970 ;
        RECT 185.465 2066.570 186.065 2066.970 ;
      LAYER met4 ;
        RECT 186.465 2066.730 191.115 2205.270 ;
      LAYER met4 ;
        RECT 191.515 2204.000 192.115 2205.670 ;
        RECT 180.615 2066.330 186.065 2066.570 ;
        RECT 191.515 2066.330 192.115 2066.970 ;
      LAYER met4 ;
        RECT 192.515 2066.730 197.965 2205.270 ;
        RECT 3390.035 2151.730 3395.485 2300.270 ;
      LAYER met4 ;
        RECT 3395.885 2299.000 3396.485 2300.670 ;
        RECT 3401.935 2300.365 3407.385 2300.670 ;
        RECT 3401.935 2299.000 3402.535 2300.365 ;
        RECT 3406.785 2299.000 3407.385 2300.365 ;
        RECT 3395.885 2151.330 3396.485 2152.035 ;
        RECT 3401.935 2151.635 3402.535 2152.035 ;
        RECT 3406.785 2151.635 3407.385 2152.035 ;
      LAYER met4 ;
        RECT 3407.785 2151.730 3412.435 2300.270 ;
      LAYER met4 ;
        RECT 3412.835 2299.000 3413.435 2300.670 ;
        RECT 3413.800 2288.065 3413.835 2299.065 ;
        RECT 3401.935 2151.330 3407.385 2151.635 ;
        RECT 3412.835 2151.330 3413.435 2152.035 ;
      LAYER met4 ;
        RECT 3413.835 2151.730 3418.485 2300.270 ;
      LAYER met4 ;
        RECT 3418.885 2299.000 3419.485 2300.670 ;
        RECT 3418.885 2151.330 3419.485 2152.035 ;
      LAYER met4 ;
        RECT 3419.885 2151.730 3423.335 2300.270 ;
      LAYER met4 ;
        RECT 3423.735 2299.000 3424.335 2300.670 ;
        RECT 3423.735 2151.330 3424.335 2152.035 ;
      LAYER met4 ;
        RECT 3424.735 2151.730 3428.185 2300.270 ;
      LAYER met4 ;
        RECT 3428.585 2299.000 3429.185 2300.670 ;
        RECT 3428.585 2151.330 3429.185 2152.035 ;
      LAYER met4 ;
        RECT 3429.585 2151.730 3434.235 2300.270 ;
      LAYER met4 ;
        RECT 3434.635 2299.000 3435.335 2300.670 ;
        RECT 3434.635 2151.330 3435.335 2152.035 ;
      LAYER met4 ;
        RECT 3435.735 2151.730 3436.065 2771.910 ;
        RECT 3436.365 2766.855 3439.345 2990.535 ;
      LAYER met4 ;
        RECT 3439.745 2966.670 3440.725 2990.935 ;
      LAYER met4 ;
        RECT 3439.645 2965.000 3440.825 2966.270 ;
      LAYER met4 ;
        RECT 3439.645 2819.000 3440.825 2965.000 ;
      LAYER met4 ;
        RECT 3439.645 2817.730 3440.825 2819.000 ;
      LAYER met4 ;
        RECT 3439.745 2782.160 3440.725 2817.330 ;
      LAYER met4 ;
        RECT 3441.125 2782.560 3444.105 3006.240 ;
      LAYER met4 ;
        RECT 3444.505 2998.310 3588.000 3006.640 ;
      LAYER met4 ;
        RECT 3444.405 2816.390 3444.735 2997.910 ;
      LAYER met4 ;
        RECT 3445.135 2966.670 3588.000 2998.310 ;
        RECT 3445.135 2966.030 3445.835 2966.670 ;
        RECT 3445.135 2819.000 3445.835 2965.000 ;
        RECT 3445.135 2817.330 3445.835 2818.035 ;
      LAYER met4 ;
        RECT 3446.235 2817.730 3450.685 2966.270 ;
      LAYER met4 ;
        RECT 3451.085 2966.030 3451.685 2966.670 ;
        RECT 3451.085 2819.000 3451.685 2965.000 ;
        RECT 3451.085 2817.330 3451.685 2818.035 ;
      LAYER met4 ;
        RECT 3452.085 2817.730 3456.535 2966.270 ;
      LAYER met4 ;
        RECT 3456.935 2966.030 3457.635 2966.670 ;
        RECT 3456.935 2819.000 3457.635 2965.000 ;
        RECT 3456.935 2817.330 3457.635 2818.035 ;
      LAYER met4 ;
        RECT 3458.035 2817.730 3483.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2966.030 3563.385 2966.670 ;
      LAYER met4 ;
        RECT 3563.785 2965.000 3588.000 2966.270 ;
      LAYER met4 ;
        RECT 3483.400 2819.000 3588.000 2965.000 ;
        RECT 3483.400 2817.330 3563.385 2818.035 ;
      LAYER met4 ;
        RECT 3563.785 2817.730 3588.000 2819.000 ;
      LAYER met4 ;
        RECT 3445.135 2815.990 3588.000 2817.330 ;
        RECT 3444.505 2782.160 3588.000 2815.990 ;
        RECT 3439.745 2780.640 3588.000 2782.160 ;
        RECT 3439.745 2766.455 3440.725 2780.640 ;
        RECT 3436.465 2764.935 3440.725 2766.455 ;
        RECT 3390.035 2079.670 3435.965 2151.330 ;
        RECT 198.365 2066.330 199.465 2066.970 ;
        RECT 152.665 2034.690 199.465 2066.330 ;
        RECT 152.035 1991.010 199.465 2034.690 ;
        RECT 147.275 1824.545 151.535 1826.065 ;
        RECT 147.275 1810.360 148.255 1824.545 ;
        RECT 0.000 1808.840 148.255 1810.360 ;
        RECT 0.000 1775.010 143.495 1808.840 ;
        RECT 0.000 1773.670 142.865 1775.010 ;
      LAYER met4 ;
        RECT 0.000 1772.000 24.215 1773.270 ;
      LAYER met4 ;
        RECT 24.615 1772.965 104.600 1773.670 ;
        RECT 0.000 1636.000 104.600 1772.000 ;
      LAYER met4 ;
        RECT 0.000 1634.730 24.215 1636.000 ;
      LAYER met4 ;
        RECT 24.615 1634.330 104.600 1634.970 ;
      LAYER met4 ;
        RECT 105.000 1634.730 129.965 1773.270 ;
      LAYER met4 ;
        RECT 130.365 1772.965 131.065 1773.670 ;
        RECT 130.365 1636.000 131.065 1772.000 ;
        RECT 130.365 1634.330 131.065 1634.970 ;
      LAYER met4 ;
        RECT 131.465 1634.730 135.915 1773.270 ;
      LAYER met4 ;
        RECT 136.315 1772.965 136.915 1773.670 ;
        RECT 136.315 1636.000 136.915 1772.000 ;
        RECT 136.315 1634.330 136.915 1634.970 ;
      LAYER met4 ;
        RECT 137.315 1634.730 141.765 1773.270 ;
      LAYER met4 ;
        RECT 142.165 1772.965 142.865 1773.670 ;
        RECT 142.165 1636.000 142.865 1772.000 ;
        RECT 142.165 1634.330 142.865 1634.970 ;
        RECT 0.000 1602.690 142.865 1634.330 ;
      LAYER met4 ;
        RECT 143.265 1603.090 143.595 1774.610 ;
      LAYER met4 ;
        RECT 0.000 1594.360 143.495 1602.690 ;
      LAYER met4 ;
        RECT 143.895 1594.760 146.875 1808.440 ;
      LAYER met4 ;
        RECT 147.275 1773.670 148.255 1808.840 ;
      LAYER met4 ;
        RECT 147.175 1772.000 148.355 1773.270 ;
      LAYER met4 ;
        RECT 147.175 1636.000 148.355 1772.000 ;
      LAYER met4 ;
        RECT 147.175 1634.730 148.355 1636.000 ;
      LAYER met4 ;
        RECT 147.275 1610.065 148.255 1634.330 ;
      LAYER met4 ;
        RECT 148.655 1610.465 151.635 1824.145 ;
        RECT 151.935 1819.090 152.265 1990.610 ;
      LAYER met4 ;
        RECT 152.665 1989.670 199.465 1991.010 ;
        RECT 152.665 1988.965 153.365 1989.670 ;
        RECT 152.665 1850.330 153.365 1850.970 ;
      LAYER met4 ;
        RECT 153.765 1850.730 158.415 1989.270 ;
      LAYER met4 ;
        RECT 158.815 1988.965 159.415 1989.670 ;
        RECT 158.815 1850.330 159.415 1850.970 ;
      LAYER met4 ;
        RECT 159.815 1850.730 163.265 1989.270 ;
      LAYER met4 ;
        RECT 163.665 1988.965 164.265 1989.670 ;
        RECT 163.665 1850.330 164.265 1850.970 ;
      LAYER met4 ;
        RECT 164.665 1850.730 168.115 1989.270 ;
      LAYER met4 ;
        RECT 168.515 1988.965 169.115 1989.670 ;
        RECT 168.515 1850.330 169.115 1850.970 ;
      LAYER met4 ;
        RECT 169.515 1850.730 174.165 1989.270 ;
      LAYER met4 ;
        RECT 174.565 1988.965 175.165 1989.670 ;
        RECT 180.615 1989.365 186.065 1989.670 ;
        RECT 174.565 1850.330 175.165 1850.970 ;
      LAYER met4 ;
        RECT 175.565 1850.730 180.215 1989.270 ;
      LAYER met4 ;
        RECT 180.615 1988.965 181.215 1989.365 ;
        RECT 185.465 1988.965 186.065 1989.365 ;
      LAYER met4 ;
        RECT 181.615 1850.970 185.065 1988.965 ;
      LAYER met4 ;
        RECT 180.615 1850.570 181.215 1850.970 ;
        RECT 185.465 1850.570 186.065 1850.970 ;
      LAYER met4 ;
        RECT 186.465 1850.730 191.115 1989.270 ;
      LAYER met4 ;
        RECT 191.515 1988.965 192.115 1989.670 ;
        RECT 180.615 1850.330 186.065 1850.570 ;
        RECT 191.515 1850.330 192.115 1850.970 ;
      LAYER met4 ;
        RECT 192.515 1850.730 197.965 1989.270 ;
      LAYER met4 ;
        RECT 198.365 1988.965 199.465 1989.670 ;
        RECT 3388.535 1931.330 3389.635 1932.035 ;
      LAYER met4 ;
        RECT 3390.035 1931.730 3395.485 2079.270 ;
      LAYER met4 ;
        RECT 3395.885 2078.965 3396.485 2079.670 ;
        RECT 3401.935 2079.365 3407.385 2079.670 ;
        RECT 3395.885 1931.330 3396.485 1932.035 ;
      LAYER met4 ;
        RECT 3396.885 1931.730 3401.535 2079.270 ;
      LAYER met4 ;
        RECT 3401.935 2078.965 3402.535 2079.365 ;
        RECT 3406.785 2078.965 3407.385 2079.365 ;
      LAYER met4 ;
        RECT 3402.935 1932.035 3406.385 2078.965 ;
      LAYER met4 ;
        RECT 3401.935 1931.635 3402.535 1932.035 ;
        RECT 3406.785 1931.635 3407.385 1932.035 ;
      LAYER met4 ;
        RECT 3407.785 1931.730 3412.435 2079.270 ;
      LAYER met4 ;
        RECT 3412.835 2078.965 3413.435 2079.670 ;
        RECT 3401.935 1931.330 3407.385 1931.635 ;
        RECT 3412.835 1931.330 3413.435 1932.035 ;
      LAYER met4 ;
        RECT 3413.835 1931.730 3418.485 2079.270 ;
      LAYER met4 ;
        RECT 3418.885 2078.965 3419.485 2079.670 ;
        RECT 3418.885 1931.330 3419.485 1932.035 ;
      LAYER met4 ;
        RECT 3419.885 1931.730 3423.335 2079.270 ;
      LAYER met4 ;
        RECT 3423.735 2078.965 3424.335 2079.670 ;
        RECT 3423.735 1931.330 3424.335 1932.035 ;
      LAYER met4 ;
        RECT 3424.735 1931.730 3428.185 2079.270 ;
      LAYER met4 ;
        RECT 3428.585 2078.965 3429.185 2079.670 ;
        RECT 3428.585 1931.330 3429.185 1932.035 ;
      LAYER met4 ;
        RECT 3429.585 1931.730 3434.235 2079.270 ;
      LAYER met4 ;
        RECT 3434.635 2078.965 3435.335 2079.670 ;
        RECT 3434.635 1931.330 3435.335 1932.035 ;
        RECT 3388.535 1929.990 3435.335 1931.330 ;
      LAYER met4 ;
        RECT 3435.735 1930.390 3436.065 2079.270 ;
      LAYER met4 ;
        RECT 3388.535 1886.310 3435.965 1929.990 ;
        RECT 3388.535 1854.670 3435.335 1886.310 ;
        RECT 3388.535 1854.030 3389.635 1854.670 ;
        RECT 198.365 1850.330 199.465 1850.970 ;
        RECT 152.665 1818.690 199.465 1850.330 ;
        RECT 152.035 1775.010 199.465 1818.690 ;
        RECT 147.275 1608.545 151.535 1610.065 ;
        RECT 147.275 1594.360 148.255 1608.545 ;
        RECT 0.000 1592.840 148.255 1594.360 ;
        RECT 0.000 1559.010 143.495 1592.840 ;
        RECT 0.000 1557.670 142.865 1559.010 ;
      LAYER met4 ;
        RECT 0.000 1556.000 24.215 1557.270 ;
      LAYER met4 ;
        RECT 24.615 1556.965 104.600 1557.670 ;
        RECT 0.000 1420.000 104.600 1556.000 ;
      LAYER met4 ;
        RECT 0.000 1418.730 24.215 1420.000 ;
      LAYER met4 ;
        RECT 24.615 1418.330 104.600 1418.970 ;
      LAYER met4 ;
        RECT 105.000 1418.730 129.965 1557.270 ;
      LAYER met4 ;
        RECT 130.365 1556.965 131.065 1557.670 ;
        RECT 130.365 1420.000 131.065 1556.000 ;
        RECT 130.365 1418.330 131.065 1418.970 ;
      LAYER met4 ;
        RECT 131.465 1418.730 135.915 1557.270 ;
      LAYER met4 ;
        RECT 136.315 1556.965 136.915 1557.670 ;
        RECT 136.315 1420.000 136.915 1556.000 ;
        RECT 136.315 1418.330 136.915 1418.970 ;
      LAYER met4 ;
        RECT 137.315 1418.730 141.765 1557.270 ;
      LAYER met4 ;
        RECT 142.165 1556.965 142.865 1557.670 ;
        RECT 142.165 1420.000 142.865 1556.000 ;
        RECT 142.165 1418.330 142.865 1418.970 ;
        RECT 0.000 1386.690 142.865 1418.330 ;
      LAYER met4 ;
        RECT 143.265 1387.090 143.595 1558.610 ;
      LAYER met4 ;
        RECT 0.000 1378.360 143.495 1386.690 ;
      LAYER met4 ;
        RECT 143.895 1378.760 146.875 1592.440 ;
      LAYER met4 ;
        RECT 147.275 1557.670 148.255 1592.840 ;
      LAYER met4 ;
        RECT 147.175 1556.000 148.355 1557.270 ;
      LAYER met4 ;
        RECT 147.175 1420.000 148.355 1556.000 ;
      LAYER met4 ;
        RECT 147.175 1418.730 148.355 1420.000 ;
      LAYER met4 ;
        RECT 147.275 1394.065 148.255 1418.330 ;
      LAYER met4 ;
        RECT 148.655 1394.465 151.635 1608.145 ;
        RECT 151.935 1603.090 152.265 1774.610 ;
      LAYER met4 ;
        RECT 152.665 1773.670 199.465 1775.010 ;
        RECT 152.665 1772.965 153.365 1773.670 ;
        RECT 152.665 1634.330 153.365 1634.970 ;
      LAYER met4 ;
        RECT 153.765 1634.730 158.415 1773.270 ;
      LAYER met4 ;
        RECT 158.815 1772.965 159.415 1773.670 ;
        RECT 158.815 1634.330 159.415 1634.970 ;
      LAYER met4 ;
        RECT 159.815 1634.730 163.265 1773.270 ;
      LAYER met4 ;
        RECT 163.665 1772.965 164.265 1773.670 ;
        RECT 163.665 1634.330 164.265 1634.970 ;
      LAYER met4 ;
        RECT 164.665 1634.730 168.115 1773.270 ;
      LAYER met4 ;
        RECT 168.515 1772.965 169.115 1773.670 ;
        RECT 168.515 1634.330 169.115 1634.970 ;
      LAYER met4 ;
        RECT 169.515 1634.730 174.165 1773.270 ;
      LAYER met4 ;
        RECT 174.565 1772.965 175.165 1773.670 ;
        RECT 180.615 1773.365 186.065 1773.670 ;
        RECT 174.565 1634.330 175.165 1634.970 ;
      LAYER met4 ;
        RECT 175.565 1634.730 180.215 1773.270 ;
      LAYER met4 ;
        RECT 180.615 1772.965 181.215 1773.365 ;
        RECT 185.465 1772.965 186.065 1773.365 ;
      LAYER met4 ;
        RECT 181.615 1634.970 185.065 1772.965 ;
      LAYER met4 ;
        RECT 180.615 1634.570 181.215 1634.970 ;
        RECT 185.465 1634.570 186.065 1634.970 ;
      LAYER met4 ;
        RECT 186.465 1634.730 191.115 1773.270 ;
      LAYER met4 ;
        RECT 191.515 1772.965 192.115 1773.670 ;
        RECT 180.615 1634.330 186.065 1634.570 ;
        RECT 191.515 1634.330 192.115 1634.970 ;
      LAYER met4 ;
        RECT 192.515 1634.730 197.965 1773.270 ;
      LAYER met4 ;
        RECT 198.365 1772.965 199.465 1773.670 ;
        RECT 3388.535 1705.330 3389.635 1706.035 ;
      LAYER met4 ;
        RECT 3390.035 1705.730 3395.485 1854.270 ;
      LAYER met4 ;
        RECT 3395.885 1854.030 3396.485 1854.670 ;
        RECT 3401.935 1854.430 3407.385 1854.670 ;
        RECT 3395.885 1705.330 3396.485 1706.035 ;
      LAYER met4 ;
        RECT 3396.885 1705.730 3401.535 1854.270 ;
      LAYER met4 ;
        RECT 3401.935 1854.030 3402.535 1854.430 ;
        RECT 3406.785 1854.030 3407.385 1854.430 ;
      LAYER met4 ;
        RECT 3402.935 1706.035 3406.385 1854.030 ;
      LAYER met4 ;
        RECT 3401.935 1705.635 3402.535 1706.035 ;
        RECT 3406.785 1705.635 3407.385 1706.035 ;
      LAYER met4 ;
        RECT 3407.785 1705.730 3412.435 1854.270 ;
      LAYER met4 ;
        RECT 3412.835 1854.030 3413.435 1854.670 ;
        RECT 3401.935 1705.330 3407.385 1705.635 ;
        RECT 3412.835 1705.330 3413.435 1706.035 ;
      LAYER met4 ;
        RECT 3413.835 1705.730 3418.485 1854.270 ;
      LAYER met4 ;
        RECT 3418.885 1854.030 3419.485 1854.670 ;
        RECT 3418.885 1705.330 3419.485 1706.035 ;
      LAYER met4 ;
        RECT 3419.885 1705.730 3423.335 1854.270 ;
      LAYER met4 ;
        RECT 3423.735 1854.030 3424.335 1854.670 ;
        RECT 3423.735 1705.330 3424.335 1706.035 ;
      LAYER met4 ;
        RECT 3424.735 1705.730 3428.185 1854.270 ;
      LAYER met4 ;
        RECT 3428.585 1854.030 3429.185 1854.670 ;
        RECT 3428.585 1705.330 3429.185 1706.035 ;
      LAYER met4 ;
        RECT 3429.585 1705.730 3434.235 1854.270 ;
      LAYER met4 ;
        RECT 3434.635 1854.030 3435.335 1854.670 ;
        RECT 3434.635 1705.330 3435.335 1706.035 ;
        RECT 3388.535 1703.990 3435.335 1705.330 ;
      LAYER met4 ;
        RECT 3435.735 1704.390 3436.065 1885.910 ;
        RECT 3436.365 1880.855 3439.345 2764.535 ;
      LAYER met4 ;
        RECT 3439.745 2740.670 3440.725 2764.935 ;
      LAYER met4 ;
        RECT 3439.645 2739.000 3440.825 2740.270 ;
      LAYER met4 ;
        RECT 3439.645 2594.000 3440.825 2739.000 ;
      LAYER met4 ;
        RECT 3439.645 2592.730 3440.825 2594.000 ;
      LAYER met4 ;
        RECT 3439.745 2520.670 3440.725 2592.330 ;
      LAYER met4 ;
        RECT 3439.645 2519.000 3440.825 2520.270 ;
      LAYER met4 ;
        RECT 3439.645 2374.000 3440.825 2519.000 ;
      LAYER met4 ;
        RECT 3439.645 2372.730 3440.825 2374.000 ;
      LAYER met4 ;
        RECT 3439.745 2300.670 3440.725 2372.330 ;
      LAYER met4 ;
        RECT 3439.645 2299.000 3440.825 2300.270 ;
      LAYER met4 ;
        RECT 3439.645 2153.000 3440.825 2299.000 ;
      LAYER met4 ;
        RECT 3439.645 2151.730 3440.825 2153.000 ;
      LAYER met4 ;
        RECT 3439.745 2079.670 3440.725 2151.330 ;
      LAYER met4 ;
        RECT 3439.645 2078.000 3440.825 2079.270 ;
      LAYER met4 ;
        RECT 3439.645 1933.000 3440.825 2078.000 ;
      LAYER met4 ;
        RECT 3439.645 1931.730 3440.825 1933.000 ;
      LAYER met4 ;
        RECT 3439.745 1896.160 3440.725 1931.330 ;
      LAYER met4 ;
        RECT 3441.125 1896.560 3444.105 2780.240 ;
      LAYER met4 ;
        RECT 3444.505 2772.310 3588.000 2780.640 ;
        RECT 3445.135 2740.670 3588.000 2772.310 ;
        RECT 3445.135 2740.030 3445.835 2740.670 ;
        RECT 3445.135 2594.000 3445.835 2739.000 ;
        RECT 3445.135 2592.330 3445.835 2593.035 ;
      LAYER met4 ;
        RECT 3446.235 2592.730 3450.685 2740.270 ;
      LAYER met4 ;
        RECT 3451.085 2740.030 3451.685 2740.670 ;
        RECT 3451.085 2594.000 3451.685 2739.000 ;
        RECT 3451.085 2592.330 3451.685 2593.035 ;
      LAYER met4 ;
        RECT 3452.085 2592.730 3456.535 2740.270 ;
      LAYER met4 ;
        RECT 3456.935 2740.030 3457.635 2740.670 ;
        RECT 3456.935 2594.000 3457.635 2739.000 ;
        RECT 3456.935 2592.330 3457.635 2593.035 ;
      LAYER met4 ;
        RECT 3458.035 2592.730 3483.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2740.030 3563.385 2740.670 ;
      LAYER met4 ;
        RECT 3563.785 2739.000 3588.000 2740.270 ;
      LAYER met4 ;
        RECT 3483.400 2594.000 3588.000 2739.000 ;
        RECT 3483.400 2592.330 3563.385 2593.035 ;
      LAYER met4 ;
        RECT 3563.785 2592.730 3588.000 2594.000 ;
      LAYER met4 ;
        RECT 3445.135 2520.670 3588.000 2592.330 ;
        RECT 3445.135 2519.965 3445.835 2520.670 ;
        RECT 3445.135 2372.330 3445.835 2519.000 ;
      LAYER met4 ;
        RECT 3446.235 2372.730 3450.685 2520.270 ;
      LAYER met4 ;
        RECT 3451.085 2519.965 3451.685 2520.670 ;
        RECT 3451.085 2372.330 3451.685 2519.000 ;
      LAYER met4 ;
        RECT 3452.085 2372.730 3456.535 2520.270 ;
      LAYER met4 ;
        RECT 3456.935 2519.965 3457.635 2520.670 ;
        RECT 3456.935 2372.330 3457.635 2519.000 ;
      LAYER met4 ;
        RECT 3458.035 2372.730 3483.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2519.965 3563.385 2520.670 ;
      LAYER met4 ;
        RECT 3563.785 2519.000 3588.000 2520.270 ;
      LAYER met4 ;
        RECT 3483.400 2374.000 3588.000 2519.000 ;
        RECT 3483.400 2372.330 3563.385 2374.000 ;
      LAYER met4 ;
        RECT 3563.785 2372.730 3588.000 2374.000 ;
      LAYER met4 ;
        RECT 3445.135 2300.670 3588.000 2372.330 ;
        RECT 3445.135 2153.000 3445.835 2300.670 ;
        RECT 3445.135 2151.330 3445.835 2152.035 ;
      LAYER met4 ;
        RECT 3446.235 2151.730 3450.685 2300.270 ;
      LAYER met4 ;
        RECT 3451.085 2153.000 3451.685 2300.670 ;
        RECT 3451.085 2151.330 3451.685 2152.035 ;
      LAYER met4 ;
        RECT 3452.085 2151.730 3456.535 2300.270 ;
      LAYER met4 ;
        RECT 3456.935 2153.000 3457.635 2300.670 ;
        RECT 3456.935 2151.330 3457.635 2152.035 ;
      LAYER met4 ;
        RECT 3458.035 2151.730 3483.000 2300.270 ;
      LAYER met4 ;
        RECT 3483.400 2299.000 3563.385 2300.670 ;
        RECT 3563.750 2299.000 3563.785 2299.215 ;
      LAYER met4 ;
        RECT 3563.785 2299.000 3588.000 2300.270 ;
      LAYER met4 ;
        RECT 3483.400 2153.000 3588.000 2299.000 ;
        RECT 3483.400 2151.330 3563.385 2152.035 ;
      LAYER met4 ;
        RECT 3563.785 2151.730 3588.000 2153.000 ;
      LAYER met4 ;
        RECT 3444.505 2079.670 3588.000 2151.330 ;
      LAYER met4 ;
        RECT 3444.405 1930.390 3444.735 2079.270 ;
      LAYER met4 ;
        RECT 3445.135 2078.965 3445.835 2079.670 ;
        RECT 3445.135 1933.000 3445.835 2078.000 ;
        RECT 3445.135 1931.330 3445.835 1932.035 ;
      LAYER met4 ;
        RECT 3446.235 1931.730 3450.685 2079.270 ;
      LAYER met4 ;
        RECT 3451.085 2078.965 3451.685 2079.670 ;
        RECT 3451.085 1933.000 3451.685 2078.000 ;
        RECT 3451.085 1931.330 3451.685 1932.035 ;
      LAYER met4 ;
        RECT 3452.085 1931.730 3456.535 2079.270 ;
      LAYER met4 ;
        RECT 3456.935 2078.965 3457.635 2079.670 ;
        RECT 3456.935 1933.000 3457.635 2078.000 ;
        RECT 3456.935 1931.330 3457.635 1932.035 ;
      LAYER met4 ;
        RECT 3458.035 1931.730 3483.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 2078.965 3563.385 2079.670 ;
      LAYER met4 ;
        RECT 3563.785 2078.000 3588.000 2079.270 ;
      LAYER met4 ;
        RECT 3483.400 1933.000 3588.000 2078.000 ;
        RECT 3483.400 1931.330 3563.385 1932.035 ;
      LAYER met4 ;
        RECT 3563.785 1931.730 3588.000 1933.000 ;
      LAYER met4 ;
        RECT 3445.135 1929.990 3588.000 1931.330 ;
        RECT 3444.505 1896.160 3588.000 1929.990 ;
        RECT 3439.745 1894.640 3588.000 1896.160 ;
        RECT 3439.745 1880.455 3440.725 1894.640 ;
        RECT 3436.465 1878.935 3440.725 1880.455 ;
        RECT 3388.535 1660.310 3435.965 1703.990 ;
        RECT 198.365 1634.330 199.465 1634.970 ;
        RECT 152.665 1602.690 199.465 1634.330 ;
        RECT 3388.535 1628.670 3435.335 1660.310 ;
        RECT 3388.535 1628.030 3389.635 1628.670 ;
        RECT 152.035 1559.010 199.465 1602.690 ;
        RECT 147.275 1392.545 151.535 1394.065 ;
        RECT 147.275 1378.360 148.255 1392.545 ;
        RECT 0.000 1376.840 148.255 1378.360 ;
        RECT 0.000 1343.010 143.495 1376.840 ;
        RECT 0.000 1341.670 142.865 1343.010 ;
      LAYER met4 ;
        RECT 0.000 1340.000 24.215 1341.270 ;
      LAYER met4 ;
        RECT 24.615 1340.965 104.600 1341.670 ;
        RECT 0.000 1204.000 104.600 1340.000 ;
      LAYER met4 ;
        RECT 0.000 1202.730 24.215 1204.000 ;
      LAYER met4 ;
        RECT 24.615 1202.330 104.600 1202.970 ;
      LAYER met4 ;
        RECT 105.000 1202.730 129.965 1341.270 ;
      LAYER met4 ;
        RECT 130.365 1340.965 131.065 1341.670 ;
        RECT 130.365 1204.000 131.065 1340.000 ;
        RECT 130.365 1202.330 131.065 1202.970 ;
      LAYER met4 ;
        RECT 131.465 1202.730 135.915 1341.270 ;
      LAYER met4 ;
        RECT 136.315 1340.965 136.915 1341.670 ;
        RECT 136.315 1204.000 136.915 1340.000 ;
        RECT 136.315 1202.330 136.915 1202.970 ;
      LAYER met4 ;
        RECT 137.315 1202.730 141.765 1341.270 ;
      LAYER met4 ;
        RECT 142.165 1340.965 142.865 1341.670 ;
        RECT 142.165 1204.000 142.865 1340.000 ;
        RECT 142.165 1202.330 142.865 1202.970 ;
        RECT 0.000 1170.690 142.865 1202.330 ;
      LAYER met4 ;
        RECT 143.265 1171.090 143.595 1342.610 ;
      LAYER met4 ;
        RECT 0.000 1162.360 143.495 1170.690 ;
      LAYER met4 ;
        RECT 143.895 1162.760 146.875 1376.440 ;
      LAYER met4 ;
        RECT 147.275 1341.670 148.255 1376.840 ;
      LAYER met4 ;
        RECT 147.175 1340.000 148.355 1341.270 ;
      LAYER met4 ;
        RECT 147.175 1204.000 148.355 1340.000 ;
      LAYER met4 ;
        RECT 147.175 1202.730 148.355 1204.000 ;
      LAYER met4 ;
        RECT 147.275 1178.065 148.255 1202.330 ;
      LAYER met4 ;
        RECT 148.655 1178.465 151.635 1392.145 ;
        RECT 151.935 1387.090 152.265 1558.610 ;
      LAYER met4 ;
        RECT 152.665 1557.670 199.465 1559.010 ;
        RECT 152.665 1556.965 153.365 1557.670 ;
        RECT 152.665 1418.330 153.365 1418.970 ;
      LAYER met4 ;
        RECT 153.765 1418.730 158.415 1557.270 ;
      LAYER met4 ;
        RECT 158.815 1556.965 159.415 1557.670 ;
        RECT 158.815 1418.330 159.415 1418.970 ;
      LAYER met4 ;
        RECT 159.815 1418.730 163.265 1557.270 ;
      LAYER met4 ;
        RECT 163.665 1556.965 164.265 1557.670 ;
        RECT 163.665 1418.330 164.265 1418.970 ;
      LAYER met4 ;
        RECT 164.665 1418.730 168.115 1557.270 ;
      LAYER met4 ;
        RECT 168.515 1556.965 169.115 1557.670 ;
        RECT 168.515 1418.330 169.115 1418.970 ;
      LAYER met4 ;
        RECT 169.515 1418.730 174.165 1557.270 ;
      LAYER met4 ;
        RECT 174.565 1556.965 175.165 1557.670 ;
        RECT 180.615 1557.365 186.065 1557.670 ;
        RECT 174.565 1418.330 175.165 1418.970 ;
      LAYER met4 ;
        RECT 175.565 1418.730 180.215 1557.270 ;
      LAYER met4 ;
        RECT 180.615 1556.965 181.215 1557.365 ;
        RECT 185.465 1556.965 186.065 1557.365 ;
      LAYER met4 ;
        RECT 181.615 1418.970 185.065 1556.965 ;
      LAYER met4 ;
        RECT 180.615 1418.570 181.215 1418.970 ;
        RECT 185.465 1418.570 186.065 1418.970 ;
      LAYER met4 ;
        RECT 186.465 1418.730 191.115 1557.270 ;
      LAYER met4 ;
        RECT 191.515 1556.965 192.115 1557.670 ;
        RECT 180.615 1418.330 186.065 1418.570 ;
        RECT 191.515 1418.330 192.115 1418.970 ;
      LAYER met4 ;
        RECT 192.515 1418.730 197.965 1557.270 ;
      LAYER met4 ;
        RECT 198.365 1556.965 199.465 1557.670 ;
        RECT 3388.535 1480.330 3389.635 1481.035 ;
      LAYER met4 ;
        RECT 3390.035 1480.730 3395.485 1628.270 ;
      LAYER met4 ;
        RECT 3395.885 1628.030 3396.485 1628.670 ;
        RECT 3401.935 1628.430 3407.385 1628.670 ;
        RECT 3395.885 1480.330 3396.485 1481.035 ;
      LAYER met4 ;
        RECT 3396.885 1480.730 3401.535 1628.270 ;
      LAYER met4 ;
        RECT 3401.935 1628.030 3402.535 1628.430 ;
        RECT 3406.785 1628.030 3407.385 1628.430 ;
      LAYER met4 ;
        RECT 3402.935 1481.035 3406.385 1628.030 ;
      LAYER met4 ;
        RECT 3401.935 1480.635 3402.535 1481.035 ;
        RECT 3406.785 1480.635 3407.385 1481.035 ;
      LAYER met4 ;
        RECT 3407.785 1480.730 3412.435 1628.270 ;
      LAYER met4 ;
        RECT 3412.835 1628.030 3413.435 1628.670 ;
        RECT 3401.935 1480.330 3407.385 1480.635 ;
        RECT 3412.835 1480.330 3413.435 1481.035 ;
      LAYER met4 ;
        RECT 3413.835 1480.730 3418.485 1628.270 ;
      LAYER met4 ;
        RECT 3418.885 1628.030 3419.485 1628.670 ;
        RECT 3418.885 1480.330 3419.485 1481.035 ;
      LAYER met4 ;
        RECT 3419.885 1480.730 3423.335 1628.270 ;
      LAYER met4 ;
        RECT 3423.735 1628.030 3424.335 1628.670 ;
        RECT 3423.735 1480.330 3424.335 1481.035 ;
      LAYER met4 ;
        RECT 3424.735 1480.730 3428.185 1628.270 ;
      LAYER met4 ;
        RECT 3428.585 1628.030 3429.185 1628.670 ;
        RECT 3428.585 1480.330 3429.185 1481.035 ;
      LAYER met4 ;
        RECT 3429.585 1480.730 3434.235 1628.270 ;
      LAYER met4 ;
        RECT 3434.635 1628.030 3435.335 1628.670 ;
        RECT 3434.635 1480.330 3435.335 1481.035 ;
        RECT 3388.535 1478.990 3435.335 1480.330 ;
      LAYER met4 ;
        RECT 3435.735 1479.390 3436.065 1659.910 ;
        RECT 3436.365 1654.855 3439.345 1878.535 ;
      LAYER met4 ;
        RECT 3439.745 1854.670 3440.725 1878.935 ;
      LAYER met4 ;
        RECT 3439.645 1853.000 3440.825 1854.270 ;
      LAYER met4 ;
        RECT 3439.645 1707.000 3440.825 1853.000 ;
      LAYER met4 ;
        RECT 3439.645 1705.730 3440.825 1707.000 ;
      LAYER met4 ;
        RECT 3439.745 1670.160 3440.725 1705.330 ;
      LAYER met4 ;
        RECT 3441.125 1670.560 3444.105 1894.240 ;
      LAYER met4 ;
        RECT 3444.505 1886.310 3588.000 1894.640 ;
      LAYER met4 ;
        RECT 3444.405 1704.390 3444.735 1885.910 ;
      LAYER met4 ;
        RECT 3445.135 1854.670 3588.000 1886.310 ;
        RECT 3445.135 1854.030 3445.835 1854.670 ;
        RECT 3445.135 1707.000 3445.835 1853.000 ;
        RECT 3445.135 1705.330 3445.835 1706.035 ;
      LAYER met4 ;
        RECT 3446.235 1705.730 3450.685 1854.270 ;
      LAYER met4 ;
        RECT 3451.085 1854.030 3451.685 1854.670 ;
        RECT 3451.085 1707.000 3451.685 1853.000 ;
        RECT 3451.085 1705.330 3451.685 1706.035 ;
      LAYER met4 ;
        RECT 3452.085 1705.730 3456.535 1854.270 ;
      LAYER met4 ;
        RECT 3456.935 1854.030 3457.635 1854.670 ;
        RECT 3456.935 1707.000 3457.635 1853.000 ;
        RECT 3456.935 1705.330 3457.635 1706.035 ;
      LAYER met4 ;
        RECT 3458.035 1705.730 3483.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1854.030 3563.385 1854.670 ;
      LAYER met4 ;
        RECT 3563.785 1853.000 3588.000 1854.270 ;
      LAYER met4 ;
        RECT 3483.400 1707.000 3588.000 1853.000 ;
        RECT 3483.400 1705.330 3563.385 1706.035 ;
      LAYER met4 ;
        RECT 3563.785 1705.730 3588.000 1707.000 ;
      LAYER met4 ;
        RECT 3445.135 1703.990 3588.000 1705.330 ;
        RECT 3444.505 1670.160 3588.000 1703.990 ;
        RECT 3439.745 1668.640 3588.000 1670.160 ;
        RECT 3439.745 1654.455 3440.725 1668.640 ;
        RECT 3436.465 1652.935 3440.725 1654.455 ;
        RECT 3388.535 1435.310 3435.965 1478.990 ;
        RECT 198.365 1418.330 199.465 1418.970 ;
        RECT 152.665 1386.690 199.465 1418.330 ;
        RECT 3388.535 1403.670 3435.335 1435.310 ;
        RECT 3388.535 1403.030 3389.635 1403.670 ;
        RECT 152.035 1343.010 199.465 1386.690 ;
        RECT 147.275 1176.545 151.535 1178.065 ;
        RECT 147.275 1162.360 148.255 1176.545 ;
        RECT 0.000 1160.840 148.255 1162.360 ;
        RECT 0.000 1127.010 143.495 1160.840 ;
        RECT 0.000 1125.670 142.865 1127.010 ;
      LAYER met4 ;
        RECT 0.000 1124.000 24.215 1125.270 ;
      LAYER met4 ;
        RECT 24.615 1124.965 104.600 1125.670 ;
        RECT 0.000 988.000 104.600 1124.000 ;
      LAYER met4 ;
        RECT 0.000 986.730 24.215 988.000 ;
      LAYER met4 ;
        RECT 24.615 986.330 104.600 986.970 ;
      LAYER met4 ;
        RECT 105.000 986.730 129.965 1125.270 ;
      LAYER met4 ;
        RECT 130.365 1124.965 131.065 1125.670 ;
        RECT 130.365 988.000 131.065 1124.000 ;
        RECT 130.365 986.330 131.065 986.970 ;
      LAYER met4 ;
        RECT 131.465 986.730 135.915 1125.270 ;
      LAYER met4 ;
        RECT 136.315 1124.965 136.915 1125.670 ;
        RECT 136.315 988.000 136.915 1124.000 ;
        RECT 136.315 986.330 136.915 986.970 ;
      LAYER met4 ;
        RECT 137.315 986.730 141.765 1125.270 ;
      LAYER met4 ;
        RECT 142.165 1124.965 142.865 1125.670 ;
        RECT 142.165 988.000 142.865 1124.000 ;
        RECT 142.165 986.330 142.865 986.970 ;
        RECT 0.000 954.690 142.865 986.330 ;
      LAYER met4 ;
        RECT 143.265 955.090 143.595 1126.610 ;
      LAYER met4 ;
        RECT 0.000 946.360 143.495 954.690 ;
      LAYER met4 ;
        RECT 143.895 946.760 146.875 1160.440 ;
      LAYER met4 ;
        RECT 147.275 1125.670 148.255 1160.840 ;
      LAYER met4 ;
        RECT 147.175 1124.000 148.355 1125.270 ;
      LAYER met4 ;
        RECT 147.175 988.000 148.355 1124.000 ;
      LAYER met4 ;
        RECT 147.175 986.730 148.355 988.000 ;
      LAYER met4 ;
        RECT 147.275 962.065 148.255 986.330 ;
      LAYER met4 ;
        RECT 148.655 962.465 151.635 1176.145 ;
        RECT 151.935 1171.090 152.265 1342.610 ;
      LAYER met4 ;
        RECT 152.665 1341.670 199.465 1343.010 ;
        RECT 152.665 1340.965 153.365 1341.670 ;
        RECT 152.665 1202.330 153.365 1202.970 ;
      LAYER met4 ;
        RECT 153.765 1202.730 158.415 1341.270 ;
      LAYER met4 ;
        RECT 158.815 1340.965 159.415 1341.670 ;
        RECT 158.815 1202.330 159.415 1202.970 ;
      LAYER met4 ;
        RECT 159.815 1202.730 163.265 1341.270 ;
      LAYER met4 ;
        RECT 163.665 1340.965 164.265 1341.670 ;
        RECT 163.665 1202.330 164.265 1202.970 ;
      LAYER met4 ;
        RECT 164.665 1202.730 168.115 1341.270 ;
      LAYER met4 ;
        RECT 168.515 1340.965 169.115 1341.670 ;
        RECT 168.515 1202.330 169.115 1202.970 ;
      LAYER met4 ;
        RECT 169.515 1202.730 174.165 1341.270 ;
      LAYER met4 ;
        RECT 174.565 1340.965 175.165 1341.670 ;
        RECT 180.615 1341.365 186.065 1341.670 ;
        RECT 174.565 1202.330 175.165 1202.970 ;
      LAYER met4 ;
        RECT 175.565 1202.730 180.215 1341.270 ;
      LAYER met4 ;
        RECT 180.615 1340.965 181.215 1341.365 ;
        RECT 185.465 1340.965 186.065 1341.365 ;
      LAYER met4 ;
        RECT 181.615 1202.970 185.065 1340.965 ;
      LAYER met4 ;
        RECT 180.615 1202.570 181.215 1202.970 ;
        RECT 185.465 1202.570 186.065 1202.970 ;
      LAYER met4 ;
        RECT 186.465 1202.730 191.115 1341.270 ;
      LAYER met4 ;
        RECT 191.515 1340.965 192.115 1341.670 ;
        RECT 180.615 1202.330 186.065 1202.570 ;
        RECT 191.515 1202.330 192.115 1202.970 ;
      LAYER met4 ;
        RECT 192.515 1202.730 197.965 1341.270 ;
      LAYER met4 ;
        RECT 198.365 1340.965 199.465 1341.670 ;
        RECT 3388.535 1255.330 3389.635 1256.035 ;
      LAYER met4 ;
        RECT 3390.035 1255.730 3395.485 1403.270 ;
      LAYER met4 ;
        RECT 3395.885 1403.030 3396.485 1403.670 ;
        RECT 3401.935 1403.430 3407.385 1403.670 ;
        RECT 3395.885 1255.330 3396.485 1256.035 ;
      LAYER met4 ;
        RECT 3396.885 1255.730 3401.535 1403.270 ;
      LAYER met4 ;
        RECT 3401.935 1403.030 3402.535 1403.430 ;
        RECT 3406.785 1403.030 3407.385 1403.430 ;
      LAYER met4 ;
        RECT 3402.935 1256.035 3406.385 1403.030 ;
      LAYER met4 ;
        RECT 3401.935 1255.635 3402.535 1256.035 ;
        RECT 3406.785 1255.635 3407.385 1256.035 ;
      LAYER met4 ;
        RECT 3407.785 1255.730 3412.435 1403.270 ;
      LAYER met4 ;
        RECT 3412.835 1403.030 3413.435 1403.670 ;
        RECT 3401.935 1255.330 3407.385 1255.635 ;
        RECT 3412.835 1255.330 3413.435 1256.035 ;
      LAYER met4 ;
        RECT 3413.835 1255.730 3418.485 1403.270 ;
      LAYER met4 ;
        RECT 3418.885 1403.030 3419.485 1403.670 ;
        RECT 3418.885 1255.330 3419.485 1256.035 ;
      LAYER met4 ;
        RECT 3419.885 1255.730 3423.335 1403.270 ;
      LAYER met4 ;
        RECT 3423.735 1403.030 3424.335 1403.670 ;
        RECT 3423.735 1255.330 3424.335 1256.035 ;
      LAYER met4 ;
        RECT 3424.735 1255.730 3428.185 1403.270 ;
      LAYER met4 ;
        RECT 3428.585 1403.030 3429.185 1403.670 ;
        RECT 3428.585 1255.330 3429.185 1256.035 ;
      LAYER met4 ;
        RECT 3429.585 1255.730 3434.235 1403.270 ;
      LAYER met4 ;
        RECT 3434.635 1403.030 3435.335 1403.670 ;
        RECT 3434.635 1255.330 3435.335 1256.035 ;
        RECT 3388.535 1253.990 3435.335 1255.330 ;
      LAYER met4 ;
        RECT 3435.735 1254.390 3436.065 1434.910 ;
        RECT 3436.365 1429.855 3439.345 1652.535 ;
      LAYER met4 ;
        RECT 3439.745 1628.670 3440.725 1652.935 ;
      LAYER met4 ;
        RECT 3439.645 1627.000 3440.825 1628.270 ;
      LAYER met4 ;
        RECT 3439.645 1482.000 3440.825 1627.000 ;
      LAYER met4 ;
        RECT 3439.645 1480.730 3440.825 1482.000 ;
      LAYER met4 ;
        RECT 3439.745 1445.160 3440.725 1480.330 ;
      LAYER met4 ;
        RECT 3441.125 1445.560 3444.105 1668.240 ;
      LAYER met4 ;
        RECT 3444.505 1660.310 3588.000 1668.640 ;
      LAYER met4 ;
        RECT 3444.405 1479.390 3444.735 1659.910 ;
      LAYER met4 ;
        RECT 3445.135 1628.670 3588.000 1660.310 ;
        RECT 3445.135 1628.030 3445.835 1628.670 ;
        RECT 3445.135 1482.000 3445.835 1627.000 ;
        RECT 3445.135 1480.330 3445.835 1481.035 ;
      LAYER met4 ;
        RECT 3446.235 1480.730 3450.685 1628.270 ;
      LAYER met4 ;
        RECT 3451.085 1628.030 3451.685 1628.670 ;
        RECT 3451.085 1482.000 3451.685 1627.000 ;
        RECT 3451.085 1480.330 3451.685 1481.035 ;
      LAYER met4 ;
        RECT 3452.085 1480.730 3456.535 1628.270 ;
      LAYER met4 ;
        RECT 3456.935 1628.030 3457.635 1628.670 ;
        RECT 3456.935 1482.000 3457.635 1627.000 ;
        RECT 3456.935 1480.330 3457.635 1481.035 ;
      LAYER met4 ;
        RECT 3458.035 1480.730 3483.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1628.030 3563.385 1628.670 ;
      LAYER met4 ;
        RECT 3563.785 1627.000 3588.000 1628.270 ;
      LAYER met4 ;
        RECT 3483.400 1482.000 3588.000 1627.000 ;
        RECT 3483.400 1480.330 3563.385 1481.035 ;
      LAYER met4 ;
        RECT 3563.785 1480.730 3588.000 1482.000 ;
      LAYER met4 ;
        RECT 3445.135 1478.990 3588.000 1480.330 ;
        RECT 3444.505 1445.160 3588.000 1478.990 ;
        RECT 3439.745 1443.640 3588.000 1445.160 ;
        RECT 3439.745 1429.455 3440.725 1443.640 ;
        RECT 3436.465 1427.935 3440.725 1429.455 ;
        RECT 3388.535 1210.310 3435.965 1253.990 ;
        RECT 198.365 1202.330 199.465 1202.970 ;
        RECT 152.665 1170.690 199.465 1202.330 ;
        RECT 3388.535 1178.670 3435.335 1210.310 ;
        RECT 3388.535 1178.030 3389.635 1178.670 ;
        RECT 152.035 1127.010 199.465 1170.690 ;
        RECT 147.275 960.545 151.535 962.065 ;
        RECT 147.275 946.360 148.255 960.545 ;
        RECT 0.000 944.840 148.255 946.360 ;
        RECT 0.000 911.010 143.495 944.840 ;
        RECT 0.000 909.670 142.865 911.010 ;
      LAYER met4 ;
        RECT 0.000 908.000 24.215 909.270 ;
      LAYER met4 ;
        RECT 24.615 908.965 104.600 909.670 ;
        RECT 0.000 767.000 104.600 908.000 ;
        RECT 0.000 762.000 24.215 767.000 ;
        RECT 0.000 626.000 104.600 762.000 ;
      LAYER met4 ;
        RECT 0.000 624.730 24.215 626.000 ;
      LAYER met4 ;
        RECT 24.615 624.330 104.600 625.035 ;
      LAYER met4 ;
        RECT 105.000 624.730 129.965 909.270 ;
      LAYER met4 ;
        RECT 130.365 908.965 131.065 909.670 ;
        RECT 130.365 767.000 131.065 908.000 ;
        RECT 130.365 626.000 131.065 762.000 ;
        RECT 130.365 624.330 131.065 625.035 ;
      LAYER met4 ;
        RECT 131.465 624.730 135.915 909.270 ;
      LAYER met4 ;
        RECT 136.315 908.965 136.915 909.670 ;
        RECT 136.315 767.000 136.915 908.000 ;
        RECT 136.315 626.000 136.915 762.000 ;
        RECT 136.315 624.330 136.915 625.035 ;
      LAYER met4 ;
        RECT 137.315 624.730 141.765 909.270 ;
      LAYER met4 ;
        RECT 142.165 908.965 142.865 909.670 ;
        RECT 142.165 767.000 142.865 908.000 ;
      LAYER met4 ;
        RECT 143.265 767.000 143.595 910.610 ;
      LAYER met4 ;
        RECT 142.165 626.000 142.865 762.000 ;
        RECT 142.165 624.330 142.865 625.035 ;
        RECT 0.000 552.670 142.865 624.330 ;
      LAYER met4 ;
        RECT 0.000 551.000 24.215 552.270 ;
      LAYER met4 ;
        RECT 24.615 551.965 104.600 552.670 ;
        RECT 0.000 415.000 104.600 551.000 ;
      LAYER met4 ;
        RECT 0.000 413.730 24.215 415.000 ;
      LAYER met4 ;
        RECT 24.615 413.330 104.600 415.000 ;
      LAYER met4 ;
        RECT 105.000 413.730 129.965 552.270 ;
      LAYER met4 ;
        RECT 130.365 551.965 131.065 552.670 ;
        RECT 130.365 413.330 131.065 551.000 ;
      LAYER met4 ;
        RECT 131.465 413.730 135.915 552.270 ;
      LAYER met4 ;
        RECT 136.315 551.965 136.915 552.670 ;
        RECT 136.315 413.330 136.915 551.000 ;
      LAYER met4 ;
        RECT 137.315 413.730 141.765 552.270 ;
      LAYER met4 ;
        RECT 142.165 551.965 142.865 552.670 ;
        RECT 142.165 413.330 142.865 551.000 ;
        RECT 0.000 341.670 142.865 413.330 ;
      LAYER met4 ;
        RECT 0.000 340.000 24.215 341.270 ;
      LAYER met4 ;
        RECT 24.615 340.965 104.600 341.670 ;
        RECT 0.000 204.000 104.600 340.000 ;
      LAYER met4 ;
        RECT 0.000 202.730 24.215 204.000 ;
      LAYER met4 ;
        RECT 24.615 202.330 104.600 202.745 ;
        RECT 0.000 201.745 104.600 202.330 ;
      LAYER met4 ;
        RECT 105.000 202.145 129.965 341.270 ;
      LAYER met4 ;
        RECT 130.365 340.965 131.065 341.670 ;
        RECT 130.365 204.000 131.065 340.000 ;
        RECT 130.365 202.330 131.065 202.745 ;
      LAYER met4 ;
        RECT 131.465 202.730 135.915 341.270 ;
      LAYER met4 ;
        RECT 136.315 340.965 136.915 341.670 ;
        RECT 136.315 204.000 136.915 340.000 ;
        RECT 136.315 202.330 136.915 202.745 ;
      LAYER met4 ;
        RECT 137.315 202.730 141.765 341.270 ;
      LAYER met4 ;
        RECT 142.165 340.965 142.865 341.670 ;
        RECT 142.165 204.000 142.865 340.000 ;
        RECT 142.165 202.330 142.865 202.745 ;
        RECT 130.365 201.745 142.865 202.330 ;
        RECT 0.000 176.425 142.865 201.745 ;
      LAYER met4 ;
        RECT 143.265 176.825 143.595 762.000 ;
        RECT 143.895 177.090 146.875 944.440 ;
      LAYER met4 ;
        RECT 147.275 909.670 148.255 944.840 ;
      LAYER met4 ;
        RECT 147.175 908.000 148.355 909.270 ;
      LAYER met4 ;
        RECT 147.175 767.000 148.355 908.000 ;
        RECT 147.175 626.000 148.355 762.000 ;
      LAYER met4 ;
        RECT 147.175 624.730 148.355 626.000 ;
      LAYER met4 ;
        RECT 147.275 552.670 148.255 624.330 ;
      LAYER met4 ;
        RECT 147.175 551.000 148.355 552.270 ;
      LAYER met4 ;
        RECT 147.175 415.000 148.355 551.000 ;
      LAYER met4 ;
        RECT 147.175 413.730 148.355 415.000 ;
      LAYER met4 ;
        RECT 147.275 341.670 148.255 413.330 ;
      LAYER met4 ;
        RECT 147.175 340.000 148.355 341.270 ;
      LAYER met4 ;
        RECT 147.175 204.000 148.355 340.000 ;
      LAYER met4 ;
        RECT 147.175 182.445 148.355 204.000 ;
        RECT 148.655 183.125 151.635 960.145 ;
        RECT 151.935 955.090 152.265 1126.610 ;
      LAYER met4 ;
        RECT 152.665 1125.670 199.465 1127.010 ;
        RECT 152.665 1124.965 153.365 1125.670 ;
        RECT 152.665 986.330 153.365 986.970 ;
      LAYER met4 ;
        RECT 153.765 986.730 158.415 1125.270 ;
      LAYER met4 ;
        RECT 158.815 1124.965 159.415 1125.670 ;
        RECT 158.815 986.330 159.415 986.970 ;
      LAYER met4 ;
        RECT 159.815 986.730 163.265 1125.270 ;
      LAYER met4 ;
        RECT 163.665 1124.965 164.265 1125.670 ;
        RECT 163.665 986.330 164.265 986.970 ;
      LAYER met4 ;
        RECT 164.665 986.730 168.115 1125.270 ;
      LAYER met4 ;
        RECT 168.515 1124.965 169.115 1125.670 ;
        RECT 168.515 986.330 169.115 986.970 ;
      LAYER met4 ;
        RECT 169.515 986.730 174.165 1125.270 ;
      LAYER met4 ;
        RECT 174.565 1124.965 175.165 1125.670 ;
        RECT 180.615 1125.365 186.065 1125.670 ;
        RECT 174.565 986.330 175.165 986.970 ;
      LAYER met4 ;
        RECT 175.565 986.730 180.215 1125.270 ;
      LAYER met4 ;
        RECT 180.615 1124.965 181.215 1125.365 ;
        RECT 185.465 1124.965 186.065 1125.365 ;
      LAYER met4 ;
        RECT 181.615 986.970 185.065 1124.965 ;
      LAYER met4 ;
        RECT 180.615 986.570 181.215 986.970 ;
        RECT 185.465 986.570 186.065 986.970 ;
      LAYER met4 ;
        RECT 186.465 986.730 191.115 1125.270 ;
      LAYER met4 ;
        RECT 191.515 1124.965 192.115 1125.670 ;
        RECT 180.615 986.330 186.065 986.570 ;
        RECT 191.515 986.330 192.115 986.970 ;
      LAYER met4 ;
        RECT 192.515 986.730 197.965 1125.270 ;
      LAYER met4 ;
        RECT 198.365 1124.965 199.465 1125.670 ;
        RECT 3388.535 1029.330 3389.635 1030.035 ;
      LAYER met4 ;
        RECT 3390.035 1029.730 3395.485 1178.270 ;
      LAYER met4 ;
        RECT 3395.885 1178.030 3396.485 1178.670 ;
        RECT 3401.935 1178.430 3407.385 1178.670 ;
        RECT 3395.885 1029.330 3396.485 1030.035 ;
      LAYER met4 ;
        RECT 3396.885 1029.730 3401.535 1178.270 ;
      LAYER met4 ;
        RECT 3401.935 1178.030 3402.535 1178.430 ;
        RECT 3406.785 1178.030 3407.385 1178.430 ;
      LAYER met4 ;
        RECT 3402.935 1030.035 3406.385 1178.030 ;
      LAYER met4 ;
        RECT 3401.935 1029.635 3402.535 1030.035 ;
        RECT 3406.785 1029.635 3407.385 1030.035 ;
      LAYER met4 ;
        RECT 3407.785 1029.730 3412.435 1178.270 ;
      LAYER met4 ;
        RECT 3412.835 1178.030 3413.435 1178.670 ;
        RECT 3401.935 1029.330 3407.385 1029.635 ;
        RECT 3412.835 1029.330 3413.435 1030.035 ;
      LAYER met4 ;
        RECT 3413.835 1029.730 3418.485 1178.270 ;
      LAYER met4 ;
        RECT 3418.885 1178.030 3419.485 1178.670 ;
        RECT 3418.885 1029.330 3419.485 1030.035 ;
      LAYER met4 ;
        RECT 3419.885 1029.730 3423.335 1178.270 ;
      LAYER met4 ;
        RECT 3423.735 1178.030 3424.335 1178.670 ;
        RECT 3423.735 1029.330 3424.335 1030.035 ;
      LAYER met4 ;
        RECT 3424.735 1029.730 3428.185 1178.270 ;
      LAYER met4 ;
        RECT 3428.585 1178.030 3429.185 1178.670 ;
        RECT 3428.585 1029.330 3429.185 1030.035 ;
      LAYER met4 ;
        RECT 3429.585 1029.730 3434.235 1178.270 ;
      LAYER met4 ;
        RECT 3434.635 1178.030 3435.335 1178.670 ;
        RECT 3434.635 1029.330 3435.335 1030.035 ;
        RECT 3388.535 1027.990 3435.335 1029.330 ;
      LAYER met4 ;
        RECT 3435.735 1028.390 3436.065 1209.910 ;
        RECT 3436.365 1204.855 3439.345 1427.535 ;
      LAYER met4 ;
        RECT 3439.745 1403.670 3440.725 1427.935 ;
      LAYER met4 ;
        RECT 3439.645 1402.000 3440.825 1403.270 ;
      LAYER met4 ;
        RECT 3439.645 1257.000 3440.825 1402.000 ;
      LAYER met4 ;
        RECT 3439.645 1255.730 3440.825 1257.000 ;
      LAYER met4 ;
        RECT 3439.745 1220.160 3440.725 1255.330 ;
      LAYER met4 ;
        RECT 3441.125 1220.560 3444.105 1443.240 ;
      LAYER met4 ;
        RECT 3444.505 1435.310 3588.000 1443.640 ;
      LAYER met4 ;
        RECT 3444.405 1254.390 3444.735 1434.910 ;
      LAYER met4 ;
        RECT 3445.135 1403.670 3588.000 1435.310 ;
        RECT 3445.135 1403.030 3445.835 1403.670 ;
        RECT 3445.135 1257.000 3445.835 1402.000 ;
        RECT 3445.135 1255.330 3445.835 1256.035 ;
      LAYER met4 ;
        RECT 3446.235 1255.730 3450.685 1403.270 ;
      LAYER met4 ;
        RECT 3451.085 1403.030 3451.685 1403.670 ;
        RECT 3451.085 1257.000 3451.685 1402.000 ;
        RECT 3451.085 1255.330 3451.685 1256.035 ;
      LAYER met4 ;
        RECT 3452.085 1255.730 3456.535 1403.270 ;
      LAYER met4 ;
        RECT 3456.935 1403.030 3457.635 1403.670 ;
        RECT 3456.935 1257.000 3457.635 1402.000 ;
        RECT 3456.935 1255.330 3457.635 1256.035 ;
      LAYER met4 ;
        RECT 3458.035 1255.730 3483.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1403.030 3563.385 1403.670 ;
      LAYER met4 ;
        RECT 3563.785 1402.000 3588.000 1403.270 ;
      LAYER met4 ;
        RECT 3483.400 1257.000 3588.000 1402.000 ;
        RECT 3483.400 1255.330 3563.385 1256.035 ;
      LAYER met4 ;
        RECT 3563.785 1255.730 3588.000 1257.000 ;
      LAYER met4 ;
        RECT 3445.135 1253.990 3588.000 1255.330 ;
        RECT 3444.505 1220.160 3588.000 1253.990 ;
        RECT 3439.745 1218.640 3588.000 1220.160 ;
        RECT 3439.745 1204.455 3440.725 1218.640 ;
        RECT 3436.465 1202.935 3440.725 1204.455 ;
        RECT 198.365 986.330 199.465 986.970 ;
        RECT 152.665 954.690 199.465 986.330 ;
        RECT 152.035 911.010 199.465 954.690 ;
        RECT 3388.535 984.310 3435.965 1027.990 ;
        RECT 3388.535 952.670 3435.335 984.310 ;
        RECT 3388.535 952.030 3389.635 952.670 ;
      LAYER met4 ;
        RECT 151.935 767.000 152.265 910.610 ;
      LAYER met4 ;
        RECT 152.665 909.670 199.465 911.010 ;
        RECT 152.665 908.965 153.365 909.670 ;
      LAYER met4 ;
        RECT 153.765 772.000 158.415 909.270 ;
      LAYER met4 ;
        RECT 158.815 908.965 159.415 909.670 ;
      LAYER met4 ;
        RECT 159.815 767.000 163.265 909.270 ;
      LAYER met4 ;
        RECT 163.665 908.965 164.265 909.670 ;
        RECT 148.755 182.045 151.535 182.725 ;
        RECT 147.275 180.025 151.535 182.045 ;
      LAYER met4 ;
        RECT 151.935 180.425 152.265 762.000 ;
      LAYER met4 ;
        RECT 152.665 624.330 153.365 625.035 ;
      LAYER met4 ;
        RECT 153.765 624.730 158.415 767.000 ;
      LAYER met4 ;
        RECT 158.815 624.330 159.415 625.035 ;
      LAYER met4 ;
        RECT 159.815 624.730 163.265 762.000 ;
      LAYER met4 ;
        RECT 163.665 624.330 164.265 625.035 ;
      LAYER met4 ;
        RECT 164.665 624.730 168.115 909.270 ;
      LAYER met4 ;
        RECT 168.515 908.965 169.115 909.670 ;
        RECT 168.515 624.330 169.115 625.035 ;
      LAYER met4 ;
        RECT 169.515 624.730 174.165 909.270 ;
      LAYER met4 ;
        RECT 174.565 908.965 175.165 909.670 ;
        RECT 180.615 909.365 186.065 909.670 ;
        RECT 174.565 624.330 175.165 625.035 ;
      LAYER met4 ;
        RECT 175.565 624.730 180.215 909.270 ;
      LAYER met4 ;
        RECT 180.615 908.965 181.215 909.365 ;
        RECT 185.465 908.965 186.065 909.365 ;
      LAYER met4 ;
        RECT 181.615 767.000 185.065 908.965 ;
        RECT 186.465 772.000 191.115 909.270 ;
      LAYER met4 ;
        RECT 191.515 908.965 192.115 909.670 ;
      LAYER met4 ;
        RECT 181.615 625.035 185.065 762.000 ;
      LAYER met4 ;
        RECT 180.615 624.635 181.215 625.035 ;
        RECT 185.465 624.635 186.065 625.035 ;
      LAYER met4 ;
        RECT 186.465 624.730 191.115 767.000 ;
      LAYER met4 ;
        RECT 180.615 624.330 186.065 624.635 ;
        RECT 191.515 624.330 192.115 625.035 ;
      LAYER met4 ;
        RECT 192.515 624.730 197.965 909.270 ;
      LAYER met4 ;
        RECT 198.365 908.965 199.465 909.670 ;
        RECT 3388.535 804.330 3389.635 805.035 ;
      LAYER met4 ;
        RECT 3390.035 804.730 3395.485 952.270 ;
      LAYER met4 ;
        RECT 3395.885 952.030 3396.485 952.670 ;
        RECT 3401.935 952.430 3407.385 952.670 ;
        RECT 3395.885 804.330 3396.485 805.035 ;
      LAYER met4 ;
        RECT 3396.885 804.730 3401.535 952.270 ;
      LAYER met4 ;
        RECT 3401.935 952.030 3402.535 952.430 ;
        RECT 3406.785 952.030 3407.385 952.430 ;
      LAYER met4 ;
        RECT 3402.935 805.035 3406.385 952.030 ;
      LAYER met4 ;
        RECT 3401.935 804.635 3402.535 805.035 ;
        RECT 3406.785 804.635 3407.385 805.035 ;
      LAYER met4 ;
        RECT 3407.785 804.730 3412.435 952.270 ;
      LAYER met4 ;
        RECT 3412.835 952.030 3413.435 952.670 ;
        RECT 3401.935 804.330 3407.385 804.635 ;
        RECT 3412.835 804.330 3413.435 805.035 ;
      LAYER met4 ;
        RECT 3413.835 804.730 3418.485 952.270 ;
      LAYER met4 ;
        RECT 3418.885 952.030 3419.485 952.670 ;
        RECT 3418.885 804.330 3419.485 805.035 ;
      LAYER met4 ;
        RECT 3419.885 804.730 3423.335 952.270 ;
      LAYER met4 ;
        RECT 3423.735 952.030 3424.335 952.670 ;
        RECT 3423.735 804.330 3424.335 805.035 ;
      LAYER met4 ;
        RECT 3424.735 804.730 3428.185 952.270 ;
      LAYER met4 ;
        RECT 3428.585 952.030 3429.185 952.670 ;
        RECT 3428.585 804.330 3429.185 805.035 ;
      LAYER met4 ;
        RECT 3429.585 804.730 3434.235 952.270 ;
      LAYER met4 ;
        RECT 3434.635 952.030 3435.335 952.670 ;
        RECT 3434.635 804.330 3435.335 805.035 ;
        RECT 3388.535 802.990 3435.335 804.330 ;
      LAYER met4 ;
        RECT 3435.735 803.390 3436.065 983.910 ;
        RECT 3436.365 978.855 3439.345 1202.535 ;
      LAYER met4 ;
        RECT 3439.745 1178.670 3440.725 1202.935 ;
      LAYER met4 ;
        RECT 3439.645 1177.000 3440.825 1178.270 ;
      LAYER met4 ;
        RECT 3439.645 1031.000 3440.825 1177.000 ;
      LAYER met4 ;
        RECT 3439.645 1029.730 3440.825 1031.000 ;
      LAYER met4 ;
        RECT 3439.745 994.160 3440.725 1029.330 ;
      LAYER met4 ;
        RECT 3441.125 994.560 3444.105 1218.240 ;
      LAYER met4 ;
        RECT 3444.505 1210.310 3588.000 1218.640 ;
      LAYER met4 ;
        RECT 3444.405 1028.390 3444.735 1209.910 ;
      LAYER met4 ;
        RECT 3445.135 1178.670 3588.000 1210.310 ;
        RECT 3445.135 1178.030 3445.835 1178.670 ;
        RECT 3445.135 1031.000 3445.835 1177.000 ;
        RECT 3445.135 1029.330 3445.835 1030.035 ;
      LAYER met4 ;
        RECT 3446.235 1029.730 3450.685 1178.270 ;
      LAYER met4 ;
        RECT 3451.085 1178.030 3451.685 1178.670 ;
        RECT 3451.085 1031.000 3451.685 1177.000 ;
        RECT 3451.085 1029.330 3451.685 1030.035 ;
      LAYER met4 ;
        RECT 3452.085 1029.730 3456.535 1178.270 ;
      LAYER met4 ;
        RECT 3456.935 1178.030 3457.635 1178.670 ;
        RECT 3456.935 1031.000 3457.635 1177.000 ;
        RECT 3456.935 1029.330 3457.635 1030.035 ;
      LAYER met4 ;
        RECT 3458.035 1029.730 3483.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1178.030 3563.385 1178.670 ;
      LAYER met4 ;
        RECT 3563.785 1177.000 3588.000 1178.270 ;
      LAYER met4 ;
        RECT 3483.400 1031.000 3588.000 1177.000 ;
        RECT 3483.400 1029.330 3563.385 1030.035 ;
      LAYER met4 ;
        RECT 3563.785 1029.730 3588.000 1031.000 ;
      LAYER met4 ;
        RECT 3445.135 1027.990 3588.000 1029.330 ;
        RECT 3444.505 994.160 3588.000 1027.990 ;
        RECT 3439.745 992.640 3588.000 994.160 ;
        RECT 3439.745 978.455 3440.725 992.640 ;
        RECT 3436.465 976.935 3440.725 978.455 ;
        RECT 3388.535 759.310 3435.965 802.990 ;
        RECT 3388.535 727.670 3435.335 759.310 ;
        RECT 3388.535 727.030 3389.635 727.670 ;
        RECT 152.665 552.670 197.965 624.330 ;
        RECT 3388.535 578.330 3389.635 579.035 ;
      LAYER met4 ;
        RECT 3390.035 578.730 3395.485 727.270 ;
      LAYER met4 ;
        RECT 3395.885 727.030 3396.485 727.670 ;
        RECT 3401.935 727.430 3407.385 727.670 ;
        RECT 3395.885 578.330 3396.485 579.035 ;
      LAYER met4 ;
        RECT 3396.885 578.730 3401.535 727.270 ;
      LAYER met4 ;
        RECT 3401.935 727.030 3402.535 727.430 ;
        RECT 3406.785 727.030 3407.385 727.430 ;
      LAYER met4 ;
        RECT 3402.935 579.035 3406.385 727.030 ;
      LAYER met4 ;
        RECT 3401.935 578.635 3402.535 579.035 ;
        RECT 3406.785 578.635 3407.385 579.035 ;
      LAYER met4 ;
        RECT 3407.785 578.730 3412.435 727.270 ;
      LAYER met4 ;
        RECT 3412.835 727.030 3413.435 727.670 ;
        RECT 3401.935 578.330 3407.385 578.635 ;
        RECT 3412.835 578.330 3413.435 579.035 ;
      LAYER met4 ;
        RECT 3413.835 578.730 3418.485 727.270 ;
      LAYER met4 ;
        RECT 3418.885 727.030 3419.485 727.670 ;
        RECT 3418.885 578.330 3419.485 579.035 ;
      LAYER met4 ;
        RECT 3419.885 578.730 3423.335 727.270 ;
      LAYER met4 ;
        RECT 3423.735 727.030 3424.335 727.670 ;
        RECT 3423.735 578.330 3424.335 579.035 ;
      LAYER met4 ;
        RECT 3424.735 578.730 3428.185 727.270 ;
      LAYER met4 ;
        RECT 3428.585 727.030 3429.185 727.670 ;
        RECT 3428.585 578.330 3429.185 579.035 ;
      LAYER met4 ;
        RECT 3429.585 578.730 3434.235 727.270 ;
      LAYER met4 ;
        RECT 3434.635 727.030 3435.335 727.670 ;
        RECT 3434.635 578.330 3435.335 579.035 ;
        RECT 3388.535 576.990 3435.335 578.330 ;
      LAYER met4 ;
        RECT 3435.735 577.390 3436.065 758.910 ;
        RECT 3436.365 753.855 3439.345 976.535 ;
      LAYER met4 ;
        RECT 3439.745 952.670 3440.725 976.935 ;
      LAYER met4 ;
        RECT 3439.645 951.000 3440.825 952.270 ;
      LAYER met4 ;
        RECT 3439.645 806.000 3440.825 951.000 ;
      LAYER met4 ;
        RECT 3439.645 804.730 3440.825 806.000 ;
      LAYER met4 ;
        RECT 3439.745 769.160 3440.725 804.330 ;
      LAYER met4 ;
        RECT 3441.125 769.560 3444.105 992.240 ;
      LAYER met4 ;
        RECT 3444.505 984.310 3588.000 992.640 ;
      LAYER met4 ;
        RECT 3444.405 803.390 3444.735 983.910 ;
      LAYER met4 ;
        RECT 3445.135 952.670 3588.000 984.310 ;
        RECT 3445.135 952.030 3445.835 952.670 ;
        RECT 3445.135 806.000 3445.835 951.000 ;
        RECT 3445.135 804.330 3445.835 805.035 ;
      LAYER met4 ;
        RECT 3446.235 804.730 3450.685 952.270 ;
      LAYER met4 ;
        RECT 3451.085 952.030 3451.685 952.670 ;
        RECT 3451.085 806.000 3451.685 951.000 ;
        RECT 3451.085 804.330 3451.685 805.035 ;
      LAYER met4 ;
        RECT 3452.085 804.730 3456.535 952.270 ;
      LAYER met4 ;
        RECT 3456.935 952.030 3457.635 952.670 ;
        RECT 3456.935 806.000 3457.635 951.000 ;
        RECT 3456.935 804.330 3457.635 805.035 ;
      LAYER met4 ;
        RECT 3458.035 804.730 3483.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 952.030 3563.385 952.670 ;
      LAYER met4 ;
        RECT 3563.785 951.000 3588.000 952.270 ;
      LAYER met4 ;
        RECT 3483.400 806.000 3588.000 951.000 ;
        RECT 3483.400 804.330 3563.385 805.035 ;
      LAYER met4 ;
        RECT 3563.785 804.730 3588.000 806.000 ;
      LAYER met4 ;
        RECT 3445.135 802.990 3588.000 804.330 ;
        RECT 3444.505 769.160 3588.000 802.990 ;
        RECT 3439.745 767.640 3588.000 769.160 ;
        RECT 3439.745 753.455 3440.725 767.640 ;
        RECT 3436.465 751.935 3440.725 753.455 ;
        RECT 152.665 551.965 153.365 552.670 ;
        RECT 152.665 413.330 153.365 415.000 ;
      LAYER met4 ;
        RECT 153.765 413.730 158.415 552.270 ;
      LAYER met4 ;
        RECT 158.815 551.965 159.415 552.670 ;
        RECT 158.815 413.330 159.415 415.000 ;
      LAYER met4 ;
        RECT 159.815 413.730 163.265 552.270 ;
      LAYER met4 ;
        RECT 163.665 551.965 164.265 552.670 ;
        RECT 163.665 413.330 164.265 415.000 ;
      LAYER met4 ;
        RECT 164.665 413.730 168.115 552.270 ;
      LAYER met4 ;
        RECT 168.515 551.965 169.115 552.670 ;
        RECT 168.515 413.330 169.115 415.000 ;
      LAYER met4 ;
        RECT 169.515 413.730 174.165 552.270 ;
      LAYER met4 ;
        RECT 174.565 551.965 175.165 552.670 ;
        RECT 180.615 552.365 186.065 552.670 ;
        RECT 174.565 413.330 175.165 415.000 ;
      LAYER met4 ;
        RECT 175.565 413.730 180.215 552.270 ;
      LAYER met4 ;
        RECT 180.615 551.965 181.215 552.365 ;
        RECT 185.465 551.965 186.065 552.365 ;
        RECT 180.615 413.635 181.215 415.000 ;
      LAYER met4 ;
        RECT 181.615 414.035 185.065 551.965 ;
      LAYER met4 ;
        RECT 185.465 413.635 186.065 415.000 ;
      LAYER met4 ;
        RECT 186.465 413.730 191.115 552.270 ;
      LAYER met4 ;
        RECT 191.515 551.965 192.115 552.670 ;
        RECT 180.615 413.330 186.065 413.635 ;
        RECT 191.515 413.330 192.115 415.000 ;
      LAYER met4 ;
        RECT 192.515 413.730 197.965 552.270 ;
      LAYER met4 ;
        RECT 3388.535 533.310 3435.965 576.990 ;
        RECT 3388.535 501.670 3435.335 533.310 ;
        RECT 3388.535 501.030 3389.635 501.670 ;
        RECT 152.665 341.670 197.965 413.330 ;
        RECT 152.665 340.965 153.365 341.670 ;
        RECT 152.665 202.330 153.365 202.745 ;
      LAYER met4 ;
        RECT 153.765 202.730 158.415 341.270 ;
      LAYER met4 ;
        RECT 158.815 340.965 159.415 341.670 ;
        RECT 158.815 202.330 159.415 202.745 ;
      LAYER met4 ;
        RECT 159.815 202.730 163.265 341.270 ;
      LAYER met4 ;
        RECT 163.665 340.965 164.265 341.670 ;
        RECT 163.665 202.330 164.265 202.745 ;
      LAYER met4 ;
        RECT 164.665 202.730 168.115 341.270 ;
      LAYER met4 ;
        RECT 168.515 340.965 169.115 341.670 ;
        RECT 168.515 202.330 169.115 202.745 ;
      LAYER met4 ;
        RECT 169.515 202.730 174.165 341.270 ;
      LAYER met4 ;
        RECT 174.565 340.965 175.165 341.670 ;
        RECT 180.615 341.365 186.065 341.670 ;
        RECT 174.565 202.330 175.165 202.745 ;
      LAYER met4 ;
        RECT 175.565 202.730 180.215 341.270 ;
      LAYER met4 ;
        RECT 180.615 340.965 181.215 341.365 ;
        RECT 185.465 340.965 186.065 341.365 ;
      LAYER met4 ;
        RECT 181.615 202.745 185.065 340.965 ;
      LAYER met4 ;
        RECT 180.615 202.345 181.215 202.745 ;
        RECT 185.465 202.345 186.065 202.745 ;
      LAYER met4 ;
        RECT 186.465 202.730 191.115 341.270 ;
      LAYER met4 ;
        RECT 191.515 340.965 192.115 341.670 ;
        RECT 180.615 202.330 186.065 202.345 ;
        RECT 191.515 202.330 192.115 202.745 ;
      LAYER met4 ;
        RECT 192.515 202.730 197.965 341.270 ;
      LAYER met4 ;
        RECT 198.365 202.330 200.000 202.745 ;
        RECT 152.665 198.365 200.000 202.330 ;
        RECT 933.030 198.365 1011.035 199.465 ;
        RECT 1476.030 198.365 1554.035 199.465 ;
        RECT 1750.030 198.365 1828.035 199.465 ;
        RECT 2024.030 198.365 2102.035 199.465 ;
        RECT 2298.030 198.365 2376.035 199.465 ;
        RECT 2572.030 198.365 2650.035 199.465 ;
        RECT 3385.255 198.365 3389.635 200.000 ;
        RECT 152.665 192.115 197.250 198.365 ;
      LAYER met4 ;
        RECT 197.650 192.515 395.270 197.965 ;
      LAYER met4 ;
        RECT 395.670 192.115 467.330 197.965 ;
      LAYER met4 ;
        RECT 467.730 192.515 664.270 197.965 ;
      LAYER met4 ;
        RECT 664.670 192.115 736.330 197.965 ;
      LAYER met4 ;
        RECT 736.730 192.515 933.270 197.965 ;
      LAYER met4 ;
        RECT 933.670 192.115 1010.330 198.365 ;
      LAYER met4 ;
        RECT 1010.730 192.515 1207.270 197.965 ;
      LAYER met4 ;
        RECT 1207.670 192.115 1279.330 197.965 ;
      LAYER met4 ;
        RECT 1279.730 192.515 1476.270 197.965 ;
      LAYER met4 ;
        RECT 1476.670 192.115 1553.330 198.365 ;
      LAYER met4 ;
        RECT 1553.730 192.515 1750.270 197.965 ;
      LAYER met4 ;
        RECT 1750.670 192.115 1827.330 198.365 ;
      LAYER met4 ;
        RECT 1827.730 192.515 2024.270 197.965 ;
      LAYER met4 ;
        RECT 2024.670 192.115 2101.330 198.365 ;
      LAYER met4 ;
        RECT 2101.730 192.515 2298.270 197.965 ;
      LAYER met4 ;
        RECT 2298.670 192.115 2375.330 198.365 ;
      LAYER met4 ;
        RECT 2375.730 192.515 2572.270 197.965 ;
      LAYER met4 ;
        RECT 2572.670 192.115 2649.330 198.365 ;
      LAYER met4 ;
        RECT 2649.730 192.515 2846.270 197.965 ;
      LAYER met4 ;
        RECT 2846.670 192.115 2918.330 197.965 ;
      LAYER met4 ;
        RECT 2918.730 192.515 3115.270 197.965 ;
      LAYER met4 ;
        RECT 3115.670 192.115 3187.330 197.965 ;
      LAYER met4 ;
        RECT 3187.730 192.515 3385.270 197.965 ;
      LAYER met4 ;
        RECT 3385.670 197.250 3389.635 198.365 ;
      LAYER met4 ;
        RECT 3390.035 197.650 3395.485 501.270 ;
      LAYER met4 ;
        RECT 3395.885 501.030 3396.485 501.670 ;
        RECT 3401.935 501.430 3407.385 501.670 ;
      LAYER met4 ;
        RECT 3396.885 355.000 3401.535 501.270 ;
      LAYER met4 ;
        RECT 3401.935 501.030 3402.535 501.430 ;
        RECT 3406.785 501.030 3407.385 501.430 ;
      LAYER met4 ;
        RECT 3402.935 350.000 3406.385 501.030 ;
      LAYER met4 ;
        RECT 3395.885 197.250 3396.485 200.000 ;
        RECT 3385.670 195.815 3396.485 197.250 ;
      LAYER met4 ;
        RECT 3396.885 196.215 3401.535 350.000 ;
      LAYER met4 ;
        RECT 3401.935 198.130 3402.535 200.000 ;
      LAYER met4 ;
        RECT 3402.935 198.530 3406.385 345.000 ;
      LAYER met4 ;
        RECT 3406.785 198.130 3407.385 200.000 ;
      LAYER met4 ;
        RECT 3407.785 198.475 3412.435 501.270 ;
      LAYER met4 ;
        RECT 3412.835 501.030 3413.435 501.670 ;
        RECT 3401.935 198.075 3407.385 198.130 ;
        RECT 3412.835 198.075 3413.435 200.000 ;
      LAYER met4 ;
        RECT 3413.835 198.400 3418.485 501.270 ;
      LAYER met4 ;
        RECT 3418.885 501.030 3419.485 501.670 ;
        RECT 3401.935 198.000 3413.435 198.075 ;
        RECT 3418.885 198.215 3419.485 200.000 ;
      LAYER met4 ;
        RECT 3419.885 198.615 3423.335 501.270 ;
      LAYER met4 ;
        RECT 3423.735 501.030 3424.335 501.670 ;
      LAYER met4 ;
        RECT 3424.735 350.000 3428.185 501.270 ;
      LAYER met4 ;
        RECT 3428.585 501.030 3429.185 501.670 ;
      LAYER met4 ;
        RECT 3429.585 355.000 3434.235 501.270 ;
      LAYER met4 ;
        RECT 3434.635 501.030 3435.335 501.670 ;
      LAYER met4 ;
        RECT 3435.735 350.000 3436.065 532.910 ;
        RECT 3436.365 527.855 3439.345 751.535 ;
      LAYER met4 ;
        RECT 3439.745 727.670 3440.725 751.935 ;
      LAYER met4 ;
        RECT 3439.645 726.000 3440.825 727.270 ;
      LAYER met4 ;
        RECT 3439.645 580.000 3440.825 726.000 ;
      LAYER met4 ;
        RECT 3439.645 578.730 3440.825 580.000 ;
      LAYER met4 ;
        RECT 3439.745 543.160 3440.725 578.330 ;
      LAYER met4 ;
        RECT 3441.125 543.560 3444.105 767.240 ;
      LAYER met4 ;
        RECT 3444.505 759.310 3588.000 767.640 ;
      LAYER met4 ;
        RECT 3444.405 577.390 3444.735 758.910 ;
      LAYER met4 ;
        RECT 3445.135 727.670 3588.000 759.310 ;
        RECT 3445.135 727.030 3445.835 727.670 ;
        RECT 3445.135 580.000 3445.835 726.000 ;
        RECT 3445.135 578.330 3445.835 579.035 ;
      LAYER met4 ;
        RECT 3446.235 578.730 3450.685 727.270 ;
      LAYER met4 ;
        RECT 3451.085 727.030 3451.685 727.670 ;
        RECT 3451.085 580.000 3451.685 726.000 ;
        RECT 3451.085 578.330 3451.685 579.035 ;
      LAYER met4 ;
        RECT 3452.085 578.730 3456.535 727.270 ;
      LAYER met4 ;
        RECT 3456.935 727.030 3457.635 727.670 ;
        RECT 3456.935 580.000 3457.635 726.000 ;
        RECT 3456.935 578.330 3457.635 579.035 ;
      LAYER met4 ;
        RECT 3458.035 578.730 3483.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 727.030 3563.385 727.670 ;
      LAYER met4 ;
        RECT 3563.785 726.000 3588.000 727.270 ;
      LAYER met4 ;
        RECT 3483.400 580.000 3588.000 726.000 ;
        RECT 3483.400 578.330 3563.385 579.035 ;
      LAYER met4 ;
        RECT 3563.785 578.730 3588.000 580.000 ;
      LAYER met4 ;
        RECT 3445.135 576.990 3588.000 578.330 ;
        RECT 3444.505 543.160 3588.000 576.990 ;
        RECT 3439.745 541.640 3588.000 543.160 ;
        RECT 3439.745 527.455 3440.725 541.640 ;
        RECT 3436.465 525.935 3440.725 527.455 ;
        RECT 3423.735 198.265 3424.335 200.000 ;
      LAYER met4 ;
        RECT 3424.735 198.665 3428.185 345.000 ;
      LAYER met4 ;
        RECT 3428.585 198.265 3429.185 200.000 ;
      LAYER met4 ;
        RECT 3429.585 198.525 3434.235 350.000 ;
      LAYER met4 ;
        RECT 3423.735 198.215 3429.185 198.265 ;
        RECT 3418.885 198.125 3429.185 198.215 ;
        RECT 3434.635 198.125 3435.335 200.000 ;
        RECT 3418.885 198.000 3435.335 198.125 ;
        RECT 3401.935 195.815 3435.335 198.000 ;
        RECT 3385.670 192.115 3435.335 195.815 ;
        RECT 152.665 191.515 200.000 192.115 ;
        RECT 394.965 191.515 468.035 192.115 ;
        RECT 663.965 191.515 737.035 192.115 ;
        RECT 933.030 191.515 1011.035 192.115 ;
        RECT 1206.000 191.515 1280.035 192.115 ;
        RECT 1476.030 191.515 1554.035 192.115 ;
        RECT 1750.030 191.515 1828.035 192.115 ;
        RECT 2024.030 191.515 2102.035 192.115 ;
        RECT 2298.030 191.515 2376.035 192.115 ;
        RECT 2572.030 191.515 2650.035 192.115 ;
        RECT 2845.965 191.515 2919.035 192.115 ;
        RECT 3114.965 191.515 3188.035 192.115 ;
        RECT 3385.255 191.515 3435.335 192.115 ;
        RECT 152.665 186.065 195.815 191.515 ;
      LAYER met4 ;
        RECT 196.215 186.465 395.270 191.115 ;
      LAYER met4 ;
        RECT 395.670 186.065 467.330 191.515 ;
      LAYER met4 ;
        RECT 467.730 186.465 664.270 191.115 ;
      LAYER met4 ;
        RECT 664.670 186.065 736.330 191.515 ;
      LAYER met4 ;
        RECT 736.730 186.465 933.270 191.115 ;
      LAYER met4 ;
        RECT 933.670 186.065 1010.330 191.515 ;
      LAYER met4 ;
        RECT 1010.730 186.465 1207.270 191.115 ;
      LAYER met4 ;
        RECT 1207.670 186.065 1279.330 191.515 ;
      LAYER met4 ;
        RECT 1279.730 186.465 1476.270 191.115 ;
      LAYER met4 ;
        RECT 1476.670 186.065 1553.330 191.515 ;
      LAYER met4 ;
        RECT 1553.730 186.465 1750.270 191.115 ;
      LAYER met4 ;
        RECT 1750.670 186.065 1827.330 191.515 ;
      LAYER met4 ;
        RECT 1827.730 186.465 2024.270 191.115 ;
      LAYER met4 ;
        RECT 2024.670 186.065 2101.330 191.515 ;
      LAYER met4 ;
        RECT 2101.730 186.465 2298.270 191.115 ;
      LAYER met4 ;
        RECT 2298.670 186.065 2375.330 191.515 ;
      LAYER met4 ;
        RECT 2375.730 186.465 2572.270 191.115 ;
      LAYER met4 ;
        RECT 2572.670 186.065 2649.330 191.515 ;
      LAYER met4 ;
        RECT 2649.730 186.465 2846.270 191.115 ;
      LAYER met4 ;
        RECT 2846.670 186.065 2918.330 191.515 ;
      LAYER met4 ;
        RECT 2918.730 186.465 3115.270 191.115 ;
      LAYER met4 ;
        RECT 3115.670 186.065 3187.330 191.515 ;
      LAYER met4 ;
        RECT 3187.730 186.465 3385.270 191.115 ;
      LAYER met4 ;
        RECT 3385.670 186.065 3435.335 191.515 ;
        RECT 152.665 185.465 200.000 186.065 ;
        RECT 394.965 185.465 468.035 186.065 ;
        RECT 663.965 185.465 737.035 186.065 ;
        RECT 933.030 185.465 1011.035 186.065 ;
        RECT 1206.000 185.465 1280.035 186.065 ;
        RECT 1476.030 185.465 1554.035 186.065 ;
        RECT 1750.030 185.465 1828.035 186.065 ;
        RECT 2024.030 185.465 2102.035 186.065 ;
        RECT 2298.030 185.465 2376.035 186.065 ;
        RECT 2572.030 185.465 2650.035 186.065 ;
        RECT 2845.965 185.465 2919.035 186.065 ;
        RECT 3114.965 185.465 3188.035 186.065 ;
        RECT 3385.255 185.465 3435.335 186.065 ;
        RECT 152.665 181.215 198.130 185.465 ;
      LAYER met4 ;
        RECT 198.530 181.615 394.965 185.065 ;
      LAYER met4 ;
        RECT 395.365 181.215 467.635 185.465 ;
        RECT 664.365 181.215 736.635 185.465 ;
      LAYER met4 ;
        RECT 737.035 181.615 933.030 185.065 ;
      LAYER met4 ;
        RECT 933.430 181.215 1010.635 185.465 ;
      LAYER met4 ;
        RECT 1011.035 181.615 1206.965 185.065 ;
      LAYER met4 ;
        RECT 1207.365 181.215 1279.635 185.465 ;
      LAYER met4 ;
        RECT 1280.035 181.615 1476.030 185.065 ;
      LAYER met4 ;
        RECT 1476.430 181.215 1553.635 185.465 ;
      LAYER met4 ;
        RECT 1554.035 181.615 1750.030 185.065 ;
      LAYER met4 ;
        RECT 1750.430 181.215 1827.635 185.465 ;
      LAYER met4 ;
        RECT 1828.035 181.615 2024.030 185.065 ;
      LAYER met4 ;
        RECT 2024.430 181.215 2101.635 185.465 ;
      LAYER met4 ;
        RECT 2102.035 181.615 2298.030 185.065 ;
      LAYER met4 ;
        RECT 2298.430 181.215 2375.635 185.465 ;
      LAYER met4 ;
        RECT 2376.035 181.615 2572.030 185.065 ;
      LAYER met4 ;
        RECT 2572.430 181.215 2649.635 185.465 ;
      LAYER met4 ;
        RECT 2650.035 181.615 2845.965 185.065 ;
      LAYER met4 ;
        RECT 2846.365 181.215 2918.635 185.465 ;
      LAYER met4 ;
        RECT 2919.035 181.615 3114.965 185.065 ;
      LAYER met4 ;
        RECT 3115.365 181.215 3187.635 185.465 ;
      LAYER met4 ;
        RECT 3188.035 181.615 3385.255 185.065 ;
      LAYER met4 ;
        RECT 3385.655 181.215 3435.335 185.465 ;
        RECT 152.665 180.615 200.000 181.215 ;
        RECT 394.965 180.615 468.035 181.215 ;
        RECT 663.965 180.615 737.035 181.215 ;
        RECT 933.030 180.615 1011.035 181.215 ;
        RECT 1206.000 180.615 1280.035 181.215 ;
        RECT 1476.030 180.615 1554.035 181.215 ;
        RECT 1750.030 180.615 1828.035 181.215 ;
        RECT 2024.030 180.615 2102.035 181.215 ;
        RECT 2298.030 180.615 2376.035 181.215 ;
        RECT 2572.030 180.615 2650.035 181.215 ;
        RECT 2845.965 180.615 2919.035 181.215 ;
        RECT 3114.965 180.615 3188.035 181.215 ;
        RECT 3385.255 180.615 3435.335 181.215 ;
        RECT 152.665 180.025 198.075 180.615 ;
        RECT 147.275 176.690 198.075 180.025 ;
        RECT 143.995 176.425 198.075 176.690 ;
        RECT 0.000 175.165 198.075 176.425 ;
      LAYER met4 ;
        RECT 198.475 175.565 395.270 180.215 ;
      LAYER met4 ;
        RECT 395.670 175.165 467.330 180.615 ;
      LAYER met4 ;
        RECT 467.730 175.565 664.270 180.215 ;
      LAYER met4 ;
        RECT 664.670 175.165 736.330 180.615 ;
      LAYER met4 ;
        RECT 736.730 175.565 933.270 180.215 ;
      LAYER met4 ;
        RECT 933.670 175.165 1010.330 180.615 ;
      LAYER met4 ;
        RECT 1010.730 175.565 1207.270 180.215 ;
      LAYER met4 ;
        RECT 1207.670 175.165 1279.330 180.615 ;
      LAYER met4 ;
        RECT 1279.730 175.565 1476.270 180.215 ;
      LAYER met4 ;
        RECT 1476.670 175.165 1553.330 180.615 ;
      LAYER met4 ;
        RECT 1553.730 175.565 1750.270 180.215 ;
      LAYER met4 ;
        RECT 1750.670 175.165 1827.330 180.615 ;
      LAYER met4 ;
        RECT 1827.730 175.565 2024.270 180.215 ;
      LAYER met4 ;
        RECT 2024.670 175.165 2101.330 180.615 ;
      LAYER met4 ;
        RECT 2101.730 175.565 2298.270 180.215 ;
      LAYER met4 ;
        RECT 2298.670 175.165 2375.330 180.615 ;
      LAYER met4 ;
        RECT 2375.730 175.565 2572.270 180.215 ;
      LAYER met4 ;
        RECT 2572.670 175.165 2649.330 180.615 ;
      LAYER met4 ;
        RECT 2649.730 175.565 2846.270 180.215 ;
      LAYER met4 ;
        RECT 2846.670 175.165 2918.330 180.615 ;
      LAYER met4 ;
        RECT 2918.730 175.565 3115.270 180.215 ;
      LAYER met4 ;
        RECT 3115.670 175.165 3187.330 180.615 ;
      LAYER met4 ;
        RECT 3187.730 175.565 3385.270 180.215 ;
      LAYER met4 ;
        RECT 3385.670 180.025 3435.335 180.615 ;
      LAYER met4 ;
        RECT 3435.735 180.425 3436.065 345.000 ;
      LAYER met4 ;
        RECT 3385.670 178.665 3435.965 180.025 ;
      LAYER met4 ;
        RECT 3436.365 179.065 3439.345 525.535 ;
      LAYER met4 ;
        RECT 3439.745 501.670 3440.725 525.935 ;
      LAYER met4 ;
        RECT 3439.645 500.000 3440.825 501.270 ;
      LAYER met4 ;
        RECT 3439.645 350.000 3440.825 500.000 ;
        RECT 3439.645 200.000 3440.825 345.000 ;
        RECT 3385.670 178.050 3439.245 178.665 ;
      LAYER met4 ;
        RECT 3439.645 178.450 3440.825 200.000 ;
      LAYER met4 ;
        RECT 3385.670 176.690 3440.725 178.050 ;
      LAYER met4 ;
        RECT 3441.125 177.090 3444.105 541.240 ;
      LAYER met4 ;
        RECT 3444.505 533.310 3588.000 541.640 ;
      LAYER met4 ;
        RECT 3444.405 350.000 3444.735 532.910 ;
      LAYER met4 ;
        RECT 3445.135 501.670 3588.000 533.310 ;
        RECT 3445.135 501.030 3445.835 501.670 ;
        RECT 3445.135 350.000 3445.835 500.000 ;
      LAYER met4 ;
        RECT 3444.405 176.825 3444.735 345.000 ;
      LAYER met4 ;
        RECT 3445.135 197.975 3445.835 345.000 ;
      LAYER met4 ;
        RECT 3446.235 198.375 3450.685 501.270 ;
      LAYER met4 ;
        RECT 3451.085 501.030 3451.685 501.670 ;
        RECT 3451.085 350.000 3451.685 500.000 ;
        RECT 3451.085 198.120 3451.685 345.000 ;
      LAYER met4 ;
        RECT 3452.085 198.520 3456.535 501.270 ;
      LAYER met4 ;
        RECT 3456.935 501.030 3457.635 501.670 ;
        RECT 3456.935 350.000 3457.635 500.000 ;
        RECT 3456.935 198.120 3457.635 345.000 ;
        RECT 3451.085 197.975 3457.635 198.120 ;
        RECT 3445.135 196.955 3457.635 197.975 ;
      LAYER met4 ;
        RECT 3458.035 197.355 3483.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 501.030 3563.385 501.670 ;
      LAYER met4 ;
        RECT 3563.785 500.000 3588.000 501.270 ;
      LAYER met4 ;
        RECT 3483.400 350.000 3588.000 500.000 ;
        RECT 3563.785 345.000 3588.000 350.000 ;
        RECT 3483.400 200.000 3588.000 345.000 ;
        RECT 3483.400 198.165 3563.385 200.000 ;
      LAYER met4 ;
        RECT 3563.785 198.565 3588.000 200.000 ;
      LAYER met4 ;
        RECT 3483.400 196.955 3588.000 198.165 ;
        RECT 3385.670 176.425 3444.005 176.690 ;
        RECT 3445.135 176.425 3588.000 196.955 ;
        RECT 3385.670 175.165 3588.000 176.425 ;
        RECT 0.000 174.565 200.000 175.165 ;
        RECT 394.965 174.565 468.035 175.165 ;
        RECT 663.965 174.565 737.035 175.165 ;
        RECT 933.030 174.565 1011.035 175.165 ;
        RECT 1206.000 174.565 1280.035 175.165 ;
        RECT 1476.030 174.565 1554.035 175.165 ;
        RECT 1750.030 174.565 1828.035 175.165 ;
        RECT 2024.030 174.565 2102.035 175.165 ;
        RECT 2298.030 174.565 2376.035 175.165 ;
        RECT 2572.030 174.565 2650.035 175.165 ;
        RECT 2845.965 174.565 2919.035 175.165 ;
        RECT 3114.965 174.565 3188.035 175.165 ;
        RECT 3385.255 174.565 3588.000 175.165 ;
        RECT 0.000 169.115 198.000 174.565 ;
      LAYER met4 ;
        RECT 198.400 169.515 395.270 174.165 ;
      LAYER met4 ;
        RECT 395.670 169.115 467.330 174.565 ;
      LAYER met4 ;
        RECT 467.730 169.515 664.270 174.165 ;
      LAYER met4 ;
        RECT 664.670 169.115 736.330 174.565 ;
      LAYER met4 ;
        RECT 736.730 169.515 933.270 174.165 ;
      LAYER met4 ;
        RECT 933.670 169.115 1010.330 174.565 ;
      LAYER met4 ;
        RECT 1010.730 169.515 1207.270 174.165 ;
      LAYER met4 ;
        RECT 1207.670 169.115 1279.330 174.565 ;
      LAYER met4 ;
        RECT 1279.730 169.515 1476.270 174.165 ;
      LAYER met4 ;
        RECT 1476.670 169.115 1553.330 174.565 ;
      LAYER met4 ;
        RECT 1553.730 169.515 1750.270 174.165 ;
      LAYER met4 ;
        RECT 1750.670 169.115 1827.330 174.565 ;
      LAYER met4 ;
        RECT 1827.730 169.515 2024.270 174.165 ;
      LAYER met4 ;
        RECT 2024.670 169.115 2101.330 174.565 ;
      LAYER met4 ;
        RECT 2101.730 169.515 2298.270 174.165 ;
      LAYER met4 ;
        RECT 2298.670 169.115 2375.330 174.565 ;
      LAYER met4 ;
        RECT 2375.730 169.515 2572.270 174.165 ;
      LAYER met4 ;
        RECT 2572.670 169.115 2649.330 174.565 ;
      LAYER met4 ;
        RECT 2649.730 169.515 2846.270 174.165 ;
      LAYER met4 ;
        RECT 2846.670 169.115 2918.330 174.565 ;
      LAYER met4 ;
        RECT 2918.730 169.515 3115.270 174.165 ;
      LAYER met4 ;
        RECT 3115.670 169.115 3187.330 174.565 ;
      LAYER met4 ;
        RECT 3187.730 169.515 3385.270 174.165 ;
      LAYER met4 ;
        RECT 3385.670 169.115 3588.000 174.565 ;
        RECT 0.000 168.515 200.000 169.115 ;
        RECT 394.965 168.515 468.035 169.115 ;
        RECT 663.965 168.515 737.035 169.115 ;
        RECT 933.030 168.515 1011.035 169.115 ;
        RECT 1206.000 168.515 1280.035 169.115 ;
        RECT 1476.030 168.515 1554.035 169.115 ;
        RECT 1750.030 168.515 1828.035 169.115 ;
        RECT 2024.030 168.515 2102.035 169.115 ;
        RECT 2298.030 168.515 2376.035 169.115 ;
        RECT 2572.030 168.515 2650.035 169.115 ;
        RECT 2845.965 168.515 2919.035 169.115 ;
        RECT 3114.965 168.515 3188.035 169.115 ;
        RECT 3385.255 168.515 3588.000 169.115 ;
        RECT 0.000 164.265 198.215 168.515 ;
      LAYER met4 ;
        RECT 198.615 164.665 395.270 168.115 ;
      LAYER met4 ;
        RECT 395.670 164.265 467.330 168.515 ;
      LAYER met4 ;
        RECT 467.730 164.665 664.270 168.115 ;
      LAYER met4 ;
        RECT 664.670 164.265 736.330 168.515 ;
      LAYER met4 ;
        RECT 736.730 164.665 933.270 168.115 ;
      LAYER met4 ;
        RECT 933.670 164.265 1010.330 168.515 ;
      LAYER met4 ;
        RECT 1010.730 164.665 1207.270 168.115 ;
      LAYER met4 ;
        RECT 1207.670 164.265 1279.330 168.515 ;
      LAYER met4 ;
        RECT 1279.730 164.665 1476.270 168.115 ;
      LAYER met4 ;
        RECT 1476.670 164.265 1553.330 168.515 ;
      LAYER met4 ;
        RECT 1553.730 164.665 1750.270 168.115 ;
      LAYER met4 ;
        RECT 1750.670 164.265 1827.330 168.515 ;
      LAYER met4 ;
        RECT 1827.730 164.665 2024.270 168.115 ;
      LAYER met4 ;
        RECT 2024.670 164.265 2101.330 168.515 ;
      LAYER met4 ;
        RECT 2101.730 164.665 2298.270 168.115 ;
      LAYER met4 ;
        RECT 2298.670 164.265 2375.330 168.515 ;
      LAYER met4 ;
        RECT 2375.730 164.665 2572.270 168.115 ;
      LAYER met4 ;
        RECT 2572.670 164.265 2649.330 168.515 ;
      LAYER met4 ;
        RECT 2649.730 164.665 2846.270 168.115 ;
      LAYER met4 ;
        RECT 2846.670 164.265 2918.330 168.515 ;
      LAYER met4 ;
        RECT 2918.730 164.665 3115.270 168.115 ;
      LAYER met4 ;
        RECT 3115.670 164.265 3187.330 168.515 ;
      LAYER met4 ;
        RECT 3187.730 164.665 3385.270 168.115 ;
      LAYER met4 ;
        RECT 3385.670 164.265 3588.000 168.515 ;
        RECT 0.000 163.665 200.000 164.265 ;
        RECT 394.965 163.665 468.035 164.265 ;
        RECT 663.965 163.665 737.035 164.265 ;
        RECT 933.030 163.665 1011.035 164.265 ;
        RECT 1206.000 163.665 1280.035 164.265 ;
        RECT 1476.030 163.665 1554.035 164.265 ;
        RECT 1750.030 163.665 1828.035 164.265 ;
        RECT 2024.030 163.665 2102.035 164.265 ;
        RECT 2298.030 163.665 2376.035 164.265 ;
        RECT 2572.030 163.665 2650.035 164.265 ;
        RECT 2845.965 163.665 2919.035 164.265 ;
        RECT 3114.965 163.665 3188.035 164.265 ;
        RECT 3385.255 163.665 3588.000 164.265 ;
        RECT 0.000 159.415 198.265 163.665 ;
      LAYER met4 ;
        RECT 198.665 159.815 395.270 163.265 ;
      LAYER met4 ;
        RECT 395.670 159.415 467.330 163.665 ;
      LAYER met4 ;
        RECT 467.730 159.815 664.270 163.265 ;
      LAYER met4 ;
        RECT 664.670 159.415 736.330 163.665 ;
      LAYER met4 ;
        RECT 736.730 159.815 933.270 163.265 ;
      LAYER met4 ;
        RECT 933.670 159.415 1010.330 163.665 ;
      LAYER met4 ;
        RECT 1010.730 159.815 1207.270 163.265 ;
      LAYER met4 ;
        RECT 1207.670 159.415 1279.330 163.665 ;
      LAYER met4 ;
        RECT 1279.730 159.815 1476.270 163.265 ;
      LAYER met4 ;
        RECT 1476.670 159.415 1553.330 163.665 ;
      LAYER met4 ;
        RECT 1553.730 159.815 1750.270 163.265 ;
      LAYER met4 ;
        RECT 1750.670 159.415 1827.330 163.665 ;
      LAYER met4 ;
        RECT 1827.730 159.815 2024.270 163.265 ;
      LAYER met4 ;
        RECT 2024.670 159.415 2101.330 163.665 ;
      LAYER met4 ;
        RECT 2101.730 159.815 2298.270 163.265 ;
      LAYER met4 ;
        RECT 2298.670 159.415 2375.330 163.665 ;
      LAYER met4 ;
        RECT 2375.730 159.815 2572.270 163.265 ;
      LAYER met4 ;
        RECT 2572.670 159.415 2649.330 163.665 ;
      LAYER met4 ;
        RECT 2649.730 159.815 2846.270 163.265 ;
      LAYER met4 ;
        RECT 2846.670 159.415 2918.330 163.665 ;
      LAYER met4 ;
        RECT 2918.730 159.815 3115.270 163.265 ;
      LAYER met4 ;
        RECT 3115.670 159.415 3187.330 163.665 ;
      LAYER met4 ;
        RECT 3187.730 159.815 3385.270 163.265 ;
      LAYER met4 ;
        RECT 3385.670 159.415 3588.000 163.665 ;
        RECT 0.000 158.815 200.000 159.415 ;
        RECT 394.965 158.815 468.035 159.415 ;
        RECT 663.965 158.815 737.035 159.415 ;
        RECT 933.030 158.815 1011.035 159.415 ;
        RECT 1206.000 158.815 1280.035 159.415 ;
        RECT 1476.030 158.815 1554.035 159.415 ;
        RECT 1750.030 158.815 1828.035 159.415 ;
        RECT 2024.030 158.815 2102.035 159.415 ;
        RECT 2298.030 158.815 2376.035 159.415 ;
        RECT 2572.030 158.815 2650.035 159.415 ;
        RECT 2845.965 158.815 2919.035 159.415 ;
        RECT 3114.965 158.815 3188.035 159.415 ;
        RECT 3385.255 158.815 3588.000 159.415 ;
        RECT 0.000 153.365 198.125 158.815 ;
      LAYER met4 ;
        RECT 198.525 153.765 395.270 158.415 ;
      LAYER met4 ;
        RECT 395.670 153.365 467.330 158.815 ;
        RECT 664.670 158.770 736.330 158.815 ;
        RECT 664.745 153.410 736.330 158.770 ;
      LAYER met4 ;
        RECT 736.730 153.765 933.270 158.415 ;
      LAYER met4 ;
        RECT 664.670 153.365 736.330 153.410 ;
        RECT 933.670 153.365 1010.330 158.815 ;
      LAYER met4 ;
        RECT 1010.730 153.765 1207.270 158.415 ;
      LAYER met4 ;
        RECT 1207.670 153.365 1279.330 158.815 ;
      LAYER met4 ;
        RECT 1279.730 153.765 1476.270 158.415 ;
      LAYER met4 ;
        RECT 1476.670 153.365 1553.330 158.815 ;
      LAYER met4 ;
        RECT 1553.730 153.765 1750.270 158.415 ;
      LAYER met4 ;
        RECT 1750.670 153.365 1827.330 158.815 ;
      LAYER met4 ;
        RECT 1827.730 153.765 2024.270 158.415 ;
      LAYER met4 ;
        RECT 2024.670 153.365 2101.330 158.815 ;
      LAYER met4 ;
        RECT 2101.730 153.765 2298.270 158.415 ;
      LAYER met4 ;
        RECT 2298.670 153.365 2375.330 158.815 ;
      LAYER met4 ;
        RECT 2375.730 153.765 2572.270 158.415 ;
      LAYER met4 ;
        RECT 2572.670 153.365 2649.330 158.815 ;
      LAYER met4 ;
        RECT 2649.730 153.765 2846.270 158.415 ;
      LAYER met4 ;
        RECT 2846.670 153.365 2918.330 158.815 ;
      LAYER met4 ;
        RECT 2918.730 153.765 3115.270 158.415 ;
      LAYER met4 ;
        RECT 3115.670 153.365 3187.330 158.815 ;
      LAYER met4 ;
        RECT 3187.730 153.765 3385.270 158.415 ;
      LAYER met4 ;
        RECT 3385.670 153.365 3588.000 158.815 ;
        RECT 0.000 152.665 200.000 153.365 ;
        RECT 394.965 152.665 468.035 153.365 ;
        RECT 663.965 152.665 737.035 153.365 ;
        RECT 933.030 152.665 1011.035 153.365 ;
        RECT 1206.000 152.665 1280.035 153.365 ;
        RECT 1476.030 152.665 1554.035 153.365 ;
        RECT 1750.030 152.665 1828.035 153.365 ;
        RECT 2024.030 152.665 2102.035 153.365 ;
        RECT 2298.030 152.665 2376.035 153.365 ;
        RECT 2572.030 152.665 2650.035 153.365 ;
        RECT 2845.965 152.665 2919.035 153.365 ;
        RECT 3114.965 152.665 3188.035 153.365 ;
        RECT 3385.255 152.665 3588.000 153.365 ;
        RECT 0.000 152.035 180.025 152.665 ;
        RECT 0.000 148.755 178.665 152.035 ;
      LAYER met4 ;
        RECT 180.425 151.935 395.270 152.265 ;
      LAYER met4 ;
        RECT 395.670 152.035 467.330 152.665 ;
      LAYER met4 ;
        RECT 467.730 151.935 964.910 152.265 ;
      LAYER met4 ;
        RECT 965.310 152.035 1008.990 152.665 ;
      LAYER met4 ;
        RECT 1009.390 151.935 1507.910 152.265 ;
      LAYER met4 ;
        RECT 1508.310 152.035 1551.990 152.665 ;
      LAYER met4 ;
        RECT 1552.390 151.935 1781.910 152.265 ;
      LAYER met4 ;
        RECT 1782.310 152.035 1825.990 152.665 ;
      LAYER met4 ;
        RECT 1826.390 151.935 2055.910 152.265 ;
      LAYER met4 ;
        RECT 2056.310 152.035 2099.990 152.665 ;
      LAYER met4 ;
        RECT 2100.390 151.935 2329.910 152.265 ;
      LAYER met4 ;
        RECT 2330.310 152.035 2373.990 152.665 ;
      LAYER met4 ;
        RECT 2374.390 151.935 2603.910 152.265 ;
      LAYER met4 ;
        RECT 2604.310 152.035 2647.990 152.665 ;
      LAYER met4 ;
        RECT 2648.390 151.935 3407.575 152.265 ;
      LAYER met4 ;
        RECT 0.000 147.275 178.050 148.755 ;
      LAYER met4 ;
        RECT 179.065 148.655 957.535 151.635 ;
      LAYER met4 ;
        RECT 0.000 143.995 176.690 147.275 ;
      LAYER met4 ;
        RECT 178.450 147.175 200.000 148.355 ;
      LAYER met4 ;
        RECT 200.000 147.175 394.000 148.355 ;
      LAYER met4 ;
        RECT 394.000 147.175 395.270 148.355 ;
      LAYER met4 ;
        RECT 395.670 147.275 467.330 148.255 ;
      LAYER met4 ;
        RECT 467.730 147.175 469.000 148.355 ;
      LAYER met4 ;
        RECT 469.000 147.175 663.000 148.355 ;
      LAYER met4 ;
        RECT 663.000 147.175 664.270 148.355 ;
      LAYER met4 ;
        RECT 664.670 147.275 736.330 148.255 ;
      LAYER met4 ;
        RECT 736.730 147.175 738.000 148.355 ;
      LAYER met4 ;
        RECT 738.000 147.175 932.000 148.355 ;
      LAYER met4 ;
        RECT 932.000 147.175 933.270 148.355 ;
      LAYER met4 ;
        RECT 957.935 148.255 959.455 151.535 ;
      LAYER met4 ;
        RECT 959.855 148.655 1500.535 151.635 ;
      LAYER met4 ;
        RECT 933.670 147.275 1010.330 148.255 ;
        RECT 0.000 142.865 176.425 143.995 ;
      LAYER met4 ;
        RECT 177.090 143.895 973.240 146.875 ;
        RECT 176.825 143.265 395.270 143.595 ;
      LAYER met4 ;
        RECT 973.640 143.495 975.160 147.275 ;
      LAYER met4 ;
        RECT 1010.730 147.175 1012.000 148.355 ;
      LAYER met4 ;
        RECT 1012.000 147.175 1206.000 148.355 ;
      LAYER met4 ;
        RECT 1206.000 147.175 1207.270 148.355 ;
      LAYER met4 ;
        RECT 1207.670 147.275 1279.330 148.255 ;
      LAYER met4 ;
        RECT 1279.730 147.175 1281.000 148.355 ;
      LAYER met4 ;
        RECT 1281.000 147.175 1475.000 148.355 ;
      LAYER met4 ;
        RECT 1475.000 147.175 1476.270 148.355 ;
      LAYER met4 ;
        RECT 1500.935 148.255 1502.455 151.535 ;
      LAYER met4 ;
        RECT 1502.855 148.655 1774.535 151.635 ;
      LAYER met4 ;
        RECT 1476.670 147.275 1553.330 148.255 ;
      LAYER met4 ;
        RECT 975.560 143.895 1516.240 146.875 ;
      LAYER met4 ;
        RECT 395.670 142.865 467.330 143.495 ;
        RECT 965.310 142.865 1008.990 143.495 ;
      LAYER met4 ;
        RECT 1009.390 143.265 1507.910 143.595 ;
      LAYER met4 ;
        RECT 1516.640 143.495 1518.160 147.275 ;
      LAYER met4 ;
        RECT 1553.730 147.175 1555.000 148.355 ;
      LAYER met4 ;
        RECT 1555.000 147.175 1749.000 148.355 ;
      LAYER met4 ;
        RECT 1749.000 147.175 1750.270 148.355 ;
      LAYER met4 ;
        RECT 1774.935 148.255 1776.455 151.535 ;
      LAYER met4 ;
        RECT 1776.855 148.655 2048.535 151.635 ;
      LAYER met4 ;
        RECT 1750.670 147.275 1827.330 148.255 ;
      LAYER met4 ;
        RECT 1518.560 143.895 1790.240 146.875 ;
      LAYER met4 ;
        RECT 1508.310 142.865 1551.990 143.495 ;
      LAYER met4 ;
        RECT 1552.390 143.265 1781.910 143.595 ;
      LAYER met4 ;
        RECT 1790.640 143.495 1792.160 147.275 ;
      LAYER met4 ;
        RECT 1827.730 147.175 1829.000 148.355 ;
      LAYER met4 ;
        RECT 1829.000 147.175 2023.000 148.355 ;
      LAYER met4 ;
        RECT 2023.000 147.175 2024.270 148.355 ;
      LAYER met4 ;
        RECT 2048.935 148.255 2050.455 151.535 ;
      LAYER met4 ;
        RECT 2050.855 148.655 2322.535 151.635 ;
      LAYER met4 ;
        RECT 2024.670 147.275 2101.330 148.255 ;
      LAYER met4 ;
        RECT 1792.560 143.895 2064.240 146.875 ;
      LAYER met4 ;
        RECT 1782.310 142.865 1825.990 143.495 ;
      LAYER met4 ;
        RECT 1826.390 143.265 2055.910 143.595 ;
      LAYER met4 ;
        RECT 2064.640 143.495 2066.160 147.275 ;
      LAYER met4 ;
        RECT 2101.730 147.175 2103.000 148.355 ;
      LAYER met4 ;
        RECT 2103.000 147.175 2297.000 148.355 ;
      LAYER met4 ;
        RECT 2297.000 147.175 2298.270 148.355 ;
      LAYER met4 ;
        RECT 2322.935 148.255 2324.455 151.535 ;
      LAYER met4 ;
        RECT 2324.855 148.655 2596.535 151.635 ;
      LAYER met4 ;
        RECT 2298.670 147.275 2375.330 148.255 ;
      LAYER met4 ;
        RECT 2066.560 143.895 2338.240 146.875 ;
      LAYER met4 ;
        RECT 2056.310 142.865 2099.990 143.495 ;
      LAYER met4 ;
        RECT 2100.390 143.265 2329.910 143.595 ;
      LAYER met4 ;
        RECT 2338.640 143.495 2340.160 147.275 ;
      LAYER met4 ;
        RECT 2375.730 147.175 2377.000 148.355 ;
      LAYER met4 ;
        RECT 2377.000 147.175 2571.000 148.355 ;
      LAYER met4 ;
        RECT 2571.000 147.175 2572.270 148.355 ;
      LAYER met4 ;
        RECT 2596.935 148.255 2598.455 151.535 ;
      LAYER met4 ;
        RECT 2598.855 148.655 3404.875 151.635 ;
      LAYER met4 ;
        RECT 3407.975 151.535 3588.000 152.665 ;
        RECT 3405.275 148.755 3588.000 151.535 ;
        RECT 2572.670 147.275 2649.330 148.255 ;
      LAYER met4 ;
        RECT 2340.560 143.895 2612.240 146.875 ;
      LAYER met4 ;
        RECT 2330.310 142.865 2373.990 143.495 ;
      LAYER met4 ;
        RECT 2374.390 143.265 2603.910 143.595 ;
      LAYER met4 ;
        RECT 2612.640 143.495 2614.160 147.275 ;
      LAYER met4 ;
        RECT 2649.730 147.175 2651.000 148.355 ;
      LAYER met4 ;
        RECT 2651.000 147.175 2845.000 148.355 ;
      LAYER met4 ;
        RECT 2845.000 147.175 2846.270 148.355 ;
      LAYER met4 ;
        RECT 2846.670 147.275 2918.330 148.255 ;
      LAYER met4 ;
        RECT 2918.730 147.175 2920.000 148.355 ;
      LAYER met4 ;
        RECT 2920.000 147.175 3114.000 148.355 ;
      LAYER met4 ;
        RECT 3114.000 147.175 3115.270 148.355 ;
      LAYER met4 ;
        RECT 3115.670 147.275 3187.330 148.255 ;
      LAYER met4 ;
        RECT 3187.730 147.175 3189.000 148.355 ;
      LAYER met4 ;
        RECT 3189.000 147.175 3384.000 148.355 ;
      LAYER met4 ;
        RECT 3384.000 147.175 3405.555 148.355 ;
      LAYER met4 ;
        RECT 3405.955 147.275 3588.000 148.755 ;
      LAYER met4 ;
        RECT 2614.560 143.895 3410.910 146.875 ;
      LAYER met4 ;
        RECT 3411.310 143.995 3588.000 147.275 ;
        RECT 2604.310 142.865 2647.990 143.495 ;
      LAYER met4 ;
        RECT 2648.390 143.265 3411.175 143.595 ;
      LAYER met4 ;
        RECT 3411.575 142.865 3588.000 143.995 ;
        RECT 0.000 142.165 394.000 142.865 ;
        RECT 394.965 142.165 468.035 142.865 ;
        RECT 469.000 142.165 663.000 142.865 ;
        RECT 663.965 142.165 737.035 142.865 ;
        RECT 738.000 142.165 932.000 142.865 ;
        RECT 933.030 142.165 1011.035 142.865 ;
        RECT 1012.000 142.165 1280.035 142.865 ;
        RECT 1281.000 142.165 1475.000 142.865 ;
        RECT 1476.030 142.165 1554.035 142.865 ;
        RECT 1555.000 142.165 1749.000 142.865 ;
        RECT 1750.030 142.165 1828.035 142.865 ;
        RECT 1829.000 142.165 2023.000 142.865 ;
        RECT 2024.030 142.165 2102.035 142.865 ;
        RECT 2103.000 142.165 2297.000 142.865 ;
        RECT 2298.030 142.165 2376.035 142.865 ;
        RECT 2377.000 142.165 2571.000 142.865 ;
        RECT 2572.030 142.165 2650.035 142.865 ;
        RECT 2651.000 142.165 2845.000 142.865 ;
        RECT 2845.965 142.165 2919.035 142.865 ;
        RECT 2920.000 142.165 3114.000 142.865 ;
        RECT 3114.965 142.165 3188.035 142.865 ;
        RECT 3189.000 142.165 3384.000 142.865 ;
        RECT 3385.255 142.165 3588.000 142.865 ;
        RECT 0.000 136.915 197.975 142.165 ;
      LAYER met4 ;
        RECT 198.375 137.315 395.270 141.765 ;
      LAYER met4 ;
        RECT 395.670 136.915 467.330 142.165 ;
      LAYER met4 ;
        RECT 467.730 137.315 664.270 141.765 ;
      LAYER met4 ;
        RECT 664.670 136.915 736.330 142.165 ;
      LAYER met4 ;
        RECT 736.730 137.315 933.270 141.765 ;
      LAYER met4 ;
        RECT 933.670 136.915 1010.330 142.165 ;
      LAYER met4 ;
        RECT 1010.730 137.315 1207.270 141.765 ;
      LAYER met4 ;
        RECT 1207.670 136.915 1279.330 142.165 ;
      LAYER met4 ;
        RECT 1279.730 137.315 1476.270 141.765 ;
      LAYER met4 ;
        RECT 1476.670 136.915 1553.330 142.165 ;
      LAYER met4 ;
        RECT 1553.730 137.315 1750.270 141.765 ;
      LAYER met4 ;
        RECT 1750.670 136.915 1827.330 142.165 ;
      LAYER met4 ;
        RECT 1827.730 137.315 2024.270 141.765 ;
      LAYER met4 ;
        RECT 2024.670 136.915 2101.330 142.165 ;
      LAYER met4 ;
        RECT 2101.730 137.315 2298.270 141.765 ;
      LAYER met4 ;
        RECT 2298.670 136.915 2375.330 142.165 ;
      LAYER met4 ;
        RECT 2375.730 137.315 2572.270 141.765 ;
      LAYER met4 ;
        RECT 2572.670 136.915 2649.330 142.165 ;
      LAYER met4 ;
        RECT 2649.730 137.315 2846.270 141.765 ;
      LAYER met4 ;
        RECT 2846.670 136.915 2918.330 142.165 ;
      LAYER met4 ;
        RECT 2918.730 137.315 3115.270 141.765 ;
      LAYER met4 ;
        RECT 3115.670 136.915 3187.330 142.165 ;
      LAYER met4 ;
        RECT 3187.730 137.315 3385.270 141.765 ;
      LAYER met4 ;
        RECT 3385.670 136.915 3588.000 142.165 ;
        RECT 0.000 136.315 394.000 136.915 ;
        RECT 394.965 136.315 468.035 136.915 ;
        RECT 469.000 136.315 663.000 136.915 ;
        RECT 663.965 136.315 737.035 136.915 ;
        RECT 738.000 136.315 932.000 136.915 ;
        RECT 933.030 136.315 1011.035 136.915 ;
        RECT 1012.000 136.315 1280.035 136.915 ;
        RECT 1281.000 136.315 1475.000 136.915 ;
        RECT 1476.030 136.315 1554.035 136.915 ;
        RECT 1555.000 136.315 1749.000 136.915 ;
        RECT 1750.030 136.315 1828.035 136.915 ;
        RECT 1829.000 136.315 2023.000 136.915 ;
        RECT 2024.030 136.315 2102.035 136.915 ;
        RECT 2103.000 136.315 2297.000 136.915 ;
        RECT 2298.030 136.315 2376.035 136.915 ;
        RECT 2377.000 136.315 2571.000 136.915 ;
        RECT 2572.030 136.315 2650.035 136.915 ;
        RECT 2651.000 136.315 2845.000 136.915 ;
        RECT 2845.965 136.315 2919.035 136.915 ;
        RECT 2920.000 136.315 3114.000 136.915 ;
        RECT 3114.965 136.315 3188.035 136.915 ;
        RECT 3189.000 136.315 3384.000 136.915 ;
        RECT 3385.255 136.315 3588.000 136.915 ;
        RECT 0.000 131.065 198.120 136.315 ;
      LAYER met4 ;
        RECT 198.520 131.465 395.270 135.915 ;
      LAYER met4 ;
        RECT 395.670 131.065 467.330 136.315 ;
      LAYER met4 ;
        RECT 467.730 131.465 664.270 135.915 ;
      LAYER met4 ;
        RECT 664.670 131.065 736.330 136.315 ;
      LAYER met4 ;
        RECT 736.730 131.465 933.270 135.915 ;
      LAYER met4 ;
        RECT 933.670 131.065 1010.330 136.315 ;
      LAYER met4 ;
        RECT 1010.730 131.465 1207.270 135.915 ;
      LAYER met4 ;
        RECT 1207.670 131.065 1279.330 136.315 ;
      LAYER met4 ;
        RECT 1279.730 131.465 1476.270 135.915 ;
      LAYER met4 ;
        RECT 1476.670 131.065 1553.330 136.315 ;
      LAYER met4 ;
        RECT 1553.730 131.465 1750.270 135.915 ;
      LAYER met4 ;
        RECT 1750.670 131.065 1827.330 136.315 ;
      LAYER met4 ;
        RECT 1827.730 131.465 2024.270 135.915 ;
      LAYER met4 ;
        RECT 2024.670 131.065 2101.330 136.315 ;
      LAYER met4 ;
        RECT 2101.730 131.465 2298.270 135.915 ;
      LAYER met4 ;
        RECT 2298.670 131.065 2375.330 136.315 ;
      LAYER met4 ;
        RECT 2375.730 131.465 2572.270 135.915 ;
      LAYER met4 ;
        RECT 2572.670 131.065 2649.330 136.315 ;
      LAYER met4 ;
        RECT 2649.730 131.465 2846.270 135.915 ;
      LAYER met4 ;
        RECT 2846.670 131.065 2918.330 136.315 ;
      LAYER met4 ;
        RECT 2918.730 131.465 3115.270 135.915 ;
      LAYER met4 ;
        RECT 3115.670 131.065 3187.330 136.315 ;
      LAYER met4 ;
        RECT 3187.730 131.465 3385.270 135.915 ;
      LAYER met4 ;
        RECT 3385.670 131.065 3588.000 136.315 ;
        RECT 0.000 130.365 394.000 131.065 ;
        RECT 394.965 130.365 468.035 131.065 ;
        RECT 469.000 130.365 663.000 131.065 ;
        RECT 663.965 130.365 737.035 131.065 ;
        RECT 738.000 130.365 932.000 131.065 ;
        RECT 933.030 130.365 1011.035 131.065 ;
        RECT 1012.000 130.365 1280.035 131.065 ;
        RECT 1281.000 130.365 1475.000 131.065 ;
        RECT 1476.030 130.365 1554.035 131.065 ;
        RECT 1555.000 130.365 1749.000 131.065 ;
        RECT 1750.030 130.365 1828.035 131.065 ;
        RECT 1829.000 130.365 2023.000 131.065 ;
        RECT 2024.030 130.365 2102.035 131.065 ;
        RECT 2103.000 130.365 2297.000 131.065 ;
        RECT 2298.030 130.365 2376.035 131.065 ;
        RECT 2377.000 130.365 2571.000 131.065 ;
        RECT 2572.030 130.365 2650.035 131.065 ;
        RECT 2651.000 130.365 2845.000 131.065 ;
        RECT 2845.965 130.365 2919.035 131.065 ;
        RECT 2920.000 130.365 3114.000 131.065 ;
        RECT 3114.965 130.365 3188.035 131.065 ;
        RECT 3189.000 130.365 3384.000 131.065 ;
        RECT 3385.255 130.365 3588.000 131.065 ;
        RECT 0.000 104.600 196.955 130.365 ;
      LAYER met4 ;
        RECT 197.355 105.000 395.270 129.965 ;
      LAYER met4 ;
        RECT 395.670 104.600 467.330 130.365 ;
      LAYER met4 ;
        RECT 467.730 105.000 664.270 129.965 ;
      LAYER met4 ;
        RECT 664.670 104.600 736.330 130.365 ;
      LAYER met4 ;
        RECT 736.730 105.000 933.270 129.965 ;
      LAYER met4 ;
        RECT 933.670 104.600 1010.330 130.365 ;
      LAYER met4 ;
        RECT 1010.730 105.000 1207.270 129.965 ;
      LAYER met4 ;
        RECT 1207.670 104.600 1279.330 130.365 ;
      LAYER met4 ;
        RECT 1279.730 105.000 1476.270 129.965 ;
      LAYER met4 ;
        RECT 1476.670 104.600 1553.330 130.365 ;
      LAYER met4 ;
        RECT 1553.730 105.000 1750.270 129.965 ;
      LAYER met4 ;
        RECT 1750.670 104.600 1827.330 130.365 ;
      LAYER met4 ;
        RECT 1827.730 105.000 2024.270 129.965 ;
      LAYER met4 ;
        RECT 2024.670 104.600 2101.330 130.365 ;
      LAYER met4 ;
        RECT 2101.730 105.000 2298.270 129.965 ;
      LAYER met4 ;
        RECT 2298.670 104.600 2375.330 130.365 ;
      LAYER met4 ;
        RECT 2375.730 105.000 2572.270 129.965 ;
      LAYER met4 ;
        RECT 2572.670 104.600 2649.330 130.365 ;
      LAYER met4 ;
        RECT 2649.730 105.000 2846.270 129.965 ;
      LAYER met4 ;
        RECT 2846.670 104.600 2918.330 130.365 ;
      LAYER met4 ;
        RECT 2918.730 105.000 3115.270 129.965 ;
      LAYER met4 ;
        RECT 3115.670 104.600 3187.330 130.365 ;
      LAYER met4 ;
        RECT 3187.730 105.000 3385.855 129.965 ;
      LAYER met4 ;
        RECT 3386.255 104.600 3588.000 130.365 ;
        RECT 0.000 24.615 394.000 104.600 ;
        RECT 394.965 24.615 468.035 104.600 ;
        RECT 0.000 0.000 198.165 24.615 ;
      LAYER met4 ;
        RECT 198.565 0.000 200.000 24.215 ;
      LAYER met4 ;
        RECT 200.000 0.000 394.000 24.615 ;
      LAYER met4 ;
        RECT 394.000 0.000 395.270 24.215 ;
      LAYER met4 ;
        RECT 395.670 0.000 467.330 24.615 ;
      LAYER met4 ;
        RECT 467.730 0.000 469.000 24.215 ;
      LAYER met4 ;
        RECT 469.000 0.000 663.000 104.600 ;
        RECT 663.965 24.615 737.035 104.600 ;
      LAYER met4 ;
        RECT 663.000 0.000 664.270 24.215 ;
      LAYER met4 ;
        RECT 664.670 0.000 736.330 24.615 ;
      LAYER met4 ;
        RECT 736.730 0.000 738.000 24.215 ;
      LAYER met4 ;
        RECT 738.000 0.000 932.000 104.600 ;
        RECT 933.030 24.615 1011.035 104.600 ;
        RECT 1012.000 24.615 1280.035 104.600 ;
      LAYER met4 ;
        RECT 932.000 0.000 933.270 24.215 ;
      LAYER met4 ;
        RECT 933.670 0.000 1010.330 24.615 ;
      LAYER met4 ;
        RECT 1010.730 0.000 1012.000 24.215 ;
      LAYER met4 ;
        RECT 1012.000 0.000 1206.000 24.615 ;
      LAYER met4 ;
        RECT 1206.000 0.000 1207.270 24.215 ;
      LAYER met4 ;
        RECT 1207.670 0.000 1279.330 24.615 ;
      LAYER met4 ;
        RECT 1279.730 0.000 1281.000 24.215 ;
      LAYER met4 ;
        RECT 1281.000 0.000 1475.000 104.600 ;
        RECT 1476.030 24.615 1554.035 104.600 ;
      LAYER met4 ;
        RECT 1475.000 0.000 1476.270 24.215 ;
      LAYER met4 ;
        RECT 1476.670 0.000 1553.330 24.615 ;
      LAYER met4 ;
        RECT 1553.730 0.000 1555.000 24.215 ;
      LAYER met4 ;
        RECT 1555.000 0.000 1749.000 104.600 ;
        RECT 1750.030 24.615 1828.035 104.600 ;
      LAYER met4 ;
        RECT 1749.000 0.000 1750.270 24.215 ;
      LAYER met4 ;
        RECT 1750.670 0.000 1827.330 24.615 ;
      LAYER met4 ;
        RECT 1827.730 0.000 1829.000 24.215 ;
      LAYER met4 ;
        RECT 1829.000 0.000 2023.000 104.600 ;
        RECT 2024.030 24.615 2102.035 104.600 ;
      LAYER met4 ;
        RECT 2023.000 0.000 2024.270 24.215 ;
      LAYER met4 ;
        RECT 2024.670 0.000 2101.330 24.615 ;
      LAYER met4 ;
        RECT 2101.730 0.000 2103.000 24.215 ;
      LAYER met4 ;
        RECT 2103.000 0.000 2297.000 104.600 ;
        RECT 2298.030 24.615 2376.035 104.600 ;
      LAYER met4 ;
        RECT 2297.000 0.000 2298.270 24.215 ;
      LAYER met4 ;
        RECT 2298.670 0.000 2375.330 24.615 ;
      LAYER met4 ;
        RECT 2375.730 0.000 2377.000 24.215 ;
      LAYER met4 ;
        RECT 2377.000 0.000 2571.000 104.600 ;
        RECT 2572.030 24.615 2650.035 104.600 ;
      LAYER met4 ;
        RECT 2571.000 0.000 2572.270 24.215 ;
      LAYER met4 ;
        RECT 2572.670 0.000 2649.330 24.615 ;
      LAYER met4 ;
        RECT 2649.730 0.000 2651.000 24.215 ;
      LAYER met4 ;
        RECT 2651.000 0.000 2845.000 104.600 ;
        RECT 2845.965 24.615 2919.035 104.600 ;
      LAYER met4 ;
        RECT 2845.000 0.000 2846.270 24.215 ;
      LAYER met4 ;
        RECT 2846.670 0.000 2918.330 24.615 ;
      LAYER met4 ;
        RECT 2918.730 0.000 2920.000 24.215 ;
      LAYER met4 ;
        RECT 2920.000 0.000 3114.000 104.600 ;
        RECT 3114.965 24.615 3188.035 104.600 ;
      LAYER met4 ;
        RECT 3114.000 0.000 3115.270 24.215 ;
      LAYER met4 ;
        RECT 3115.670 0.000 3187.330 24.615 ;
      LAYER met4 ;
        RECT 3187.730 0.000 3189.000 24.215 ;
      LAYER met4 ;
        RECT 3189.000 0.000 3384.000 104.600 ;
        RECT 3385.255 24.615 3588.000 104.600 ;
      LAYER met4 ;
        RECT 3384.000 0.000 3385.270 24.215 ;
      LAYER met4 ;
        RECT 3385.670 0.000 3588.000 24.615 ;
      LAYER met5 ;
        RECT 0.000 5084.585 204.000 5188.000 ;
      LAYER met5 ;
        RECT 204.000 5163.785 381.000 5188.000 ;
      LAYER met5 ;
        RECT 381.000 5156.610 461.000 5188.000 ;
      LAYER met5 ;
        RECT 461.000 5163.785 638.000 5188.000 ;
      LAYER met5 ;
        RECT 381.000 5090.960 390.500 5156.610 ;
        RECT 456.400 5090.960 461.000 5156.610 ;
        RECT 381.000 5084.585 461.000 5090.960 ;
        RECT 638.000 5156.610 718.000 5188.000 ;
      LAYER met5 ;
        RECT 718.000 5163.785 895.000 5188.000 ;
      LAYER met5 ;
        RECT 638.000 5090.960 647.500 5156.610 ;
        RECT 713.400 5090.960 718.000 5156.610 ;
        RECT 638.000 5084.585 718.000 5090.960 ;
        RECT 895.000 5156.610 975.000 5188.000 ;
      LAYER met5 ;
        RECT 975.000 5163.785 1152.000 5188.000 ;
      LAYER met5 ;
        RECT 895.000 5090.960 904.500 5156.610 ;
        RECT 970.400 5090.960 975.000 5156.610 ;
        RECT 895.000 5084.585 975.000 5090.960 ;
        RECT 1152.000 5156.610 1232.000 5188.000 ;
      LAYER met5 ;
        RECT 1232.000 5163.785 1410.000 5188.000 ;
      LAYER met5 ;
        RECT 1152.000 5090.960 1161.500 5156.610 ;
        RECT 1227.400 5090.960 1232.000 5156.610 ;
        RECT 1152.000 5084.585 1232.000 5090.960 ;
        RECT 1410.000 5156.610 1490.000 5188.000 ;
      LAYER met5 ;
        RECT 1490.000 5163.785 1667.000 5188.000 ;
      LAYER met5 ;
        RECT 1410.000 5090.960 1419.500 5156.610 ;
        RECT 1485.400 5090.960 1490.000 5156.610 ;
        RECT 1410.000 5084.585 1490.000 5090.960 ;
        RECT 1667.000 5155.545 1742.000 5188.000 ;
      LAYER met5 ;
        RECT 1742.000 5163.785 1919.000 5188.000 ;
      LAYER met5 ;
        RECT 1667.000 5091.520 1672.450 5155.545 ;
        RECT 1736.490 5091.520 1742.000 5155.545 ;
        RECT 1667.000 5084.585 1742.000 5091.520 ;
        RECT 1919.000 5156.610 1999.000 5188.000 ;
      LAYER met5 ;
        RECT 1999.000 5163.785 2364.000 5188.000 ;
      LAYER met5 ;
        RECT 1919.000 5090.960 1928.500 5156.610 ;
        RECT 1994.400 5090.960 1999.000 5156.610 ;
        RECT 1919.000 5084.585 1999.000 5090.960 ;
        RECT 2364.000 5156.610 2444.000 5188.000 ;
      LAYER met5 ;
        RECT 2444.000 5163.785 2621.000 5188.000 ;
      LAYER met5 ;
        RECT 2364.000 5090.960 2373.500 5156.610 ;
        RECT 2439.400 5090.960 2444.000 5156.610 ;
        RECT 2364.000 5084.585 2444.000 5090.960 ;
        RECT 2621.000 5156.610 2701.000 5188.000 ;
      LAYER met5 ;
        RECT 2701.000 5163.785 2878.000 5188.000 ;
      LAYER met5 ;
        RECT 2621.000 5090.960 2630.500 5156.610 ;
        RECT 2696.400 5090.960 2701.000 5156.610 ;
        RECT 2621.000 5084.585 2701.000 5090.960 ;
        RECT 2878.000 5155.545 2953.000 5188.000 ;
      LAYER met5 ;
        RECT 2953.000 5163.785 3130.000 5188.000 ;
      LAYER met5 ;
        RECT 2878.000 5091.520 2883.450 5155.545 ;
        RECT 2947.490 5091.520 2953.000 5155.545 ;
        RECT 2878.000 5084.585 2953.000 5091.520 ;
        RECT 3130.000 5156.610 3210.000 5188.000 ;
      LAYER met5 ;
        RECT 3210.000 5163.785 3388.000 5188.000 ;
      LAYER met5 ;
        RECT 3130.000 5090.960 3139.500 5156.610 ;
        RECT 3205.400 5090.960 3210.000 5156.610 ;
        RECT 3130.000 5084.585 3210.000 5090.960 ;
        RECT 3388.000 5084.585 3588.000 5188.000 ;
        RECT 0.000 5056.435 200.545 5084.585 ;
      LAYER met5 ;
        RECT 202.145 5058.035 382.270 5082.985 ;
      LAYER met5 ;
        RECT 0.000 5046.335 201.130 5056.435 ;
      LAYER met5 ;
        RECT 202.730 5052.185 382.270 5056.435 ;
        RECT 202.730 5046.335 382.270 5050.585 ;
      LAYER met5 ;
        RECT 0.000 5034.135 175.245 5046.335 ;
      LAYER met5 ;
        RECT 176.845 5035.735 382.270 5044.735 ;
      LAYER met5 ;
        RECT 0.000 5012.755 201.130 5034.135 ;
      LAYER met5 ;
        RECT 202.730 5029.685 382.270 5034.135 ;
        RECT 202.730 5024.840 382.270 5028.085 ;
        RECT 204.000 5024.835 381.000 5024.840 ;
        RECT 202.730 5019.985 382.270 5023.235 ;
        RECT 202.730 5013.935 382.270 5018.385 ;
      LAYER met5 ;
        RECT 0.000 4992.245 141.665 5012.755 ;
        RECT 0.000 4988.000 103.415 4992.245 ;
        RECT 131.565 4991.225 141.665 4992.245 ;
        RECT 131.565 4991.080 135.815 4991.225 ;
      LAYER met5 ;
        RECT 0.000 4851.000 24.215 4988.000 ;
      LAYER met5 ;
        RECT 0.000 4848.130 103.415 4851.000 ;
      LAYER met5 ;
        RECT 105.015 4849.730 129.965 4990.645 ;
        RECT 131.565 4849.730 135.815 4989.480 ;
        RECT 137.415 4849.730 141.665 4989.625 ;
        RECT 143.265 4849.730 152.265 5011.155 ;
      LAYER met5 ;
        RECT 153.865 5006.285 201.130 5012.755 ;
      LAYER met5 ;
        RECT 202.730 5007.885 382.270 5012.335 ;
      LAYER met5 ;
        RECT 383.870 5006.285 458.130 5084.585 ;
      LAYER met5 ;
        RECT 459.730 5058.035 639.270 5082.985 ;
        RECT 459.730 5052.185 639.270 5056.435 ;
        RECT 459.730 5046.335 639.270 5050.585 ;
        RECT 459.730 5035.735 639.270 5044.735 ;
        RECT 459.730 5029.685 639.270 5034.135 ;
        RECT 459.730 5024.840 639.270 5028.085 ;
        RECT 461.000 5024.835 638.000 5024.840 ;
        RECT 459.730 5019.985 639.270 5023.235 ;
        RECT 459.730 5013.935 639.270 5018.385 ;
        RECT 459.730 5007.885 639.270 5012.335 ;
      LAYER met5 ;
        RECT 640.870 5006.285 715.130 5084.585 ;
      LAYER met5 ;
        RECT 716.730 5058.035 896.270 5082.985 ;
        RECT 716.730 5052.185 896.270 5056.435 ;
        RECT 716.730 5046.335 896.270 5050.585 ;
        RECT 716.730 5035.735 896.270 5044.735 ;
        RECT 716.730 5029.685 896.270 5034.135 ;
        RECT 716.730 5024.840 896.270 5028.085 ;
        RECT 718.000 5024.835 895.000 5024.840 ;
        RECT 716.730 5019.985 896.270 5023.235 ;
        RECT 716.730 5013.935 896.270 5018.385 ;
        RECT 716.730 5007.885 896.270 5012.335 ;
      LAYER met5 ;
        RECT 897.870 5006.285 972.130 5084.585 ;
      LAYER met5 ;
        RECT 973.730 5058.035 1153.270 5082.985 ;
        RECT 973.730 5052.185 1153.270 5056.435 ;
        RECT 973.730 5046.335 1153.270 5050.585 ;
        RECT 973.730 5035.735 1153.270 5044.735 ;
        RECT 973.730 5029.685 1153.270 5034.135 ;
        RECT 973.730 5024.840 1153.270 5028.085 ;
        RECT 975.000 5024.835 1152.000 5024.840 ;
        RECT 973.730 5019.985 1153.270 5023.235 ;
        RECT 973.730 5013.935 1153.270 5018.385 ;
        RECT 973.730 5007.885 1153.270 5012.335 ;
      LAYER met5 ;
        RECT 1154.870 5006.285 1229.130 5084.585 ;
      LAYER met5 ;
        RECT 1230.730 5058.035 1411.270 5082.985 ;
        RECT 1230.730 5052.185 1411.270 5056.435 ;
        RECT 1230.730 5046.335 1411.270 5050.585 ;
        RECT 1230.730 5035.735 1411.270 5044.735 ;
        RECT 1230.730 5029.685 1411.270 5034.135 ;
        RECT 1230.730 5024.840 1411.270 5028.085 ;
        RECT 1232.000 5024.835 1410.000 5024.840 ;
        RECT 1230.730 5019.985 1411.270 5023.235 ;
        RECT 1230.730 5013.935 1411.270 5018.385 ;
        RECT 1230.730 5007.885 1411.270 5012.335 ;
      LAYER met5 ;
        RECT 1412.870 5006.285 1487.130 5084.585 ;
      LAYER met5 ;
        RECT 1488.730 5058.035 1668.270 5082.985 ;
        RECT 1488.730 5052.185 1668.270 5056.435 ;
        RECT 1488.730 5046.335 1668.270 5050.585 ;
        RECT 1488.730 5035.735 1668.270 5044.735 ;
        RECT 1488.730 5029.685 1668.270 5034.135 ;
        RECT 1488.730 5024.840 1668.270 5028.085 ;
      LAYER met5 ;
        RECT 1669.870 5024.840 1739.130 5084.585 ;
      LAYER met5 ;
        RECT 1740.730 5058.035 1920.270 5082.985 ;
        RECT 1740.730 5052.185 1920.270 5056.435 ;
        RECT 1740.730 5046.335 1920.270 5050.585 ;
        RECT 1740.730 5035.735 1742.000 5044.735 ;
        RECT 1747.000 5035.735 1920.270 5044.735 ;
        RECT 1740.730 5029.685 1747.000 5034.135 ;
        RECT 1752.000 5029.685 1920.270 5034.135 ;
        RECT 1740.730 5024.840 1742.000 5028.085 ;
        RECT 1490.000 5024.835 1667.000 5024.840 ;
      LAYER met5 ;
        RECT 1667.000 5024.835 1742.000 5024.840 ;
      LAYER met5 ;
        RECT 1747.000 5024.840 1920.270 5028.085 ;
        RECT 1747.000 5024.835 1919.000 5024.840 ;
        RECT 1488.730 5019.985 1668.270 5023.235 ;
        RECT 1488.730 5013.935 1668.270 5018.385 ;
        RECT 1488.730 5007.885 1668.270 5012.335 ;
      LAYER met5 ;
        RECT 1669.870 5006.285 1739.130 5024.835 ;
      LAYER met5 ;
        RECT 1740.730 5019.985 1920.270 5023.235 ;
        RECT 1740.730 5013.935 1920.270 5018.385 ;
        RECT 1740.730 5007.885 1920.270 5012.335 ;
      LAYER met5 ;
        RECT 1921.870 5006.285 1996.130 5084.585 ;
      LAYER met5 ;
        RECT 1997.730 5058.035 2365.270 5082.985 ;
        RECT 1997.730 5052.185 2365.270 5056.435 ;
        RECT 1997.730 5046.335 2365.270 5050.585 ;
        RECT 1997.730 5035.735 2365.270 5044.735 ;
        RECT 1997.730 5029.685 2365.270 5034.135 ;
        RECT 1997.730 5024.840 2365.270 5028.085 ;
        RECT 1999.000 5024.835 2364.000 5024.840 ;
        RECT 1997.730 5019.985 2365.270 5023.235 ;
        RECT 1997.730 5013.935 2365.270 5018.385 ;
        RECT 1997.730 5007.885 2365.270 5012.335 ;
      LAYER met5 ;
        RECT 2366.870 5006.285 2441.130 5084.585 ;
      LAYER met5 ;
        RECT 2442.730 5058.035 2622.270 5082.985 ;
        RECT 2442.730 5052.185 2622.270 5056.435 ;
        RECT 2442.730 5046.335 2622.270 5050.585 ;
        RECT 2442.730 5035.735 2622.270 5044.735 ;
        RECT 2442.730 5029.685 2622.270 5034.135 ;
        RECT 2442.730 5024.840 2622.270 5028.085 ;
        RECT 2444.000 5024.835 2621.000 5024.840 ;
        RECT 2442.730 5019.985 2622.270 5023.235 ;
        RECT 2442.730 5013.935 2622.270 5018.385 ;
        RECT 2442.730 5007.885 2622.270 5012.335 ;
      LAYER met5 ;
        RECT 2623.870 5006.285 2698.130 5084.585 ;
      LAYER met5 ;
        RECT 2699.730 5058.035 2879.270 5082.985 ;
        RECT 2699.730 5052.185 2879.270 5056.435 ;
        RECT 2699.730 5046.335 2879.270 5050.585 ;
        RECT 2699.730 5035.735 2879.270 5044.735 ;
        RECT 2699.730 5029.685 2879.270 5034.135 ;
        RECT 2699.730 5024.840 2879.270 5028.085 ;
      LAYER met5 ;
        RECT 2880.870 5024.840 2950.130 5084.585 ;
      LAYER met5 ;
        RECT 2951.730 5058.035 3131.270 5082.985 ;
        RECT 2951.730 5052.185 3131.270 5056.435 ;
        RECT 2951.730 5046.335 3131.270 5050.585 ;
        RECT 2951.730 5035.735 3131.270 5044.735 ;
        RECT 2951.730 5029.685 3131.270 5034.135 ;
        RECT 2951.730 5024.840 3131.270 5028.085 ;
        RECT 2701.000 5024.835 2878.000 5024.840 ;
      LAYER met5 ;
        RECT 2878.000 5024.835 2953.000 5024.840 ;
      LAYER met5 ;
        RECT 2953.000 5024.835 3130.000 5024.840 ;
        RECT 2699.730 5019.985 2879.270 5023.235 ;
        RECT 2699.730 5013.935 2879.270 5018.385 ;
        RECT 2699.730 5007.885 2879.270 5012.335 ;
      LAYER met5 ;
        RECT 2880.870 5006.285 2950.130 5024.835 ;
      LAYER met5 ;
        RECT 2951.730 5019.985 3131.270 5023.235 ;
        RECT 2951.730 5013.935 3131.270 5018.385 ;
        RECT 2951.730 5007.885 3131.270 5012.335 ;
      LAYER met5 ;
        RECT 3132.870 5006.285 3207.130 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5058.035 3390.645 5082.985 ;
      LAYER met5 ;
        RECT 3392.245 5056.435 3588.000 5084.585 ;
      LAYER met5 ;
        RECT 3208.730 5052.185 3389.480 5056.435 ;
      LAYER met5 ;
        RECT 3391.080 5052.185 3588.000 5056.435 ;
      LAYER met5 ;
        RECT 3208.730 5046.335 3389.625 5050.585 ;
      LAYER met5 ;
        RECT 3391.225 5046.335 3588.000 5052.185 ;
      LAYER met5 ;
        RECT 3208.730 5035.735 3411.155 5044.735 ;
      LAYER met5 ;
        RECT 3412.755 5034.135 3588.000 5046.335 ;
      LAYER met5 ;
        RECT 3208.730 5029.685 3389.475 5034.135 ;
      LAYER met5 ;
        RECT 3391.075 5028.085 3588.000 5034.135 ;
      LAYER met5 ;
        RECT 3208.730 5024.840 3389.335 5028.085 ;
        RECT 3210.000 5024.835 3389.335 5024.840 ;
      LAYER met5 ;
        RECT 3390.935 5024.835 3588.000 5028.085 ;
      LAYER met5 ;
        RECT 3208.730 5019.985 3389.385 5023.235 ;
      LAYER met5 ;
        RECT 3390.985 5019.985 3588.000 5024.835 ;
      LAYER met5 ;
        RECT 3208.730 5013.935 3389.600 5018.385 ;
      LAYER met5 ;
        RECT 3391.200 5012.755 3588.000 5019.985 ;
        RECT 3391.200 5012.335 3434.135 5012.755 ;
      LAYER met5 ;
        RECT 3208.730 5007.885 3389.525 5012.335 ;
      LAYER met5 ;
        RECT 3391.125 5006.285 3434.135 5012.335 ;
        RECT 153.865 5003.035 201.145 5006.285 ;
      LAYER met5 ;
        RECT 202.745 5003.035 381.965 5006.285 ;
      LAYER met5 ;
        RECT 383.565 5003.035 458.370 5006.285 ;
      LAYER met5 ;
        RECT 459.970 5003.035 638.965 5006.285 ;
      LAYER met5 ;
        RECT 640.565 5003.035 715.370 5006.285 ;
      LAYER met5 ;
        RECT 716.970 5003.035 895.965 5006.285 ;
      LAYER met5 ;
        RECT 897.565 5003.035 972.370 5006.285 ;
      LAYER met5 ;
        RECT 973.970 5003.035 1152.965 5006.285 ;
      LAYER met5 ;
        RECT 1154.565 5003.035 1229.370 5006.285 ;
      LAYER met5 ;
        RECT 1230.970 5003.035 1410.965 5006.285 ;
      LAYER met5 ;
        RECT 1412.565 5003.035 1487.370 5006.285 ;
      LAYER met5 ;
        RECT 1488.970 5003.035 1667.965 5006.285 ;
      LAYER met5 ;
        RECT 1669.565 5003.035 1739.435 5006.285 ;
      LAYER met5 ;
        RECT 1741.035 5003.035 1742.000 5006.285 ;
        RECT 1747.000 5003.035 1919.965 5006.285 ;
      LAYER met5 ;
        RECT 1921.565 5003.035 1996.370 5006.285 ;
      LAYER met5 ;
        RECT 1997.970 5003.035 2364.965 5006.285 ;
      LAYER met5 ;
        RECT 2366.565 5003.035 2441.370 5006.285 ;
      LAYER met5 ;
        RECT 2442.970 5003.035 2621.965 5006.285 ;
      LAYER met5 ;
        RECT 2623.565 5003.035 2698.370 5006.285 ;
      LAYER met5 ;
        RECT 2699.970 5003.035 2878.965 5006.285 ;
      LAYER met5 ;
        RECT 2880.565 5003.035 2950.435 5006.285 ;
      LAYER met5 ;
        RECT 2952.035 5003.035 3130.965 5006.285 ;
      LAYER met5 ;
        RECT 3132.565 5003.035 3207.370 5006.285 ;
      LAYER met5 ;
        RECT 3208.970 5003.035 3389.470 5006.285 ;
      LAYER met5 ;
        RECT 3391.070 5003.035 3434.135 5006.285 ;
        RECT 153.865 4993.385 201.130 5003.035 ;
      LAYER met5 ;
        RECT 202.730 4996.985 382.270 5001.435 ;
      LAYER met5 ;
        RECT 153.865 4991.200 184.965 4993.385 ;
        RECT 192.615 4991.950 201.130 4993.385 ;
        RECT 153.865 4991.075 168.015 4991.200 ;
        RECT 175.665 4991.125 184.965 4991.200 ;
        RECT 159.915 4990.985 168.015 4991.075 ;
        RECT 181.715 4991.070 184.965 4991.125 ;
        RECT 159.915 4990.935 163.165 4990.985 ;
      LAYER met5 ;
        RECT 153.865 4849.730 158.315 4989.475 ;
        RECT 159.915 4851.000 163.165 4989.335 ;
        RECT 159.915 4849.730 163.160 4851.000 ;
        RECT 164.765 4849.730 168.015 4989.385 ;
        RECT 169.615 4849.730 174.065 4989.600 ;
        RECT 175.665 4849.730 180.115 4989.525 ;
        RECT 181.715 4849.970 184.965 4989.470 ;
        RECT 186.565 4849.730 191.015 4991.785 ;
        RECT 192.615 4849.730 197.865 4990.350 ;
      LAYER met5 ;
        RECT 199.465 4988.535 201.130 4991.950 ;
      LAYER met5 ;
        RECT 202.730 4990.135 382.270 4995.385 ;
      LAYER met5 ;
        RECT 383.870 4990.135 458.130 5003.035 ;
      LAYER met5 ;
        RECT 459.730 4996.985 639.270 5001.435 ;
        RECT 459.730 4990.135 639.270 4995.385 ;
      LAYER met5 ;
        RECT 640.870 4990.135 715.130 5003.035 ;
      LAYER met5 ;
        RECT 716.730 4996.985 896.270 5001.435 ;
        RECT 716.730 4990.135 896.270 4995.385 ;
      LAYER met5 ;
        RECT 897.870 4990.135 972.130 5003.035 ;
      LAYER met5 ;
        RECT 973.730 4996.985 1153.270 5001.435 ;
        RECT 973.730 4990.135 1153.270 4995.385 ;
      LAYER met5 ;
        RECT 1154.870 4990.135 1229.130 5003.035 ;
      LAYER met5 ;
        RECT 1230.730 4996.985 1411.270 5001.435 ;
        RECT 1230.730 4990.135 1411.270 4995.385 ;
      LAYER met5 ;
        RECT 1412.870 4990.135 1487.130 5003.035 ;
      LAYER met5 ;
        RECT 1488.730 4996.985 1668.270 5001.435 ;
        RECT 1488.730 4990.135 1668.270 4995.385 ;
      LAYER met5 ;
        RECT 1669.870 4990.135 1739.130 5003.035 ;
      LAYER met5 ;
        RECT 1740.730 4996.985 1747.000 5001.435 ;
        RECT 1752.000 4996.985 1920.270 5001.435 ;
        RECT 1740.730 4990.135 1920.270 4995.385 ;
      LAYER met5 ;
        RECT 1921.870 4990.135 1996.130 5003.035 ;
      LAYER met5 ;
        RECT 1997.730 4996.985 2365.270 5001.435 ;
        RECT 1997.730 4990.135 2365.270 4995.385 ;
      LAYER met5 ;
        RECT 2366.870 4990.135 2441.130 5003.035 ;
      LAYER met5 ;
        RECT 2442.730 4996.985 2622.270 5001.435 ;
        RECT 2442.730 4990.135 2622.270 4995.385 ;
      LAYER met5 ;
        RECT 2623.870 4990.135 2698.130 5003.035 ;
      LAYER met5 ;
        RECT 2699.730 4996.985 2879.270 5001.435 ;
        RECT 2699.730 4990.135 2879.270 4995.385 ;
      LAYER met5 ;
        RECT 2880.870 4990.135 2950.130 5003.035 ;
      LAYER met5 ;
        RECT 2951.730 4996.985 3131.270 5001.435 ;
        RECT 2951.730 4990.135 3131.270 4995.385 ;
      LAYER met5 ;
        RECT 3132.870 4990.135 3207.130 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4996.985 3391.785 5001.435 ;
      LAYER met5 ;
        RECT 3393.385 4995.385 3434.135 5003.035 ;
      LAYER met5 ;
        RECT 3208.730 4990.135 3390.350 4995.385 ;
      LAYER met5 ;
        RECT 3391.950 4988.535 3434.135 4995.385 ;
        RECT 199.465 4988.000 204.000 4988.535 ;
        RECT 3388.000 4986.870 3434.135 4988.535 ;
        RECT 3388.000 4984.000 3388.535 4986.870 ;
        RECT 3403.035 4986.855 3406.285 4986.870 ;
        RECT 181.715 4848.130 184.965 4848.370 ;
        RECT 0.000 4846.400 197.865 4848.130 ;
        RECT 0.000 4780.500 31.390 4846.400 ;
        RECT 97.040 4780.500 197.865 4846.400 ;
      LAYER met5 ;
        RECT 3390.135 4836.730 3395.385 4985.270 ;
        RECT 3396.985 4836.730 3401.435 4985.270 ;
        RECT 3403.035 4837.035 3406.285 4985.255 ;
        RECT 3407.885 4836.730 3412.335 4985.270 ;
        RECT 3413.935 4836.730 3418.385 4985.270 ;
        RECT 3419.985 4836.730 3423.235 4985.270 ;
        RECT 3424.840 4984.000 3428.085 4985.270 ;
        RECT 3424.835 4838.000 3428.085 4984.000 ;
        RECT 3424.840 4836.730 3428.085 4838.000 ;
        RECT 3429.685 4836.730 3434.135 4985.270 ;
        RECT 3435.735 4836.730 3444.735 5011.155 ;
      LAYER met5 ;
        RECT 3446.335 4987.455 3588.000 5012.755 ;
        RECT 3446.335 4986.870 3456.435 4987.455 ;
      LAYER met5 ;
        RECT 3446.335 4836.730 3450.585 4985.270 ;
        RECT 3452.185 4836.730 3456.435 4985.270 ;
        RECT 3458.035 4836.730 3482.985 4985.855 ;
      LAYER met5 ;
        RECT 3484.585 4984.000 3588.000 4987.455 ;
      LAYER met5 ;
        RECT 3563.785 4838.000 3588.000 4984.000 ;
      LAYER met5 ;
        RECT 3403.035 4835.130 3406.285 4835.435 ;
        RECT 3484.585 4835.130 3588.000 4838.000 ;
        RECT 0.000 4773.870 197.865 4780.500 ;
        RECT 3390.135 4828.500 3588.000 4835.130 ;
        RECT 0.000 4771.000 103.415 4773.870 ;
        RECT 181.715 4773.565 184.965 4773.870 ;
      LAYER met5 ;
        RECT 0.000 4635.000 24.215 4771.000 ;
      LAYER met5 ;
        RECT 0.000 4632.130 103.415 4635.000 ;
      LAYER met5 ;
        RECT 105.015 4633.730 129.965 4772.270 ;
        RECT 131.565 4633.730 135.815 4772.270 ;
        RECT 137.415 4633.730 141.665 4772.270 ;
        RECT 143.265 4633.730 152.265 4772.270 ;
        RECT 153.865 4633.730 158.315 4772.270 ;
        RECT 159.915 4771.000 163.160 4772.270 ;
        RECT 159.915 4635.000 163.165 4771.000 ;
        RECT 159.915 4633.730 163.160 4635.000 ;
        RECT 164.765 4633.730 168.015 4772.270 ;
        RECT 169.615 4633.730 174.065 4772.270 ;
        RECT 175.665 4633.730 180.115 4772.270 ;
        RECT 181.715 4634.035 184.965 4771.965 ;
        RECT 186.565 4633.730 191.015 4772.270 ;
        RECT 192.615 4633.730 197.865 4772.270 ;
      LAYER met5 ;
        RECT 3390.135 4762.600 3490.960 4828.500 ;
        RECT 3556.610 4762.600 3588.000 4828.500 ;
        RECT 3390.135 4760.870 3588.000 4762.600 ;
        RECT 3403.035 4760.630 3406.285 4760.870 ;
        RECT 181.715 4632.130 184.965 4632.435 ;
        RECT 0.000 4626.270 197.865 4632.130 ;
        RECT 0.000 4568.670 29.235 4626.270 ;
        RECT 99.700 4568.670 197.865 4626.270 ;
      LAYER met5 ;
        RECT 3390.135 4611.730 3395.385 4759.270 ;
        RECT 3396.985 4611.730 3401.435 4759.270 ;
        RECT 3403.035 4612.035 3406.285 4759.030 ;
        RECT 3407.885 4611.730 3412.335 4759.270 ;
        RECT 3413.935 4611.730 3418.385 4759.270 ;
        RECT 3419.985 4611.730 3423.235 4759.270 ;
        RECT 3424.840 4758.000 3428.085 4759.270 ;
        RECT 3424.835 4613.000 3428.085 4758.000 ;
        RECT 3424.840 4611.730 3428.085 4613.000 ;
        RECT 3429.685 4611.730 3434.135 4759.270 ;
        RECT 3435.735 4611.730 3444.735 4759.270 ;
        RECT 3446.335 4611.730 3450.585 4759.270 ;
        RECT 3452.185 4611.730 3456.435 4759.270 ;
        RECT 3458.035 4611.730 3482.985 4759.270 ;
      LAYER met5 ;
        RECT 3484.585 4758.000 3588.000 4760.870 ;
      LAYER met5 ;
        RECT 3563.785 4613.000 3588.000 4758.000 ;
      LAYER met5 ;
        RECT 3403.035 4610.130 3406.285 4610.435 ;
        RECT 3484.585 4610.130 3588.000 4613.000 ;
        RECT 0.000 4562.870 197.865 4568.670 ;
        RECT 3390.135 4604.330 3588.000 4610.130 ;
        RECT 0.000 4560.000 103.415 4562.870 ;
        RECT 181.715 4562.565 184.965 4562.870 ;
      LAYER met5 ;
        RECT 0.000 4424.000 24.215 4560.000 ;
      LAYER met5 ;
        RECT 0.000 4421.130 103.415 4424.000 ;
      LAYER met5 ;
        RECT 105.015 4422.730 129.965 4561.270 ;
        RECT 131.565 4422.730 135.815 4561.270 ;
        RECT 137.415 4422.730 141.665 4561.270 ;
        RECT 143.265 4422.730 152.265 4561.270 ;
        RECT 153.865 4422.730 158.315 4561.270 ;
        RECT 159.915 4560.000 163.160 4561.270 ;
        RECT 159.915 4424.000 163.165 4560.000 ;
        RECT 159.915 4422.730 163.160 4424.000 ;
      LAYER met5 ;
        RECT 163.160 4421.130 163.165 4424.000 ;
      LAYER met5 ;
        RECT 164.765 4422.730 168.015 4561.270 ;
        RECT 169.615 4422.730 174.065 4561.270 ;
        RECT 175.665 4422.730 180.115 4561.270 ;
        RECT 181.715 4423.035 184.965 4560.965 ;
        RECT 186.565 4422.730 191.015 4561.270 ;
        RECT 192.615 4422.730 197.865 4561.270 ;
      LAYER met5 ;
        RECT 3390.135 4546.730 3488.300 4604.330 ;
        RECT 3558.765 4546.730 3588.000 4604.330 ;
        RECT 3390.135 4540.870 3588.000 4546.730 ;
        RECT 3403.035 4540.565 3406.285 4540.870 ;
        RECT 181.715 4421.130 184.965 4421.435 ;
        RECT 0.000 4418.490 197.865 4421.130 ;
        RECT 0.000 4354.450 32.455 4418.490 ;
        RECT 96.480 4354.450 197.865 4418.490 ;
      LAYER met5 ;
        RECT 3390.135 4390.730 3395.385 4539.270 ;
        RECT 3396.985 4390.730 3401.435 4539.270 ;
        RECT 3403.035 4391.035 3406.285 4538.965 ;
        RECT 3407.885 4390.730 3412.335 4539.270 ;
        RECT 3413.935 4390.730 3418.385 4539.270 ;
        RECT 3419.985 4390.730 3423.235 4539.270 ;
        RECT 3424.840 4538.000 3428.085 4539.270 ;
        RECT 3424.835 4392.000 3428.085 4538.000 ;
        RECT 3424.840 4390.730 3428.085 4392.000 ;
        RECT 3429.685 4390.730 3434.135 4539.270 ;
        RECT 3435.735 4390.730 3444.735 4539.270 ;
        RECT 3446.335 4390.730 3450.585 4539.270 ;
        RECT 3452.185 4390.730 3456.435 4539.270 ;
        RECT 3458.035 4390.730 3482.985 4539.270 ;
      LAYER met5 ;
        RECT 3484.585 4538.000 3588.000 4540.870 ;
      LAYER met5 ;
        RECT 3563.785 4392.000 3588.000 4538.000 ;
      LAYER met5 ;
        RECT 3403.035 4389.130 3406.285 4389.435 ;
        RECT 3484.585 4389.130 3588.000 4392.000 ;
        RECT 0.000 4351.870 197.865 4354.450 ;
        RECT 3390.135 4382.500 3588.000 4389.130 ;
        RECT 0.000 4349.000 103.415 4351.870 ;
      LAYER met5 ;
        RECT 0.000 4213.000 24.215 4349.000 ;
      LAYER met5 ;
        RECT 0.000 4210.130 103.415 4213.000 ;
      LAYER met5 ;
        RECT 105.015 4211.730 129.965 4350.270 ;
        RECT 131.565 4211.730 135.815 4350.270 ;
        RECT 137.415 4211.730 141.665 4350.270 ;
        RECT 143.265 4211.730 152.265 4350.270 ;
        RECT 153.865 4211.730 158.315 4350.270 ;
        RECT 159.915 4349.000 163.160 4350.270 ;
      LAYER met5 ;
        RECT 163.160 4349.000 163.165 4351.870 ;
        RECT 181.715 4351.565 184.965 4351.870 ;
      LAYER met5 ;
        RECT 159.915 4213.000 163.165 4349.000 ;
        RECT 159.915 4211.730 163.160 4213.000 ;
      LAYER met5 ;
        RECT 163.160 4210.130 163.165 4213.000 ;
      LAYER met5 ;
        RECT 164.765 4211.730 168.015 4350.270 ;
        RECT 169.615 4211.730 174.065 4350.270 ;
        RECT 175.665 4211.730 180.115 4350.270 ;
        RECT 181.715 4212.035 184.965 4349.965 ;
        RECT 186.565 4211.730 191.015 4350.270 ;
        RECT 192.615 4211.730 197.865 4350.270 ;
      LAYER met5 ;
        RECT 3390.135 4316.600 3490.960 4382.500 ;
        RECT 3556.610 4316.600 3588.000 4382.500 ;
        RECT 3390.135 4314.870 3588.000 4316.600 ;
        RECT 3403.035 4314.630 3406.285 4314.870 ;
        RECT 181.715 4210.130 184.965 4210.435 ;
        RECT 0.000 4207.490 197.865 4210.130 ;
        RECT 0.000 4143.450 32.455 4207.490 ;
        RECT 96.480 4143.450 197.865 4207.490 ;
      LAYER met5 ;
        RECT 3390.135 4165.730 3395.385 4313.270 ;
        RECT 3396.985 4165.730 3401.435 4313.270 ;
        RECT 3403.035 4166.035 3406.285 4313.030 ;
        RECT 3407.885 4165.730 3412.335 4313.270 ;
        RECT 3413.935 4165.730 3418.385 4313.270 ;
        RECT 3419.985 4165.730 3423.235 4313.270 ;
        RECT 3424.840 4312.000 3428.085 4313.270 ;
        RECT 3424.835 4167.000 3428.085 4312.000 ;
      LAYER met5 ;
        RECT 3403.035 4164.130 3406.285 4164.435 ;
        RECT 3424.835 4164.130 3424.840 4167.000 ;
      LAYER met5 ;
        RECT 3424.840 4165.730 3428.085 4167.000 ;
        RECT 3429.685 4165.730 3434.135 4313.270 ;
        RECT 3435.735 4165.730 3444.735 4313.270 ;
        RECT 3446.335 4165.730 3450.585 4313.270 ;
        RECT 3452.185 4165.730 3456.435 4313.270 ;
        RECT 3458.035 4165.730 3482.985 4313.270 ;
      LAYER met5 ;
        RECT 3484.585 4312.000 3588.000 4314.870 ;
      LAYER met5 ;
        RECT 3563.785 4167.000 3588.000 4312.000 ;
      LAYER met5 ;
        RECT 3484.585 4164.130 3588.000 4167.000 ;
        RECT 0.000 4140.870 197.865 4143.450 ;
        RECT 3390.135 4161.550 3588.000 4164.130 ;
        RECT 0.000 4138.000 103.415 4140.870 ;
      LAYER met5 ;
        RECT 0.000 4002.000 24.215 4138.000 ;
      LAYER met5 ;
        RECT 0.000 3999.130 103.415 4002.000 ;
      LAYER met5 ;
        RECT 105.015 4000.730 129.965 4139.270 ;
        RECT 131.565 4000.730 135.815 4139.270 ;
        RECT 137.415 4000.730 141.665 4139.270 ;
        RECT 143.265 4000.730 152.265 4139.270 ;
        RECT 153.865 4000.730 158.315 4139.270 ;
        RECT 159.915 4138.000 163.160 4139.270 ;
      LAYER met5 ;
        RECT 163.160 4138.000 163.165 4140.870 ;
        RECT 181.715 4140.565 184.965 4140.870 ;
      LAYER met5 ;
        RECT 159.915 4002.000 163.165 4138.000 ;
        RECT 159.915 4000.730 163.160 4002.000 ;
        RECT 164.765 4000.730 168.015 4139.270 ;
        RECT 169.615 4000.730 174.065 4139.270 ;
        RECT 175.665 4000.730 180.115 4139.270 ;
        RECT 181.715 4000.970 184.965 4138.965 ;
        RECT 186.565 4000.730 191.015 4139.270 ;
        RECT 192.615 4000.730 197.865 4139.270 ;
      LAYER met5 ;
        RECT 3390.135 4097.510 3491.520 4161.550 ;
        RECT 3555.545 4097.510 3588.000 4161.550 ;
        RECT 3390.135 4094.870 3588.000 4097.510 ;
        RECT 3403.035 4094.565 3406.285 4094.870 ;
        RECT 181.715 3999.130 184.965 3999.370 ;
        RECT 0.000 3997.400 197.865 3999.130 ;
        RECT 0.000 3931.500 31.390 3997.400 ;
        RECT 97.040 3931.500 197.865 3997.400 ;
      LAYER met5 ;
        RECT 3390.135 3944.730 3395.385 4093.270 ;
        RECT 3396.985 3944.730 3401.435 4093.270 ;
        RECT 3403.035 3945.035 3406.285 4092.965 ;
        RECT 3407.885 3944.730 3412.335 4093.270 ;
        RECT 3413.935 3944.730 3418.385 4093.270 ;
        RECT 3419.985 3944.730 3423.235 4093.270 ;
      LAYER met5 ;
        RECT 3424.835 4092.000 3424.840 4094.870 ;
      LAYER met5 ;
        RECT 3424.840 4092.000 3428.085 4093.270 ;
        RECT 3424.835 3946.000 3428.085 4092.000 ;
        RECT 3424.840 3944.730 3428.085 3946.000 ;
        RECT 3429.685 3944.730 3434.135 4093.270 ;
        RECT 3435.735 3944.730 3444.735 4093.270 ;
        RECT 3446.335 3944.730 3450.585 4093.270 ;
        RECT 3452.185 3944.730 3456.435 4093.270 ;
        RECT 3458.035 3944.730 3482.985 4093.270 ;
      LAYER met5 ;
        RECT 3484.585 4092.000 3588.000 4094.870 ;
      LAYER met5 ;
        RECT 3563.785 3946.000 3588.000 4092.000 ;
      LAYER met5 ;
        RECT 3403.035 3943.130 3406.285 3943.435 ;
        RECT 3484.585 3943.130 3588.000 3946.000 ;
        RECT 0.000 3924.870 197.865 3931.500 ;
        RECT 3390.135 3936.500 3588.000 3943.130 ;
        RECT 0.000 3922.000 103.415 3924.870 ;
        RECT 181.715 3924.565 184.965 3924.870 ;
      LAYER met5 ;
        RECT 0.000 3786.000 24.215 3922.000 ;
      LAYER met5 ;
        RECT 0.000 3783.130 103.415 3786.000 ;
      LAYER met5 ;
        RECT 105.015 3784.730 129.965 3923.270 ;
        RECT 131.565 3784.730 135.815 3923.270 ;
        RECT 137.415 3784.730 141.665 3923.270 ;
        RECT 143.265 3784.730 152.265 3923.270 ;
        RECT 153.865 3784.730 158.315 3923.270 ;
        RECT 159.915 3922.000 163.160 3923.270 ;
        RECT 159.915 3786.000 163.165 3922.000 ;
        RECT 159.915 3784.730 163.160 3786.000 ;
        RECT 164.765 3784.730 168.015 3923.270 ;
        RECT 169.615 3784.730 174.065 3923.270 ;
        RECT 175.665 3784.730 180.115 3923.270 ;
        RECT 181.715 3784.970 184.965 3922.965 ;
        RECT 186.565 3784.730 191.015 3923.270 ;
        RECT 192.615 3784.730 197.865 3923.270 ;
      LAYER met5 ;
        RECT 3390.135 3870.600 3490.960 3936.500 ;
        RECT 3556.610 3870.600 3588.000 3936.500 ;
        RECT 3390.135 3868.870 3588.000 3870.600 ;
        RECT 3403.035 3868.630 3406.285 3868.870 ;
        RECT 181.715 3783.130 184.965 3783.370 ;
        RECT 0.000 3781.400 197.865 3783.130 ;
        RECT 0.000 3715.500 31.390 3781.400 ;
        RECT 97.040 3715.500 197.865 3781.400 ;
      LAYER met5 ;
        RECT 3390.135 3719.730 3395.385 3867.270 ;
        RECT 3396.985 3719.730 3401.435 3867.270 ;
        RECT 3403.035 3720.035 3406.285 3867.030 ;
        RECT 3407.885 3719.730 3412.335 3867.270 ;
        RECT 3413.935 3719.730 3418.385 3867.270 ;
        RECT 3419.985 3719.730 3423.235 3867.270 ;
        RECT 3424.840 3866.000 3428.085 3867.270 ;
        RECT 3424.835 3721.000 3428.085 3866.000 ;
        RECT 3424.840 3719.730 3428.085 3721.000 ;
        RECT 3429.685 3719.730 3434.135 3867.270 ;
        RECT 3435.735 3719.730 3444.735 3867.270 ;
        RECT 3446.335 3719.730 3450.585 3867.270 ;
        RECT 3452.185 3719.730 3456.435 3867.270 ;
        RECT 3458.035 3719.730 3482.985 3867.270 ;
      LAYER met5 ;
        RECT 3484.585 3866.000 3588.000 3868.870 ;
      LAYER met5 ;
        RECT 3563.785 3721.000 3588.000 3866.000 ;
      LAYER met5 ;
        RECT 3403.035 3718.130 3406.285 3718.435 ;
        RECT 3484.585 3718.130 3588.000 3721.000 ;
        RECT 0.000 3708.870 197.865 3715.500 ;
        RECT 3390.135 3711.500 3588.000 3718.130 ;
        RECT 0.000 3706.000 103.415 3708.870 ;
        RECT 181.715 3708.565 184.965 3708.870 ;
      LAYER met5 ;
        RECT 0.000 3570.000 24.215 3706.000 ;
      LAYER met5 ;
        RECT 0.000 3567.130 103.415 3570.000 ;
      LAYER met5 ;
        RECT 105.015 3568.730 129.965 3707.270 ;
        RECT 131.565 3568.730 135.815 3707.270 ;
        RECT 137.415 3568.730 141.665 3707.270 ;
        RECT 143.265 3568.730 152.265 3707.270 ;
        RECT 153.865 3568.730 158.315 3707.270 ;
        RECT 159.915 3706.000 163.160 3707.270 ;
        RECT 159.915 3570.000 163.165 3706.000 ;
        RECT 159.915 3568.730 163.160 3570.000 ;
        RECT 164.765 3568.730 168.015 3707.270 ;
        RECT 169.615 3568.730 174.065 3707.270 ;
        RECT 175.665 3568.730 180.115 3707.270 ;
        RECT 181.715 3568.970 184.965 3706.965 ;
        RECT 186.565 3568.730 191.015 3707.270 ;
        RECT 192.615 3568.730 197.865 3707.270 ;
      LAYER met5 ;
        RECT 3390.135 3645.600 3490.960 3711.500 ;
        RECT 3556.610 3645.600 3588.000 3711.500 ;
        RECT 3390.135 3643.870 3588.000 3645.600 ;
        RECT 3403.035 3643.630 3406.285 3643.870 ;
        RECT 181.715 3567.130 184.965 3567.370 ;
        RECT 0.000 3565.400 197.865 3567.130 ;
        RECT 0.000 3499.500 31.390 3565.400 ;
        RECT 97.040 3499.500 197.865 3565.400 ;
        RECT 0.000 3492.870 197.865 3499.500 ;
      LAYER met5 ;
        RECT 3390.135 3494.730 3395.385 3642.270 ;
        RECT 3396.985 3494.730 3401.435 3642.270 ;
        RECT 3403.035 3495.035 3406.285 3642.030 ;
        RECT 3407.885 3494.730 3412.335 3642.270 ;
        RECT 3413.935 3494.730 3418.385 3642.270 ;
        RECT 3419.985 3494.730 3423.235 3642.270 ;
        RECT 3424.840 3641.000 3428.085 3642.270 ;
        RECT 3424.835 3496.000 3428.085 3641.000 ;
        RECT 3424.840 3494.730 3428.085 3496.000 ;
        RECT 3429.685 3494.730 3434.135 3642.270 ;
        RECT 3435.735 3494.730 3444.735 3642.270 ;
        RECT 3446.335 3494.730 3450.585 3642.270 ;
        RECT 3452.185 3494.730 3456.435 3642.270 ;
        RECT 3458.035 3494.730 3482.985 3642.270 ;
      LAYER met5 ;
        RECT 3484.585 3641.000 3588.000 3643.870 ;
      LAYER met5 ;
        RECT 3563.785 3496.000 3588.000 3641.000 ;
      LAYER met5 ;
        RECT 3403.035 3493.130 3406.285 3493.435 ;
        RECT 3484.585 3493.130 3588.000 3496.000 ;
        RECT 0.000 3490.000 103.415 3492.870 ;
        RECT 181.715 3492.565 184.965 3492.870 ;
      LAYER met5 ;
        RECT 0.000 3354.000 24.215 3490.000 ;
      LAYER met5 ;
        RECT 0.000 3351.130 103.415 3354.000 ;
      LAYER met5 ;
        RECT 105.015 3352.730 129.965 3491.270 ;
        RECT 131.565 3352.730 135.815 3491.270 ;
        RECT 137.415 3352.730 141.665 3491.270 ;
        RECT 143.265 3352.730 152.265 3491.270 ;
        RECT 153.865 3352.730 158.315 3491.270 ;
        RECT 159.915 3490.000 163.160 3491.270 ;
        RECT 159.915 3354.000 163.165 3490.000 ;
        RECT 159.915 3352.730 163.160 3354.000 ;
        RECT 164.765 3352.730 168.015 3491.270 ;
        RECT 169.615 3352.730 174.065 3491.270 ;
        RECT 175.665 3352.730 180.115 3491.270 ;
        RECT 181.715 3352.970 184.965 3490.965 ;
        RECT 186.565 3352.730 191.015 3491.270 ;
        RECT 192.615 3352.730 197.865 3491.270 ;
      LAYER met5 ;
        RECT 3390.135 3486.500 3588.000 3493.130 ;
        RECT 3390.135 3420.600 3490.960 3486.500 ;
        RECT 3556.610 3420.600 3588.000 3486.500 ;
        RECT 3390.135 3418.870 3588.000 3420.600 ;
        RECT 3403.035 3418.630 3406.285 3418.870 ;
        RECT 181.715 3351.130 184.965 3351.370 ;
        RECT 0.000 3349.400 197.865 3351.130 ;
        RECT 0.000 3283.500 31.390 3349.400 ;
        RECT 97.040 3283.500 197.865 3349.400 ;
        RECT 0.000 3276.870 197.865 3283.500 ;
        RECT 0.000 3274.000 103.415 3276.870 ;
        RECT 181.715 3276.565 184.965 3276.870 ;
      LAYER met5 ;
        RECT 0.000 3138.000 24.215 3274.000 ;
      LAYER met5 ;
        RECT 0.000 3135.130 103.415 3138.000 ;
      LAYER met5 ;
        RECT 105.015 3136.730 129.965 3275.270 ;
        RECT 131.565 3136.730 135.815 3275.270 ;
        RECT 137.415 3136.730 141.665 3275.270 ;
        RECT 143.265 3136.730 152.265 3275.270 ;
        RECT 153.865 3136.730 158.315 3275.270 ;
        RECT 159.915 3274.000 163.160 3275.270 ;
        RECT 159.915 3138.000 163.165 3274.000 ;
        RECT 159.915 3136.730 163.160 3138.000 ;
        RECT 164.765 3136.730 168.015 3275.270 ;
        RECT 169.615 3136.730 174.065 3275.270 ;
        RECT 175.665 3136.730 180.115 3275.270 ;
        RECT 181.715 3136.970 184.965 3274.965 ;
        RECT 186.565 3136.730 191.015 3275.270 ;
        RECT 192.615 3136.730 197.865 3275.270 ;
        RECT 3390.135 3268.730 3395.385 3417.270 ;
        RECT 3396.985 3268.730 3401.435 3417.270 ;
        RECT 3403.035 3269.035 3406.285 3417.030 ;
        RECT 3407.885 3268.730 3412.335 3417.270 ;
        RECT 3413.935 3268.730 3418.385 3417.270 ;
        RECT 3419.985 3268.730 3423.235 3417.270 ;
        RECT 3424.840 3416.000 3428.085 3417.270 ;
        RECT 3424.835 3270.000 3428.085 3416.000 ;
        RECT 3424.840 3268.730 3428.085 3270.000 ;
        RECT 3429.685 3268.730 3434.135 3417.270 ;
        RECT 3435.735 3268.730 3444.735 3417.270 ;
        RECT 3446.335 3268.730 3450.585 3417.270 ;
        RECT 3452.185 3268.730 3456.435 3417.270 ;
        RECT 3458.035 3268.730 3482.985 3417.270 ;
      LAYER met5 ;
        RECT 3484.585 3416.000 3588.000 3418.870 ;
      LAYER met5 ;
        RECT 3563.785 3270.000 3588.000 3416.000 ;
      LAYER met5 ;
        RECT 3403.035 3267.130 3406.285 3267.435 ;
        RECT 3484.585 3267.130 3588.000 3270.000 ;
        RECT 3390.135 3260.500 3588.000 3267.130 ;
        RECT 3390.135 3194.600 3490.960 3260.500 ;
        RECT 3556.610 3194.600 3588.000 3260.500 ;
        RECT 3390.135 3192.870 3588.000 3194.600 ;
        RECT 3403.035 3192.630 3406.285 3192.870 ;
        RECT 181.715 3135.130 184.965 3135.370 ;
        RECT 0.000 3133.400 197.865 3135.130 ;
        RECT 0.000 3067.500 31.390 3133.400 ;
        RECT 97.040 3067.500 197.865 3133.400 ;
        RECT 0.000 3060.870 197.865 3067.500 ;
        RECT 0.000 3058.000 103.415 3060.870 ;
        RECT 181.715 3060.565 184.965 3060.870 ;
      LAYER met5 ;
        RECT 0.000 2922.000 24.215 3058.000 ;
      LAYER met5 ;
        RECT 0.000 2919.130 103.415 2922.000 ;
      LAYER met5 ;
        RECT 105.015 2920.730 129.965 3059.270 ;
        RECT 131.565 2920.730 135.815 3059.270 ;
        RECT 137.415 2920.730 141.665 3059.270 ;
        RECT 143.265 2920.730 152.265 3059.270 ;
        RECT 153.865 2920.730 158.315 3059.270 ;
        RECT 159.915 3058.000 163.160 3059.270 ;
        RECT 159.915 2922.000 163.165 3058.000 ;
        RECT 159.915 2920.730 163.160 2922.000 ;
        RECT 164.765 2920.730 168.015 3059.270 ;
        RECT 169.615 2920.730 174.065 3059.270 ;
        RECT 175.665 2920.730 180.115 3059.270 ;
        RECT 181.715 2920.970 184.965 3058.965 ;
        RECT 186.565 2920.730 191.015 3059.270 ;
        RECT 192.615 2920.730 197.865 3059.270 ;
        RECT 3390.135 3043.730 3395.385 3191.270 ;
        RECT 3396.985 3043.730 3401.435 3191.270 ;
        RECT 3403.035 3044.035 3406.285 3191.030 ;
        RECT 3407.885 3043.730 3412.335 3191.270 ;
        RECT 3413.935 3043.730 3418.385 3191.270 ;
        RECT 3419.985 3043.730 3423.235 3191.270 ;
        RECT 3424.840 3190.000 3428.085 3191.270 ;
        RECT 3424.835 3045.000 3428.085 3190.000 ;
        RECT 3424.840 3043.730 3428.085 3045.000 ;
        RECT 3429.685 3043.730 3434.135 3191.270 ;
        RECT 3435.735 3043.730 3444.735 3191.270 ;
        RECT 3446.335 3043.730 3450.585 3191.270 ;
        RECT 3452.185 3043.730 3456.435 3191.270 ;
        RECT 3458.035 3043.730 3482.985 3191.270 ;
      LAYER met5 ;
        RECT 3484.585 3190.000 3588.000 3192.870 ;
      LAYER met5 ;
        RECT 3563.785 3045.000 3588.000 3190.000 ;
      LAYER met5 ;
        RECT 3403.035 3042.130 3406.285 3042.435 ;
        RECT 3484.585 3042.130 3588.000 3045.000 ;
        RECT 3390.135 3035.500 3588.000 3042.130 ;
        RECT 3390.135 2969.600 3490.960 3035.500 ;
        RECT 3556.610 2969.600 3588.000 3035.500 ;
        RECT 3390.135 2967.870 3588.000 2969.600 ;
        RECT 3403.035 2967.630 3406.285 2967.870 ;
        RECT 181.715 2919.130 184.965 2919.370 ;
        RECT 0.000 2917.400 197.865 2919.130 ;
        RECT 0.000 2851.500 31.390 2917.400 ;
        RECT 97.040 2851.500 197.865 2917.400 ;
        RECT 0.000 2844.870 197.865 2851.500 ;
        RECT 0.000 2842.000 103.415 2844.870 ;
        RECT 181.715 2844.565 184.965 2844.870 ;
      LAYER met5 ;
        RECT 0.000 2706.000 24.215 2842.000 ;
      LAYER met5 ;
        RECT 0.000 2703.130 103.415 2706.000 ;
      LAYER met5 ;
        RECT 105.015 2704.730 129.965 2843.270 ;
        RECT 131.565 2704.730 135.815 2843.270 ;
        RECT 137.415 2704.730 141.665 2843.270 ;
        RECT 143.265 2704.730 152.265 2843.270 ;
        RECT 153.865 2704.730 158.315 2843.270 ;
        RECT 159.915 2842.000 163.160 2843.270 ;
        RECT 159.915 2706.000 163.165 2842.000 ;
        RECT 159.915 2704.730 163.160 2706.000 ;
        RECT 164.765 2704.730 168.015 2843.270 ;
        RECT 169.615 2704.730 174.065 2843.270 ;
        RECT 175.665 2704.730 180.115 2843.270 ;
        RECT 181.715 2704.970 184.965 2842.965 ;
        RECT 186.565 2704.730 191.015 2843.270 ;
        RECT 192.615 2704.730 197.865 2843.270 ;
        RECT 3390.135 2817.730 3395.385 2966.270 ;
        RECT 3396.985 2817.730 3401.435 2966.270 ;
        RECT 3403.035 2818.035 3406.285 2966.030 ;
        RECT 3407.885 2817.730 3412.335 2966.270 ;
        RECT 3413.935 2817.730 3418.385 2966.270 ;
        RECT 3419.985 2817.730 3423.235 2966.270 ;
        RECT 3424.840 2965.000 3428.085 2966.270 ;
        RECT 3424.835 2819.000 3428.085 2965.000 ;
        RECT 3424.840 2817.730 3428.085 2819.000 ;
        RECT 3429.685 2817.730 3434.135 2966.270 ;
        RECT 3435.735 2817.730 3444.735 2966.270 ;
        RECT 3446.335 2817.730 3450.585 2966.270 ;
        RECT 3452.185 2817.730 3456.435 2966.270 ;
        RECT 3458.035 2817.730 3482.985 2966.270 ;
      LAYER met5 ;
        RECT 3484.585 2965.000 3588.000 2967.870 ;
      LAYER met5 ;
        RECT 3563.785 2819.000 3588.000 2965.000 ;
      LAYER met5 ;
        RECT 3403.035 2816.130 3406.285 2816.435 ;
        RECT 3484.585 2816.130 3588.000 2819.000 ;
        RECT 3390.135 2809.500 3588.000 2816.130 ;
        RECT 3390.135 2743.600 3490.960 2809.500 ;
        RECT 3556.610 2743.600 3588.000 2809.500 ;
        RECT 3390.135 2741.870 3588.000 2743.600 ;
        RECT 3403.035 2741.630 3406.285 2741.870 ;
        RECT 181.715 2703.130 184.965 2703.370 ;
        RECT 0.000 2701.400 197.865 2703.130 ;
        RECT 0.000 2635.500 31.390 2701.400 ;
        RECT 97.040 2635.500 197.865 2701.400 ;
        RECT 0.000 2628.870 197.865 2635.500 ;
        RECT 0.000 2626.000 103.415 2628.870 ;
        RECT 181.715 2628.565 184.965 2628.870 ;
      LAYER met5 ;
        RECT 0.000 2490.000 24.215 2626.000 ;
      LAYER met5 ;
        RECT 0.000 2487.130 103.415 2490.000 ;
      LAYER met5 ;
        RECT 105.015 2488.730 129.965 2627.270 ;
        RECT 131.565 2488.730 135.815 2627.270 ;
        RECT 137.415 2488.730 141.665 2627.270 ;
        RECT 143.265 2488.730 152.265 2627.270 ;
        RECT 153.865 2488.730 158.315 2627.270 ;
        RECT 159.915 2626.000 163.160 2627.270 ;
        RECT 159.915 2490.000 163.165 2626.000 ;
        RECT 159.915 2488.730 163.160 2490.000 ;
      LAYER met5 ;
        RECT 163.160 2487.130 163.165 2490.000 ;
      LAYER met5 ;
        RECT 164.765 2488.730 168.015 2627.270 ;
        RECT 169.615 2488.730 174.065 2627.270 ;
        RECT 175.665 2488.730 180.115 2627.270 ;
        RECT 181.715 2489.035 184.965 2626.965 ;
        RECT 186.565 2488.730 191.015 2627.270 ;
        RECT 192.615 2488.730 197.865 2627.270 ;
        RECT 3390.135 2592.730 3395.385 2740.270 ;
        RECT 3396.985 2592.730 3401.435 2740.270 ;
        RECT 3403.035 2593.035 3406.285 2740.030 ;
        RECT 3407.885 2592.730 3412.335 2740.270 ;
        RECT 3413.935 2592.730 3418.385 2740.270 ;
        RECT 3419.985 2592.730 3423.235 2740.270 ;
        RECT 3424.840 2739.000 3428.085 2740.270 ;
        RECT 3424.835 2594.000 3428.085 2739.000 ;
      LAYER met5 ;
        RECT 3403.035 2591.130 3406.285 2591.435 ;
        RECT 3424.835 2591.130 3424.840 2594.000 ;
      LAYER met5 ;
        RECT 3424.840 2592.730 3428.085 2594.000 ;
        RECT 3429.685 2592.730 3434.135 2740.270 ;
        RECT 3435.735 2592.730 3444.735 2740.270 ;
        RECT 3446.335 2592.730 3450.585 2740.270 ;
        RECT 3452.185 2592.730 3456.435 2740.270 ;
        RECT 3458.035 2592.730 3482.985 2740.270 ;
      LAYER met5 ;
        RECT 3484.585 2739.000 3588.000 2741.870 ;
      LAYER met5 ;
        RECT 3563.785 2594.000 3588.000 2739.000 ;
      LAYER met5 ;
        RECT 3484.585 2591.130 3588.000 2594.000 ;
        RECT 3390.135 2588.550 3588.000 2591.130 ;
        RECT 3390.135 2524.510 3491.520 2588.550 ;
        RECT 3555.545 2524.510 3588.000 2588.550 ;
        RECT 3390.135 2521.870 3588.000 2524.510 ;
        RECT 3403.035 2521.565 3406.285 2521.870 ;
        RECT 181.715 2487.130 184.965 2487.435 ;
        RECT 0.000 2484.490 197.865 2487.130 ;
        RECT 0.000 2420.450 32.455 2484.490 ;
        RECT 96.480 2420.450 197.865 2484.490 ;
        RECT 0.000 2417.870 197.865 2420.450 ;
        RECT 0.000 2415.000 103.415 2417.870 ;
      LAYER met5 ;
        RECT 0.000 2279.000 24.215 2415.000 ;
      LAYER met5 ;
        RECT 0.000 2276.130 103.415 2279.000 ;
      LAYER met5 ;
        RECT 105.015 2277.730 129.965 2416.270 ;
        RECT 131.565 2277.730 135.815 2416.270 ;
        RECT 137.415 2277.730 141.665 2416.270 ;
        RECT 143.265 2277.730 152.265 2416.270 ;
        RECT 153.865 2277.730 158.315 2416.270 ;
        RECT 159.915 2415.000 163.160 2416.270 ;
      LAYER met5 ;
        RECT 163.160 2415.000 163.165 2417.870 ;
        RECT 181.715 2417.565 184.965 2417.870 ;
      LAYER met5 ;
        RECT 159.915 2279.000 163.165 2415.000 ;
        RECT 159.915 2277.730 163.160 2279.000 ;
        RECT 164.765 2277.730 168.015 2416.270 ;
        RECT 169.615 2277.730 174.065 2416.270 ;
        RECT 175.665 2277.730 180.115 2416.270 ;
        RECT 181.715 2278.035 184.965 2415.965 ;
        RECT 186.565 2277.730 191.015 2416.270 ;
        RECT 192.615 2277.730 197.865 2416.270 ;
        RECT 3390.135 2372.730 3395.385 2520.270 ;
        RECT 3396.985 2372.730 3401.435 2520.270 ;
        RECT 3403.035 2373.035 3406.285 2519.965 ;
        RECT 3407.885 2372.730 3412.335 2520.270 ;
        RECT 3413.935 2372.730 3418.385 2520.270 ;
        RECT 3419.985 2372.730 3423.235 2520.270 ;
      LAYER met5 ;
        RECT 3424.835 2519.000 3424.840 2521.870 ;
      LAYER met5 ;
        RECT 3424.840 2519.000 3428.085 2520.270 ;
        RECT 3424.835 2374.000 3428.085 2519.000 ;
        RECT 3424.840 2372.730 3428.085 2374.000 ;
        RECT 3429.685 2372.730 3434.135 2520.270 ;
        RECT 3435.735 2372.730 3444.735 2520.270 ;
        RECT 3446.335 2372.730 3450.585 2520.270 ;
        RECT 3452.185 2372.730 3456.435 2520.270 ;
        RECT 3458.035 2372.730 3482.985 2520.270 ;
      LAYER met5 ;
        RECT 3484.585 2519.000 3588.000 2521.870 ;
      LAYER met5 ;
        RECT 3563.785 2374.000 3588.000 2519.000 ;
      LAYER met5 ;
        RECT 3403.035 2371.130 3406.285 2371.435 ;
        RECT 3484.585 2371.130 3588.000 2374.000 ;
        RECT 3390.135 2365.330 3588.000 2371.130 ;
        RECT 3390.135 2307.730 3488.300 2365.330 ;
        RECT 3558.765 2307.730 3588.000 2365.330 ;
        RECT 3390.135 2301.870 3588.000 2307.730 ;
        RECT 3403.035 2301.565 3406.285 2301.870 ;
        RECT 181.715 2276.130 184.965 2276.435 ;
        RECT 0.000 2270.270 197.865 2276.130 ;
        RECT 0.000 2212.670 29.235 2270.270 ;
        RECT 99.700 2212.670 197.865 2270.270 ;
        RECT 0.000 2206.870 197.865 2212.670 ;
        RECT 0.000 2204.000 103.415 2206.870 ;
        RECT 181.715 2206.565 184.965 2206.870 ;
      LAYER met5 ;
        RECT 0.000 2068.000 24.215 2204.000 ;
      LAYER met5 ;
        RECT 0.000 2065.130 103.415 2068.000 ;
      LAYER met5 ;
        RECT 105.015 2066.730 129.965 2205.270 ;
        RECT 131.565 2066.730 135.815 2205.270 ;
        RECT 137.415 2066.730 141.665 2205.270 ;
        RECT 143.265 2066.730 152.265 2205.270 ;
        RECT 153.865 2066.730 158.315 2205.270 ;
        RECT 159.915 2204.000 163.160 2205.270 ;
        RECT 159.915 2068.000 163.165 2204.000 ;
        RECT 159.915 2066.730 163.160 2068.000 ;
        RECT 164.765 2066.730 168.015 2205.270 ;
        RECT 169.615 2066.730 174.065 2205.270 ;
        RECT 175.665 2066.730 180.115 2205.270 ;
        RECT 181.715 2066.970 184.965 2204.965 ;
        RECT 186.565 2066.730 191.015 2205.270 ;
        RECT 192.615 2066.730 197.865 2205.270 ;
        RECT 3390.135 2151.730 3395.385 2300.270 ;
        RECT 3396.985 2151.730 3401.435 2300.270 ;
        RECT 3403.035 2152.035 3406.285 2299.965 ;
        RECT 3407.885 2151.730 3412.335 2300.270 ;
        RECT 3413.935 2151.730 3418.385 2300.270 ;
        RECT 3419.985 2151.730 3423.235 2300.270 ;
        RECT 3424.840 2299.000 3428.085 2300.270 ;
        RECT 3424.835 2153.000 3428.085 2299.000 ;
      LAYER met5 ;
        RECT 3403.035 2150.130 3406.285 2150.435 ;
        RECT 3424.835 2150.130 3424.840 2153.000 ;
      LAYER met5 ;
        RECT 3424.840 2151.730 3428.085 2153.000 ;
        RECT 3429.685 2151.730 3434.135 2300.270 ;
        RECT 3435.735 2151.730 3444.735 2300.270 ;
        RECT 3446.335 2151.730 3450.585 2300.270 ;
        RECT 3452.185 2151.730 3456.435 2300.270 ;
        RECT 3458.035 2151.730 3482.985 2300.270 ;
      LAYER met5 ;
        RECT 3484.585 2299.000 3588.000 2301.870 ;
      LAYER met5 ;
        RECT 3563.785 2153.000 3588.000 2299.000 ;
      LAYER met5 ;
        RECT 3484.585 2150.130 3588.000 2153.000 ;
        RECT 3390.135 2147.550 3588.000 2150.130 ;
        RECT 3390.135 2083.510 3491.520 2147.550 ;
        RECT 3555.545 2083.510 3588.000 2147.550 ;
        RECT 3390.135 2080.870 3588.000 2083.510 ;
        RECT 3403.035 2080.565 3406.285 2080.870 ;
        RECT 181.715 2065.130 184.965 2065.370 ;
        RECT 0.000 2063.400 197.865 2065.130 ;
        RECT 0.000 1997.500 31.390 2063.400 ;
        RECT 97.040 1997.500 197.865 2063.400 ;
        RECT 0.000 1990.870 197.865 1997.500 ;
        RECT 0.000 1988.000 103.415 1990.870 ;
        RECT 181.715 1990.565 184.965 1990.870 ;
      LAYER met5 ;
        RECT 0.000 1852.000 24.215 1988.000 ;
      LAYER met5 ;
        RECT 0.000 1849.130 103.415 1852.000 ;
      LAYER met5 ;
        RECT 105.015 1850.730 129.965 1989.270 ;
        RECT 131.565 1850.730 135.815 1989.270 ;
        RECT 137.415 1850.730 141.665 1989.270 ;
        RECT 143.265 1850.730 152.265 1989.270 ;
        RECT 153.865 1850.730 158.315 1989.270 ;
        RECT 159.915 1988.000 163.160 1989.270 ;
        RECT 159.915 1852.000 163.165 1988.000 ;
        RECT 159.915 1850.730 163.160 1852.000 ;
        RECT 164.765 1850.730 168.015 1989.270 ;
        RECT 169.615 1850.730 174.065 1989.270 ;
        RECT 175.665 1850.730 180.115 1989.270 ;
        RECT 181.715 1850.970 184.965 1988.965 ;
        RECT 186.565 1850.730 191.015 1989.270 ;
        RECT 192.615 1850.730 197.865 1989.270 ;
        RECT 3390.135 1931.730 3395.385 2079.270 ;
        RECT 3396.985 1931.730 3401.435 2079.270 ;
        RECT 3403.035 1932.035 3406.285 2078.965 ;
        RECT 3407.885 1931.730 3412.335 2079.270 ;
        RECT 3413.935 1931.730 3418.385 2079.270 ;
        RECT 3419.985 1931.730 3423.235 2079.270 ;
      LAYER met5 ;
        RECT 3424.835 2078.000 3424.840 2080.870 ;
      LAYER met5 ;
        RECT 3424.840 2078.000 3428.085 2079.270 ;
        RECT 3424.835 1933.000 3428.085 2078.000 ;
        RECT 3424.840 1931.730 3428.085 1933.000 ;
        RECT 3429.685 1931.730 3434.135 2079.270 ;
        RECT 3435.735 1931.730 3444.735 2079.270 ;
        RECT 3446.335 1931.730 3450.585 2079.270 ;
        RECT 3452.185 1931.730 3456.435 2079.270 ;
        RECT 3458.035 1931.730 3482.985 2079.270 ;
      LAYER met5 ;
        RECT 3484.585 2078.000 3588.000 2080.870 ;
      LAYER met5 ;
        RECT 3563.785 1933.000 3588.000 2078.000 ;
      LAYER met5 ;
        RECT 3403.035 1930.130 3406.285 1930.435 ;
        RECT 3484.585 1930.130 3588.000 1933.000 ;
        RECT 3390.135 1923.500 3588.000 1930.130 ;
        RECT 3390.135 1857.600 3490.960 1923.500 ;
        RECT 3556.610 1857.600 3588.000 1923.500 ;
        RECT 3390.135 1855.870 3588.000 1857.600 ;
        RECT 3403.035 1855.630 3406.285 1855.870 ;
        RECT 181.715 1849.130 184.965 1849.370 ;
        RECT 0.000 1847.400 197.865 1849.130 ;
        RECT 0.000 1781.500 31.390 1847.400 ;
        RECT 97.040 1781.500 197.865 1847.400 ;
        RECT 0.000 1774.870 197.865 1781.500 ;
        RECT 0.000 1772.000 103.415 1774.870 ;
        RECT 181.715 1774.565 184.965 1774.870 ;
      LAYER met5 ;
        RECT 0.000 1636.000 24.215 1772.000 ;
      LAYER met5 ;
        RECT 0.000 1633.130 103.415 1636.000 ;
      LAYER met5 ;
        RECT 105.015 1634.730 129.965 1773.270 ;
        RECT 131.565 1634.730 135.815 1773.270 ;
        RECT 137.415 1634.730 141.665 1773.270 ;
        RECT 143.265 1634.730 152.265 1773.270 ;
        RECT 153.865 1634.730 158.315 1773.270 ;
        RECT 159.915 1772.000 163.160 1773.270 ;
        RECT 159.915 1636.000 163.165 1772.000 ;
        RECT 159.915 1634.730 163.160 1636.000 ;
        RECT 164.765 1634.730 168.015 1773.270 ;
        RECT 169.615 1634.730 174.065 1773.270 ;
        RECT 175.665 1634.730 180.115 1773.270 ;
        RECT 181.715 1634.970 184.965 1772.965 ;
        RECT 186.565 1634.730 191.015 1773.270 ;
        RECT 192.615 1634.730 197.865 1773.270 ;
        RECT 3390.135 1705.730 3395.385 1854.270 ;
        RECT 3396.985 1705.730 3401.435 1854.270 ;
        RECT 3403.035 1706.035 3406.285 1854.030 ;
        RECT 3407.885 1705.730 3412.335 1854.270 ;
        RECT 3413.935 1705.730 3418.385 1854.270 ;
        RECT 3419.985 1705.730 3423.235 1854.270 ;
        RECT 3424.840 1853.000 3428.085 1854.270 ;
        RECT 3424.835 1707.000 3428.085 1853.000 ;
        RECT 3424.840 1705.730 3428.085 1707.000 ;
        RECT 3429.685 1705.730 3434.135 1854.270 ;
        RECT 3435.735 1705.730 3444.735 1854.270 ;
        RECT 3446.335 1705.730 3450.585 1854.270 ;
        RECT 3452.185 1705.730 3456.435 1854.270 ;
        RECT 3458.035 1705.730 3482.985 1854.270 ;
      LAYER met5 ;
        RECT 3484.585 1853.000 3588.000 1855.870 ;
      LAYER met5 ;
        RECT 3563.785 1707.000 3588.000 1853.000 ;
      LAYER met5 ;
        RECT 3403.035 1704.130 3406.285 1704.435 ;
        RECT 3484.585 1704.130 3588.000 1707.000 ;
        RECT 3390.135 1697.500 3588.000 1704.130 ;
        RECT 181.715 1633.130 184.965 1633.370 ;
        RECT 0.000 1631.400 197.865 1633.130 ;
        RECT 0.000 1565.500 31.390 1631.400 ;
        RECT 97.040 1565.500 197.865 1631.400 ;
        RECT 3390.135 1631.600 3490.960 1697.500 ;
        RECT 3556.610 1631.600 3588.000 1697.500 ;
        RECT 3390.135 1629.870 3588.000 1631.600 ;
        RECT 3403.035 1629.630 3406.285 1629.870 ;
        RECT 0.000 1558.870 197.865 1565.500 ;
        RECT 0.000 1556.000 103.415 1558.870 ;
        RECT 181.715 1558.565 184.965 1558.870 ;
      LAYER met5 ;
        RECT 0.000 1420.000 24.215 1556.000 ;
      LAYER met5 ;
        RECT 0.000 1417.130 103.415 1420.000 ;
      LAYER met5 ;
        RECT 105.015 1418.730 129.965 1557.270 ;
        RECT 131.565 1418.730 135.815 1557.270 ;
        RECT 137.415 1418.730 141.665 1557.270 ;
        RECT 143.265 1418.730 152.265 1557.270 ;
        RECT 153.865 1418.730 158.315 1557.270 ;
        RECT 159.915 1556.000 163.160 1557.270 ;
        RECT 159.915 1420.000 163.165 1556.000 ;
        RECT 159.915 1418.730 163.160 1420.000 ;
        RECT 164.765 1418.730 168.015 1557.270 ;
        RECT 169.615 1418.730 174.065 1557.270 ;
        RECT 175.665 1418.730 180.115 1557.270 ;
        RECT 181.715 1418.970 184.965 1556.965 ;
        RECT 186.565 1418.730 191.015 1557.270 ;
        RECT 192.615 1418.730 197.865 1557.270 ;
        RECT 3390.135 1480.730 3395.385 1628.270 ;
        RECT 3396.985 1480.730 3401.435 1628.270 ;
        RECT 3403.035 1481.035 3406.285 1628.030 ;
        RECT 3407.885 1480.730 3412.335 1628.270 ;
        RECT 3413.935 1480.730 3418.385 1628.270 ;
        RECT 3419.985 1480.730 3423.235 1628.270 ;
        RECT 3424.840 1627.000 3428.085 1628.270 ;
        RECT 3424.835 1482.000 3428.085 1627.000 ;
        RECT 3424.840 1480.730 3428.085 1482.000 ;
        RECT 3429.685 1480.730 3434.135 1628.270 ;
        RECT 3435.735 1480.730 3444.735 1628.270 ;
        RECT 3446.335 1480.730 3450.585 1628.270 ;
        RECT 3452.185 1480.730 3456.435 1628.270 ;
        RECT 3458.035 1480.730 3482.985 1628.270 ;
      LAYER met5 ;
        RECT 3484.585 1627.000 3588.000 1629.870 ;
      LAYER met5 ;
        RECT 3563.785 1482.000 3588.000 1627.000 ;
      LAYER met5 ;
        RECT 3403.035 1479.130 3406.285 1479.435 ;
        RECT 3484.585 1479.130 3588.000 1482.000 ;
        RECT 3390.135 1472.500 3588.000 1479.130 ;
        RECT 181.715 1417.130 184.965 1417.370 ;
        RECT 0.000 1415.400 197.865 1417.130 ;
        RECT 0.000 1349.500 31.390 1415.400 ;
        RECT 97.040 1349.500 197.865 1415.400 ;
        RECT 3390.135 1406.600 3490.960 1472.500 ;
        RECT 3556.610 1406.600 3588.000 1472.500 ;
        RECT 3390.135 1404.870 3588.000 1406.600 ;
        RECT 3403.035 1404.630 3406.285 1404.870 ;
        RECT 0.000 1342.870 197.865 1349.500 ;
        RECT 0.000 1340.000 103.415 1342.870 ;
        RECT 181.715 1342.565 184.965 1342.870 ;
      LAYER met5 ;
        RECT 0.000 1204.000 24.215 1340.000 ;
      LAYER met5 ;
        RECT 0.000 1201.130 103.415 1204.000 ;
      LAYER met5 ;
        RECT 105.015 1202.730 129.965 1341.270 ;
        RECT 131.565 1202.730 135.815 1341.270 ;
        RECT 137.415 1202.730 141.665 1341.270 ;
        RECT 143.265 1202.730 152.265 1341.270 ;
        RECT 153.865 1202.730 158.315 1341.270 ;
        RECT 159.915 1340.000 163.160 1341.270 ;
        RECT 159.915 1204.000 163.165 1340.000 ;
        RECT 159.915 1202.730 163.160 1204.000 ;
        RECT 164.765 1202.730 168.015 1341.270 ;
        RECT 169.615 1202.730 174.065 1341.270 ;
        RECT 175.665 1202.730 180.115 1341.270 ;
        RECT 181.715 1202.970 184.965 1340.965 ;
        RECT 186.565 1202.730 191.015 1341.270 ;
        RECT 192.615 1202.730 197.865 1341.270 ;
        RECT 3390.135 1255.730 3395.385 1403.270 ;
        RECT 3396.985 1255.730 3401.435 1403.270 ;
        RECT 3403.035 1256.035 3406.285 1403.030 ;
        RECT 3407.885 1255.730 3412.335 1403.270 ;
        RECT 3413.935 1255.730 3418.385 1403.270 ;
        RECT 3419.985 1255.730 3423.235 1403.270 ;
        RECT 3424.840 1402.000 3428.085 1403.270 ;
        RECT 3424.835 1257.000 3428.085 1402.000 ;
        RECT 3424.840 1255.730 3428.085 1257.000 ;
        RECT 3429.685 1255.730 3434.135 1403.270 ;
        RECT 3435.735 1255.730 3444.735 1403.270 ;
        RECT 3446.335 1255.730 3450.585 1403.270 ;
        RECT 3452.185 1255.730 3456.435 1403.270 ;
        RECT 3458.035 1255.730 3482.985 1403.270 ;
      LAYER met5 ;
        RECT 3484.585 1402.000 3588.000 1404.870 ;
      LAYER met5 ;
        RECT 3563.785 1257.000 3588.000 1402.000 ;
      LAYER met5 ;
        RECT 3403.035 1254.130 3406.285 1254.435 ;
        RECT 3484.585 1254.130 3588.000 1257.000 ;
        RECT 3390.135 1247.500 3588.000 1254.130 ;
        RECT 181.715 1201.130 184.965 1201.370 ;
        RECT 0.000 1199.400 197.865 1201.130 ;
        RECT 0.000 1133.500 31.390 1199.400 ;
        RECT 97.040 1133.500 197.865 1199.400 ;
        RECT 3390.135 1181.600 3490.960 1247.500 ;
        RECT 3556.610 1181.600 3588.000 1247.500 ;
        RECT 3390.135 1179.870 3588.000 1181.600 ;
        RECT 3403.035 1179.630 3406.285 1179.870 ;
        RECT 0.000 1126.870 197.865 1133.500 ;
        RECT 0.000 1124.000 103.415 1126.870 ;
        RECT 181.715 1126.565 184.965 1126.870 ;
      LAYER met5 ;
        RECT 0.000 988.000 24.215 1124.000 ;
      LAYER met5 ;
        RECT 0.000 985.130 103.415 988.000 ;
      LAYER met5 ;
        RECT 105.015 986.730 129.965 1125.270 ;
        RECT 131.565 986.730 135.815 1125.270 ;
        RECT 137.415 986.730 141.665 1125.270 ;
        RECT 143.265 986.730 152.265 1125.270 ;
        RECT 153.865 986.730 158.315 1125.270 ;
        RECT 159.915 1124.000 163.160 1125.270 ;
        RECT 159.915 988.000 163.165 1124.000 ;
        RECT 159.915 986.730 163.160 988.000 ;
        RECT 164.765 986.730 168.015 1125.270 ;
        RECT 169.615 986.730 174.065 1125.270 ;
        RECT 175.665 986.730 180.115 1125.270 ;
        RECT 181.715 986.970 184.965 1124.965 ;
        RECT 186.565 986.730 191.015 1125.270 ;
        RECT 192.615 986.730 197.865 1125.270 ;
        RECT 3390.135 1029.730 3395.385 1178.270 ;
        RECT 3396.985 1029.730 3401.435 1178.270 ;
        RECT 3403.035 1030.035 3406.285 1178.030 ;
        RECT 3407.885 1029.730 3412.335 1178.270 ;
        RECT 3413.935 1029.730 3418.385 1178.270 ;
        RECT 3419.985 1029.730 3423.235 1178.270 ;
        RECT 3424.840 1177.000 3428.085 1178.270 ;
        RECT 3424.835 1031.000 3428.085 1177.000 ;
        RECT 3424.840 1029.730 3428.085 1031.000 ;
        RECT 3429.685 1029.730 3434.135 1178.270 ;
        RECT 3435.735 1029.730 3444.735 1178.270 ;
        RECT 3446.335 1029.730 3450.585 1178.270 ;
        RECT 3452.185 1029.730 3456.435 1178.270 ;
        RECT 3458.035 1029.730 3482.985 1178.270 ;
      LAYER met5 ;
        RECT 3484.585 1177.000 3588.000 1179.870 ;
      LAYER met5 ;
        RECT 3563.785 1031.000 3588.000 1177.000 ;
      LAYER met5 ;
        RECT 3403.035 1028.130 3406.285 1028.435 ;
        RECT 3484.585 1028.130 3588.000 1031.000 ;
        RECT 3390.135 1021.500 3588.000 1028.130 ;
        RECT 181.715 985.130 184.965 985.370 ;
        RECT 0.000 983.400 197.865 985.130 ;
        RECT 0.000 917.500 31.390 983.400 ;
        RECT 97.040 917.500 197.865 983.400 ;
        RECT 3390.135 955.600 3490.960 1021.500 ;
        RECT 3556.610 955.600 3588.000 1021.500 ;
        RECT 3390.135 953.870 3588.000 955.600 ;
        RECT 3403.035 953.630 3406.285 953.870 ;
        RECT 0.000 910.870 197.865 917.500 ;
        RECT 0.000 908.000 103.415 910.870 ;
        RECT 181.715 910.565 184.965 910.870 ;
      LAYER met5 ;
        RECT 0.000 626.000 24.215 908.000 ;
      LAYER met5 ;
        RECT 0.000 623.130 103.415 626.000 ;
      LAYER met5 ;
        RECT 105.015 624.730 129.965 909.270 ;
        RECT 131.565 624.730 135.815 909.270 ;
        RECT 137.415 624.730 141.665 909.270 ;
        RECT 143.265 767.000 152.265 909.270 ;
        RECT 153.865 772.000 158.315 909.270 ;
        RECT 159.915 908.000 163.160 909.270 ;
        RECT 159.915 767.000 163.165 908.000 ;
        RECT 143.265 624.730 152.265 762.000 ;
        RECT 153.865 624.730 158.315 767.000 ;
        RECT 159.915 626.000 163.165 762.000 ;
        RECT 159.915 624.730 163.160 626.000 ;
      LAYER met5 ;
        RECT 163.160 623.130 163.165 626.000 ;
      LAYER met5 ;
        RECT 164.765 624.730 168.015 909.270 ;
        RECT 169.615 624.730 174.065 909.270 ;
        RECT 175.665 624.730 180.115 909.270 ;
        RECT 181.715 767.000 184.965 908.965 ;
        RECT 186.565 772.000 191.015 909.270 ;
        RECT 181.715 625.035 184.965 762.000 ;
        RECT 186.565 624.730 191.015 767.000 ;
        RECT 192.615 624.730 197.865 909.270 ;
        RECT 3390.135 804.730 3395.385 952.270 ;
        RECT 3396.985 804.730 3401.435 952.270 ;
        RECT 3403.035 805.035 3406.285 952.030 ;
        RECT 3407.885 804.730 3412.335 952.270 ;
        RECT 3413.935 804.730 3418.385 952.270 ;
        RECT 3419.985 804.730 3423.235 952.270 ;
        RECT 3424.840 951.000 3428.085 952.270 ;
        RECT 3424.835 806.000 3428.085 951.000 ;
        RECT 3424.840 804.730 3428.085 806.000 ;
        RECT 3429.685 804.730 3434.135 952.270 ;
        RECT 3435.735 804.730 3444.735 952.270 ;
        RECT 3446.335 804.730 3450.585 952.270 ;
        RECT 3452.185 804.730 3456.435 952.270 ;
        RECT 3458.035 804.730 3482.985 952.270 ;
      LAYER met5 ;
        RECT 3484.585 951.000 3588.000 953.870 ;
      LAYER met5 ;
        RECT 3563.785 806.000 3588.000 951.000 ;
      LAYER met5 ;
        RECT 3403.035 803.130 3406.285 803.435 ;
        RECT 3484.585 803.130 3588.000 806.000 ;
        RECT 3390.135 796.500 3588.000 803.130 ;
        RECT 3390.135 730.600 3490.960 796.500 ;
        RECT 3556.610 730.600 3588.000 796.500 ;
        RECT 3390.135 728.870 3588.000 730.600 ;
        RECT 3403.035 728.630 3406.285 728.870 ;
        RECT 181.715 623.130 184.965 623.435 ;
        RECT 0.000 620.490 197.865 623.130 ;
        RECT 0.000 556.450 32.455 620.490 ;
        RECT 96.480 556.450 197.865 620.490 ;
      LAYER met5 ;
        RECT 3390.135 578.730 3395.385 727.270 ;
        RECT 3396.985 578.730 3401.435 727.270 ;
        RECT 3403.035 579.035 3406.285 727.030 ;
        RECT 3407.885 578.730 3412.335 727.270 ;
        RECT 3413.935 578.730 3418.385 727.270 ;
        RECT 3419.985 578.730 3423.235 727.270 ;
        RECT 3424.840 726.000 3428.085 727.270 ;
        RECT 3424.835 580.000 3428.085 726.000 ;
        RECT 3424.840 578.730 3428.085 580.000 ;
        RECT 3429.685 578.730 3434.135 727.270 ;
        RECT 3435.735 578.730 3444.735 727.270 ;
        RECT 3446.335 578.730 3450.585 727.270 ;
        RECT 3452.185 578.730 3456.435 727.270 ;
        RECT 3458.035 578.730 3482.985 727.270 ;
      LAYER met5 ;
        RECT 3484.585 726.000 3588.000 728.870 ;
      LAYER met5 ;
        RECT 3563.785 580.000 3588.000 726.000 ;
      LAYER met5 ;
        RECT 3403.035 577.130 3406.285 577.435 ;
        RECT 3484.585 577.130 3588.000 580.000 ;
        RECT 0.000 553.870 197.865 556.450 ;
        RECT 3390.135 570.500 3588.000 577.130 ;
        RECT 0.000 551.000 103.415 553.870 ;
      LAYER met5 ;
        RECT 0.000 415.000 24.215 551.000 ;
      LAYER met5 ;
        RECT 0.000 412.130 103.415 415.000 ;
      LAYER met5 ;
        RECT 105.015 413.730 129.965 552.270 ;
        RECT 131.565 413.730 135.815 552.270 ;
        RECT 137.415 413.730 141.665 552.270 ;
        RECT 143.265 413.730 152.265 552.270 ;
        RECT 153.865 413.730 158.315 552.270 ;
        RECT 159.915 551.000 163.160 552.270 ;
      LAYER met5 ;
        RECT 163.160 551.000 163.165 553.870 ;
        RECT 181.715 553.565 184.965 553.870 ;
      LAYER met5 ;
        RECT 159.915 415.000 163.165 551.000 ;
        RECT 159.915 413.730 163.160 415.000 ;
      LAYER met5 ;
        RECT 163.160 412.130 163.165 415.000 ;
      LAYER met5 ;
        RECT 164.765 413.730 168.015 552.270 ;
        RECT 169.615 413.730 174.065 552.270 ;
        RECT 175.665 413.730 180.115 552.270 ;
        RECT 181.715 414.035 184.965 551.965 ;
        RECT 186.565 413.730 191.015 552.270 ;
        RECT 192.615 413.730 197.865 552.270 ;
      LAYER met5 ;
        RECT 3390.135 504.600 3490.960 570.500 ;
        RECT 3556.610 504.600 3588.000 570.500 ;
        RECT 3390.135 502.870 3588.000 504.600 ;
        RECT 3403.035 502.630 3406.285 502.870 ;
        RECT 181.715 412.130 184.965 412.435 ;
        RECT 0.000 406.270 197.865 412.130 ;
        RECT 0.000 348.670 29.235 406.270 ;
        RECT 99.700 348.670 197.865 406.270 ;
        RECT 0.000 342.870 197.865 348.670 ;
        RECT 0.000 340.000 103.415 342.870 ;
      LAYER met5 ;
        RECT 0.000 204.000 24.215 340.000 ;
      LAYER met5 ;
        RECT 0.000 200.545 103.415 204.000 ;
      LAYER met5 ;
        RECT 105.015 202.145 129.965 341.270 ;
        RECT 131.565 202.730 135.815 341.270 ;
        RECT 137.415 202.730 141.665 341.270 ;
      LAYER met5 ;
        RECT 131.565 200.545 141.665 201.130 ;
        RECT 0.000 175.245 141.665 200.545 ;
      LAYER met5 ;
        RECT 143.265 176.845 152.265 341.270 ;
        RECT 153.865 202.730 158.315 341.270 ;
        RECT 159.915 340.000 163.160 341.270 ;
      LAYER met5 ;
        RECT 163.160 340.000 163.165 342.870 ;
        RECT 181.715 342.565 184.965 342.870 ;
      LAYER met5 ;
        RECT 159.915 204.000 163.165 340.000 ;
        RECT 159.915 202.730 163.160 204.000 ;
        RECT 164.765 202.730 168.015 341.270 ;
        RECT 169.615 202.730 174.065 341.270 ;
        RECT 175.665 202.730 180.115 341.270 ;
        RECT 181.715 202.745 184.965 340.965 ;
        RECT 186.565 202.730 191.015 341.270 ;
        RECT 192.615 202.730 197.865 341.270 ;
      LAYER met5 ;
        RECT 181.715 201.130 184.965 201.145 ;
        RECT 199.465 201.130 200.000 204.000 ;
        RECT 153.865 199.465 200.000 201.130 ;
        RECT 3384.000 199.465 3388.535 200.000 ;
        RECT 153.865 192.615 196.050 199.465 ;
      LAYER met5 ;
        RECT 197.650 192.615 395.270 197.865 ;
      LAYER met5 ;
        RECT 153.865 184.965 194.615 192.615 ;
      LAYER met5 ;
        RECT 237.000 191.015 357.000 192.615 ;
        RECT 196.215 186.565 395.270 191.015 ;
      LAYER met5 ;
        RECT 396.870 184.965 466.130 197.865 ;
      LAYER met5 ;
        RECT 467.730 192.615 664.270 197.865 ;
        RECT 506.000 191.015 626.000 192.615 ;
        RECT 467.730 186.565 664.270 191.015 ;
      LAYER met5 ;
        RECT 665.870 184.965 735.130 197.865 ;
      LAYER met5 ;
        RECT 736.730 192.615 933.270 197.865 ;
        RECT 775.000 191.015 895.000 192.615 ;
        RECT 736.730 186.565 933.270 191.015 ;
      LAYER met5 ;
        RECT 934.870 184.965 1009.130 197.865 ;
      LAYER met5 ;
        RECT 1010.730 192.615 1207.270 197.865 ;
        RECT 1049.000 191.015 1169.000 192.615 ;
        RECT 1010.730 186.565 1207.270 191.015 ;
      LAYER met5 ;
        RECT 1208.870 184.965 1278.130 197.865 ;
      LAYER met5 ;
        RECT 1279.730 192.615 1476.270 197.865 ;
        RECT 1318.000 191.015 1438.000 192.615 ;
        RECT 1279.730 186.565 1476.270 191.015 ;
      LAYER met5 ;
        RECT 1477.870 184.965 1552.130 197.865 ;
      LAYER met5 ;
        RECT 1553.730 192.615 1750.270 197.865 ;
        RECT 1592.000 191.015 1712.000 192.615 ;
        RECT 1553.730 186.565 1750.270 191.015 ;
      LAYER met5 ;
        RECT 1751.870 184.965 1826.130 197.865 ;
      LAYER met5 ;
        RECT 1827.730 192.615 2024.270 197.865 ;
        RECT 1866.000 191.015 1986.000 192.615 ;
        RECT 1827.730 186.565 2024.270 191.015 ;
      LAYER met5 ;
        RECT 2025.870 184.965 2100.130 197.865 ;
      LAYER met5 ;
        RECT 2101.730 192.615 2298.270 197.865 ;
        RECT 2140.000 191.015 2260.000 192.615 ;
        RECT 2101.730 186.565 2298.270 191.015 ;
      LAYER met5 ;
        RECT 2299.870 184.965 2374.130 197.865 ;
      LAYER met5 ;
        RECT 2375.730 192.615 2572.270 197.865 ;
        RECT 2414.000 191.015 2534.000 192.615 ;
        RECT 2375.730 186.565 2572.270 191.015 ;
      LAYER met5 ;
        RECT 2573.870 184.965 2648.130 197.865 ;
      LAYER met5 ;
        RECT 2649.730 192.615 2846.270 197.865 ;
        RECT 2688.000 191.015 2808.000 192.615 ;
        RECT 2649.730 186.565 2846.270 191.015 ;
      LAYER met5 ;
        RECT 2847.870 184.965 2917.130 197.865 ;
      LAYER met5 ;
        RECT 2918.730 192.615 3115.270 197.865 ;
        RECT 2957.000 191.015 3077.000 192.615 ;
        RECT 2918.730 186.565 3115.270 191.015 ;
      LAYER met5 ;
        RECT 3116.870 184.965 3186.130 197.865 ;
      LAYER met5 ;
        RECT 3187.730 192.615 3385.270 197.865 ;
      LAYER met5 ;
        RECT 3386.870 196.050 3388.535 199.465 ;
      LAYER met5 ;
        RECT 3390.135 197.650 3395.385 501.270 ;
        RECT 3396.985 355.000 3401.435 501.270 ;
        RECT 3403.035 350.000 3406.285 501.030 ;
        RECT 3396.985 196.215 3401.435 350.000 ;
        RECT 3403.035 198.530 3406.285 345.000 ;
        RECT 3407.885 198.475 3412.335 501.270 ;
        RECT 3413.935 198.400 3418.385 501.270 ;
        RECT 3419.985 198.615 3423.235 501.270 ;
        RECT 3424.840 500.000 3428.085 501.270 ;
        RECT 3424.835 350.000 3428.085 500.000 ;
        RECT 3429.685 355.000 3434.135 501.270 ;
        RECT 3435.735 350.000 3444.735 501.270 ;
        RECT 3424.835 198.665 3428.085 345.000 ;
        RECT 3429.685 198.525 3434.135 350.000 ;
      LAYER met5 ;
        RECT 3424.835 197.015 3428.085 197.065 ;
        RECT 3403.035 196.875 3406.285 196.930 ;
        RECT 3419.985 196.925 3428.085 197.015 ;
        RECT 3403.035 196.800 3412.335 196.875 ;
        RECT 3419.985 196.800 3434.135 196.925 ;
        RECT 3386.870 194.615 3395.385 196.050 ;
        RECT 3403.035 194.615 3434.135 196.800 ;
      LAYER met5 ;
        RECT 3226.000 191.015 3346.000 192.615 ;
        RECT 3187.730 186.565 3385.270 191.015 ;
      LAYER met5 ;
        RECT 3386.870 184.965 3434.135 194.615 ;
        RECT 153.865 181.715 196.930 184.965 ;
      LAYER met5 ;
        RECT 198.530 181.715 394.965 184.965 ;
      LAYER met5 ;
        RECT 396.565 181.715 466.435 184.965 ;
      LAYER met5 ;
        RECT 468.035 181.715 663.965 184.965 ;
      LAYER met5 ;
        RECT 665.565 181.715 735.435 184.965 ;
      LAYER met5 ;
        RECT 737.035 181.715 933.030 184.965 ;
      LAYER met5 ;
        RECT 934.630 181.715 1009.435 184.965 ;
      LAYER met5 ;
        RECT 1011.035 181.715 1206.965 184.965 ;
      LAYER met5 ;
        RECT 1208.565 181.715 1278.435 184.965 ;
      LAYER met5 ;
        RECT 1280.035 181.715 1476.030 184.965 ;
      LAYER met5 ;
        RECT 1477.630 181.715 1552.435 184.965 ;
      LAYER met5 ;
        RECT 1554.035 181.715 1750.030 184.965 ;
      LAYER met5 ;
        RECT 1751.630 181.715 1826.435 184.965 ;
      LAYER met5 ;
        RECT 1828.035 181.715 2024.030 184.965 ;
      LAYER met5 ;
        RECT 2025.630 181.715 2100.435 184.965 ;
      LAYER met5 ;
        RECT 2102.035 181.715 2298.030 184.965 ;
      LAYER met5 ;
        RECT 2299.630 181.715 2374.435 184.965 ;
      LAYER met5 ;
        RECT 2376.035 181.715 2572.030 184.965 ;
      LAYER met5 ;
        RECT 2573.630 181.715 2648.435 184.965 ;
      LAYER met5 ;
        RECT 2650.035 181.715 2845.965 184.965 ;
      LAYER met5 ;
        RECT 2847.565 181.715 2917.435 184.965 ;
      LAYER met5 ;
        RECT 2919.035 181.715 3114.965 184.965 ;
      LAYER met5 ;
        RECT 3116.565 181.715 3186.435 184.965 ;
      LAYER met5 ;
        RECT 3188.035 181.715 3385.255 184.965 ;
      LAYER met5 ;
        RECT 3386.855 181.715 3434.135 184.965 ;
        RECT 153.865 175.665 196.875 181.715 ;
      LAYER met5 ;
        RECT 198.475 175.665 395.270 180.115 ;
      LAYER met5 ;
        RECT 153.865 175.245 196.800 175.665 ;
        RECT 0.000 168.015 196.800 175.245 ;
      LAYER met5 ;
        RECT 198.400 169.615 395.270 174.065 ;
      LAYER met5 ;
        RECT 0.000 163.165 197.015 168.015 ;
      LAYER met5 ;
        RECT 198.615 164.765 395.270 168.015 ;
      LAYER met5 ;
        RECT 396.870 163.165 466.130 181.715 ;
      LAYER met5 ;
        RECT 467.730 175.665 664.270 180.115 ;
        RECT 467.730 169.615 664.270 174.065 ;
        RECT 467.730 164.765 664.270 168.015 ;
      LAYER met5 ;
        RECT 0.000 159.915 197.065 163.165 ;
      LAYER met5 ;
        RECT 198.665 163.160 394.000 163.165 ;
      LAYER met5 ;
        RECT 394.000 163.160 469.000 163.165 ;
      LAYER met5 ;
        RECT 469.000 163.160 663.000 163.165 ;
        RECT 198.665 159.915 395.270 163.160 ;
      LAYER met5 ;
        RECT 0.000 153.865 196.925 159.915 ;
      LAYER met5 ;
        RECT 198.525 153.865 395.270 158.315 ;
      LAYER met5 ;
        RECT 0.000 141.665 175.245 153.865 ;
      LAYER met5 ;
        RECT 176.845 143.265 395.270 152.265 ;
      LAYER met5 ;
        RECT 0.000 135.815 196.775 141.665 ;
      LAYER met5 ;
        RECT 198.375 137.415 395.270 141.665 ;
      LAYER met5 ;
        RECT 0.000 131.565 196.920 135.815 ;
      LAYER met5 ;
        RECT 198.520 131.565 395.270 135.815 ;
      LAYER met5 ;
        RECT 0.000 103.415 195.755 131.565 ;
      LAYER met5 ;
        RECT 197.355 105.015 395.270 129.965 ;
      LAYER met5 ;
        RECT 396.870 103.415 466.130 163.160 ;
      LAYER met5 ;
        RECT 467.730 159.915 664.270 163.160 ;
        RECT 467.730 153.865 664.270 158.315 ;
        RECT 467.730 143.265 664.270 152.265 ;
        RECT 467.730 137.415 664.270 141.665 ;
        RECT 467.730 131.565 664.270 135.815 ;
        RECT 467.730 105.015 664.270 129.965 ;
      LAYER met5 ;
        RECT 665.870 103.415 735.130 181.715 ;
      LAYER met5 ;
        RECT 736.730 175.665 933.270 180.115 ;
        RECT 736.730 169.615 933.270 174.065 ;
        RECT 736.730 164.765 933.270 168.015 ;
        RECT 738.000 163.160 932.000 163.165 ;
        RECT 736.730 159.915 933.270 163.160 ;
        RECT 736.730 153.865 933.270 158.315 ;
        RECT 736.730 143.265 933.270 152.265 ;
        RECT 736.730 137.415 933.270 141.665 ;
        RECT 736.730 131.565 933.270 135.815 ;
        RECT 736.730 105.015 933.270 129.965 ;
      LAYER met5 ;
        RECT 934.870 103.415 1009.130 181.715 ;
      LAYER met5 ;
        RECT 1010.730 175.665 1207.270 180.115 ;
        RECT 1010.730 169.615 1207.270 174.065 ;
        RECT 1010.730 164.765 1207.270 168.015 ;
      LAYER met5 ;
        RECT 1208.870 163.165 1278.130 181.715 ;
      LAYER met5 ;
        RECT 1279.730 175.665 1476.270 180.115 ;
        RECT 1279.730 169.615 1476.270 174.065 ;
        RECT 1279.730 164.765 1476.270 168.015 ;
        RECT 1012.000 163.160 1206.000 163.165 ;
      LAYER met5 ;
        RECT 1206.000 163.160 1281.000 163.165 ;
      LAYER met5 ;
        RECT 1281.000 163.160 1475.000 163.165 ;
        RECT 1010.730 159.915 1207.270 163.160 ;
        RECT 1010.730 153.865 1207.270 158.315 ;
        RECT 1010.730 143.265 1207.270 152.265 ;
        RECT 1010.730 137.415 1207.270 141.665 ;
        RECT 1010.730 131.565 1207.270 135.815 ;
        RECT 1010.730 105.015 1207.270 129.965 ;
      LAYER met5 ;
        RECT 1208.870 103.415 1278.130 163.160 ;
      LAYER met5 ;
        RECT 1279.730 159.915 1476.270 163.160 ;
        RECT 1279.730 153.865 1476.270 158.315 ;
        RECT 1279.730 143.265 1476.270 152.265 ;
        RECT 1279.730 137.415 1476.270 141.665 ;
        RECT 1279.730 131.565 1476.270 135.815 ;
        RECT 1279.730 105.015 1476.270 129.965 ;
      LAYER met5 ;
        RECT 1477.870 103.415 1552.130 181.715 ;
      LAYER met5 ;
        RECT 1553.730 175.665 1750.270 180.115 ;
        RECT 1553.730 169.615 1750.270 174.065 ;
        RECT 1553.730 164.765 1750.270 168.015 ;
        RECT 1555.000 163.160 1749.000 163.165 ;
        RECT 1553.730 159.915 1750.270 163.160 ;
        RECT 1553.730 153.865 1750.270 158.315 ;
        RECT 1553.730 143.265 1750.270 152.265 ;
        RECT 1553.730 137.415 1750.270 141.665 ;
        RECT 1553.730 131.565 1750.270 135.815 ;
        RECT 1553.730 105.015 1750.270 129.965 ;
      LAYER met5 ;
        RECT 1751.870 103.415 1826.130 181.715 ;
      LAYER met5 ;
        RECT 1827.730 175.665 2024.270 180.115 ;
        RECT 1827.730 169.615 2024.270 174.065 ;
        RECT 1827.730 164.765 2024.270 168.015 ;
        RECT 1829.000 163.160 2023.000 163.165 ;
        RECT 1827.730 159.915 2024.270 163.160 ;
        RECT 1827.730 153.865 2024.270 158.315 ;
        RECT 1827.730 143.265 2024.270 152.265 ;
        RECT 1827.730 137.415 2024.270 141.665 ;
        RECT 1827.730 131.565 2024.270 135.815 ;
        RECT 1827.730 105.015 2024.270 129.965 ;
      LAYER met5 ;
        RECT 2025.870 103.415 2100.130 181.715 ;
      LAYER met5 ;
        RECT 2101.730 175.665 2298.270 180.115 ;
        RECT 2101.730 169.615 2298.270 174.065 ;
        RECT 2101.730 164.765 2298.270 168.015 ;
        RECT 2103.000 163.160 2297.000 163.165 ;
        RECT 2101.730 159.915 2298.270 163.160 ;
        RECT 2101.730 153.865 2298.270 158.315 ;
        RECT 2101.730 143.265 2298.270 152.265 ;
        RECT 2101.730 137.415 2298.270 141.665 ;
        RECT 2101.730 131.565 2298.270 135.815 ;
        RECT 2101.730 105.015 2298.270 129.965 ;
      LAYER met5 ;
        RECT 2299.870 103.415 2374.130 181.715 ;
      LAYER met5 ;
        RECT 2375.730 175.665 2572.270 180.115 ;
        RECT 2375.730 169.615 2572.270 174.065 ;
        RECT 2375.730 164.765 2572.270 168.015 ;
        RECT 2377.000 163.160 2571.000 163.165 ;
        RECT 2375.730 159.915 2572.270 163.160 ;
        RECT 2375.730 153.865 2572.270 158.315 ;
        RECT 2375.730 143.265 2572.270 152.265 ;
        RECT 2375.730 137.415 2572.270 141.665 ;
        RECT 2375.730 131.565 2572.270 135.815 ;
        RECT 2375.730 105.015 2572.270 129.965 ;
      LAYER met5 ;
        RECT 2573.870 103.415 2648.130 181.715 ;
      LAYER met5 ;
        RECT 2649.730 175.665 2846.270 180.115 ;
        RECT 2649.730 169.615 2846.270 174.065 ;
        RECT 2649.730 164.765 2846.270 168.015 ;
      LAYER met5 ;
        RECT 2847.870 163.165 2917.130 181.715 ;
      LAYER met5 ;
        RECT 2918.730 175.665 3115.270 180.115 ;
        RECT 2918.730 169.615 3115.270 174.065 ;
        RECT 2918.730 164.765 3115.270 168.015 ;
      LAYER met5 ;
        RECT 3116.870 163.165 3186.130 181.715 ;
      LAYER met5 ;
        RECT 3187.730 175.665 3385.270 180.115 ;
      LAYER met5 ;
        RECT 3386.870 175.245 3434.135 181.715 ;
      LAYER met5 ;
        RECT 3435.735 176.845 3444.735 345.000 ;
        RECT 3446.335 198.375 3450.585 501.270 ;
        RECT 3452.185 198.520 3456.435 501.270 ;
        RECT 3458.035 197.355 3482.985 501.270 ;
      LAYER met5 ;
        RECT 3484.585 500.000 3588.000 502.870 ;
      LAYER met5 ;
        RECT 3563.785 200.000 3588.000 500.000 ;
      LAYER met5 ;
        RECT 3452.185 196.775 3456.435 196.920 ;
        RECT 3446.335 195.755 3456.435 196.775 ;
        RECT 3484.585 195.755 3588.000 200.000 ;
        RECT 3446.335 175.245 3588.000 195.755 ;
      LAYER met5 ;
        RECT 3187.730 169.615 3385.270 174.065 ;
        RECT 3187.730 164.765 3385.270 168.015 ;
        RECT 2651.000 163.160 2845.000 163.165 ;
      LAYER met5 ;
        RECT 2845.000 163.160 2920.000 163.165 ;
      LAYER met5 ;
        RECT 2920.000 163.160 3114.000 163.165 ;
      LAYER met5 ;
        RECT 3114.000 163.160 3189.000 163.165 ;
      LAYER met5 ;
        RECT 3189.000 163.160 3384.000 163.165 ;
        RECT 2649.730 159.915 2846.270 163.160 ;
        RECT 2649.730 153.865 2846.270 158.315 ;
        RECT 2649.730 143.265 2846.270 152.265 ;
        RECT 2649.730 137.415 2846.270 141.665 ;
        RECT 2649.730 131.565 2846.270 135.815 ;
        RECT 2649.730 105.015 2846.270 129.965 ;
      LAYER met5 ;
        RECT 2847.870 103.415 2917.130 163.160 ;
      LAYER met5 ;
        RECT 2918.730 159.915 3115.270 163.160 ;
        RECT 2918.730 153.865 3115.270 158.315 ;
        RECT 2918.730 143.265 3115.270 152.265 ;
        RECT 2918.730 137.415 3115.270 141.665 ;
        RECT 2918.730 131.565 3115.270 135.815 ;
        RECT 2918.730 105.015 3115.270 129.965 ;
      LAYER met5 ;
        RECT 3116.870 103.415 3186.130 163.160 ;
      LAYER met5 ;
        RECT 3187.730 159.915 3385.270 163.160 ;
        RECT 3187.730 153.865 3385.270 158.315 ;
      LAYER met5 ;
        RECT 3386.870 153.865 3588.000 175.245 ;
      LAYER met5 ;
        RECT 3187.730 143.265 3411.155 152.265 ;
      LAYER met5 ;
        RECT 3412.755 141.665 3588.000 153.865 ;
      LAYER met5 ;
        RECT 3187.730 137.415 3385.270 141.665 ;
        RECT 3187.730 131.565 3385.270 135.815 ;
      LAYER met5 ;
        RECT 3386.870 131.565 3588.000 141.665 ;
      LAYER met5 ;
        RECT 3187.730 105.015 3385.855 129.965 ;
      LAYER met5 ;
        RECT 3387.455 103.415 3588.000 131.565 ;
        RECT 0.000 0.000 200.000 103.415 ;
        RECT 394.000 96.480 469.000 103.415 ;
        RECT 394.000 32.455 399.510 96.480 ;
        RECT 463.550 32.455 469.000 96.480 ;
      LAYER met5 ;
        RECT 200.000 0.000 394.000 24.215 ;
      LAYER met5 ;
        RECT 394.000 0.000 469.000 32.455 ;
        RECT 663.000 93.145 738.000 103.415 ;
        RECT 663.000 34.115 681.965 93.145 ;
        RECT 722.350 34.115 738.000 93.145 ;
        RECT 663.000 25.815 738.000 34.115 ;
        RECT 932.000 97.040 1012.000 103.415 ;
        RECT 932.000 31.390 936.600 97.040 ;
        RECT 1002.500 31.390 1012.000 97.040 ;
      LAYER met5 ;
        RECT 469.000 0.000 664.270 24.215 ;
      LAYER met5 ;
        RECT 665.870 0.000 735.130 25.815 ;
      LAYER met5 ;
        RECT 736.730 0.000 932.000 24.215 ;
      LAYER met5 ;
        RECT 932.000 0.000 1012.000 31.390 ;
        RECT 1206.000 99.700 1281.000 103.415 ;
        RECT 1206.000 29.235 1214.730 99.700 ;
        RECT 1272.330 29.235 1281.000 99.700 ;
      LAYER met5 ;
        RECT 1012.000 0.000 1206.000 24.215 ;
      LAYER met5 ;
        RECT 1206.000 0.000 1281.000 29.235 ;
        RECT 1475.000 97.040 1555.000 103.415 ;
        RECT 1475.000 31.390 1479.600 97.040 ;
        RECT 1545.500 31.390 1555.000 97.040 ;
      LAYER met5 ;
        RECT 1281.000 0.000 1475.000 24.215 ;
      LAYER met5 ;
        RECT 1475.000 0.000 1555.000 31.390 ;
        RECT 1749.000 97.040 1829.000 103.415 ;
        RECT 1749.000 31.390 1753.600 97.040 ;
        RECT 1819.500 31.390 1829.000 97.040 ;
      LAYER met5 ;
        RECT 1555.000 0.000 1749.000 24.215 ;
      LAYER met5 ;
        RECT 1749.000 0.000 1829.000 31.390 ;
        RECT 2023.000 97.040 2103.000 103.415 ;
        RECT 2023.000 31.390 2027.600 97.040 ;
        RECT 2093.500 31.390 2103.000 97.040 ;
      LAYER met5 ;
        RECT 1829.000 0.000 2023.000 24.215 ;
      LAYER met5 ;
        RECT 2023.000 0.000 2103.000 31.390 ;
        RECT 2297.000 97.040 2377.000 103.415 ;
        RECT 2297.000 31.390 2301.600 97.040 ;
        RECT 2367.500 31.390 2377.000 97.040 ;
      LAYER met5 ;
        RECT 2103.000 0.000 2297.000 24.215 ;
      LAYER met5 ;
        RECT 2297.000 0.000 2377.000 31.390 ;
        RECT 2571.000 97.040 2651.000 103.415 ;
        RECT 2571.000 31.390 2575.600 97.040 ;
        RECT 2641.500 31.390 2651.000 97.040 ;
      LAYER met5 ;
        RECT 2377.000 0.000 2571.000 24.215 ;
      LAYER met5 ;
        RECT 2571.000 0.000 2651.000 31.390 ;
        RECT 2845.000 96.480 2920.000 103.415 ;
        RECT 2845.000 32.455 2850.510 96.480 ;
        RECT 2914.550 32.455 2920.000 96.480 ;
      LAYER met5 ;
        RECT 2651.000 0.000 2845.000 24.215 ;
      LAYER met5 ;
        RECT 2845.000 0.000 2920.000 32.455 ;
        RECT 3114.000 96.480 3189.000 103.415 ;
        RECT 3114.000 32.455 3119.510 96.480 ;
        RECT 3183.550 32.455 3189.000 96.480 ;
      LAYER met5 ;
        RECT 2920.000 0.000 3114.000 24.215 ;
      LAYER met5 ;
        RECT 3114.000 0.000 3189.000 32.455 ;
      LAYER met5 ;
        RECT 3189.000 0.000 3384.000 24.215 ;
      LAYER met5 ;
        RECT 3384.000 0.000 3588.000 103.415 ;
  END
END chip_io
END LIBRARY

