magic
tech sky130A
magscale 1 2
timestamp 1606523612
<< checkpaint >>
rect -1260 -1260 6192 6260
<< locali >>
rect 3937 2052 3971 2610
<< viali >>
rect 1057 2610 1091 2644
rect 2785 2610 2819 2644
rect 3937 2610 3971 2644
rect 289 2240 323 2274
rect 1633 2092 1667 2126
rect 3937 2018 3971 2052
rect 4321 2018 4355 2052
rect 3265 1870 3299 1904
<< metal1 >>
rect 1906 4155 1912 4207
rect 1964 4195 1970 4207
rect 4210 4195 4216 4207
rect 1964 4167 4216 4195
rect 1964 4155 1970 4167
rect 4210 4155 4216 4167
rect 4268 4155 4274 4207
rect 66 4096 4866 4121
rect 66 4044 745 4096
rect 797 4044 809 4096
rect 861 4044 873 4096
rect 925 4044 937 4096
rect 989 4044 2348 4096
rect 2400 4044 2412 4096
rect 2464 4044 2476 4096
rect 2528 4044 2540 4096
rect 2592 4044 3950 4096
rect 4002 4044 4014 4096
rect 4066 4044 4078 4096
rect 4130 4044 4142 4096
rect 4194 4044 4866 4096
rect 66 4019 4866 4044
rect 66 3282 4866 3307
rect 66 3230 1546 3282
rect 1598 3230 1610 3282
rect 1662 3230 1674 3282
rect 1726 3230 1738 3282
rect 1790 3230 3149 3282
rect 3201 3230 3213 3282
rect 3265 3230 3277 3282
rect 3329 3230 3341 3282
rect 3393 3230 4866 3282
rect 66 3205 4866 3230
rect 274 2601 280 2653
rect 332 2641 338 2653
rect 1045 2644 1103 2650
rect 1045 2641 1057 2644
rect 332 2613 1057 2641
rect 332 2601 338 2613
rect 1045 2610 1057 2613
rect 1091 2610 1103 2644
rect 1045 2604 1103 2610
rect 2773 2644 2831 2650
rect 2773 2610 2785 2644
rect 2819 2641 2831 2644
rect 3925 2644 3983 2650
rect 3925 2641 3937 2644
rect 2819 2613 3937 2641
rect 2819 2610 2831 2613
rect 2773 2604 2831 2610
rect 3925 2610 3937 2613
rect 3971 2610 3983 2644
rect 3925 2604 3983 2610
rect 66 2468 4866 2493
rect 66 2416 745 2468
rect 797 2416 809 2468
rect 861 2416 873 2468
rect 925 2416 937 2468
rect 989 2416 2348 2468
rect 2400 2416 2412 2468
rect 2464 2416 2476 2468
rect 2528 2416 2540 2468
rect 2592 2416 3950 2468
rect 4002 2416 4014 2468
rect 4066 2416 4078 2468
rect 4130 2416 4142 2468
rect 4194 2416 4866 2468
rect 66 2391 4866 2416
rect 274 2271 280 2283
rect 235 2243 280 2271
rect 274 2231 280 2243
rect 332 2231 338 2283
rect 1621 2126 1679 2132
rect 1621 2092 1633 2126
rect 1667 2123 1679 2126
rect 1906 2123 1912 2135
rect 1667 2095 1912 2123
rect 1667 2092 1679 2095
rect 1621 2086 1679 2092
rect 1906 2083 1912 2095
rect 1964 2083 1970 2135
rect 3925 2052 3983 2058
rect 3925 2018 3937 2052
rect 3971 2049 3983 2052
rect 4309 2052 4367 2058
rect 4309 2049 4321 2052
rect 3971 2021 4321 2049
rect 3971 2018 3983 2021
rect 3925 2012 3983 2018
rect 4309 2018 4321 2021
rect 4355 2018 4367 2052
rect 4309 2012 4367 2018
rect 562 1861 568 1913
rect 620 1901 626 1913
rect 3253 1904 3311 1910
rect 3253 1901 3265 1904
rect 620 1873 3265 1901
rect 620 1861 626 1873
rect 3253 1870 3265 1873
rect 3299 1870 3311 1904
rect 3253 1864 3311 1870
rect 66 1654 4866 1679
rect 66 1602 1546 1654
rect 1598 1602 1610 1654
rect 1662 1602 1674 1654
rect 1726 1602 1738 1654
rect 1790 1602 3149 1654
rect 3201 1602 3213 1654
rect 3265 1602 3277 1654
rect 3329 1602 3341 1654
rect 3393 1602 4866 1654
rect 66 1577 4866 1602
rect 66 840 4866 865
rect 66 788 745 840
rect 797 788 809 840
rect 861 788 873 840
rect 925 788 937 840
rect 989 788 2348 840
rect 2400 788 2412 840
rect 2464 788 2476 840
rect 2528 788 2540 840
rect 2592 788 3950 840
rect 4002 788 4014 840
rect 4066 788 4078 840
rect 4130 788 4142 840
rect 4194 788 4866 840
rect 66 763 4866 788
<< via1 >>
rect 1912 4155 1964 4207
rect 4216 4155 4268 4207
rect 745 4044 797 4096
rect 809 4044 861 4096
rect 873 4044 925 4096
rect 937 4044 989 4096
rect 2348 4044 2400 4096
rect 2412 4044 2464 4096
rect 2476 4044 2528 4096
rect 2540 4044 2592 4096
rect 3950 4044 4002 4096
rect 4014 4044 4066 4096
rect 4078 4044 4130 4096
rect 4142 4044 4194 4096
rect 1546 3230 1598 3282
rect 1610 3230 1662 3282
rect 1674 3230 1726 3282
rect 1738 3230 1790 3282
rect 3149 3230 3201 3282
rect 3213 3230 3265 3282
rect 3277 3230 3329 3282
rect 3341 3230 3393 3282
rect 280 2601 332 2653
rect 745 2416 797 2468
rect 809 2416 861 2468
rect 873 2416 925 2468
rect 937 2416 989 2468
rect 2348 2416 2400 2468
rect 2412 2416 2464 2468
rect 2476 2416 2528 2468
rect 2540 2416 2592 2468
rect 3950 2416 4002 2468
rect 4014 2416 4066 2468
rect 4078 2416 4130 2468
rect 4142 2416 4194 2468
rect 280 2274 332 2283
rect 280 2240 289 2274
rect 289 2240 323 2274
rect 323 2240 332 2274
rect 280 2231 332 2240
rect 1912 2083 1964 2135
rect 568 1861 620 1913
rect 1546 1602 1598 1654
rect 1610 1602 1662 1654
rect 1674 1602 1726 1654
rect 1738 1602 1790 1654
rect 3149 1602 3201 1654
rect 3213 1602 3265 1654
rect 3277 1602 3329 1654
rect 3341 1602 3393 1654
rect 745 788 797 840
rect 809 788 861 840
rect 873 788 925 840
rect 937 788 989 840
rect 2348 788 2400 840
rect 2412 788 2464 840
rect 2476 788 2528 840
rect 2540 788 2592 840
rect 3950 788 4002 840
rect 4014 788 4066 840
rect 4078 788 4130 840
rect 4142 788 4194 840
<< metal2 >>
rect 1912 4207 1964 4213
rect 4214 4207 4270 5000
rect 4214 4200 4216 4207
rect 1912 4149 1964 4155
rect 4268 4200 4270 4207
rect 4216 4149 4268 4155
rect 719 4098 1015 4121
rect 775 4096 799 4098
rect 855 4096 879 4098
rect 935 4096 959 4098
rect 797 4044 799 4096
rect 861 4044 873 4096
rect 935 4044 937 4096
rect 775 4042 799 4044
rect 855 4042 879 4044
rect 935 4042 959 4044
rect 719 4019 1015 4042
rect 1520 3284 1816 3307
rect 1576 3282 1600 3284
rect 1656 3282 1680 3284
rect 1736 3282 1760 3284
rect 1598 3230 1600 3282
rect 1662 3230 1674 3282
rect 1736 3230 1738 3282
rect 1576 3228 1600 3230
rect 1656 3228 1680 3230
rect 1736 3228 1760 3230
rect 1520 3205 1816 3228
rect 280 2653 332 2659
rect 280 2595 332 2601
rect 292 2289 320 2595
rect 719 2470 1015 2493
rect 775 2468 799 2470
rect 855 2468 879 2470
rect 935 2468 959 2470
rect 797 2416 799 2468
rect 861 2416 873 2468
rect 935 2416 937 2468
rect 775 2414 799 2416
rect 855 2414 879 2416
rect 935 2414 959 2416
rect 719 2391 1015 2414
rect 280 2283 332 2289
rect 280 2225 332 2231
rect 1924 2141 1952 4149
rect 2322 4098 2618 4121
rect 2378 4096 2402 4098
rect 2458 4096 2482 4098
rect 2538 4096 2562 4098
rect 2400 4044 2402 4096
rect 2464 4044 2476 4096
rect 2538 4044 2540 4096
rect 2378 4042 2402 4044
rect 2458 4042 2482 4044
rect 2538 4042 2562 4044
rect 2322 4019 2618 4042
rect 3924 4098 4220 4121
rect 3980 4096 4004 4098
rect 4060 4096 4084 4098
rect 4140 4096 4164 4098
rect 4002 4044 4004 4096
rect 4066 4044 4078 4096
rect 4140 4044 4142 4096
rect 3980 4042 4004 4044
rect 4060 4042 4084 4044
rect 4140 4042 4164 4044
rect 3924 4019 4220 4042
rect 3123 3284 3419 3307
rect 3179 3282 3203 3284
rect 3259 3282 3283 3284
rect 3339 3282 3363 3284
rect 3201 3230 3203 3282
rect 3265 3230 3277 3282
rect 3339 3230 3341 3282
rect 3179 3228 3203 3230
rect 3259 3228 3283 3230
rect 3339 3228 3363 3230
rect 3123 3205 3419 3228
rect 2322 2470 2618 2493
rect 2378 2468 2402 2470
rect 2458 2468 2482 2470
rect 2538 2468 2562 2470
rect 2400 2416 2402 2468
rect 2464 2416 2476 2468
rect 2538 2416 2540 2468
rect 2378 2414 2402 2416
rect 2458 2414 2482 2416
rect 2538 2414 2562 2416
rect 2322 2391 2618 2414
rect 3924 2470 4220 2493
rect 3980 2468 4004 2470
rect 4060 2468 4084 2470
rect 4140 2468 4164 2470
rect 4002 2416 4004 2468
rect 4066 2416 4078 2468
rect 4140 2416 4142 2468
rect 3980 2414 4004 2416
rect 4060 2414 4084 2416
rect 4140 2414 4164 2416
rect 3924 2391 4220 2414
rect 1912 2135 1964 2141
rect 1912 2077 1964 2083
rect 568 1913 620 1919
rect 568 1855 620 1861
rect 580 800 608 1855
rect 1520 1656 1816 1679
rect 1576 1654 1600 1656
rect 1656 1654 1680 1656
rect 1736 1654 1760 1656
rect 1598 1602 1600 1654
rect 1662 1602 1674 1654
rect 1736 1602 1738 1654
rect 1576 1600 1600 1602
rect 1656 1600 1680 1602
rect 1736 1600 1760 1602
rect 1520 1577 1816 1600
rect 3123 1656 3419 1679
rect 3179 1654 3203 1656
rect 3259 1654 3283 1656
rect 3339 1654 3363 1656
rect 3201 1602 3203 1654
rect 3265 1602 3277 1654
rect 3339 1602 3341 1654
rect 3179 1600 3203 1602
rect 3259 1600 3283 1602
rect 3339 1600 3363 1602
rect 3123 1577 3419 1600
rect 719 842 1015 865
rect 775 840 799 842
rect 855 840 879 842
rect 935 840 959 842
rect 566 0 622 800
rect 797 788 799 840
rect 861 788 873 840
rect 935 788 937 840
rect 775 786 799 788
rect 855 786 879 788
rect 935 786 959 788
rect 719 763 1015 786
rect 2322 842 2618 865
rect 2378 840 2402 842
rect 2458 840 2482 842
rect 2538 840 2562 842
rect 2400 788 2402 840
rect 2464 788 2476 840
rect 2538 788 2540 840
rect 2378 786 2402 788
rect 2458 786 2482 788
rect 2538 786 2562 788
rect 2322 763 2618 786
rect 3924 842 4220 865
rect 3980 840 4004 842
rect 4060 840 4084 842
rect 4140 840 4164 842
rect 4002 788 4004 840
rect 4066 788 4078 840
rect 4140 788 4142 840
rect 3980 786 4004 788
rect 4060 786 4084 788
rect 4140 786 4164 788
rect 3924 763 4220 786
<< via2 >>
rect 719 4096 775 4098
rect 799 4096 855 4098
rect 879 4096 935 4098
rect 959 4096 1015 4098
rect 719 4044 745 4096
rect 745 4044 775 4096
rect 799 4044 809 4096
rect 809 4044 855 4096
rect 879 4044 925 4096
rect 925 4044 935 4096
rect 959 4044 989 4096
rect 989 4044 1015 4096
rect 719 4042 775 4044
rect 799 4042 855 4044
rect 879 4042 935 4044
rect 959 4042 1015 4044
rect 1520 3282 1576 3284
rect 1600 3282 1656 3284
rect 1680 3282 1736 3284
rect 1760 3282 1816 3284
rect 1520 3230 1546 3282
rect 1546 3230 1576 3282
rect 1600 3230 1610 3282
rect 1610 3230 1656 3282
rect 1680 3230 1726 3282
rect 1726 3230 1736 3282
rect 1760 3230 1790 3282
rect 1790 3230 1816 3282
rect 1520 3228 1576 3230
rect 1600 3228 1656 3230
rect 1680 3228 1736 3230
rect 1760 3228 1816 3230
rect 719 2468 775 2470
rect 799 2468 855 2470
rect 879 2468 935 2470
rect 959 2468 1015 2470
rect 719 2416 745 2468
rect 745 2416 775 2468
rect 799 2416 809 2468
rect 809 2416 855 2468
rect 879 2416 925 2468
rect 925 2416 935 2468
rect 959 2416 989 2468
rect 989 2416 1015 2468
rect 719 2414 775 2416
rect 799 2414 855 2416
rect 879 2414 935 2416
rect 959 2414 1015 2416
rect 2322 4096 2378 4098
rect 2402 4096 2458 4098
rect 2482 4096 2538 4098
rect 2562 4096 2618 4098
rect 2322 4044 2348 4096
rect 2348 4044 2378 4096
rect 2402 4044 2412 4096
rect 2412 4044 2458 4096
rect 2482 4044 2528 4096
rect 2528 4044 2538 4096
rect 2562 4044 2592 4096
rect 2592 4044 2618 4096
rect 2322 4042 2378 4044
rect 2402 4042 2458 4044
rect 2482 4042 2538 4044
rect 2562 4042 2618 4044
rect 3924 4096 3980 4098
rect 4004 4096 4060 4098
rect 4084 4096 4140 4098
rect 4164 4096 4220 4098
rect 3924 4044 3950 4096
rect 3950 4044 3980 4096
rect 4004 4044 4014 4096
rect 4014 4044 4060 4096
rect 4084 4044 4130 4096
rect 4130 4044 4140 4096
rect 4164 4044 4194 4096
rect 4194 4044 4220 4096
rect 3924 4042 3980 4044
rect 4004 4042 4060 4044
rect 4084 4042 4140 4044
rect 4164 4042 4220 4044
rect 3123 3282 3179 3284
rect 3203 3282 3259 3284
rect 3283 3282 3339 3284
rect 3363 3282 3419 3284
rect 3123 3230 3149 3282
rect 3149 3230 3179 3282
rect 3203 3230 3213 3282
rect 3213 3230 3259 3282
rect 3283 3230 3329 3282
rect 3329 3230 3339 3282
rect 3363 3230 3393 3282
rect 3393 3230 3419 3282
rect 3123 3228 3179 3230
rect 3203 3228 3259 3230
rect 3283 3228 3339 3230
rect 3363 3228 3419 3230
rect 2322 2468 2378 2470
rect 2402 2468 2458 2470
rect 2482 2468 2538 2470
rect 2562 2468 2618 2470
rect 2322 2416 2348 2468
rect 2348 2416 2378 2468
rect 2402 2416 2412 2468
rect 2412 2416 2458 2468
rect 2482 2416 2528 2468
rect 2528 2416 2538 2468
rect 2562 2416 2592 2468
rect 2592 2416 2618 2468
rect 2322 2414 2378 2416
rect 2402 2414 2458 2416
rect 2482 2414 2538 2416
rect 2562 2414 2618 2416
rect 3924 2468 3980 2470
rect 4004 2468 4060 2470
rect 4084 2468 4140 2470
rect 4164 2468 4220 2470
rect 3924 2416 3950 2468
rect 3950 2416 3980 2468
rect 4004 2416 4014 2468
rect 4014 2416 4060 2468
rect 4084 2416 4130 2468
rect 4130 2416 4140 2468
rect 4164 2416 4194 2468
rect 4194 2416 4220 2468
rect 3924 2414 3980 2416
rect 4004 2414 4060 2416
rect 4084 2414 4140 2416
rect 4164 2414 4220 2416
rect 1520 1654 1576 1656
rect 1600 1654 1656 1656
rect 1680 1654 1736 1656
rect 1760 1654 1816 1656
rect 1520 1602 1546 1654
rect 1546 1602 1576 1654
rect 1600 1602 1610 1654
rect 1610 1602 1656 1654
rect 1680 1602 1726 1654
rect 1726 1602 1736 1654
rect 1760 1602 1790 1654
rect 1790 1602 1816 1654
rect 1520 1600 1576 1602
rect 1600 1600 1656 1602
rect 1680 1600 1736 1602
rect 1760 1600 1816 1602
rect 3123 1654 3179 1656
rect 3203 1654 3259 1656
rect 3283 1654 3339 1656
rect 3363 1654 3419 1656
rect 3123 1602 3149 1654
rect 3149 1602 3179 1654
rect 3203 1602 3213 1654
rect 3213 1602 3259 1654
rect 3283 1602 3329 1654
rect 3329 1602 3339 1654
rect 3363 1602 3393 1654
rect 3393 1602 3419 1654
rect 3123 1600 3179 1602
rect 3203 1600 3259 1602
rect 3283 1600 3339 1602
rect 3363 1600 3419 1602
rect 719 840 775 842
rect 799 840 855 842
rect 879 840 935 842
rect 959 840 1015 842
rect 719 788 745 840
rect 745 788 775 840
rect 799 788 809 840
rect 809 788 855 840
rect 879 788 925 840
rect 925 788 935 840
rect 959 788 989 840
rect 989 788 1015 840
rect 719 786 775 788
rect 799 786 855 788
rect 879 786 935 788
rect 959 786 1015 788
rect 2322 840 2378 842
rect 2402 840 2458 842
rect 2482 840 2538 842
rect 2562 840 2618 842
rect 2322 788 2348 840
rect 2348 788 2378 840
rect 2402 788 2412 840
rect 2412 788 2458 840
rect 2482 788 2528 840
rect 2528 788 2538 840
rect 2562 788 2592 840
rect 2592 788 2618 840
rect 2322 786 2378 788
rect 2402 786 2458 788
rect 2482 786 2538 788
rect 2562 786 2618 788
rect 3924 840 3980 842
rect 4004 840 4060 842
rect 4084 840 4140 842
rect 4164 840 4220 842
rect 3924 788 3950 840
rect 3950 788 3980 840
rect 4004 788 4014 840
rect 4014 788 4060 840
rect 4084 788 4130 840
rect 4130 788 4140 840
rect 4164 788 4194 840
rect 4194 788 4220 840
rect 3924 786 3980 788
rect 4004 786 4060 788
rect 4084 786 4140 788
rect 4164 786 4220 788
<< metal3 >>
rect 707 4102 1027 4103
rect 707 4038 715 4102
rect 779 4038 795 4102
rect 859 4038 875 4102
rect 939 4038 955 4102
rect 1019 4038 1027 4102
rect 707 4037 1027 4038
rect 2310 4102 2630 4103
rect 2310 4038 2318 4102
rect 2382 4038 2398 4102
rect 2462 4038 2478 4102
rect 2542 4038 2558 4102
rect 2622 4038 2630 4102
rect 2310 4037 2630 4038
rect 3912 4102 4232 4103
rect 3912 4038 3920 4102
rect 3984 4038 4000 4102
rect 4064 4038 4080 4102
rect 4144 4038 4160 4102
rect 4224 4038 4232 4102
rect 3912 4037 4232 4038
rect 1508 3288 1828 3289
rect 1508 3224 1516 3288
rect 1580 3224 1596 3288
rect 1660 3224 1676 3288
rect 1740 3224 1756 3288
rect 1820 3224 1828 3288
rect 1508 3223 1828 3224
rect 3111 3288 3431 3289
rect 3111 3224 3119 3288
rect 3183 3224 3199 3288
rect 3263 3224 3279 3288
rect 3343 3224 3359 3288
rect 3423 3224 3431 3288
rect 3111 3223 3431 3224
rect 707 2474 1027 2475
rect 707 2410 715 2474
rect 779 2410 795 2474
rect 859 2410 875 2474
rect 939 2410 955 2474
rect 1019 2410 1027 2474
rect 707 2409 1027 2410
rect 2310 2474 2630 2475
rect 2310 2410 2318 2474
rect 2382 2410 2398 2474
rect 2462 2410 2478 2474
rect 2542 2410 2558 2474
rect 2622 2410 2630 2474
rect 2310 2409 2630 2410
rect 3912 2474 4232 2475
rect 3912 2410 3920 2474
rect 3984 2410 4000 2474
rect 4064 2410 4080 2474
rect 4144 2410 4160 2474
rect 4224 2410 4232 2474
rect 3912 2409 4232 2410
rect 1508 1660 1828 1661
rect 1508 1596 1516 1660
rect 1580 1596 1596 1660
rect 1660 1596 1676 1660
rect 1740 1596 1756 1660
rect 1820 1596 1828 1660
rect 1508 1595 1828 1596
rect 3111 1660 3431 1661
rect 3111 1596 3119 1660
rect 3183 1596 3199 1660
rect 3263 1596 3279 1660
rect 3343 1596 3359 1660
rect 3423 1596 3431 1660
rect 3111 1595 3431 1596
rect 707 846 1027 847
rect 707 782 715 846
rect 779 782 795 846
rect 859 782 875 846
rect 939 782 955 846
rect 1019 782 1027 846
rect 707 781 1027 782
rect 2310 846 2630 847
rect 2310 782 2318 846
rect 2382 782 2398 846
rect 2462 782 2478 846
rect 2542 782 2558 846
rect 2622 782 2630 846
rect 2310 781 2630 782
rect 3912 846 4232 847
rect 3912 782 3920 846
rect 3984 782 4000 846
rect 4064 782 4080 846
rect 4144 782 4160 846
rect 4224 782 4232 846
rect 3912 781 4232 782
<< via3 >>
rect 715 4098 779 4102
rect 715 4042 719 4098
rect 719 4042 775 4098
rect 775 4042 779 4098
rect 715 4038 779 4042
rect 795 4098 859 4102
rect 795 4042 799 4098
rect 799 4042 855 4098
rect 855 4042 859 4098
rect 795 4038 859 4042
rect 875 4098 939 4102
rect 875 4042 879 4098
rect 879 4042 935 4098
rect 935 4042 939 4098
rect 875 4038 939 4042
rect 955 4098 1019 4102
rect 955 4042 959 4098
rect 959 4042 1015 4098
rect 1015 4042 1019 4098
rect 955 4038 1019 4042
rect 2318 4098 2382 4102
rect 2318 4042 2322 4098
rect 2322 4042 2378 4098
rect 2378 4042 2382 4098
rect 2318 4038 2382 4042
rect 2398 4098 2462 4102
rect 2398 4042 2402 4098
rect 2402 4042 2458 4098
rect 2458 4042 2462 4098
rect 2398 4038 2462 4042
rect 2478 4098 2542 4102
rect 2478 4042 2482 4098
rect 2482 4042 2538 4098
rect 2538 4042 2542 4098
rect 2478 4038 2542 4042
rect 2558 4098 2622 4102
rect 2558 4042 2562 4098
rect 2562 4042 2618 4098
rect 2618 4042 2622 4098
rect 2558 4038 2622 4042
rect 3920 4098 3984 4102
rect 3920 4042 3924 4098
rect 3924 4042 3980 4098
rect 3980 4042 3984 4098
rect 3920 4038 3984 4042
rect 4000 4098 4064 4102
rect 4000 4042 4004 4098
rect 4004 4042 4060 4098
rect 4060 4042 4064 4098
rect 4000 4038 4064 4042
rect 4080 4098 4144 4102
rect 4080 4042 4084 4098
rect 4084 4042 4140 4098
rect 4140 4042 4144 4098
rect 4080 4038 4144 4042
rect 4160 4098 4224 4102
rect 4160 4042 4164 4098
rect 4164 4042 4220 4098
rect 4220 4042 4224 4098
rect 4160 4038 4224 4042
rect 1516 3284 1580 3288
rect 1516 3228 1520 3284
rect 1520 3228 1576 3284
rect 1576 3228 1580 3284
rect 1516 3224 1580 3228
rect 1596 3284 1660 3288
rect 1596 3228 1600 3284
rect 1600 3228 1656 3284
rect 1656 3228 1660 3284
rect 1596 3224 1660 3228
rect 1676 3284 1740 3288
rect 1676 3228 1680 3284
rect 1680 3228 1736 3284
rect 1736 3228 1740 3284
rect 1676 3224 1740 3228
rect 1756 3284 1820 3288
rect 1756 3228 1760 3284
rect 1760 3228 1816 3284
rect 1816 3228 1820 3284
rect 1756 3224 1820 3228
rect 3119 3284 3183 3288
rect 3119 3228 3123 3284
rect 3123 3228 3179 3284
rect 3179 3228 3183 3284
rect 3119 3224 3183 3228
rect 3199 3284 3263 3288
rect 3199 3228 3203 3284
rect 3203 3228 3259 3284
rect 3259 3228 3263 3284
rect 3199 3224 3263 3228
rect 3279 3284 3343 3288
rect 3279 3228 3283 3284
rect 3283 3228 3339 3284
rect 3339 3228 3343 3284
rect 3279 3224 3343 3228
rect 3359 3284 3423 3288
rect 3359 3228 3363 3284
rect 3363 3228 3419 3284
rect 3419 3228 3423 3284
rect 3359 3224 3423 3228
rect 715 2470 779 2474
rect 715 2414 719 2470
rect 719 2414 775 2470
rect 775 2414 779 2470
rect 715 2410 779 2414
rect 795 2470 859 2474
rect 795 2414 799 2470
rect 799 2414 855 2470
rect 855 2414 859 2470
rect 795 2410 859 2414
rect 875 2470 939 2474
rect 875 2414 879 2470
rect 879 2414 935 2470
rect 935 2414 939 2470
rect 875 2410 939 2414
rect 955 2470 1019 2474
rect 955 2414 959 2470
rect 959 2414 1015 2470
rect 1015 2414 1019 2470
rect 955 2410 1019 2414
rect 2318 2470 2382 2474
rect 2318 2414 2322 2470
rect 2322 2414 2378 2470
rect 2378 2414 2382 2470
rect 2318 2410 2382 2414
rect 2398 2470 2462 2474
rect 2398 2414 2402 2470
rect 2402 2414 2458 2470
rect 2458 2414 2462 2470
rect 2398 2410 2462 2414
rect 2478 2470 2542 2474
rect 2478 2414 2482 2470
rect 2482 2414 2538 2470
rect 2538 2414 2542 2470
rect 2478 2410 2542 2414
rect 2558 2470 2622 2474
rect 2558 2414 2562 2470
rect 2562 2414 2618 2470
rect 2618 2414 2622 2470
rect 2558 2410 2622 2414
rect 3920 2470 3984 2474
rect 3920 2414 3924 2470
rect 3924 2414 3980 2470
rect 3980 2414 3984 2470
rect 3920 2410 3984 2414
rect 4000 2470 4064 2474
rect 4000 2414 4004 2470
rect 4004 2414 4060 2470
rect 4060 2414 4064 2470
rect 4000 2410 4064 2414
rect 4080 2470 4144 2474
rect 4080 2414 4084 2470
rect 4084 2414 4140 2470
rect 4140 2414 4144 2470
rect 4080 2410 4144 2414
rect 4160 2470 4224 2474
rect 4160 2414 4164 2470
rect 4164 2414 4220 2470
rect 4220 2414 4224 2470
rect 4160 2410 4224 2414
rect 1516 1656 1580 1660
rect 1516 1600 1520 1656
rect 1520 1600 1576 1656
rect 1576 1600 1580 1656
rect 1516 1596 1580 1600
rect 1596 1656 1660 1660
rect 1596 1600 1600 1656
rect 1600 1600 1656 1656
rect 1656 1600 1660 1656
rect 1596 1596 1660 1600
rect 1676 1656 1740 1660
rect 1676 1600 1680 1656
rect 1680 1600 1736 1656
rect 1736 1600 1740 1656
rect 1676 1596 1740 1600
rect 1756 1656 1820 1660
rect 1756 1600 1760 1656
rect 1760 1600 1816 1656
rect 1816 1600 1820 1656
rect 1756 1596 1820 1600
rect 3119 1656 3183 1660
rect 3119 1600 3123 1656
rect 3123 1600 3179 1656
rect 3179 1600 3183 1656
rect 3119 1596 3183 1600
rect 3199 1656 3263 1660
rect 3199 1600 3203 1656
rect 3203 1600 3259 1656
rect 3259 1600 3263 1656
rect 3199 1596 3263 1600
rect 3279 1656 3343 1660
rect 3279 1600 3283 1656
rect 3283 1600 3339 1656
rect 3339 1600 3343 1656
rect 3279 1596 3343 1600
rect 3359 1656 3423 1660
rect 3359 1600 3363 1656
rect 3363 1600 3419 1656
rect 3419 1600 3423 1656
rect 3359 1596 3423 1600
rect 715 842 779 846
rect 715 786 719 842
rect 719 786 775 842
rect 775 786 779 842
rect 715 782 779 786
rect 795 842 859 846
rect 795 786 799 842
rect 799 786 855 842
rect 855 786 859 842
rect 795 782 859 786
rect 875 842 939 846
rect 875 786 879 842
rect 879 786 935 842
rect 935 786 939 842
rect 875 782 939 786
rect 955 842 1019 846
rect 955 786 959 842
rect 959 786 1015 842
rect 1015 786 1019 842
rect 955 782 1019 786
rect 2318 842 2382 846
rect 2318 786 2322 842
rect 2322 786 2378 842
rect 2378 786 2382 842
rect 2318 782 2382 786
rect 2398 842 2462 846
rect 2398 786 2402 842
rect 2402 786 2458 842
rect 2458 786 2462 842
rect 2398 782 2462 786
rect 2478 842 2542 846
rect 2478 786 2482 842
rect 2482 786 2538 842
rect 2538 786 2542 842
rect 2478 782 2542 786
rect 2558 842 2622 846
rect 2558 786 2562 842
rect 2562 786 2618 842
rect 2618 786 2622 842
rect 2558 782 2622 786
rect 3920 842 3984 846
rect 3920 786 3924 842
rect 3924 786 3980 842
rect 3980 786 3984 842
rect 3920 782 3984 786
rect 4000 842 4064 846
rect 4000 786 4004 842
rect 4004 786 4060 842
rect 4060 786 4064 842
rect 4000 782 4064 786
rect 4080 842 4144 846
rect 4080 786 4084 842
rect 4084 786 4140 842
rect 4140 786 4144 842
rect 4080 782 4144 786
rect 4160 842 4224 846
rect 4160 786 4164 842
rect 4164 786 4220 842
rect 4220 786 4224 842
rect 4160 782 4224 786
<< metal4 >>
rect 707 4102 1027 4121
rect 707 4038 715 4102
rect 779 4038 795 4102
rect 859 4038 875 4102
rect 939 4038 955 4102
rect 1019 4038 1027 4102
rect 707 3691 1027 4038
rect 707 3455 749 3691
rect 985 3455 1027 3691
rect 707 2567 1027 3455
rect 707 2474 749 2567
rect 985 2474 1027 2567
rect 707 2410 715 2474
rect 1019 2410 1027 2474
rect 707 2331 749 2410
rect 985 2331 1027 2410
rect 707 1443 1027 2331
rect 707 1207 749 1443
rect 985 1207 1027 1443
rect 707 846 1027 1207
rect 707 782 715 846
rect 779 782 795 846
rect 859 782 875 846
rect 939 782 955 846
rect 1019 782 1027 846
rect 707 763 1027 782
rect 1508 3288 1828 4121
rect 1508 3224 1516 3288
rect 1580 3224 1596 3288
rect 1660 3224 1676 3288
rect 1740 3224 1756 3288
rect 1820 3224 1828 3288
rect 1508 3129 1828 3224
rect 1508 2893 1550 3129
rect 1786 2893 1828 3129
rect 1508 2005 1828 2893
rect 1508 1769 1550 2005
rect 1786 1769 1828 2005
rect 1508 1660 1828 1769
rect 1508 1596 1516 1660
rect 1580 1596 1596 1660
rect 1660 1596 1676 1660
rect 1740 1596 1756 1660
rect 1820 1596 1828 1660
rect 1508 763 1828 1596
rect 2310 4102 2630 4121
rect 2310 4038 2318 4102
rect 2382 4038 2398 4102
rect 2462 4038 2478 4102
rect 2542 4038 2558 4102
rect 2622 4038 2630 4102
rect 2310 3691 2630 4038
rect 2310 3455 2352 3691
rect 2588 3455 2630 3691
rect 2310 2567 2630 3455
rect 2310 2474 2352 2567
rect 2588 2474 2630 2567
rect 2310 2410 2318 2474
rect 2622 2410 2630 2474
rect 2310 2331 2352 2410
rect 2588 2331 2630 2410
rect 2310 1443 2630 2331
rect 2310 1207 2352 1443
rect 2588 1207 2630 1443
rect 2310 846 2630 1207
rect 2310 782 2318 846
rect 2382 782 2398 846
rect 2462 782 2478 846
rect 2542 782 2558 846
rect 2622 782 2630 846
rect 2310 763 2630 782
rect 3111 3288 3431 4121
rect 3111 3224 3119 3288
rect 3183 3224 3199 3288
rect 3263 3224 3279 3288
rect 3343 3224 3359 3288
rect 3423 3224 3431 3288
rect 3111 3129 3431 3224
rect 3111 2893 3153 3129
rect 3389 2893 3431 3129
rect 3111 2005 3431 2893
rect 3111 1769 3153 2005
rect 3389 1769 3431 2005
rect 3111 1660 3431 1769
rect 3111 1596 3119 1660
rect 3183 1596 3199 1660
rect 3263 1596 3279 1660
rect 3343 1596 3359 1660
rect 3423 1596 3431 1660
rect 3111 763 3431 1596
rect 3912 4102 4232 4121
rect 3912 4038 3920 4102
rect 3984 4038 4000 4102
rect 4064 4038 4080 4102
rect 4144 4038 4160 4102
rect 4224 4038 4232 4102
rect 3912 3691 4232 4038
rect 3912 3455 3954 3691
rect 4190 3455 4232 3691
rect 3912 2567 4232 3455
rect 3912 2474 3954 2567
rect 4190 2474 4232 2567
rect 3912 2410 3920 2474
rect 4224 2410 4232 2474
rect 3912 2331 3954 2410
rect 4190 2331 4232 2410
rect 3912 1443 4232 2331
rect 3912 1207 3954 1443
rect 4190 1207 4232 1443
rect 3912 846 4232 1207
rect 3912 782 3920 846
rect 3984 782 4000 846
rect 4064 782 4080 846
rect 4144 782 4160 846
rect 4224 782 4232 846
rect 3912 763 4232 782
<< via4 >>
rect 749 3455 985 3691
rect 749 2474 985 2567
rect 749 2410 779 2474
rect 779 2410 795 2474
rect 795 2410 859 2474
rect 859 2410 875 2474
rect 875 2410 939 2474
rect 939 2410 955 2474
rect 955 2410 985 2474
rect 749 2331 985 2410
rect 749 1207 985 1443
rect 1550 2893 1786 3129
rect 1550 1769 1786 2005
rect 2352 3455 2588 3691
rect 2352 2474 2588 2567
rect 2352 2410 2382 2474
rect 2382 2410 2398 2474
rect 2398 2410 2462 2474
rect 2462 2410 2478 2474
rect 2478 2410 2542 2474
rect 2542 2410 2558 2474
rect 2558 2410 2588 2474
rect 2352 2331 2588 2410
rect 2352 1207 2588 1443
rect 3153 2893 3389 3129
rect 3153 1769 3389 2005
rect 3954 3455 4190 3691
rect 3954 2474 4190 2567
rect 3954 2410 3984 2474
rect 3984 2410 4000 2474
rect 4000 2410 4064 2474
rect 4064 2410 4080 2474
rect 4080 2410 4144 2474
rect 4144 2410 4160 2474
rect 4160 2410 4190 2474
rect 3954 2331 4190 2410
rect 3954 1207 4190 1443
<< metal5 >>
rect 66 3691 4866 3733
rect 66 3455 749 3691
rect 985 3455 2352 3691
rect 2588 3455 3954 3691
rect 4190 3455 4866 3691
rect 66 3413 4866 3455
rect 66 3129 4866 3171
rect 66 2893 1550 3129
rect 1786 2893 3153 3129
rect 3389 2893 4866 3129
rect 66 2851 4866 2893
rect 66 2567 4866 2609
rect 66 2331 749 2567
rect 985 2331 2352 2567
rect 2588 2331 3954 2567
rect 4190 2331 4866 2567
rect 66 2289 4866 2331
rect 66 2005 4866 2047
rect 66 1769 1550 2005
rect 1786 1769 3153 2005
rect 3389 1769 4866 2005
rect 66 1727 4866 1769
rect 66 1443 4866 1485
rect 66 1207 749 1443
rect 985 1207 2352 1443
rect 2588 1207 3954 1443
rect 4190 1207 4866 1443
rect 66 1165 4866 1207
use sky130_fd_sc_hvl__decap_8  FILLER_3_40
timestamp 1606523612
transform 1 0 3906 0 1 3256
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_2  FILLER_3_48
timestamp 1606523612
transform 1 0 4674 0 1 3256
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_24
timestamp 1606523612
transform 1 0 2370 0 1 3256
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_32
timestamp 1606523612
transform 1 0 3138 0 1 3256
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_0
timestamp 1606523612
transform 1 0 66 0 1 3256
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_8
timestamp 1606523612
transform 1 0 834 0 1 3256
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_3_16
timestamp 1606523612
transform 1 0 1602 0 1 3256
box -66 -23 834 897
use sky130_fd_sc_hvl__conb_1  mprj_logic_high_hvl
timestamp 1606523612
transform 1 0 4194 0 1 1628
box -66 -23 546 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_40
timestamp 1606523612
transform 1 0 3906 0 -1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_48
timestamp 1606523612
transform 1 0 4674 0 -1 1628
box -66 -23 258 897
use sky130_fd_sc_hvl__fill_2  FILLER_1_48
timestamp 1606523612
transform 1 0 4674 0 1 1628
box -66 -23 258 897
use sky130_fd_sc_hvl__decap_4  FILLER_2_43
timestamp 1606523612
transform 1 0 4194 0 -1 3256
box -66 -23 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_2_47
timestamp 1606523612
transform 1 0 4578 0 -1 3256
box -66 -23 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_49
timestamp 1606523612
transform 1 0 4770 0 -1 3256
box -66 -23 162 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  mprj_logic_high_lv
timestamp 1606523612
transform 1 0 2562 0 1 1628
box -66 -23 1698 1651
use sky130_fd_sc_hvl__decap_8  FILLER_0_24
timestamp 1606523612
transform 1 0 2370 0 -1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_32
timestamp 1606523612
transform 1 0 3138 0 -1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__conb_1  mprj2_logic_high_hvl
timestamp 1606523612
transform 1 0 66 0 1 1628
box -66 -23 546 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  mprj2_logic_high_lv
timestamp 1606523612
transform 1 0 930 0 1 1628
box -66 -23 1698 1651
use sky130_fd_sc_hvl__decap_8  FILLER_0_0
timestamp 1606523612
transform 1 0 66 0 -1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_8
timestamp 1606523612
transform 1 0 834 0 -1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_16
timestamp 1606523612
transform 1 0 1602 0 -1 1628
box -66 -23 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_5
timestamp 1606523612
transform 1 0 546 0 1 1628
box -66 -23 450 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_0
timestamp 1606523612
transform 1 0 66 0 -1 3256
box -66 -23 834 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_8
timestamp 1606523612
transform 1 0 834 0 -1 3256
box -66 -23 162 897
<< labels >>
rlabel metal2 s 4214 4200 4270 5000 4 mprj2_vdd_logic1
port 1 nsew
rlabel metal2 s 566 0 622 800 4 mprj_vdd_logic1
port 2 nsew
rlabel metal1 s 66 4019 4866 4121 4 VPWR
port 3 nsew
rlabel metal1 s 66 3205 4866 3307 4 VGND
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 4932 5000
<< end >>
