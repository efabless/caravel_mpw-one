magic
tech sky130A
magscale 1 2
timestamp 1609274408
<< obsli1 >>
rect 76168 997646 92232 1037541
rect 127568 997646 143632 1037541
rect 178968 997646 195032 1037541
rect 230368 997646 246432 1037541
rect 281968 997646 298032 1037541
rect 333614 998007 347955 1037539
rect 335813 997978 336009 998007
rect 347352 997978 347530 998007
rect 335813 997800 347530 997978
rect 383768 997646 399832 1037541
rect 472768 997646 488832 1037541
rect 524168 997646 540232 1037541
rect 575814 998007 590155 1037539
rect 578013 997978 578209 998007
rect 589552 997978 589730 998007
rect 578013 997800 589730 997978
rect 625968 997646 642032 1037541
rect 59 954168 39954 970232
rect 677646 951568 717541 967632
rect 44 912048 39396 926951
rect 678204 907649 717556 922552
rect 61 883936 39593 884371
rect 61 883746 39806 883936
rect 61 872409 39593 883746
rect 39616 872409 39806 883746
rect 61 872207 39806 872409
rect 61 872031 39593 872207
rect 61 869922 39787 872031
rect 677646 862368 717541 878432
rect 61 841730 39593 842155
rect 61 841552 39800 841730
rect 61 830209 39593 841552
rect 39622 830209 39800 841552
rect 677813 831169 717539 833278
rect 678007 830993 717539 831169
rect 61 830013 39800 830209
rect 677794 830791 717539 830993
rect 61 827814 39593 830013
rect 677794 819454 677984 830791
rect 678007 819454 717539 830791
rect 677794 819264 717539 819454
rect 678007 818829 717539 819264
rect 59 784368 39954 800432
rect 677646 773168 717541 789232
rect 59 741168 39954 757232
rect 677646 728168 717541 744232
rect 59 697968 39954 714032
rect 677646 683168 717541 699232
rect 59 654768 39954 670832
rect 677646 637968 717541 654032
rect 59 611568 39954 627632
rect 677646 592968 717541 609032
rect 59 568368 39954 584432
rect 677646 547768 717541 563832
rect 59 525168 39954 541232
rect 677813 516569 717539 518678
rect 678007 516393 717539 516569
rect 677794 516191 717539 516393
rect 677794 504854 677984 516191
rect 678007 504854 717539 516191
rect 677794 504664 717539 504854
rect 678007 504229 717539 504664
rect 61 497136 39593 497571
rect 61 496946 39806 497136
rect 61 485609 39593 496946
rect 39616 485609 39806 496946
rect 61 485407 39806 485609
rect 61 485231 39593 485407
rect 61 483122 39787 485231
rect 678204 459849 717556 474752
rect 44 440848 39396 455751
rect 678007 428187 717539 430386
rect 677800 427991 717539 428187
rect 677800 416648 677978 427991
rect 678007 416648 717539 427991
rect 677800 416470 717539 416648
rect 678007 416045 717539 416470
rect 59 397568 39954 413632
rect 677646 370568 717541 386632
rect 59 354368 39954 370432
rect 59 311168 39954 327232
rect 677646 325368 717541 341432
rect 59 267968 39954 284032
rect 677646 280368 717541 296432
rect 59 224768 39954 240832
rect 677646 235368 717541 251432
rect 59 181568 39954 197632
rect 677646 190168 717541 206232
rect 677646 145168 717541 161232
rect 61 124336 39593 124771
rect 61 124146 39806 124336
rect 61 112809 39593 124146
rect 39616 112809 39806 124146
rect 61 112607 39806 112809
rect 61 112431 39593 112607
rect 61 110322 39787 112431
rect 677646 99968 717541 116032
rect 44 68048 39396 82951
rect 79670 39622 91387 39800
rect 79670 39593 79848 39622
rect 91191 39593 91387 39622
rect 79245 61 93586 39593
rect 132600 156 147600 39963
rect 186368 59 202432 39954
rect 241249 44 256152 39396
rect 294968 59 311032 39954
rect 349768 59 365832 39954
rect 404568 59 420632 39954
rect 459368 59 475432 39954
rect 514168 59 530232 39954
rect 569870 39622 581587 39800
rect 569870 39593 570048 39622
rect 581391 39593 581587 39622
rect 623664 39616 635393 39806
rect 623664 39593 623854 39616
rect 635191 39593 635393 39616
rect 635569 39593 637678 39787
rect 569445 61 583786 39593
rect 623229 61 637678 39593
<< metal1 >>
rect 585042 992196 585048 992248
rect 585100 992236 585106 992248
rect 674742 992236 674748 992248
rect 585100 992208 674748 992236
rect 585100 992196 585106 992208
rect 674742 992196 674748 992208
rect 674800 992196 674806 992248
rect 78858 990768 78864 990820
rect 78916 990808 78922 990820
rect 130286 990808 130292 990820
rect 78916 990780 130292 990808
rect 78916 990768 78922 990780
rect 130286 990768 130292 990780
rect 130344 990768 130350 990820
rect 233050 990808 233056 990820
rect 194704 990780 233056 990808
rect 89990 990700 89996 990752
rect 90048 990740 90054 990752
rect 141418 990740 141424 990752
rect 90048 990712 141424 990740
rect 90048 990700 90054 990712
rect 141418 990700 141424 990712
rect 141476 990740 141482 990752
rect 192846 990740 192852 990752
rect 141476 990712 192852 990740
rect 141476 990700 141482 990712
rect 192846 990700 192852 990712
rect 192904 990700 192910 990752
rect 130286 990632 130292 990684
rect 130344 990672 130350 990684
rect 181714 990672 181720 990684
rect 130344 990644 181720 990672
rect 130344 990632 130350 990644
rect 181714 990632 181720 990644
rect 181772 990672 181778 990684
rect 194704 990672 194732 990780
rect 233050 990768 233056 990780
rect 233108 990808 233114 990820
rect 284662 990808 284668 990820
rect 233108 990780 284668 990808
rect 233108 990768 233114 990780
rect 284662 990768 284668 990780
rect 284720 990808 284726 990820
rect 286962 990808 286968 990820
rect 284720 990780 286968 990808
rect 284720 990768 284726 990780
rect 286962 990768 286968 990780
rect 287020 990768 287026 990820
rect 345106 990768 345112 990820
rect 345164 990808 345170 990820
rect 372522 990808 372528 990820
rect 345164 990780 372528 990808
rect 345164 990768 345170 990780
rect 372522 990768 372528 990780
rect 372580 990768 372586 990820
rect 372614 990768 372620 990820
rect 372672 990808 372678 990820
rect 372672 990780 383608 990808
rect 372672 990768 372678 990780
rect 194962 990700 194968 990752
rect 195020 990740 195026 990752
rect 244182 990740 244188 990752
rect 195020 990712 244188 990740
rect 195020 990700 195026 990712
rect 244182 990700 244188 990712
rect 244240 990740 244246 990752
rect 295794 990740 295800 990752
rect 244240 990712 295800 990740
rect 244240 990700 244246 990712
rect 295794 990700 295800 990712
rect 295852 990700 295858 990752
rect 233694 990672 233700 990684
rect 181772 990644 194732 990672
rect 195072 990644 233700 990672
rect 181772 990632 181778 990644
rect 121270 990604 121276 990616
rect 102060 990576 121276 990604
rect 102060 990536 102088 990576
rect 121270 990564 121276 990576
rect 121328 990564 121334 990616
rect 96540 990508 102088 990536
rect 96540 990264 96568 990508
rect 160186 990428 160192 990480
rect 160244 990468 160250 990480
rect 160244 990440 173940 990468
rect 160244 990428 160250 990440
rect 173912 990412 173940 990440
rect 192846 990428 192852 990480
rect 192904 990468 192910 990480
rect 194962 990468 194968 990480
rect 192904 990440 194968 990468
rect 192904 990428 192910 990440
rect 194962 990428 194968 990440
rect 195020 990428 195026 990480
rect 173894 990360 173900 990412
rect 173952 990360 173958 990412
rect 182450 990360 182456 990412
rect 182508 990400 182514 990412
rect 195072 990400 195100 990644
rect 233694 990632 233700 990644
rect 233752 990672 233758 990684
rect 285306 990672 285312 990684
rect 233752 990644 285312 990672
rect 233752 990632 233758 990644
rect 285306 990632 285312 990644
rect 285364 990672 285370 990684
rect 342162 990672 342168 990684
rect 285364 990644 342168 990672
rect 285364 990632 285370 990644
rect 342162 990632 342168 990644
rect 342220 990672 342226 990684
rect 345014 990672 345020 990684
rect 342220 990644 345020 990672
rect 342220 990632 342226 990644
rect 345014 990632 345020 990644
rect 345072 990632 345078 990684
rect 383580 990672 383608 990780
rect 397454 990768 397460 990820
rect 397512 990808 397518 990820
rect 397638 990808 397644 990820
rect 397512 990780 397644 990808
rect 397512 990768 397518 990780
rect 397638 990768 397644 990780
rect 397696 990808 397702 990820
rect 486602 990808 486608 990820
rect 397696 990780 486608 990808
rect 397696 990768 397702 990780
rect 486602 990768 486608 990780
rect 486660 990808 486666 990820
rect 538030 990808 538036 990820
rect 486660 990780 538036 990808
rect 486660 990768 486666 990780
rect 538030 990768 538036 990780
rect 538088 990808 538094 990820
rect 639782 990808 639788 990820
rect 538088 990780 639788 990808
rect 538088 990768 538094 990780
rect 639782 990768 639788 990780
rect 639840 990768 639846 990820
rect 400122 990700 400128 990752
rect 400180 990740 400186 990752
rect 419534 990740 419540 990752
rect 400180 990712 419540 990740
rect 400180 990700 400186 990712
rect 419534 990700 419540 990712
rect 419592 990700 419598 990752
rect 438762 990700 438768 990752
rect 438820 990740 438826 990752
rect 458174 990740 458180 990752
rect 438820 990712 458180 990740
rect 438820 990700 438826 990712
rect 458174 990700 458180 990712
rect 458232 990700 458238 990752
rect 477402 990700 477408 990752
rect 477460 990740 477466 990752
rect 527542 990740 527548 990752
rect 477460 990712 527548 990740
rect 477460 990700 477466 990712
rect 527542 990700 527548 990712
rect 527600 990740 527606 990752
rect 629294 990740 629300 990752
rect 527600 990712 629300 990740
rect 527600 990700 527606 990712
rect 629294 990700 629300 990712
rect 629352 990740 629358 990752
rect 631226 990740 631232 990752
rect 629352 990712 631232 990740
rect 629352 990700 629358 990712
rect 631226 990700 631232 990712
rect 631284 990700 631290 990752
rect 386414 990672 386420 990684
rect 383580 990644 386420 990672
rect 386414 990632 386420 990644
rect 386472 990632 386478 990684
rect 386506 990632 386512 990684
rect 386564 990672 386570 990684
rect 475470 990672 475476 990684
rect 386564 990644 475476 990672
rect 386564 990632 386570 990644
rect 475470 990632 475476 990644
rect 475528 990672 475534 990684
rect 526898 990672 526904 990684
rect 475528 990644 526904 990672
rect 475528 990632 475534 990644
rect 526898 990632 526904 990644
rect 526956 990672 526962 990684
rect 626534 990672 626540 990684
rect 526956 990644 626540 990672
rect 526956 990632 526962 990644
rect 626534 990632 626540 990644
rect 626592 990632 626598 990684
rect 286962 990564 286968 990616
rect 287020 990604 287026 990616
rect 386524 990604 386552 990632
rect 287020 990576 386552 990604
rect 287020 990564 287026 990576
rect 295794 990496 295800 990548
rect 295852 990536 295858 990548
rect 397454 990536 397460 990548
rect 295852 990508 397460 990536
rect 295852 990496 295858 990508
rect 397454 990496 397460 990508
rect 397512 990496 397518 990548
rect 419534 990496 419540 990548
rect 419592 990536 419598 990548
rect 438762 990536 438768 990548
rect 419592 990508 438768 990536
rect 419592 990496 419598 990508
rect 438762 990496 438768 990508
rect 438820 990496 438826 990548
rect 458174 990496 458180 990548
rect 458232 990536 458238 990548
rect 476114 990536 476120 990548
rect 458232 990508 476120 990536
rect 458232 990496 458238 990508
rect 476114 990496 476120 990508
rect 476172 990536 476178 990548
rect 477402 990536 477408 990548
rect 476172 990508 477408 990536
rect 476172 990496 476178 990508
rect 477402 990496 477408 990508
rect 477460 990496 477466 990548
rect 386414 990428 386420 990480
rect 386472 990468 386478 990480
rect 387150 990468 387156 990480
rect 386472 990440 387156 990468
rect 386472 990428 386478 990440
rect 387150 990428 387156 990440
rect 387208 990468 387214 990480
rect 400122 990468 400128 990480
rect 387208 990440 400128 990468
rect 387208 990428 387214 990440
rect 400122 990428 400128 990440
rect 400180 990428 400186 990480
rect 182508 990372 195100 990400
rect 182508 990360 182514 990372
rect 140682 990332 140688 990344
rect 135272 990304 140688 990332
rect 84396 990236 96568 990264
rect 42242 990156 42248 990208
rect 42300 990196 42306 990208
rect 78858 990196 78864 990208
rect 42300 990168 78864 990196
rect 42300 990156 42306 990168
rect 78858 990156 78864 990168
rect 78916 990156 78922 990208
rect 42334 990088 42340 990140
rect 42392 990128 42398 990140
rect 79502 990128 79508 990140
rect 42392 990100 79508 990128
rect 42392 990088 42398 990100
rect 79502 990088 79508 990100
rect 79560 990128 79566 990140
rect 84396 990128 84424 990236
rect 131022 990224 131028 990276
rect 131080 990264 131086 990276
rect 135272 990264 135300 990304
rect 140682 990292 140688 990304
rect 140740 990292 140746 990344
rect 160002 990332 160008 990344
rect 154500 990304 160008 990332
rect 131080 990236 135300 990264
rect 131080 990224 131086 990236
rect 140774 990224 140780 990276
rect 140832 990264 140838 990276
rect 154500 990264 154528 990304
rect 160002 990292 160008 990304
rect 160060 990292 160066 990344
rect 140832 990236 154528 990264
rect 140832 990224 140838 990236
rect 173894 990224 173900 990276
rect 173952 990264 173958 990276
rect 182468 990264 182496 990360
rect 173952 990236 182496 990264
rect 173952 990224 173958 990236
rect 639782 990156 639788 990208
rect 639840 990196 639846 990208
rect 673638 990196 673644 990208
rect 639840 990168 673644 990196
rect 639840 990156 639846 990168
rect 673638 990156 673644 990168
rect 673696 990156 673702 990208
rect 79560 990100 84424 990128
rect 79560 990088 79566 990100
rect 89898 990088 89904 990140
rect 89956 990088 89962 990140
rect 626534 990088 626540 990140
rect 626592 990088 626598 990140
rect 628650 990088 628656 990140
rect 628708 990088 628714 990140
rect 631226 990088 631232 990140
rect 631284 990128 631290 990140
rect 673546 990128 673552 990140
rect 631284 990100 673552 990128
rect 631284 990088 631290 990100
rect 673546 990088 673552 990100
rect 673604 990088 673610 990140
rect 42518 990020 42524 990072
rect 42576 990060 42582 990072
rect 89916 990060 89944 990088
rect 42576 990032 89944 990060
rect 626552 990060 626580 990088
rect 628668 990060 628696 990088
rect 673454 990060 673460 990072
rect 626552 990032 673460 990060
rect 42576 990020 42582 990032
rect 673454 990020 673460 990032
rect 673512 990020 673518 990072
rect 41782 968464 41788 968516
rect 41840 968504 41846 968516
rect 42518 968504 42524 968516
rect 41840 968476 42524 968504
rect 41840 968464 41846 968476
rect 42518 968464 42524 968476
rect 42576 968464 42582 968516
rect 673454 965268 673460 965320
rect 673512 965308 673518 965320
rect 675386 965308 675392 965320
rect 673512 965280 675392 965308
rect 673512 965268 673518 965280
rect 675386 965268 675392 965280
rect 675444 965268 675450 965320
rect 673546 964724 673552 964776
rect 673604 964764 673610 964776
rect 675386 964764 675392 964776
rect 673604 964736 675392 964764
rect 673604 964724 673610 964736
rect 675386 964724 675392 964736
rect 675444 964724 675450 964776
rect 41782 958060 41788 958112
rect 41840 958100 41846 958112
rect 42334 958100 42340 958112
rect 41840 958072 42340 958100
rect 41840 958060 41846 958072
rect 42334 958060 42340 958072
rect 42392 958060 42398 958112
rect 42242 957720 42248 957772
rect 42300 957720 42306 957772
rect 42260 957568 42288 957720
rect 42242 957516 42248 957568
rect 42300 957516 42306 957568
rect 673638 953300 673644 953352
rect 673696 953340 673702 953352
rect 675386 953340 675392 953352
rect 673696 953312 675392 953340
rect 673696 953300 673702 953312
rect 675386 953300 675392 953312
rect 675444 953300 675450 953352
rect 673454 875168 673460 875220
rect 673512 875208 673518 875220
rect 675386 875208 675392 875220
rect 673512 875180 675392 875208
rect 673512 875168 673518 875180
rect 675386 875168 675392 875180
rect 675444 875168 675450 875220
rect 673546 874488 673552 874540
rect 673604 874528 673610 874540
rect 675386 874528 675392 874540
rect 673604 874500 675392 874528
rect 673604 874488 673610 874500
rect 675386 874488 675392 874500
rect 675444 874488 675450 874540
rect 673638 864424 673644 864476
rect 673696 864464 673702 864476
rect 675386 864464 675392 864476
rect 673696 864436 675392 864464
rect 673696 864424 673702 864436
rect 675386 864424 675392 864436
rect 675444 864424 675450 864476
rect 675294 818320 675300 818372
rect 675352 818360 675358 818372
rect 677502 818360 677508 818372
rect 675352 818332 677508 818360
rect 675352 818320 675358 818332
rect 677502 818320 677508 818332
rect 677560 818320 677566 818372
rect 41782 797716 41788 797768
rect 41840 797756 41846 797768
rect 42518 797756 42524 797768
rect 41840 797728 42524 797756
rect 41840 797716 41846 797728
rect 42518 797716 42524 797728
rect 42576 797756 42582 797768
rect 42702 797756 42708 797768
rect 42576 797728 42708 797756
rect 42576 797716 42582 797728
rect 42702 797716 42708 797728
rect 42760 797716 42766 797768
rect 41782 787244 41788 787296
rect 41840 787284 41846 787296
rect 42610 787284 42616 787296
rect 41840 787256 42616 787284
rect 41840 787244 41846 787256
rect 42610 787244 42616 787256
rect 42668 787244 42674 787296
rect 41782 786632 41788 786684
rect 41840 786672 41846 786684
rect 42518 786672 42524 786684
rect 41840 786644 42524 786672
rect 41840 786632 41846 786644
rect 42518 786632 42524 786644
rect 42576 786632 42582 786684
rect 673454 786564 673460 786616
rect 673512 786604 673518 786616
rect 674006 786604 674012 786616
rect 673512 786576 674012 786604
rect 673512 786564 673518 786576
rect 674006 786564 674012 786576
rect 674064 786604 674070 786616
rect 675386 786604 675392 786616
rect 674064 786576 675392 786604
rect 674064 786564 674070 786576
rect 675386 786564 675392 786576
rect 675444 786564 675450 786616
rect 673546 786360 673552 786412
rect 673604 786400 673610 786412
rect 675386 786400 675392 786412
rect 673604 786372 675392 786400
rect 673604 786360 673610 786372
rect 675386 786360 675392 786372
rect 675444 786360 675450 786412
rect 675294 781600 675300 781652
rect 675352 781600 675358 781652
rect 675312 781448 675340 781600
rect 675294 781396 675300 781448
rect 675352 781396 675358 781448
rect 673454 774868 673460 774920
rect 673512 774908 673518 774920
rect 673638 774908 673644 774920
rect 673512 774880 673644 774908
rect 673512 774868 673518 774880
rect 673638 774868 673644 774880
rect 673696 774908 673702 774920
rect 675386 774908 675392 774920
rect 673696 774880 675392 774908
rect 673696 774868 673702 774880
rect 675386 774868 675392 774880
rect 675444 774868 675450 774920
rect 673730 772760 673736 772812
rect 673788 772800 673794 772812
rect 674006 772800 674012 772812
rect 673788 772772 674012 772800
rect 673788 772760 673794 772772
rect 674006 772760 674012 772772
rect 674064 772760 674070 772812
rect 42426 767320 42432 767372
rect 42484 767360 42490 767372
rect 42702 767360 42708 767372
rect 42484 767332 42708 767360
rect 42484 767320 42490 767332
rect 42702 767320 42708 767332
rect 42760 767320 42766 767372
rect 42518 758956 42524 759008
rect 42576 758996 42582 759008
rect 42794 758996 42800 759008
rect 42576 758968 42800 758996
rect 42576 758956 42582 758968
rect 42794 758956 42800 758968
rect 42852 758956 42858 759008
rect 41782 754468 41788 754520
rect 41840 754508 41846 754520
rect 42426 754508 42432 754520
rect 41840 754480 42432 754508
rect 41840 754468 41846 754480
rect 42426 754468 42432 754480
rect 42484 754468 42490 754520
rect 673730 753516 673736 753568
rect 673788 753556 673794 753568
rect 673914 753556 673920 753568
rect 673788 753528 673920 753556
rect 673788 753516 673794 753528
rect 673914 753516 673920 753528
rect 673972 753516 673978 753568
rect 42518 753448 42524 753500
rect 42576 753488 42582 753500
rect 42794 753488 42800 753500
rect 42576 753460 42800 753488
rect 42576 753448 42582 753460
rect 42794 753448 42800 753460
rect 42852 753448 42858 753500
rect 41782 744132 41788 744184
rect 41840 744172 41846 744184
rect 42334 744172 42340 744184
rect 41840 744144 42340 744172
rect 41840 744132 41846 744144
rect 42334 744132 42340 744144
rect 42392 744172 42398 744184
rect 42610 744172 42616 744184
rect 42392 744144 42616 744172
rect 42392 744132 42398 744144
rect 42610 744132 42616 744144
rect 42668 744132 42674 744184
rect 41782 743996 41788 744048
rect 41840 744036 41846 744048
rect 42518 744036 42524 744048
rect 41840 744008 42524 744036
rect 41840 743996 41846 744008
rect 42518 743996 42524 744008
rect 42576 744036 42582 744048
rect 42978 744036 42984 744048
rect 42576 744008 42984 744036
rect 42576 743996 42582 744008
rect 42978 743996 42984 744008
rect 43036 743996 43042 744048
rect 673638 741956 673644 742008
rect 673696 741996 673702 742008
rect 673914 741996 673920 742008
rect 673696 741968 673920 741996
rect 673696 741956 673702 741968
rect 673914 741956 673920 741968
rect 673972 741996 673978 742008
rect 673972 741968 675432 741996
rect 673972 741956 673978 741968
rect 675404 741940 675432 741968
rect 675386 741888 675392 741940
rect 675444 741888 675450 741940
rect 673546 740664 673552 740716
rect 673604 740704 673610 740716
rect 675386 740704 675392 740716
rect 673604 740676 675392 740704
rect 673604 740664 673610 740676
rect 675386 740664 675392 740676
rect 675444 740664 675450 740716
rect 673638 739780 673644 739832
rect 673696 739780 673702 739832
rect 673656 739696 673684 739780
rect 673638 739644 673644 739696
rect 673696 739644 673702 739696
rect 42334 739576 42340 739628
rect 42392 739616 42398 739628
rect 42610 739616 42616 739628
rect 42392 739588 42616 739616
rect 42392 739576 42398 739588
rect 42610 739576 42616 739588
rect 42668 739576 42674 739628
rect 42518 734136 42524 734188
rect 42576 734176 42582 734188
rect 42978 734176 42984 734188
rect 42576 734148 42984 734176
rect 42576 734136 42582 734148
rect 42978 734136 42984 734148
rect 43036 734136 43042 734188
rect 673454 730124 673460 730176
rect 673512 730164 673518 730176
rect 675386 730164 675392 730176
rect 673512 730136 675392 730164
rect 673512 730124 673518 730136
rect 675386 730124 675392 730136
rect 675444 730124 675450 730176
rect 42518 720332 42524 720384
rect 42576 720372 42582 720384
rect 42886 720372 42892 720384
rect 42576 720344 42892 720372
rect 42576 720332 42582 720344
rect 42886 720332 42892 720344
rect 42944 720332 42950 720384
rect 41782 711288 41788 711340
rect 41840 711328 41846 711340
rect 42426 711328 42432 711340
rect 41840 711300 42432 711328
rect 41840 711288 41846 711300
rect 42426 711288 42432 711300
rect 42484 711328 42490 711340
rect 42702 711328 42708 711340
rect 42484 711300 42708 711328
rect 42484 711288 42490 711300
rect 42702 711288 42708 711300
rect 42760 711288 42766 711340
rect 673638 701020 673644 701072
rect 673696 701060 673702 701072
rect 673822 701060 673828 701072
rect 673696 701032 673828 701060
rect 673696 701020 673702 701032
rect 673822 701020 673828 701032
rect 673880 701020 673886 701072
rect 41782 700952 41788 701004
rect 41840 700992 41846 701004
rect 42610 700992 42616 701004
rect 41840 700964 42616 700992
rect 41840 700952 41846 700964
rect 42610 700952 42616 700964
rect 42668 700952 42674 701004
rect 41782 700816 41788 700868
rect 41840 700856 41846 700868
rect 42886 700856 42892 700868
rect 41840 700828 42892 700856
rect 41840 700816 41846 700828
rect 42886 700816 42892 700828
rect 42944 700816 42950 700868
rect 675386 695920 675392 695972
rect 675444 695920 675450 695972
rect 673638 695852 673644 695904
rect 673696 695892 673702 695904
rect 675404 695892 675432 695920
rect 673696 695864 675432 695892
rect 673696 695852 673702 695864
rect 42426 695512 42432 695564
rect 42484 695552 42490 695564
rect 42886 695552 42892 695564
rect 42484 695524 42892 695552
rect 42484 695512 42490 695524
rect 42886 695512 42892 695524
rect 42944 695512 42950 695564
rect 673546 695308 673552 695360
rect 673604 695348 673610 695360
rect 675386 695348 675392 695360
rect 673604 695320 675392 695348
rect 673604 695308 673610 695320
rect 675386 695308 675392 695320
rect 675444 695308 675450 695360
rect 673454 685176 673460 685228
rect 673512 685216 673518 685228
rect 675386 685216 675392 685228
rect 673512 685188 675392 685216
rect 673512 685176 673518 685188
rect 675386 685176 675392 685188
rect 675444 685176 675450 685228
rect 42426 681640 42432 681692
rect 42484 681640 42490 681692
rect 42444 681612 42472 681640
rect 42794 681612 42800 681624
rect 42444 681584 42800 681612
rect 42794 681572 42800 681584
rect 42852 681572 42858 681624
rect 42610 678512 42616 678564
rect 42668 678552 42674 678564
rect 42978 678552 42984 678564
rect 42668 678524 42984 678552
rect 42668 678512 42674 678524
rect 42978 678512 42984 678524
rect 43036 678512 43042 678564
rect 42426 676132 42432 676184
rect 42484 676172 42490 676184
rect 42978 676172 42984 676184
rect 42484 676144 42984 676172
rect 42484 676132 42490 676144
rect 42978 676132 42984 676144
rect 43036 676132 43042 676184
rect 41782 669060 41788 669112
rect 41840 669100 41846 669112
rect 42518 669100 42524 669112
rect 41840 669072 42524 669100
rect 41840 669060 41846 669072
rect 42518 669060 42524 669072
rect 42576 669060 42582 669112
rect 41782 658656 41788 658708
rect 41840 658696 41846 658708
rect 42426 658696 42432 658708
rect 41840 658668 42432 658696
rect 41840 658656 41846 658668
rect 42426 658656 42432 658668
rect 42484 658696 42490 658708
rect 42702 658696 42708 658708
rect 42484 658668 42708 658696
rect 42484 658656 42490 658668
rect 42702 658656 42708 658668
rect 42760 658656 42766 658708
rect 41782 658044 41788 658096
rect 41840 658084 41846 658096
rect 42794 658084 42800 658096
rect 41840 658056 42800 658084
rect 41840 658044 41846 658056
rect 42794 658044 42800 658056
rect 42852 658044 42858 658096
rect 673638 651720 673644 651772
rect 673696 651760 673702 651772
rect 675386 651760 675392 651772
rect 673696 651732 675392 651760
rect 673696 651720 673702 651732
rect 675386 651720 675392 651732
rect 675444 651720 675450 651772
rect 42426 651380 42432 651432
rect 42484 651420 42490 651432
rect 42794 651420 42800 651432
rect 42484 651392 42800 651420
rect 42484 651380 42490 651392
rect 42794 651380 42800 651392
rect 42852 651380 42858 651432
rect 673546 651108 673552 651160
rect 673604 651148 673610 651160
rect 675386 651148 675392 651160
rect 673604 651120 675392 651148
rect 673604 651108 673610 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 675202 646008 675208 646060
rect 675260 646008 675266 646060
rect 675220 645776 675248 646008
rect 675294 645776 675300 645788
rect 675220 645748 675300 645776
rect 675294 645736 675300 645748
rect 675352 645736 675358 645788
rect 673454 639684 673460 639736
rect 673512 639724 673518 639736
rect 673914 639724 673920 639736
rect 673512 639696 673920 639724
rect 673512 639684 673518 639696
rect 673914 639684 673920 639696
rect 673972 639724 673978 639736
rect 675386 639724 675392 639736
rect 673972 639696 675392 639724
rect 673972 639684 673978 639696
rect 675386 639684 675392 639696
rect 675444 639684 675450 639736
rect 42518 632000 42524 632052
rect 42576 632000 42582 632052
rect 42702 632000 42708 632052
rect 42760 632040 42766 632052
rect 42978 632040 42984 632052
rect 42760 632012 42984 632040
rect 42760 632000 42766 632012
rect 42978 632000 42984 632012
rect 43036 632000 43042 632052
rect 42536 631904 42564 632000
rect 42794 631904 42800 631916
rect 42536 631876 42800 631904
rect 42794 631864 42800 631876
rect 42852 631864 42858 631916
rect 41782 624928 41788 624980
rect 41840 624968 41846 624980
rect 42794 624968 42800 624980
rect 41840 624940 42800 624968
rect 41840 624928 41846 624940
rect 42794 624928 42800 624940
rect 42852 624928 42858 624980
rect 41782 615476 41788 615528
rect 41840 615516 41846 615528
rect 42978 615516 42984 615528
rect 41840 615488 42984 615516
rect 41840 615476 41846 615488
rect 42978 615476 42984 615488
rect 43036 615476 43042 615528
rect 41782 614796 41788 614848
rect 41840 614836 41846 614848
rect 42518 614836 42524 614848
rect 41840 614808 42524 614836
rect 41840 614796 41846 614808
rect 42518 614796 42524 614808
rect 42576 614796 42582 614848
rect 42794 612824 42800 612876
rect 42852 612824 42858 612876
rect 42610 612756 42616 612808
rect 42668 612796 42674 612808
rect 42812 612796 42840 612824
rect 42668 612768 42840 612796
rect 42668 612756 42674 612768
rect 42610 612620 42616 612672
rect 42668 612660 42674 612672
rect 42794 612660 42800 612672
rect 42668 612632 42800 612660
rect 42668 612620 42674 612632
rect 42794 612620 42800 612632
rect 42852 612620 42858 612672
rect 673638 606704 673644 606756
rect 673696 606744 673702 606756
rect 675386 606744 675392 606756
rect 673696 606716 675392 606744
rect 673696 606704 673702 606716
rect 675386 606704 675392 606716
rect 675444 606704 675450 606756
rect 673546 606160 673552 606212
rect 673604 606200 673610 606212
rect 675018 606200 675024 606212
rect 673604 606172 675024 606200
rect 673604 606160 673610 606172
rect 675018 606160 675024 606172
rect 675076 606200 675082 606212
rect 675386 606200 675392 606212
rect 675076 606172 675392 606200
rect 675076 606160 675082 606172
rect 675386 606160 675392 606172
rect 675444 606160 675450 606212
rect 673638 594872 673644 594924
rect 673696 594912 673702 594924
rect 673914 594912 673920 594924
rect 673696 594884 673920 594912
rect 673696 594872 673702 594884
rect 673914 594872 673920 594884
rect 673972 594912 673978 594924
rect 675386 594912 675392 594924
rect 673972 594884 675392 594912
rect 673972 594872 673978 594884
rect 675386 594872 675392 594884
rect 675444 594872 675450 594924
rect 673730 594736 673736 594788
rect 673788 594776 673794 594788
rect 675018 594776 675024 594788
rect 673788 594748 675024 594776
rect 673788 594736 673794 594748
rect 675018 594736 675024 594748
rect 675076 594736 675082 594788
rect 675294 593376 675300 593428
rect 675352 593376 675358 593428
rect 675312 593224 675340 593376
rect 675294 593172 675300 593224
rect 675352 593172 675358 593224
rect 673546 585148 673552 585200
rect 673604 585188 673610 585200
rect 673822 585188 673828 585200
rect 673604 585160 673828 585188
rect 673604 585148 673610 585160
rect 673822 585148 673828 585160
rect 673880 585148 673886 585200
rect 41782 582632 41788 582684
rect 41840 582672 41846 582684
rect 42794 582672 42800 582684
rect 41840 582644 42800 582672
rect 41840 582632 41846 582644
rect 42794 582632 42800 582644
rect 42852 582632 42858 582684
rect 673730 575424 673736 575476
rect 673788 575464 673794 575476
rect 674374 575464 674380 575476
rect 673788 575436 674380 575464
rect 673788 575424 673794 575436
rect 674374 575424 674380 575436
rect 674432 575424 674438 575476
rect 42334 574064 42340 574116
rect 42392 574104 42398 574116
rect 42794 574104 42800 574116
rect 42392 574076 42800 574104
rect 42392 574064 42398 574076
rect 42794 574064 42800 574076
rect 42852 574064 42858 574116
rect 41782 571208 41788 571260
rect 41840 571248 41846 571260
rect 42794 571248 42800 571260
rect 41840 571220 42800 571248
rect 41840 571208 41846 571220
rect 42794 571208 42800 571220
rect 42852 571208 42858 571260
rect 41782 570664 41788 570716
rect 41840 570704 41846 570716
rect 42518 570704 42524 570716
rect 41840 570676 42524 570704
rect 41840 570664 41846 570676
rect 42518 570664 42524 570676
rect 42576 570704 42582 570716
rect 42702 570704 42708 570716
rect 42576 570676 42708 570704
rect 42576 570664 42582 570676
rect 42702 570664 42708 570676
rect 42760 570664 42766 570716
rect 673546 560532 673552 560584
rect 673604 560572 673610 560584
rect 673822 560572 673828 560584
rect 673604 560544 673828 560572
rect 673604 560532 673610 560544
rect 673822 560532 673828 560544
rect 673880 560572 673886 560584
rect 675386 560572 675392 560584
rect 673880 560544 675392 560572
rect 673880 560532 673886 560544
rect 675386 560532 675392 560544
rect 675444 560532 675450 560584
rect 674006 559920 674012 559972
rect 674064 559960 674070 559972
rect 674374 559960 674380 559972
rect 674064 559932 674380 559960
rect 674064 559920 674070 559932
rect 674374 559920 674380 559932
rect 674432 559960 674438 559972
rect 675386 559960 675392 559972
rect 674432 559932 675392 559960
rect 674432 559920 674438 559932
rect 675386 559920 675392 559932
rect 675444 559920 675450 559972
rect 42610 554752 42616 554804
rect 42668 554792 42674 554804
rect 42794 554792 42800 554804
rect 42668 554764 42800 554792
rect 42668 554752 42674 554764
rect 42794 554752 42800 554764
rect 42852 554752 42858 554804
rect 673638 550468 673644 550520
rect 673696 550508 673702 550520
rect 675386 550508 675392 550520
rect 673696 550480 675392 550508
rect 673696 550468 673702 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 673546 546388 673552 546440
rect 673604 546388 673610 546440
rect 673564 546360 673592 546388
rect 673822 546360 673828 546372
rect 673564 546332 673828 546360
rect 673822 546320 673828 546332
rect 673880 546320 673886 546372
rect 41782 539452 41788 539504
rect 41840 539492 41846 539504
rect 42518 539492 42524 539504
rect 41840 539464 42524 539492
rect 41840 539452 41846 539464
rect 42518 539452 42524 539464
rect 42576 539452 42582 539504
rect 41782 528028 41788 528080
rect 41840 528068 41846 528080
rect 42610 528068 42616 528080
rect 41840 528040 42616 528068
rect 41840 528028 41846 528040
rect 42610 528028 42616 528040
rect 42668 528028 42674 528080
rect 41782 527484 41788 527536
rect 41840 527524 41846 527536
rect 42426 527524 42432 527536
rect 41840 527496 42432 527524
rect 41840 527484 41846 527496
rect 42426 527484 42432 527496
rect 42484 527524 42490 527536
rect 42702 527524 42708 527536
rect 42484 527496 42708 527524
rect 42484 527484 42490 527496
rect 42702 527484 42708 527496
rect 42760 527484 42766 527536
rect 675294 513748 675300 513800
rect 675352 513788 675358 513800
rect 677686 513788 677692 513800
rect 675352 513760 677692 513788
rect 675352 513748 675358 513760
rect 677686 513748 677692 513760
rect 677744 513748 677750 513800
rect 673730 502324 673736 502376
rect 673788 502364 673794 502376
rect 673914 502364 673920 502376
rect 673788 502336 673920 502364
rect 673788 502324 673794 502336
rect 673914 502324 673920 502336
rect 673972 502324 673978 502376
rect 673546 498176 673552 498228
rect 673604 498216 673610 498228
rect 673822 498216 673828 498228
rect 673604 498188 673828 498216
rect 673604 498176 673610 498188
rect 673822 498176 673828 498188
rect 673880 498176 673886 498228
rect 673822 469316 673828 469328
rect 673748 469288 673828 469316
rect 673748 469192 673776 469288
rect 673822 469276 673828 469288
rect 673880 469276 673886 469328
rect 673730 469140 673736 469192
rect 673788 469140 673794 469192
rect 673730 463632 673736 463684
rect 673788 463672 673794 463684
rect 674006 463672 674012 463684
rect 673788 463644 674012 463672
rect 673788 463632 673794 463644
rect 674006 463632 674012 463644
rect 674064 463632 674070 463684
rect 673546 449556 673552 449608
rect 673604 449596 673610 449608
rect 673822 449596 673828 449608
rect 673604 449568 673828 449596
rect 673604 449556 673610 449568
rect 673822 449556 673828 449568
rect 673880 449556 673886 449608
rect 42610 444320 42616 444372
rect 42668 444360 42674 444372
rect 42794 444360 42800 444372
rect 42668 444332 42800 444360
rect 42668 444320 42674 444332
rect 42794 444320 42800 444332
rect 42852 444320 42858 444372
rect 673730 444320 673736 444372
rect 673788 444360 673794 444372
rect 674006 444360 674012 444372
rect 673788 444332 674012 444360
rect 673788 444320 673794 444332
rect 674006 444320 674012 444332
rect 674064 444320 674070 444372
rect 42702 441532 42708 441584
rect 42760 441572 42766 441584
rect 42794 441572 42800 441584
rect 42760 441544 42800 441572
rect 42760 441532 42766 441544
rect 42794 441532 42800 441544
rect 42852 441532 42858 441584
rect 674742 427796 674748 427848
rect 674800 427836 674806 427848
rect 677118 427836 677124 427848
rect 674800 427808 677124 427836
rect 674800 427796 674806 427808
rect 677118 427796 677124 427808
rect 677176 427796 677182 427848
rect 42610 422288 42616 422340
rect 42668 422328 42674 422340
rect 42702 422328 42708 422340
rect 42668 422300 42708 422328
rect 42668 422288 42674 422300
rect 42702 422288 42708 422300
rect 42760 422288 42766 422340
rect 673638 420724 673644 420776
rect 673696 420764 673702 420776
rect 673822 420764 673828 420776
rect 673696 420736 673828 420764
rect 673696 420724 673702 420736
rect 673822 420724 673828 420736
rect 673880 420724 673886 420776
rect 41782 411204 41788 411256
rect 41840 411244 41846 411256
rect 42518 411244 42524 411256
rect 41840 411216 42524 411244
rect 41840 411204 41846 411216
rect 42518 411204 42524 411216
rect 42576 411204 42582 411256
rect 42610 405696 42616 405748
rect 42668 405736 42674 405748
rect 42886 405736 42892 405748
rect 42668 405708 42892 405736
rect 42668 405696 42674 405708
rect 42886 405696 42892 405708
rect 42944 405696 42950 405748
rect 673822 401548 673828 401600
rect 673880 401588 673886 401600
rect 675294 401588 675300 401600
rect 673880 401560 675300 401588
rect 673880 401548 673886 401560
rect 675294 401548 675300 401560
rect 675352 401548 675358 401600
rect 41782 401344 41788 401396
rect 41840 401384 41846 401396
rect 42886 401384 42892 401396
rect 41840 401356 42892 401384
rect 41840 401344 41846 401356
rect 42886 401344 42892 401356
rect 42944 401344 42950 401396
rect 41782 400800 41788 400852
rect 41840 400840 41846 400852
rect 42426 400840 42432 400852
rect 41840 400812 42432 400840
rect 41840 400800 41846 400812
rect 42426 400800 42432 400812
rect 42484 400800 42490 400852
rect 42610 386316 42616 386368
rect 42668 386356 42674 386368
rect 42886 386356 42892 386368
rect 42668 386328 42892 386356
rect 42668 386316 42674 386328
rect 42886 386316 42892 386328
rect 42944 386316 42950 386368
rect 673730 384276 673736 384328
rect 673788 384316 673794 384328
rect 675386 384316 675392 384328
rect 673788 384288 675392 384316
rect 673788 384276 673794 384288
rect 675386 384276 675392 384288
rect 675444 384276 675450 384328
rect 673638 383188 673644 383240
rect 673696 383228 673702 383240
rect 675294 383228 675300 383240
rect 673696 383200 675300 383228
rect 673696 383188 673702 383200
rect 675294 383188 675300 383200
rect 675352 383188 675358 383240
rect 673546 380876 673552 380928
rect 673604 380916 673610 380928
rect 673730 380916 673736 380928
rect 673604 380888 673736 380916
rect 673604 380876 673610 380888
rect 673730 380876 673736 380888
rect 673788 380876 673794 380928
rect 42794 372580 42800 372632
rect 42852 372620 42858 372632
rect 42978 372620 42984 372632
rect 42852 372592 42984 372620
rect 42852 372580 42858 372592
rect 42978 372580 42984 372592
rect 43036 372580 43042 372632
rect 673730 372308 673736 372360
rect 673788 372348 673794 372360
rect 675386 372348 675392 372360
rect 673788 372320 675392 372348
rect 673788 372308 673794 372320
rect 675386 372308 675392 372320
rect 675444 372308 675450 372360
rect 41782 368636 41788 368688
rect 41840 368676 41846 368688
rect 42886 368676 42892 368688
rect 41840 368648 42892 368676
rect 41840 368636 41846 368648
rect 42886 368636 42892 368648
rect 42944 368636 42950 368688
rect 42518 367820 42524 367872
rect 42576 367860 42582 367872
rect 42794 367860 42800 367872
rect 42576 367832 42800 367860
rect 42576 367820 42582 367832
rect 42794 367820 42800 367832
rect 42852 367820 42858 367872
rect 41782 358232 41788 358284
rect 41840 358272 41846 358284
rect 42518 358272 42524 358284
rect 41840 358244 42524 358272
rect 41840 358232 41846 358244
rect 42518 358232 42524 358244
rect 42576 358232 42582 358284
rect 41782 357620 41788 357672
rect 41840 357660 41846 357672
rect 42426 357660 42432 357672
rect 41840 357632 42432 357660
rect 41840 357620 41846 357632
rect 42426 357620 42432 357632
rect 42484 357660 42490 357672
rect 42610 357660 42616 357672
rect 42484 357632 42616 357660
rect 42484 357620 42490 357632
rect 42610 357620 42616 357632
rect 42668 357620 42674 357672
rect 673546 338104 673552 338156
rect 673604 338144 673610 338156
rect 675386 338144 675392 338156
rect 673604 338116 675392 338144
rect 673604 338104 673610 338116
rect 675386 338104 675392 338116
rect 675444 338104 675450 338156
rect 673638 337492 673644 337544
rect 673696 337532 673702 337544
rect 675386 337532 675392 337544
rect 673696 337504 675392 337532
rect 673696 337492 673702 337504
rect 675386 337492 675392 337504
rect 675444 337492 675450 337544
rect 673730 328040 673736 328092
rect 673788 328080 673794 328092
rect 675386 328080 675392 328092
rect 673788 328052 675392 328080
rect 673788 328040 673794 328052
rect 675386 328040 675392 328052
rect 675444 328040 675450 328092
rect 41782 325456 41788 325508
rect 41840 325496 41846 325508
rect 42426 325496 42432 325508
rect 41840 325468 42432 325496
rect 41840 325456 41846 325468
rect 42426 325456 42432 325468
rect 42484 325496 42490 325508
rect 42702 325496 42708 325508
rect 42484 325468 42708 325496
rect 42484 325456 42490 325468
rect 42702 325456 42708 325468
rect 42760 325456 42766 325508
rect 42426 322872 42432 322924
rect 42484 322912 42490 322924
rect 42484 322884 42748 322912
rect 42484 322872 42490 322884
rect 42720 322856 42748 322884
rect 42610 322804 42616 322856
rect 42668 322804 42674 322856
rect 42702 322804 42708 322856
rect 42760 322804 42766 322856
rect 42628 322776 42656 322804
rect 42886 322776 42892 322788
rect 42628 322748 42892 322776
rect 42886 322736 42892 322748
rect 42944 322736 42950 322788
rect 42334 314168 42340 314220
rect 42392 314208 42398 314220
rect 42702 314208 42708 314220
rect 42392 314180 42708 314208
rect 42392 314168 42398 314180
rect 42702 314168 42708 314180
rect 42760 314168 42766 314220
rect 41782 314032 41788 314084
rect 41840 314072 41846 314084
rect 42518 314072 42524 314084
rect 41840 314044 42524 314072
rect 41840 314032 41846 314044
rect 42518 314032 42524 314044
rect 42576 314072 42582 314084
rect 42702 314072 42708 314084
rect 42576 314044 42708 314072
rect 42576 314032 42582 314044
rect 42702 314032 42708 314044
rect 42760 314032 42766 314084
rect 41782 313488 41788 313540
rect 41840 313488 41846 313540
rect 41800 313460 41828 313488
rect 42794 313460 42800 313472
rect 41800 313432 42800 313460
rect 42794 313420 42800 313432
rect 42852 313420 42858 313472
rect 673546 303560 673552 303612
rect 673604 303600 673610 303612
rect 675294 303600 675300 303612
rect 673604 303572 675300 303600
rect 673604 303560 673610 303572
rect 675294 303560 675300 303572
rect 675352 303560 675358 303612
rect 673638 293564 673644 293616
rect 673696 293604 673702 293616
rect 673914 293604 673920 293616
rect 673696 293576 673920 293604
rect 673696 293564 673702 293576
rect 673914 293564 673920 293576
rect 673972 293604 673978 293616
rect 675386 293604 675392 293616
rect 673972 293576 675392 293604
rect 673972 293564 673978 293576
rect 675386 293564 675392 293576
rect 675444 293564 675450 293616
rect 673638 293428 673644 293480
rect 673696 293468 673702 293480
rect 675294 293468 675300 293480
rect 673696 293440 675300 293468
rect 673696 293428 673702 293440
rect 675294 293428 675300 293440
rect 675352 293428 675358 293480
rect 41782 282276 41788 282328
rect 41840 282316 41846 282328
rect 42518 282316 42524 282328
rect 41840 282288 42524 282316
rect 41840 282276 41846 282288
rect 42518 282276 42524 282288
rect 42576 282276 42582 282328
rect 673730 282072 673736 282124
rect 673788 282112 673794 282124
rect 675386 282112 675392 282124
rect 673788 282084 675392 282112
rect 673788 282072 673794 282084
rect 675386 282072 675392 282084
rect 675444 282072 675450 282124
rect 41782 271872 41788 271924
rect 41840 271912 41846 271924
rect 42702 271912 42708 271924
rect 41840 271884 42708 271912
rect 41840 271872 41846 271884
rect 42702 271872 42708 271884
rect 42760 271872 42766 271924
rect 41782 271192 41788 271244
rect 41840 271232 41846 271244
rect 42518 271232 42524 271244
rect 41840 271204 42524 271232
rect 41840 271192 41846 271204
rect 42518 271192 42524 271204
rect 42576 271232 42582 271244
rect 42794 271232 42800 271244
rect 42576 271204 42800 271232
rect 42576 271192 42582 271204
rect 42794 271192 42800 271204
rect 42852 271192 42858 271244
rect 673454 264936 673460 264988
rect 673512 264976 673518 264988
rect 673638 264976 673644 264988
rect 673512 264948 673644 264976
rect 673512 264936 673518 264948
rect 673638 264936 673644 264948
rect 673696 264936 673702 264988
rect 673454 248684 673460 248736
rect 673512 248724 673518 248736
rect 675294 248724 675300 248736
rect 673512 248696 675300 248724
rect 673512 248684 673518 248696
rect 675294 248684 675300 248696
rect 675352 248684 675358 248736
rect 673638 247460 673644 247512
rect 673696 247500 673702 247512
rect 673914 247500 673920 247512
rect 673696 247472 673920 247500
rect 673696 247460 673702 247472
rect 673914 247460 673920 247472
rect 673972 247500 673978 247512
rect 675386 247500 675392 247512
rect 673972 247472 675392 247500
rect 673972 247460 673978 247472
rect 675386 247460 675392 247472
rect 675444 247460 675450 247512
rect 42334 245556 42340 245608
rect 42392 245596 42398 245608
rect 42886 245596 42892 245608
rect 42392 245568 42892 245596
rect 42392 245556 42398 245568
rect 42886 245556 42892 245568
rect 42944 245556 42950 245608
rect 42518 245488 42524 245540
rect 42576 245528 42582 245540
rect 42794 245528 42800 245540
rect 42576 245500 42800 245528
rect 42576 245488 42582 245500
rect 42794 245488 42800 245500
rect 42852 245488 42858 245540
rect 673822 243788 673828 243840
rect 673880 243828 673886 243840
rect 675294 243828 675300 243840
rect 673880 243800 675300 243828
rect 673880 243788 673886 243800
rect 675294 243788 675300 243800
rect 675352 243788 675358 243840
rect 41782 238076 41788 238128
rect 41840 238116 41846 238128
rect 42610 238116 42616 238128
rect 41840 238088 42616 238116
rect 41840 238076 41846 238088
rect 42610 238076 42616 238088
rect 42668 238116 42674 238128
rect 42886 238116 42892 238128
rect 42668 238088 42892 238116
rect 42668 238076 42674 238088
rect 42886 238076 42892 238088
rect 42944 238076 42950 238128
rect 673914 237668 673920 237720
rect 673972 237708 673978 237720
rect 675386 237708 675392 237720
rect 673972 237680 675392 237708
rect 673972 237668 673978 237680
rect 675386 237668 675392 237680
rect 675444 237668 675450 237720
rect 673914 237328 673920 237380
rect 673972 237368 673978 237380
rect 674098 237368 674104 237380
rect 673972 237340 674104 237368
rect 673972 237328 673978 237340
rect 674098 237328 674104 237340
rect 674156 237328 674162 237380
rect 42334 232840 42340 232892
rect 42392 232880 42398 232892
rect 42610 232880 42616 232892
rect 42392 232852 42616 232880
rect 42392 232840 42398 232852
rect 42610 232840 42616 232852
rect 42668 232840 42674 232892
rect 674098 231752 674104 231804
rect 674156 231792 674162 231804
rect 674282 231792 674288 231804
rect 674156 231764 674288 231792
rect 674156 231752 674162 231764
rect 674282 231752 674288 231764
rect 674340 231752 674346 231804
rect 41782 228624 41788 228676
rect 41840 228664 41846 228676
rect 42702 228664 42708 228676
rect 41840 228636 42708 228664
rect 41840 228624 41846 228636
rect 42702 228624 42708 228636
rect 42760 228624 42766 228676
rect 41782 228012 41788 228064
rect 41840 228052 41846 228064
rect 42610 228052 42616 228064
rect 41840 228024 42616 228052
rect 41840 228012 41846 228024
rect 42610 228012 42616 228024
rect 42668 228052 42674 228064
rect 42794 228052 42800 228064
rect 42668 228024 42800 228052
rect 42668 228012 42674 228024
rect 42794 228012 42800 228024
rect 42852 228012 42858 228064
rect 673822 218084 673828 218136
rect 673880 218084 673886 218136
rect 673840 218000 673868 218084
rect 673822 217948 673828 218000
rect 673880 217948 673886 218000
rect 673730 212508 673736 212560
rect 673788 212548 673794 212560
rect 673822 212548 673828 212560
rect 673788 212520 673828 212548
rect 673788 212508 673794 212520
rect 673822 212508 673828 212520
rect 673880 212508 673886 212560
rect 674006 212508 674012 212560
rect 674064 212548 674070 212560
rect 674282 212548 674288 212560
rect 674064 212520 674288 212548
rect 674064 212508 674070 212520
rect 674282 212508 674288 212520
rect 674340 212508 674346 212560
rect 42334 208360 42340 208412
rect 42392 208400 42398 208412
rect 42886 208400 42892 208412
rect 42392 208372 42892 208400
rect 42392 208360 42398 208372
rect 42886 208360 42892 208372
rect 42944 208360 42950 208412
rect 673730 203872 673736 203924
rect 673788 203912 673794 203924
rect 675386 203912 675392 203924
rect 673788 203884 675392 203912
rect 673788 203872 673794 203884
rect 675386 203872 675392 203884
rect 675444 203872 675450 203924
rect 673638 203328 673644 203380
rect 673696 203368 673702 203380
rect 675386 203368 675392 203380
rect 673696 203340 675392 203368
rect 673696 203328 673702 203340
rect 675386 203328 675392 203340
rect 675444 203328 675450 203380
rect 674006 198704 674012 198756
rect 674064 198744 674070 198756
rect 675202 198744 675208 198756
rect 674064 198716 675208 198744
rect 674064 198704 674070 198716
rect 675202 198704 675208 198716
rect 675260 198704 675266 198756
rect 41782 194896 41788 194948
rect 41840 194936 41846 194948
rect 42426 194936 42432 194948
rect 41840 194908 42432 194936
rect 41840 194896 41846 194908
rect 42426 194896 42432 194908
rect 42484 194936 42490 194948
rect 42886 194936 42892 194948
rect 42484 194908 42892 194936
rect 42484 194896 42490 194908
rect 42886 194896 42892 194908
rect 42944 194896 42950 194948
rect 674742 192108 674748 192160
rect 674800 192148 674806 192160
rect 675202 192148 675208 192160
rect 674800 192120 675208 192148
rect 674800 192108 674806 192120
rect 675202 192108 675208 192120
rect 675260 192148 675266 192160
rect 675386 192148 675392 192160
rect 675260 192120 675392 192148
rect 675260 192108 675266 192120
rect 675386 192108 675392 192120
rect 675444 192108 675450 192160
rect 41782 185444 41788 185496
rect 41840 185484 41846 185496
rect 42334 185484 42340 185496
rect 41840 185456 42340 185484
rect 41840 185444 41846 185456
rect 42334 185444 42340 185456
rect 42392 185484 42398 185496
rect 42702 185484 42708 185496
rect 42392 185456 42708 185484
rect 42392 185444 42398 185456
rect 42702 185444 42708 185456
rect 42760 185444 42766 185496
rect 42426 185308 42432 185360
rect 42484 185348 42490 185360
rect 42702 185348 42708 185360
rect 42484 185320 42708 185348
rect 42484 185308 42490 185320
rect 42702 185308 42708 185320
rect 42760 185308 42766 185360
rect 41782 184832 41788 184884
rect 41840 184872 41846 184884
rect 42426 184872 42432 184884
rect 41840 184844 42432 184872
rect 41840 184832 41846 184844
rect 42426 184832 42432 184844
rect 42484 184872 42490 184884
rect 42610 184872 42616 184884
rect 42484 184844 42616 184872
rect 42484 184832 42490 184844
rect 42610 184832 42616 184844
rect 42668 184832 42674 184884
rect 673822 173884 673828 173936
rect 673880 173924 673886 173936
rect 674742 173924 674748 173936
rect 673880 173896 674748 173924
rect 673880 173884 673886 173896
rect 674742 173884 674748 173896
rect 674800 173884 674806 173936
rect 673546 158312 673552 158364
rect 673604 158352 673610 158364
rect 675386 158352 675392 158364
rect 673604 158324 675392 158352
rect 673604 158312 673610 158324
rect 675386 158312 675392 158324
rect 675444 158312 675450 158364
rect 673454 157292 673460 157344
rect 673512 157332 673518 157344
rect 675386 157332 675392 157344
rect 673512 157304 675392 157332
rect 673512 157292 673518 157304
rect 675386 157292 675392 157304
rect 675444 157292 675450 157344
rect 42518 149064 42524 149116
rect 42576 149104 42582 149116
rect 42702 149104 42708 149116
rect 42576 149076 42708 149104
rect 42576 149064 42582 149076
rect 42702 149064 42708 149076
rect 42760 149064 42766 149116
rect 673638 147092 673644 147144
rect 673696 147132 673702 147144
rect 675018 147132 675024 147144
rect 673696 147104 675024 147132
rect 673696 147092 673702 147104
rect 675018 147092 675024 147104
rect 675076 147132 675082 147144
rect 675386 147132 675392 147144
rect 675076 147104 675392 147132
rect 675076 147092 675082 147104
rect 675386 147092 675392 147104
rect 675444 147092 675450 147144
rect 674006 140632 674012 140684
rect 674064 140672 674070 140684
rect 675018 140672 675024 140684
rect 674064 140644 675024 140672
rect 674064 140632 674070 140644
rect 675018 140632 675024 140644
rect 675076 140632 675082 140684
rect 42242 121456 42248 121508
rect 42300 121496 42306 121508
rect 44726 121496 44732 121508
rect 42300 121468 44732 121496
rect 42300 121456 42306 121468
rect 44726 121456 44732 121468
rect 44784 121456 44790 121508
rect 673822 115948 673828 116000
rect 673880 115988 673886 116000
rect 674006 115988 674012 116000
rect 673880 115960 674012 115988
rect 673880 115948 673886 115960
rect 674006 115948 674012 115960
rect 674064 115948 674070 116000
rect 42978 115880 42984 115932
rect 43036 115920 43042 115932
rect 44726 115920 44732 115932
rect 43036 115892 44732 115920
rect 43036 115880 43042 115892
rect 44726 115880 44732 115892
rect 44784 115880 44790 115932
rect 673822 115812 673828 115864
rect 673880 115852 673886 115864
rect 675018 115852 675024 115864
rect 673880 115824 675024 115852
rect 673880 115812 673886 115824
rect 675018 115812 675024 115824
rect 675076 115812 675082 115864
rect 673546 112752 673552 112804
rect 673604 112792 673610 112804
rect 675386 112792 675392 112804
rect 673604 112764 675392 112792
rect 673604 112752 673610 112764
rect 675386 112752 675392 112764
rect 675444 112752 675450 112804
rect 673454 112072 673460 112124
rect 673512 112112 673518 112124
rect 675386 112112 675392 112124
rect 673512 112084 675392 112112
rect 673512 112072 673518 112084
rect 675386 112072 675392 112084
rect 675444 112072 675450 112124
rect 42518 110440 42524 110492
rect 42576 110480 42582 110492
rect 42702 110480 42708 110492
rect 42576 110452 42708 110480
rect 42576 110440 42582 110452
rect 42702 110440 42708 110452
rect 42760 110440 42766 110492
rect 673638 102280 673644 102332
rect 673696 102320 673702 102332
rect 675018 102320 675024 102332
rect 673696 102292 675024 102320
rect 673696 102280 673702 102292
rect 675018 102280 675024 102292
rect 675076 102320 675082 102332
rect 675386 102320 675392 102332
rect 675076 102292 675392 102320
rect 675076 102280 675082 102292
rect 675386 102280 675392 102292
rect 675444 102280 675450 102332
rect 44634 82832 44640 82884
rect 44692 82832 44698 82884
rect 44652 82804 44680 82832
rect 44818 82804 44824 82816
rect 44652 82776 44824 82804
rect 44818 82764 44824 82776
rect 44876 82764 44882 82816
rect 42334 45704 42340 45756
rect 42392 45744 42398 45756
rect 140958 45744 140964 45756
rect 42392 45716 140964 45744
rect 42392 45704 42398 45716
rect 140958 45704 140964 45716
rect 141016 45704 141022 45756
rect 42426 45636 42432 45688
rect 42484 45676 42490 45688
rect 143626 45676 143632 45688
rect 42484 45648 143632 45676
rect 42484 45636 42490 45648
rect 143626 45636 143632 45648
rect 143684 45636 143690 45688
rect 42702 45568 42708 45620
rect 42760 45608 42766 45620
rect 143534 45608 143540 45620
rect 42760 45580 143540 45608
rect 42760 45568 42766 45580
rect 143534 45568 143540 45580
rect 143592 45568 143598 45620
rect 527450 45568 527456 45620
rect 527508 45608 527514 45620
rect 673546 45608 673552 45620
rect 527508 45580 673552 45608
rect 527508 45568 527514 45580
rect 673546 45568 673552 45580
rect 673604 45568 673610 45620
rect 44910 45500 44916 45552
rect 44968 45540 44974 45552
rect 195974 45540 195980 45552
rect 44968 45512 195980 45540
rect 44968 45500 44974 45512
rect 195974 45500 195980 45512
rect 196032 45500 196038 45552
rect 516318 45500 516324 45552
rect 516376 45540 516382 45552
rect 673638 45540 673644 45552
rect 516376 45512 673644 45540
rect 516376 45500 516382 45512
rect 673638 45500 673644 45512
rect 673696 45500 673702 45552
rect 405642 44752 405648 44804
rect 405700 44792 405706 44804
rect 411254 44792 411260 44804
rect 405700 44764 411260 44792
rect 405700 44752 405706 44764
rect 411254 44752 411260 44764
rect 411312 44752 411318 44804
rect 359366 44724 359372 44736
rect 342272 44696 359372 44724
rect 195974 44412 195980 44464
rect 196032 44452 196038 44464
rect 304534 44452 304540 44464
rect 196032 44424 304540 44452
rect 196032 44412 196038 44424
rect 304534 44412 304540 44424
rect 304592 44452 304598 44464
rect 342272 44452 342300 44696
rect 359366 44684 359372 44696
rect 359424 44684 359430 44736
rect 406746 44684 406752 44736
rect 406804 44724 406810 44736
rect 406804 44696 411300 44724
rect 406804 44684 406810 44696
rect 411272 44588 411300 44696
rect 425054 44684 425060 44736
rect 425112 44724 425118 44736
rect 444190 44724 444196 44736
rect 425112 44696 444196 44724
rect 425112 44684 425118 44696
rect 444190 44684 444196 44696
rect 444248 44684 444254 44736
rect 483014 44656 483020 44668
rect 473280 44628 483020 44656
rect 425054 44588 425060 44600
rect 411272 44560 425060 44588
rect 425054 44548 425060 44560
rect 425112 44548 425118 44600
rect 461486 44588 461492 44600
rect 449820 44560 461492 44588
rect 354398 44480 354404 44532
rect 354456 44520 354462 44532
rect 360562 44520 360568 44532
rect 354456 44492 360568 44520
rect 354456 44480 354462 44492
rect 360562 44480 360568 44492
rect 360620 44480 360626 44532
rect 360654 44480 360660 44532
rect 360712 44520 360718 44532
rect 386414 44520 386420 44532
rect 360712 44492 386420 44520
rect 360712 44480 360718 44492
rect 386414 44480 386420 44492
rect 386472 44480 386478 44532
rect 399662 44480 399668 44532
rect 399720 44520 399726 44532
rect 406746 44520 406752 44532
rect 399720 44492 406752 44520
rect 399720 44480 399726 44492
rect 406746 44480 406752 44492
rect 406804 44480 406810 44532
rect 411254 44480 411260 44532
rect 411312 44520 411318 44532
rect 411312 44492 414244 44520
rect 411312 44480 411318 44492
rect 414216 44464 414244 44492
rect 444282 44480 444288 44532
rect 444340 44520 444346 44532
rect 449820 44520 449848 44560
rect 461486 44548 461492 44560
rect 461544 44588 461550 44600
rect 469122 44588 469128 44600
rect 461544 44560 469128 44588
rect 461544 44548 461550 44560
rect 469122 44548 469128 44560
rect 469180 44548 469186 44600
rect 469214 44548 469220 44600
rect 469272 44588 469278 44600
rect 473280 44588 473308 44628
rect 483014 44616 483020 44628
rect 483072 44616 483078 44668
rect 469272 44560 473308 44588
rect 502260 44560 502380 44588
rect 469272 44548 469278 44560
rect 502260 44532 502288 44560
rect 444340 44492 449848 44520
rect 444340 44480 444346 44492
rect 502242 44480 502248 44532
rect 502300 44480 502306 44532
rect 502352 44520 502380 44560
rect 516318 44520 516324 44532
rect 502352 44492 516324 44520
rect 516318 44480 516324 44492
rect 516376 44480 516382 44532
rect 304592 44424 342300 44452
rect 304592 44412 304598 44424
rect 414198 44412 414204 44464
rect 414256 44452 414262 44464
rect 419810 44452 419816 44464
rect 414256 44424 419816 44452
rect 414256 44412 414262 44424
rect 419810 44412 419816 44424
rect 419868 44412 419874 44464
rect 143626 44344 143632 44396
rect 143684 44384 143690 44396
rect 145098 44384 145104 44396
rect 143684 44356 145104 44384
rect 143684 44344 143690 44356
rect 145098 44344 145104 44356
rect 145156 44384 145162 44396
rect 195330 44384 195336 44396
rect 145156 44356 195336 44384
rect 145156 44344 145162 44356
rect 195330 44344 195336 44356
rect 195388 44384 195394 44396
rect 199654 44384 199660 44396
rect 195388 44356 199660 44384
rect 195388 44344 195394 44356
rect 199654 44344 199660 44356
rect 199712 44344 199718 44396
rect 200850 44344 200856 44396
rect 200908 44384 200914 44396
rect 241330 44384 241336 44396
rect 200908 44356 241336 44384
rect 200908 44344 200914 44356
rect 241330 44344 241336 44356
rect 241388 44384 241394 44396
rect 251082 44384 251088 44396
rect 241388 44356 251088 44384
rect 241388 44344 241394 44356
rect 251082 44344 251088 44356
rect 251140 44344 251146 44396
rect 306374 44344 306380 44396
rect 306432 44384 306438 44396
rect 309410 44384 309416 44396
rect 306432 44356 309416 44384
rect 306432 44344 306438 44356
rect 309410 44344 309416 44356
rect 309468 44384 309474 44396
rect 352558 44384 352564 44396
rect 309468 44356 352564 44384
rect 309468 44344 309474 44356
rect 352558 44344 352564 44356
rect 352616 44384 352622 44396
rect 355410 44384 355416 44396
rect 352616 44356 355416 44384
rect 352616 44344 352622 44356
rect 355410 44344 355416 44356
rect 355468 44344 355474 44396
rect 359366 44344 359372 44396
rect 359424 44384 359430 44396
rect 360654 44384 360660 44396
rect 359424 44356 360660 44384
rect 359424 44344 359430 44356
rect 360654 44344 360660 44356
rect 360712 44344 360718 44396
rect 364242 44344 364248 44396
rect 364300 44384 364306 44396
rect 407390 44384 407396 44396
rect 364300 44356 407396 44384
rect 364300 44344 364306 44356
rect 407390 44344 407396 44356
rect 407448 44384 407454 44396
rect 410426 44384 410432 44396
rect 407448 44356 410432 44384
rect 407448 44344 407454 44356
rect 410426 44344 410432 44356
rect 410484 44344 410490 44396
rect 419074 44344 419080 44396
rect 419132 44384 419138 44396
rect 462130 44384 462136 44396
rect 419132 44356 462136 44384
rect 419132 44344 419138 44356
rect 462130 44344 462136 44356
rect 462188 44384 462194 44396
rect 465166 44384 465172 44396
rect 462188 44356 465172 44384
rect 462188 44344 462194 44356
rect 465166 44344 465172 44356
rect 465224 44344 465230 44396
rect 473814 44344 473820 44396
rect 473872 44384 473878 44396
rect 516962 44384 516968 44396
rect 473872 44356 516968 44384
rect 473872 44344 473878 44356
rect 516962 44344 516968 44356
rect 517020 44384 517026 44396
rect 519998 44384 520004 44396
rect 517020 44356 520004 44384
rect 517020 44344 517026 44356
rect 519998 44344 520004 44356
rect 520056 44344 520062 44396
rect 188522 44276 188528 44328
rect 188580 44316 188586 44328
rect 192846 44316 192852 44328
rect 188580 44288 192852 44316
rect 188580 44276 188586 44288
rect 192846 44276 192852 44288
rect 192904 44316 192910 44328
rect 201494 44316 201500 44328
rect 192904 44288 201500 44316
rect 192904 44276 192910 44288
rect 201494 44276 201500 44288
rect 201552 44316 201558 44328
rect 297082 44316 297088 44328
rect 201552 44288 297088 44316
rect 201552 44276 201558 44288
rect 297082 44276 297088 44288
rect 297140 44316 297146 44328
rect 299566 44316 299572 44328
rect 297140 44288 299572 44316
rect 297140 44276 297146 44288
rect 299566 44276 299572 44288
rect 299624 44316 299630 44328
rect 305730 44316 305736 44328
rect 299624 44288 305736 44316
rect 299624 44276 299630 44288
rect 305730 44276 305736 44288
rect 305788 44316 305794 44328
rect 351914 44316 351920 44328
rect 305788 44288 351920 44316
rect 305788 44276 305794 44288
rect 351914 44276 351920 44288
rect 351972 44316 351978 44328
rect 354398 44316 354404 44328
rect 351972 44288 354404 44316
rect 351972 44276 351978 44288
rect 354398 44276 354404 44288
rect 354456 44276 354462 44328
rect 358722 44316 358728 44328
rect 355520 44288 358728 44316
rect 199654 44208 199660 44260
rect 199712 44248 199718 44260
rect 303890 44248 303896 44260
rect 199712 44220 303896 44248
rect 199712 44208 199718 44220
rect 303890 44208 303896 44220
rect 303948 44248 303954 44260
rect 308214 44248 308220 44260
rect 303948 44220 308220 44248
rect 303948 44208 303954 44220
rect 308214 44208 308220 44220
rect 308272 44248 308278 44260
rect 355520 44248 355548 44288
rect 358722 44276 358728 44288
rect 358780 44276 358786 44328
rect 360562 44276 360568 44328
rect 360620 44316 360626 44328
rect 399662 44316 399668 44328
rect 360620 44288 399668 44316
rect 360620 44276 360626 44288
rect 399662 44276 399668 44288
rect 399720 44276 399726 44328
rect 413554 44316 413560 44328
rect 399772 44288 413560 44316
rect 308272 44220 355548 44248
rect 308272 44208 308278 44220
rect 355594 44208 355600 44260
rect 355652 44248 355658 44260
rect 359918 44248 359924 44260
rect 355652 44220 359924 44248
rect 355652 44208 355658 44220
rect 359918 44208 359924 44220
rect 359976 44208 359982 44260
rect 363046 44208 363052 44260
rect 363104 44248 363110 44260
rect 399772 44248 399800 44288
rect 413554 44276 413560 44288
rect 413612 44316 413618 44328
rect 417878 44316 417884 44328
rect 413612 44288 417884 44316
rect 413612 44276 413618 44288
rect 417878 44276 417884 44288
rect 417936 44316 417942 44328
rect 468294 44316 468300 44328
rect 417936 44288 468300 44316
rect 417936 44276 417942 44288
rect 468294 44276 468300 44288
rect 468352 44316 468358 44328
rect 472618 44316 472624 44328
rect 468352 44288 472624 44316
rect 468352 44276 468358 44288
rect 472618 44276 472624 44288
rect 472676 44316 472682 44328
rect 523126 44316 523132 44328
rect 472676 44288 523132 44316
rect 472676 44276 472682 44288
rect 523126 44276 523132 44288
rect 523184 44276 523190 44328
rect 363104 44220 399800 44248
rect 363104 44208 363110 44220
rect 411070 44208 411076 44260
rect 411128 44248 411134 44260
rect 419718 44248 419724 44260
rect 411128 44220 419724 44248
rect 411128 44208 411134 44220
rect 419718 44208 419724 44220
rect 419776 44208 419782 44260
rect 419810 44208 419816 44260
rect 419868 44248 419874 44260
rect 468938 44248 468944 44260
rect 419868 44220 468944 44248
rect 419868 44208 419874 44220
rect 468938 44208 468944 44220
rect 468996 44248 469002 44260
rect 523770 44248 523776 44260
rect 468996 44220 523776 44248
rect 468996 44208 469002 44220
rect 523770 44208 523776 44220
rect 523828 44208 523834 44260
rect 358722 44140 358728 44192
rect 358780 44180 358786 44192
rect 363064 44180 363092 44208
rect 358780 44152 363092 44180
rect 358780 44140 358786 44152
rect 523126 44140 523132 44192
rect 523184 44180 523190 44192
rect 527450 44180 527456 44192
rect 523184 44152 527456 44180
rect 523184 44140 523190 44152
rect 527450 44140 527456 44152
rect 527508 44140 527514 44192
rect 576762 42712 576768 42764
rect 576820 42752 576826 42764
rect 673454 42752 673460 42764
rect 576820 42724 673460 42752
rect 576820 42712 576826 42724
rect 673454 42712 673460 42724
rect 673512 42712 673518 42764
rect 251082 42032 251088 42084
rect 251140 42072 251146 42084
rect 255222 42072 255228 42084
rect 251140 42044 255228 42072
rect 251140 42032 251146 42044
rect 255222 42032 255228 42044
rect 255280 42032 255286 42084
rect 146294 41964 146300 42016
rect 146352 42004 146358 42016
rect 569126 42004 569132 42016
rect 146352 41976 569132 42004
rect 146352 41964 146358 41976
rect 569126 41964 569132 41976
rect 569184 42004 569190 42016
rect 576762 42004 576768 42016
rect 569184 41976 576768 42004
rect 569184 41964 569190 41976
rect 576762 41964 576768 41976
rect 576820 41964 576826 42016
rect 187694 41896 187700 41948
rect 187752 41936 187758 41948
rect 188430 41936 188436 41948
rect 187752 41908 188436 41936
rect 187752 41896 187758 41908
rect 188430 41896 188436 41908
rect 188488 41896 188494 41948
rect 198918 41896 198924 41948
rect 198976 41936 198982 41948
rect 307478 41936 307484 41948
rect 198976 41908 307484 41936
rect 198976 41896 198982 41908
rect 198458 41828 198464 41880
rect 198516 41868 198522 41880
rect 200114 41868 200120 41880
rect 198516 41840 200120 41868
rect 198516 41828 198522 41840
rect 200114 41828 200120 41840
rect 200172 41828 200178 41880
rect 255222 41828 255228 41880
rect 255280 41868 255286 41880
rect 297634 41868 297640 41880
rect 255280 41840 297640 41868
rect 255280 41828 255286 41840
rect 297634 41828 297640 41840
rect 297692 41868 297698 41880
rect 300670 41868 300676 41880
rect 297692 41840 300676 41868
rect 297692 41828 297698 41840
rect 300670 41828 300676 41840
rect 300728 41828 300734 41880
rect 149606 41760 149612 41812
rect 149664 41800 149670 41812
rect 187694 41800 187700 41812
rect 149664 41772 187700 41800
rect 149664 41760 149670 41772
rect 187694 41760 187700 41772
rect 187752 41760 187758 41812
rect 189258 41760 189264 41812
rect 189316 41800 189322 41812
rect 191098 41800 191104 41812
rect 189316 41772 191104 41800
rect 189316 41760 189322 41772
rect 191098 41760 191104 41772
rect 191156 41800 191162 41812
rect 192294 41800 192300 41812
rect 191156 41772 192300 41800
rect 191156 41760 191162 41772
rect 192294 41760 192300 41772
rect 192352 41800 192358 41812
rect 193582 41800 193588 41812
rect 192352 41772 193588 41800
rect 192352 41760 192358 41772
rect 193582 41760 193588 41772
rect 193640 41800 193646 41812
rect 196434 41800 196440 41812
rect 193640 41772 196440 41800
rect 193640 41760 193646 41772
rect 196434 41760 196440 41772
rect 196492 41760 196498 41812
rect 198826 41800 198832 41812
rect 198752 41772 198832 41800
rect 168282 41732 168288 41744
rect 160020 41704 168288 41732
rect 160020 41664 160048 41704
rect 168282 41692 168288 41704
rect 168340 41692 168346 41744
rect 154500 41636 160048 41664
rect 93762 41556 93768 41608
rect 93820 41596 93826 41608
rect 93820 41568 102180 41596
rect 93820 41556 93826 41568
rect 102152 41528 102180 41568
rect 121546 41556 121552 41608
rect 121604 41596 121610 41608
rect 121604 41568 135300 41596
rect 121604 41556 121610 41568
rect 121270 41528 121276 41540
rect 102152 41500 121276 41528
rect 121270 41488 121276 41500
rect 121328 41488 121334 41540
rect 135272 41528 135300 41568
rect 140866 41556 140872 41608
rect 140924 41596 140930 41608
rect 154500 41596 154528 41636
rect 140924 41568 154528 41596
rect 140924 41556 140930 41568
rect 140682 41528 140688 41540
rect 135272 41500 140688 41528
rect 140682 41488 140688 41500
rect 140740 41488 140746 41540
rect 168282 41488 168288 41540
rect 168340 41528 168346 41540
rect 198752 41528 198780 41772
rect 198826 41760 198832 41772
rect 198884 41760 198890 41812
rect 168340 41500 198780 41528
rect 168340 41488 168346 41500
rect 144638 40740 144644 40792
rect 144696 40780 144702 40792
rect 146294 40780 146300 40792
rect 144696 40752 146300 40780
rect 144696 40740 144702 40752
rect 146294 40740 146300 40752
rect 146352 40740 146358 40792
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143074 40100 143080 40112
rect 141048 40072 143080 40100
rect 141048 40060 141054 40072
rect 142586 40000 142614 40072
rect 143074 40060 143080 40072
rect 143132 40100 143138 40112
rect 144638 40100 144644 40112
rect 143132 40072 144644 40100
rect 143132 40060 143138 40072
rect 144638 40060 144644 40072
rect 144696 40060 144702 40112
rect 142573 38005 142619 40000
rect 145091 39934 145143 40000
rect 302234 41760 302240 41812
rect 302292 41800 302298 41812
rect 304994 41800 305000 41812
rect 302292 41772 305000 41800
rect 302292 41760 302298 41772
rect 304994 41760 305000 41772
rect 305052 41800 305058 41812
rect 306282 41800 306288 41812
rect 305052 41772 306288 41800
rect 305052 41760 305058 41772
rect 306282 41760 306288 41772
rect 306340 41760 306346 41812
rect 307404 41732 307432 41908
rect 307478 41896 307484 41908
rect 307536 41896 307542 41948
rect 362494 41896 362500 41948
rect 362552 41936 362558 41948
rect 367094 41936 367100 41948
rect 362552 41908 367100 41936
rect 362552 41896 362558 41908
rect 367094 41896 367100 41908
rect 367152 41896 367158 41948
rect 360010 41828 360016 41880
rect 360068 41868 360074 41880
rect 361114 41868 361120 41880
rect 360068 41840 361120 41868
rect 360068 41828 360074 41840
rect 361114 41828 361120 41840
rect 361172 41868 361178 41880
rect 363506 41868 363512 41880
rect 361172 41840 363512 41868
rect 361172 41828 361178 41840
rect 363506 41828 363512 41840
rect 363564 41828 363570 41880
rect 410518 41828 410524 41880
rect 410576 41868 410582 41880
rect 411806 41868 411812 41880
rect 410576 41840 411812 41868
rect 410576 41828 410582 41840
rect 411806 41828 411812 41840
rect 411864 41868 411870 41880
rect 414842 41868 414848 41880
rect 411864 41840 414848 41868
rect 411864 41828 411870 41840
rect 414842 41828 414848 41840
rect 414900 41868 414906 41880
rect 416130 41868 416136 41880
rect 414900 41840 416136 41868
rect 414900 41828 414906 41840
rect 416130 41828 416136 41840
rect 416188 41868 416194 41880
rect 418522 41868 418528 41880
rect 416188 41840 418528 41868
rect 416188 41828 416194 41840
rect 418522 41828 418528 41840
rect 418580 41828 418586 41880
rect 464154 41828 464160 41880
rect 464212 41868 464218 41880
rect 467190 41868 467196 41880
rect 464212 41840 467196 41868
rect 464212 41828 464218 41840
rect 467190 41828 467196 41840
rect 467248 41868 467254 41880
rect 470042 41868 470048 41880
rect 467248 41840 470048 41868
rect 467248 41828 467254 41840
rect 470042 41828 470048 41840
rect 470100 41828 470106 41880
rect 470962 41868 470968 41880
rect 470152 41840 470968 41868
rect 409322 41760 409328 41812
rect 409380 41800 409386 41812
rect 412358 41800 412364 41812
rect 409380 41772 412364 41800
rect 409380 41760 409386 41772
rect 412358 41760 412364 41772
rect 412416 41800 412422 41812
rect 415210 41800 415216 41812
rect 412416 41772 415216 41800
rect 412416 41760 412422 41772
rect 415210 41760 415216 41772
rect 415268 41760 415274 41812
rect 417050 41760 417056 41812
rect 417108 41800 417114 41812
rect 417108 41772 417280 41800
rect 417108 41760 417114 41772
rect 307404 41704 309180 41732
rect 309152 41664 309180 41704
rect 314562 41664 314568 41676
rect 309152 41636 314568 41664
rect 314562 41624 314568 41636
rect 314620 41624 314626 41676
rect 314654 41624 314660 41676
rect 314712 41664 314718 41676
rect 314712 41636 328408 41664
rect 314712 41624 314718 41636
rect 328380 41596 328408 41636
rect 386322 41624 386328 41676
rect 386380 41664 386386 41676
rect 417252 41664 417280 41772
rect 465350 41760 465356 41812
rect 465408 41800 465414 41812
rect 466362 41800 466368 41812
rect 465408 41772 466368 41800
rect 465408 41760 465414 41772
rect 466362 41760 466368 41772
rect 466420 41800 466426 41812
rect 469674 41800 469680 41812
rect 466420 41772 469680 41800
rect 466420 41760 466426 41772
rect 469674 41760 469680 41772
rect 469732 41800 469738 41812
rect 470152 41800 470180 41840
rect 470962 41828 470968 41840
rect 471020 41868 471026 41880
rect 473078 41868 473084 41880
rect 471020 41840 473084 41868
rect 471020 41828 471026 41840
rect 473078 41828 473084 41840
rect 473136 41828 473142 41880
rect 520090 41828 520096 41880
rect 520148 41868 520154 41880
rect 521194 41868 521200 41880
rect 520148 41840 521200 41868
rect 520148 41828 520154 41840
rect 521194 41828 521200 41840
rect 521252 41868 521258 41880
rect 524230 41868 524236 41880
rect 521252 41840 524236 41868
rect 521252 41828 521258 41840
rect 524230 41828 524236 41840
rect 524288 41868 524294 41880
rect 525518 41868 525524 41880
rect 524288 41840 525524 41868
rect 524288 41828 524294 41840
rect 525518 41828 525524 41840
rect 525576 41868 525582 41880
rect 527910 41868 527916 41880
rect 525576 41840 527916 41868
rect 525576 41828 525582 41840
rect 527910 41828 527916 41840
rect 527968 41828 527974 41880
rect 469732 41772 470180 41800
rect 469732 41760 469738 41772
rect 471882 41760 471888 41812
rect 471940 41800 471946 41812
rect 471940 41772 472112 41800
rect 471940 41760 471946 41772
rect 472084 41664 472112 41772
rect 526714 41760 526720 41812
rect 526772 41760 526778 41812
rect 386380 41636 391888 41664
rect 386380 41624 386386 41636
rect 349614 41596 349620 41608
rect 328380 41568 333928 41596
rect 333900 41528 333928 41568
rect 333992 41568 349620 41596
rect 333992 41528 334020 41568
rect 349614 41556 349620 41568
rect 349672 41556 349678 41608
rect 333900 41500 334020 41528
rect 391860 41460 391888 41636
rect 417252 41636 430528 41664
rect 417252 41460 417280 41636
rect 430500 41528 430528 41636
rect 472084 41636 488488 41664
rect 472084 41528 472112 41636
rect 488460 41596 488488 41636
rect 488460 41568 502380 41596
rect 430500 41500 472112 41528
rect 502352 41528 502380 41568
rect 507854 41556 507860 41608
rect 507912 41596 507918 41608
rect 507912 41568 521608 41596
rect 507912 41556 507918 41568
rect 507762 41528 507768 41540
rect 502352 41500 507768 41528
rect 507762 41488 507768 41500
rect 507820 41488 507826 41540
rect 521580 41528 521608 41568
rect 526732 41528 526760 41760
rect 521580 41500 526760 41528
rect 391860 41432 417280 41460
<< via1 >>
rect 585048 992196 585100 992248
rect 674748 992196 674800 992248
rect 78864 990768 78916 990820
rect 130292 990768 130344 990820
rect 89996 990700 90048 990752
rect 141424 990700 141476 990752
rect 192852 990700 192904 990752
rect 130292 990632 130344 990684
rect 181720 990632 181772 990684
rect 233056 990768 233108 990820
rect 284668 990768 284720 990820
rect 286968 990768 287020 990820
rect 345112 990768 345164 990820
rect 372528 990768 372580 990820
rect 372620 990768 372672 990820
rect 194968 990700 195020 990752
rect 244188 990700 244240 990752
rect 295800 990700 295852 990752
rect 121276 990564 121328 990616
rect 160192 990428 160244 990480
rect 192852 990428 192904 990480
rect 194968 990428 195020 990480
rect 173900 990360 173952 990412
rect 182456 990360 182508 990412
rect 233700 990632 233752 990684
rect 285312 990632 285364 990684
rect 342168 990632 342220 990684
rect 345020 990632 345072 990684
rect 397460 990768 397512 990820
rect 397644 990768 397696 990820
rect 486608 990768 486660 990820
rect 538036 990768 538088 990820
rect 639788 990768 639840 990820
rect 400128 990700 400180 990752
rect 419540 990700 419592 990752
rect 438768 990700 438820 990752
rect 458180 990700 458232 990752
rect 477408 990700 477460 990752
rect 527548 990700 527600 990752
rect 629300 990700 629352 990752
rect 631232 990700 631284 990752
rect 386420 990632 386472 990684
rect 386512 990632 386564 990684
rect 475476 990632 475528 990684
rect 526904 990632 526956 990684
rect 626540 990632 626592 990684
rect 286968 990564 287020 990616
rect 295800 990496 295852 990548
rect 397460 990496 397512 990548
rect 419540 990496 419592 990548
rect 438768 990496 438820 990548
rect 458180 990496 458232 990548
rect 476120 990496 476172 990548
rect 477408 990496 477460 990548
rect 386420 990428 386472 990480
rect 387156 990428 387208 990480
rect 400128 990428 400180 990480
rect 42248 990156 42300 990208
rect 78864 990156 78916 990208
rect 42340 990088 42392 990140
rect 79508 990088 79560 990140
rect 131028 990224 131080 990276
rect 140688 990292 140740 990344
rect 140780 990224 140832 990276
rect 160008 990292 160060 990344
rect 173900 990224 173952 990276
rect 639788 990156 639840 990208
rect 673644 990156 673696 990208
rect 89904 990088 89956 990140
rect 626540 990088 626592 990140
rect 628656 990088 628708 990140
rect 631232 990088 631284 990140
rect 673552 990088 673604 990140
rect 42524 990020 42576 990072
rect 673460 990020 673512 990072
rect 41788 968464 41840 968516
rect 42524 968464 42576 968516
rect 673460 965268 673512 965320
rect 675392 965268 675444 965320
rect 673552 964724 673604 964776
rect 675392 964724 675444 964776
rect 41788 958060 41840 958112
rect 42340 958060 42392 958112
rect 42248 957720 42300 957772
rect 42248 957516 42300 957568
rect 673644 953300 673696 953352
rect 675392 953300 675444 953352
rect 673460 875168 673512 875220
rect 675392 875168 675444 875220
rect 673552 874488 673604 874540
rect 675392 874488 675444 874540
rect 673644 864424 673696 864476
rect 675392 864424 675444 864476
rect 675300 818320 675352 818372
rect 677508 818320 677560 818372
rect 41788 797716 41840 797768
rect 42524 797716 42576 797768
rect 42708 797716 42760 797768
rect 41788 787244 41840 787296
rect 42616 787244 42668 787296
rect 41788 786632 41840 786684
rect 42524 786632 42576 786684
rect 673460 786564 673512 786616
rect 674012 786564 674064 786616
rect 675392 786564 675444 786616
rect 673552 786360 673604 786412
rect 675392 786360 675444 786412
rect 675300 781600 675352 781652
rect 675300 781396 675352 781448
rect 673460 774868 673512 774920
rect 673644 774868 673696 774920
rect 675392 774868 675444 774920
rect 673736 772760 673788 772812
rect 674012 772760 674064 772812
rect 42432 767320 42484 767372
rect 42708 767320 42760 767372
rect 42524 758956 42576 759008
rect 42800 758956 42852 759008
rect 41788 754468 41840 754520
rect 42432 754468 42484 754520
rect 673736 753516 673788 753568
rect 673920 753516 673972 753568
rect 42524 753448 42576 753500
rect 42800 753448 42852 753500
rect 41788 744132 41840 744184
rect 42340 744132 42392 744184
rect 42616 744132 42668 744184
rect 41788 743996 41840 744048
rect 42524 743996 42576 744048
rect 42984 743996 43036 744048
rect 673644 741956 673696 742008
rect 673920 741956 673972 742008
rect 675392 741888 675444 741940
rect 673552 740664 673604 740716
rect 675392 740664 675444 740716
rect 673644 739780 673696 739832
rect 673644 739644 673696 739696
rect 42340 739576 42392 739628
rect 42616 739576 42668 739628
rect 42524 734136 42576 734188
rect 42984 734136 43036 734188
rect 673460 730124 673512 730176
rect 675392 730124 675444 730176
rect 42524 720332 42576 720384
rect 42892 720332 42944 720384
rect 41788 711288 41840 711340
rect 42432 711288 42484 711340
rect 42708 711288 42760 711340
rect 673644 701020 673696 701072
rect 673828 701020 673880 701072
rect 41788 700952 41840 701004
rect 42616 700952 42668 701004
rect 41788 700816 41840 700868
rect 42892 700816 42944 700868
rect 675392 695920 675444 695972
rect 673644 695852 673696 695904
rect 42432 695512 42484 695564
rect 42892 695512 42944 695564
rect 673552 695308 673604 695360
rect 675392 695308 675444 695360
rect 673460 685176 673512 685228
rect 675392 685176 675444 685228
rect 42432 681640 42484 681692
rect 42800 681572 42852 681624
rect 42616 678512 42668 678564
rect 42984 678512 43036 678564
rect 42432 676132 42484 676184
rect 42984 676132 43036 676184
rect 41788 669060 41840 669112
rect 42524 669060 42576 669112
rect 41788 658656 41840 658708
rect 42432 658656 42484 658708
rect 42708 658656 42760 658708
rect 41788 658044 41840 658096
rect 42800 658044 42852 658096
rect 673644 651720 673696 651772
rect 675392 651720 675444 651772
rect 42432 651380 42484 651432
rect 42800 651380 42852 651432
rect 673552 651108 673604 651160
rect 675392 651108 675444 651160
rect 675208 646008 675260 646060
rect 675300 645736 675352 645788
rect 673460 639684 673512 639736
rect 673920 639684 673972 639736
rect 675392 639684 675444 639736
rect 42524 632000 42576 632052
rect 42708 632000 42760 632052
rect 42984 632000 43036 632052
rect 42800 631864 42852 631916
rect 41788 624928 41840 624980
rect 42800 624928 42852 624980
rect 41788 615476 41840 615528
rect 42984 615476 43036 615528
rect 41788 614796 41840 614848
rect 42524 614796 42576 614848
rect 42800 612824 42852 612876
rect 42616 612756 42668 612808
rect 42616 612620 42668 612672
rect 42800 612620 42852 612672
rect 673644 606704 673696 606756
rect 675392 606704 675444 606756
rect 673552 606160 673604 606212
rect 675024 606160 675076 606212
rect 675392 606160 675444 606212
rect 673644 594872 673696 594924
rect 673920 594872 673972 594924
rect 675392 594872 675444 594924
rect 673736 594736 673788 594788
rect 675024 594736 675076 594788
rect 675300 593376 675352 593428
rect 675300 593172 675352 593224
rect 673552 585148 673604 585200
rect 673828 585148 673880 585200
rect 41788 582632 41840 582684
rect 42800 582632 42852 582684
rect 673736 575424 673788 575476
rect 674380 575424 674432 575476
rect 42340 574064 42392 574116
rect 42800 574064 42852 574116
rect 41788 571208 41840 571260
rect 42800 571208 42852 571260
rect 41788 570664 41840 570716
rect 42524 570664 42576 570716
rect 42708 570664 42760 570716
rect 673552 560532 673604 560584
rect 673828 560532 673880 560584
rect 675392 560532 675444 560584
rect 674012 559920 674064 559972
rect 674380 559920 674432 559972
rect 675392 559920 675444 559972
rect 42616 554752 42668 554804
rect 42800 554752 42852 554804
rect 673644 550468 673696 550520
rect 675392 550468 675444 550520
rect 673552 546388 673604 546440
rect 673828 546320 673880 546372
rect 41788 539452 41840 539504
rect 42524 539452 42576 539504
rect 41788 528028 41840 528080
rect 42616 528028 42668 528080
rect 41788 527484 41840 527536
rect 42432 527484 42484 527536
rect 42708 527484 42760 527536
rect 675300 513748 675352 513800
rect 677692 513748 677744 513800
rect 673736 502324 673788 502376
rect 673920 502324 673972 502376
rect 673552 498176 673604 498228
rect 673828 498176 673880 498228
rect 673828 469276 673880 469328
rect 673736 469140 673788 469192
rect 673736 463632 673788 463684
rect 674012 463632 674064 463684
rect 673552 449556 673604 449608
rect 673828 449556 673880 449608
rect 42616 444320 42668 444372
rect 42800 444320 42852 444372
rect 673736 444320 673788 444372
rect 674012 444320 674064 444372
rect 42708 441532 42760 441584
rect 42800 441532 42852 441584
rect 674748 427796 674800 427848
rect 677124 427796 677176 427848
rect 42616 422288 42668 422340
rect 42708 422288 42760 422340
rect 673644 420724 673696 420776
rect 673828 420724 673880 420776
rect 41788 411204 41840 411256
rect 42524 411204 42576 411256
rect 42616 405696 42668 405748
rect 42892 405696 42944 405748
rect 673828 401548 673880 401600
rect 675300 401548 675352 401600
rect 41788 401344 41840 401396
rect 42892 401344 42944 401396
rect 41788 400800 41840 400852
rect 42432 400800 42484 400852
rect 42616 386316 42668 386368
rect 42892 386316 42944 386368
rect 673736 384276 673788 384328
rect 675392 384276 675444 384328
rect 673644 383188 673696 383240
rect 675300 383188 675352 383240
rect 673552 380876 673604 380928
rect 673736 380876 673788 380928
rect 42800 372580 42852 372632
rect 42984 372580 43036 372632
rect 673736 372308 673788 372360
rect 675392 372308 675444 372360
rect 41788 368636 41840 368688
rect 42892 368636 42944 368688
rect 42524 367820 42576 367872
rect 42800 367820 42852 367872
rect 41788 358232 41840 358284
rect 42524 358232 42576 358284
rect 41788 357620 41840 357672
rect 42432 357620 42484 357672
rect 42616 357620 42668 357672
rect 673552 338104 673604 338156
rect 675392 338104 675444 338156
rect 673644 337492 673696 337544
rect 675392 337492 675444 337544
rect 673736 328040 673788 328092
rect 675392 328040 675444 328092
rect 41788 325456 41840 325508
rect 42432 325456 42484 325508
rect 42708 325456 42760 325508
rect 42432 322872 42484 322924
rect 42616 322804 42668 322856
rect 42708 322804 42760 322856
rect 42892 322736 42944 322788
rect 42340 314168 42392 314220
rect 42708 314168 42760 314220
rect 41788 314032 41840 314084
rect 42524 314032 42576 314084
rect 42708 314032 42760 314084
rect 41788 313488 41840 313540
rect 42800 313420 42852 313472
rect 673552 303560 673604 303612
rect 675300 303560 675352 303612
rect 673644 293564 673696 293616
rect 673920 293564 673972 293616
rect 675392 293564 675444 293616
rect 673644 293428 673696 293480
rect 675300 293428 675352 293480
rect 41788 282276 41840 282328
rect 42524 282276 42576 282328
rect 673736 282072 673788 282124
rect 675392 282072 675444 282124
rect 41788 271872 41840 271924
rect 42708 271872 42760 271924
rect 41788 271192 41840 271244
rect 42524 271192 42576 271244
rect 42800 271192 42852 271244
rect 673460 264936 673512 264988
rect 673644 264936 673696 264988
rect 673460 248684 673512 248736
rect 675300 248684 675352 248736
rect 673644 247460 673696 247512
rect 673920 247460 673972 247512
rect 675392 247460 675444 247512
rect 42340 245556 42392 245608
rect 42892 245556 42944 245608
rect 42524 245488 42576 245540
rect 42800 245488 42852 245540
rect 673828 243788 673880 243840
rect 675300 243788 675352 243840
rect 41788 238076 41840 238128
rect 42616 238076 42668 238128
rect 42892 238076 42944 238128
rect 673920 237668 673972 237720
rect 675392 237668 675444 237720
rect 673920 237328 673972 237380
rect 674104 237328 674156 237380
rect 42340 232840 42392 232892
rect 42616 232840 42668 232892
rect 674104 231752 674156 231804
rect 674288 231752 674340 231804
rect 41788 228624 41840 228676
rect 42708 228624 42760 228676
rect 41788 228012 41840 228064
rect 42616 228012 42668 228064
rect 42800 228012 42852 228064
rect 673828 218084 673880 218136
rect 673828 217948 673880 218000
rect 673736 212508 673788 212560
rect 673828 212508 673880 212560
rect 674012 212508 674064 212560
rect 674288 212508 674340 212560
rect 42340 208360 42392 208412
rect 42892 208360 42944 208412
rect 673736 203872 673788 203924
rect 675392 203872 675444 203924
rect 673644 203328 673696 203380
rect 675392 203328 675444 203380
rect 674012 198704 674064 198756
rect 675208 198704 675260 198756
rect 41788 194896 41840 194948
rect 42432 194896 42484 194948
rect 42892 194896 42944 194948
rect 674748 192108 674800 192160
rect 675208 192108 675260 192160
rect 675392 192108 675444 192160
rect 41788 185444 41840 185496
rect 42340 185444 42392 185496
rect 42708 185444 42760 185496
rect 42432 185308 42484 185360
rect 42708 185308 42760 185360
rect 41788 184832 41840 184884
rect 42432 184832 42484 184884
rect 42616 184832 42668 184884
rect 673828 173884 673880 173936
rect 674748 173884 674800 173936
rect 673552 158312 673604 158364
rect 675392 158312 675444 158364
rect 673460 157292 673512 157344
rect 675392 157292 675444 157344
rect 42524 149064 42576 149116
rect 42708 149064 42760 149116
rect 673644 147092 673696 147144
rect 675024 147092 675076 147144
rect 675392 147092 675444 147144
rect 674012 140632 674064 140684
rect 675024 140632 675076 140684
rect 42248 121456 42300 121508
rect 44732 121456 44784 121508
rect 673828 115948 673880 116000
rect 674012 115948 674064 116000
rect 42984 115880 43036 115932
rect 44732 115880 44784 115932
rect 673828 115812 673880 115864
rect 675024 115812 675076 115864
rect 673552 112752 673604 112804
rect 675392 112752 675444 112804
rect 673460 112072 673512 112124
rect 675392 112072 675444 112124
rect 42524 110440 42576 110492
rect 42708 110440 42760 110492
rect 673644 102280 673696 102332
rect 675024 102280 675076 102332
rect 675392 102280 675444 102332
rect 44640 82832 44692 82884
rect 44824 82764 44876 82816
rect 42340 45704 42392 45756
rect 140964 45704 141016 45756
rect 42432 45636 42484 45688
rect 143632 45636 143684 45688
rect 42708 45568 42760 45620
rect 143540 45568 143592 45620
rect 527456 45568 527508 45620
rect 673552 45568 673604 45620
rect 44916 45500 44968 45552
rect 195980 45500 196032 45552
rect 516324 45500 516376 45552
rect 673644 45500 673696 45552
rect 405648 44752 405700 44804
rect 411260 44752 411312 44804
rect 195980 44412 196032 44464
rect 304540 44412 304592 44464
rect 359372 44684 359424 44736
rect 406752 44684 406804 44736
rect 425060 44684 425112 44736
rect 444196 44684 444248 44736
rect 425060 44548 425112 44600
rect 354404 44480 354456 44532
rect 360568 44480 360620 44532
rect 360660 44480 360712 44532
rect 386420 44480 386472 44532
rect 399668 44480 399720 44532
rect 406752 44480 406804 44532
rect 411260 44480 411312 44532
rect 444288 44480 444340 44532
rect 461492 44548 461544 44600
rect 469128 44548 469180 44600
rect 469220 44548 469272 44600
rect 483020 44616 483072 44668
rect 502248 44480 502300 44532
rect 516324 44480 516376 44532
rect 414204 44412 414256 44464
rect 419816 44412 419868 44464
rect 143632 44344 143684 44396
rect 145104 44344 145156 44396
rect 195336 44344 195388 44396
rect 199660 44344 199712 44396
rect 200856 44344 200908 44396
rect 241336 44344 241388 44396
rect 251088 44344 251140 44396
rect 306380 44344 306432 44396
rect 309416 44344 309468 44396
rect 352564 44344 352616 44396
rect 355416 44344 355468 44396
rect 359372 44344 359424 44396
rect 360660 44344 360712 44396
rect 364248 44344 364300 44396
rect 407396 44344 407448 44396
rect 410432 44344 410484 44396
rect 419080 44344 419132 44396
rect 462136 44344 462188 44396
rect 465172 44344 465224 44396
rect 473820 44344 473872 44396
rect 516968 44344 517020 44396
rect 520004 44344 520056 44396
rect 188528 44276 188580 44328
rect 192852 44276 192904 44328
rect 201500 44276 201552 44328
rect 297088 44276 297140 44328
rect 299572 44276 299624 44328
rect 305736 44276 305788 44328
rect 351920 44276 351972 44328
rect 354404 44276 354456 44328
rect 199660 44208 199712 44260
rect 303896 44208 303948 44260
rect 308220 44208 308272 44260
rect 358728 44276 358780 44328
rect 360568 44276 360620 44328
rect 399668 44276 399720 44328
rect 355600 44208 355652 44260
rect 359924 44208 359976 44260
rect 363052 44208 363104 44260
rect 413560 44276 413612 44328
rect 417884 44276 417936 44328
rect 468300 44276 468352 44328
rect 472624 44276 472676 44328
rect 523132 44276 523184 44328
rect 411076 44208 411128 44260
rect 419724 44208 419776 44260
rect 419816 44208 419868 44260
rect 468944 44208 468996 44260
rect 523776 44208 523828 44260
rect 358728 44140 358780 44192
rect 523132 44140 523184 44192
rect 527456 44140 527508 44192
rect 576768 42712 576820 42764
rect 673460 42712 673512 42764
rect 251088 42032 251140 42084
rect 255228 42032 255280 42084
rect 146300 41964 146352 42016
rect 569132 41964 569184 42016
rect 576768 41964 576820 42016
rect 187700 41896 187752 41948
rect 188436 41896 188488 41948
rect 198924 41896 198976 41948
rect 198464 41828 198516 41880
rect 200120 41828 200172 41880
rect 255228 41828 255280 41880
rect 297640 41828 297692 41880
rect 300676 41828 300728 41880
rect 149612 41760 149664 41812
rect 187700 41760 187752 41812
rect 189264 41760 189316 41812
rect 191104 41760 191156 41812
rect 192300 41760 192352 41812
rect 193588 41760 193640 41812
rect 196440 41760 196492 41812
rect 168288 41692 168340 41744
rect 93768 41556 93820 41608
rect 121552 41556 121604 41608
rect 121276 41488 121328 41540
rect 140872 41556 140924 41608
rect 140688 41488 140740 41540
rect 168288 41488 168340 41540
rect 198832 41760 198884 41812
rect 144644 40740 144696 40792
rect 146300 40740 146352 40792
rect 140996 40060 141048 40112
rect 143080 40060 143132 40112
rect 144644 40060 144696 40112
rect 302240 41760 302292 41812
rect 305000 41760 305052 41812
rect 306288 41760 306340 41812
rect 307484 41896 307536 41948
rect 362500 41896 362552 41948
rect 367100 41896 367152 41948
rect 360016 41828 360068 41880
rect 361120 41828 361172 41880
rect 363512 41828 363564 41880
rect 410524 41828 410576 41880
rect 411812 41828 411864 41880
rect 414848 41828 414900 41880
rect 416136 41828 416188 41880
rect 418528 41828 418580 41880
rect 464160 41828 464212 41880
rect 467196 41828 467248 41880
rect 470048 41828 470100 41880
rect 409328 41760 409380 41812
rect 412364 41760 412416 41812
rect 415216 41760 415268 41812
rect 417056 41760 417108 41812
rect 314568 41624 314620 41676
rect 314660 41624 314712 41676
rect 386328 41624 386380 41676
rect 465356 41760 465408 41812
rect 466368 41760 466420 41812
rect 469680 41760 469732 41812
rect 470968 41828 471020 41880
rect 473084 41828 473136 41880
rect 520096 41828 520148 41880
rect 521200 41828 521252 41880
rect 524236 41828 524288 41880
rect 525524 41828 525576 41880
rect 527916 41828 527968 41880
rect 471888 41760 471940 41812
rect 526720 41760 526772 41812
rect 349620 41556 349672 41608
rect 507860 41556 507912 41608
rect 507768 41488 507820 41540
<< obsm1 >>
rect 76171 996231 92229 1037600
rect 127571 996231 143629 1037600
rect 178971 996231 195029 1037600
rect 230371 996231 246429 1037600
rect 281971 996231 298029 1037600
rect 333437 998007 348124 1037545
rect 335807 997984 336070 998007
tri 336070 997984 336093 998007 sw
tri 347285 997984 347308 998007 se
rect 347308 997984 347536 998007
rect 335807 997794 347536 997984
rect 383771 996231 399829 1037600
rect 472771 996231 488829 1037600
rect 524171 996231 540229 1037600
rect 575637 998007 590324 1037545
rect 578007 997984 578270 998007
tri 578270 997984 578293 998007 sw
tri 589485 997984 589508 998007 se
rect 589508 997984 589736 998007
rect 578007 997794 589736 997984
rect 625971 996231 642029 1037600
rect 84010 995636 84074 995648
rect 91738 995636 91802 995648
rect 84010 995608 91802 995636
rect 84010 995596 84074 995608
rect 91738 995596 91802 995608
rect 238202 995636 238266 995648
rect 245930 995636 245994 995648
rect 238202 995608 245994 995636
rect 238202 995596 238266 995608
rect 245930 995596 245994 995608
rect 531958 995636 532022 995648
rect 539686 995636 539750 995648
rect 531958 995608 539750 995636
rect 531958 995596 532022 995608
rect 539686 995596 539750 995608
rect 135346 995500 135410 995512
rect 143166 995500 143230 995512
rect 135346 995472 143230 995500
rect 135346 995460 135410 995472
rect 143166 995460 143230 995472
rect 633802 995500 633866 995512
rect 641530 995500 641594 995512
rect 633802 995472 641594 995500
rect 633802 995460 633866 995472
rect 641530 995460 641594 995472
rect 289630 995296 289694 995308
rect 297634 995296 297698 995308
rect 289630 995268 297698 995296
rect 289630 995256 289694 995268
rect 297634 995256 297698 995268
rect 391474 995296 391538 995308
rect 399478 995296 399542 995308
rect 391474 995268 399542 995296
rect 391474 995256 391538 995268
rect 399478 995256 399542 995268
rect 480438 995296 480502 995308
rect 488442 995296 488506 995308
rect 480438 995268 488506 995296
rect 480438 995256 480502 995268
rect 488442 995256 488506 995268
rect 186682 990604 186746 990616
rect 194686 990604 194750 990616
rect 186682 990576 194750 990604
rect 186682 990564 186746 990576
rect 194686 990564 194750 990576
rect 0 954171 41369 970229
rect 41782 969388 41846 969400
rect 42426 969388 42490 969400
rect 41782 969360 42490 969388
rect 41782 969348 41846 969360
rect 42426 969348 42490 969360
rect 41782 962452 41846 962464
rect 42426 962452 42490 962464
rect 41782 962424 42490 962452
rect 41782 962412 41846 962424
rect 42426 962412 42490 962424
rect 676231 951571 717600 967629
rect 31928 929187 32702 929239
rect 31928 928387 40900 929187
tri 40900 928387 41700 929187 sw
rect 31928 927240 41700 928387
rect 31928 927049 32702 927240
rect 32 923313 39593 927000
rect 32 922707 39600 923313
rect 39756 922707 41700 927240
rect 32 916185 41700 922707
rect 678007 919269 717568 922576
rect 678000 918415 717568 919269
rect 32 915331 39600 916185
rect 32 912024 39593 915331
rect 675900 911893 717568 918415
rect 675900 907360 677844 911893
rect 678000 911287 717568 911893
rect 678007 907600 717568 911287
rect 684898 907360 685672 907551
rect 675900 906213 685672 907360
tri 675900 905413 676700 906213 ne
rect 676700 905413 685672 906213
rect 684898 905361 685672 905413
rect 55 883936 39593 884383
rect 55 883708 39806 883936
rect 55 872470 39593 883708
tri 39593 883685 39616 883708 ne
tri 39593 872470 39616 872493 se
rect 39616 872470 39806 883708
rect 55 872207 39806 872470
rect 55 871571 39593 872207
rect 55 870525 39774 871571
rect 55 869837 39593 870525
rect 673730 870176 673794 870188
rect 675386 870176 675450 870188
rect 673730 870148 675450 870176
rect 673730 870136 673794 870148
rect 675386 870136 675450 870148
rect 673730 863240 673794 863252
rect 675386 863240 675450 863252
rect 673730 863212 675450 863240
rect 673730 863200 673794 863212
rect 675386 863200 675450 863212
rect 676231 862371 717600 878429
rect 55 841736 39593 842324
rect 55 841508 39806 841736
rect 55 830270 39593 841508
tri 39593 841485 39616 841508 ne
tri 39593 830270 39616 830293 se
rect 39616 830270 39806 841508
rect 678007 832675 717545 833363
rect 677826 831629 717545 832675
rect 678007 830993 717545 831629
rect 55 830007 39806 830270
rect 677794 830730 717545 830993
rect 55 827637 39593 830007
rect 677794 819492 677984 830730
tri 677984 830707 678007 830730 nw
tri 677984 819492 678007 819515 sw
rect 678007 819492 717545 830730
rect 677794 819264 717545 819492
rect 678007 818817 717545 819264
rect 0 784371 41369 800429
rect 41782 799592 41846 799604
rect 42334 799592 42398 799604
rect 41782 799564 42398 799592
rect 41782 799552 41846 799564
rect 42334 799552 42398 799564
rect 41782 792588 41846 792600
rect 42334 792588 42398 792600
rect 41782 792560 42398 792588
rect 41782 792548 41846 792560
rect 42334 792548 42398 792560
rect 675202 774024 675266 774036
rect 675386 774024 675450 774036
rect 675202 773996 675450 774024
rect 675202 773984 675266 773996
rect 675386 773984 675450 773996
rect 676231 773171 717600 789229
rect 0 741171 41369 757229
rect 41782 756412 41846 756424
rect 42334 756412 42398 756424
rect 41782 756384 42398 756412
rect 41782 756372 41846 756384
rect 42334 756372 42398 756384
rect 41782 749408 41846 749420
rect 42334 749408 42398 749420
rect 41782 749380 42398 749408
rect 41782 749368 41846 749380
rect 42334 749368 42398 749380
rect 676231 728171 717600 744229
rect 0 697971 41369 714029
rect 41782 713164 41846 713176
rect 42334 713164 42398 713176
rect 41782 713136 42398 713164
rect 41782 713124 41846 713136
rect 42334 713124 42398 713136
rect 41782 706228 41846 706240
rect 42334 706228 42398 706240
rect 41782 706200 42398 706228
rect 41782 706188 41846 706200
rect 42334 706188 42398 706200
rect 676231 683171 717600 699229
rect 0 654771 41369 670829
rect 41782 669984 41846 669996
rect 42334 669984 42398 669996
rect 41782 669956 42398 669984
rect 41782 669944 41846 669956
rect 42334 669944 42398 669956
rect 41782 663048 41846 663060
rect 42334 663048 42398 663060
rect 41782 663020 42398 663048
rect 41782 663008 41846 663020
rect 42334 663008 42398 663020
rect 675202 638840 675266 638852
rect 675386 638840 675450 638852
rect 675202 638812 675450 638840
rect 675202 638800 675266 638812
rect 675386 638800 675450 638812
rect 676231 637971 717600 654029
rect 0 611571 41369 627629
rect 41782 626804 41846 626816
rect 42334 626804 42398 626816
rect 41782 626776 42398 626804
rect 41782 626764 41846 626776
rect 42334 626764 42398 626776
rect 41782 619800 41846 619812
rect 42334 619800 42398 619812
rect 41782 619772 42398 619800
rect 41782 619760 41846 619772
rect 42334 619760 42398 619772
rect 675202 600828 675266 600840
rect 675386 600828 675450 600840
rect 675202 600800 675450 600828
rect 675202 600788 675266 600800
rect 675386 600788 675450 600800
rect 676231 592971 717600 609029
rect 0 568371 41369 584429
rect 41782 583556 41846 583568
rect 42334 583556 42398 583568
rect 41782 583528 42398 583556
rect 41782 583516 41846 583528
rect 42334 583516 42398 583528
rect 41782 576620 41846 576632
rect 42334 576620 42398 576632
rect 41782 576592 42398 576620
rect 41782 576580 41846 576592
rect 42334 576580 42398 576592
rect 676231 547771 717600 563829
rect 0 525171 41369 541229
rect 41782 540376 41846 540388
rect 42334 540376 42398 540388
rect 41782 540348 42398 540376
rect 41782 540336 41846 540348
rect 42334 540336 42398 540348
rect 41782 533440 41846 533452
rect 42334 533440 42398 533452
rect 41782 533412 42398 533440
rect 41782 533400 41846 533412
rect 42334 533400 42398 533412
rect 678007 518075 717545 518763
rect 677826 517029 717545 518075
rect 678007 516393 717545 517029
rect 677794 516130 717545 516393
rect 677794 504892 677984 516130
tri 677984 516107 678007 516130 nw
tri 677984 504892 678007 504915 sw
rect 678007 504892 717545 516130
rect 677794 504664 717545 504892
rect 678007 504217 717545 504664
rect 55 497136 39593 497583
rect 55 496908 39806 497136
rect 55 485670 39593 496908
tri 39593 496885 39616 496908 ne
tri 39593 485670 39616 485693 se
rect 39616 485670 39806 496908
rect 55 485407 39806 485670
rect 55 484771 39593 485407
rect 55 483725 39774 484771
rect 55 483037 39593 483725
rect 678007 471469 717568 474776
rect 678000 470615 717568 471469
rect 675900 464093 717568 470615
rect 675900 459560 677844 464093
rect 678000 463487 717568 464093
rect 678007 459800 717568 463487
rect 684898 459560 685672 459751
rect 675900 458413 685672 459560
tri 675900 458039 676274 458413 ne
rect 676274 458039 685672 458413
rect 31928 457987 32702 458039
tri 676274 457987 676326 458039 ne
rect 676326 457987 685672 458039
rect 31928 457187 40900 457987
tri 40900 457187 41700 457987 sw
tri 676326 457613 676700 457987 ne
rect 676700 457613 685672 457987
rect 684898 457561 685672 457613
rect 31928 456040 41700 457187
rect 31928 455849 32702 456040
rect 32 452113 39593 455800
rect 32 451507 39600 452113
rect 39756 451507 41700 456040
rect 32 444985 41700 451507
rect 32 444131 39600 444985
rect 32 440824 39593 444131
rect 678007 428193 717545 430563
rect 677794 427930 717545 428193
rect 677794 416692 677984 427930
tri 677984 427907 678007 427930 nw
tri 677984 416692 678007 416715 sw
rect 678007 416692 717545 427930
rect 677794 416464 717545 416692
rect 678007 415876 717545 416464
rect 0 397571 41369 413629
rect 41782 412808 41846 412820
rect 42334 412808 42398 412820
rect 41782 412780 42398 412808
rect 41782 412768 41846 412780
rect 42334 412768 42398 412780
rect 41782 405804 41846 405816
rect 42334 405804 42398 405816
rect 41782 405776 42398 405804
rect 41782 405764 41846 405776
rect 42334 405764 42398 405776
rect 676231 370571 717600 386629
rect 0 354371 41369 370429
rect 41782 369560 41846 369572
rect 42334 369560 42398 369572
rect 41782 369532 42398 369560
rect 41782 369520 41846 369532
rect 42334 369520 42398 369532
rect 41782 362624 41846 362636
rect 42334 362624 42398 362636
rect 41782 362596 42398 362624
rect 41782 362584 41846 362596
rect 42334 362584 42398 362596
rect 0 311171 41369 327229
rect 41782 326380 41846 326392
rect 42334 326380 42398 326392
rect 41782 326352 42398 326380
rect 41782 326340 41846 326352
rect 42334 326340 42398 326352
rect 676231 325371 717600 341429
rect 41782 319444 41846 319456
rect 42334 319444 42398 319456
rect 41782 319416 42398 319444
rect 41782 319404 41846 319416
rect 42334 319404 42398 319416
rect 0 267971 41369 284029
rect 41782 283200 41846 283212
rect 42334 283200 42398 283212
rect 41782 283172 42398 283200
rect 41782 283160 41846 283172
rect 42334 283160 42398 283172
rect 676231 280371 717600 296429
rect 41782 276196 41846 276208
rect 42334 276196 42398 276208
rect 41782 276168 42398 276196
rect 41782 276156 41846 276168
rect 42334 276156 42398 276168
rect 0 224771 41369 240829
rect 41782 239952 41846 239964
rect 42334 239952 42398 239964
rect 41782 239924 42398 239952
rect 41782 239912 41846 239924
rect 42334 239912 42398 239924
rect 676231 235371 717600 251429
rect 41782 233016 41846 233028
rect 42334 233016 42398 233028
rect 41782 232988 42398 233016
rect 41782 232976 41846 232988
rect 42334 232976 42398 232988
rect 0 181571 41369 197629
rect 41782 196772 41846 196784
rect 42334 196772 42398 196784
rect 41782 196744 42398 196772
rect 41782 196732 41846 196744
rect 42334 196732 42398 196744
rect 676231 190171 717600 206229
rect 41782 189836 41846 189848
rect 42334 189836 42398 189848
rect 41782 189808 42398 189836
rect 41782 189796 41846 189808
rect 42334 189796 42398 189808
rect 676231 145171 717600 161229
rect 55 124336 39593 124783
rect 55 124108 39806 124336
rect 55 112870 39593 124108
tri 39593 124085 39616 124108 ne
tri 39593 112870 39616 112893 se
rect 39616 112870 39806 124108
rect 55 112607 39806 112870
rect 55 111971 39593 112607
rect 55 110925 39774 111971
rect 55 110237 39593 110925
rect 676231 99971 717600 116029
rect 24523 84387 40977 85187
tri 40977 84387 41777 85187 sw
rect 24523 83240 41777 84387
rect 32 79313 39593 83000
rect 32 78707 39600 79313
rect 39756 78707 41777 83240
rect 32 72185 41777 78707
rect 32 71331 39600 72185
rect 32 68024 39593 71331
rect 186682 44248 186746 44260
rect 194686 44248 194750 44260
rect 186682 44220 194750 44248
rect 186682 44208 186746 44220
rect 194686 44208 194750 44220
rect 295242 44180 295306 44192
rect 303246 44180 303310 44192
rect 295242 44152 303310 44180
rect 295242 44140 295306 44152
rect 303246 44140 303310 44152
rect 350074 44180 350138 44192
rect 358078 44180 358142 44192
rect 350074 44152 358142 44180
rect 350074 44140 350138 44152
rect 358078 44140 358142 44152
rect 404906 44180 404970 44192
rect 412910 44180 412974 44192
rect 404906 44152 412974 44180
rect 404906 44140 404970 44152
rect 412910 44140 412974 44152
rect 459646 44180 459710 44192
rect 467650 44180 467714 44192
rect 459646 44152 467714 44180
rect 459646 44140 459710 44152
rect 467650 44140 467714 44152
rect 514478 44180 514542 44192
rect 522482 44180 522546 44192
rect 514478 44152 522546 44180
rect 514478 44140 514542 44152
rect 522482 44140 522546 44152
rect 135162 40236 135226 40248
rect 143534 40236 143598 40248
rect 135162 40208 143598 40236
rect 135162 40196 135226 40208
rect 143534 40196 143598 40208
rect 132600 39878 140940 39963
rect 140996 39934 141048 40000
rect 141104 39878 141313 39963
rect 141369 39934 141499 40000
rect 141555 39878 141898 39963
rect 141954 39934 142084 40000
rect 142140 39878 142517 39963
rect 79664 39616 91393 39806
rect 79664 39593 79892 39616
tri 79892 39593 79915 39616 nw
tri 91107 39593 91130 39616 ne
rect 91130 39593 91393 39616
rect 79076 55 93763 39593
rect 132600 37949 142517 39878
rect 142675 39878 143012 39963
rect 143068 39934 143128 40000
rect 143184 39878 144517 39963
rect 144573 39934 144689 40000
rect 144745 39878 145035 39963
rect 145199 39878 147600 39963
rect 142675 37949 147600 39878
rect 132600 158 147600 37949
rect 186371 0 202429 41369
tri 239013 40977 239813 41777 se
rect 239813 40977 252015 41777
rect 239013 39756 252015 40977
rect 239013 24523 240960 39756
rect 245493 39600 252015 39756
rect 244887 39593 252869 39600
rect 241200 32 256176 39593
rect 294971 0 311029 41369
rect 349771 0 365829 41369
rect 404571 0 420629 41369
rect 459371 0 475429 41369
rect 514171 0 530229 41369
rect 569864 39616 581593 39806
rect 569864 39593 570092 39616
tri 570092 39593 570115 39616 nw
tri 581307 39593 581330 39616 ne
rect 581330 39593 581593 39616
rect 623664 39616 635393 39806
rect 623664 39593 623892 39616
tri 623892 39593 623915 39616 nw
tri 635107 39593 635130 39616 ne
rect 635130 39593 635393 39616
rect 636029 39593 637075 39774
rect 569276 55 583963 39593
rect 623217 55 637763 39593
<< metal2 >>
rect 342164 997474 342224 997483
rect 342164 997405 342224 997414
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 78889 995452 78945 995887
rect 79533 995452 79589 995887
rect 78876 995407 78945 995452
rect 79520 995407 79589 995452
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 82569 995407 82625 995887
rect 83213 995407 83269 995887
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 90021 995452 90077 995887
rect 90008 995407 90077 995452
rect 91217 995407 91273 995887
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 130289 995407 130345 995887
rect 130933 995466 130989 995887
rect 130933 995438 131068 995466
rect 130933 995407 130989 995438
rect 78876 990826 78904 995407
rect 78864 990820 78916 990826
rect 78864 990762 78916 990768
rect 78876 990214 78904 990762
rect 42248 990208 42300 990214
rect 42248 990150 42300 990156
rect 78864 990208 78916 990214
rect 78864 990150 78916 990156
rect 41713 969217 42193 969273
rect 41788 968516 41840 968522
rect 41788 968458 41840 968464
rect 41800 968077 41828 968458
rect 41713 968021 42193 968077
rect 41713 967377 42193 967433
rect 41713 966733 42193 966789
rect 41713 965537 42193 965593
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 41713 963053 42193 963109
rect 41713 962501 42193 962557
rect 41713 961213 42193 961269
rect 41713 960569 42193 960625
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 41713 958729 42193 958785
rect 41713 958177 42193 958233
rect 41788 958112 41840 958118
rect 41788 958054 41840 958060
rect 41800 957589 41828 958054
rect 42260 957778 42288 990150
rect 79520 990146 79548 995407
rect 90008 990758 90036 995407
rect 130304 990826 130332 995407
rect 130292 990820 130344 990826
rect 130292 990762 130344 990768
rect 89996 990752 90048 990758
rect 89996 990694 90048 990700
rect 90008 990162 90036 990694
rect 130304 990690 130332 990762
rect 130292 990684 130344 990690
rect 130292 990626 130344 990632
rect 121276 990616 121328 990622
rect 121276 990558 121328 990564
rect 121288 990457 121316 990558
rect 131040 990457 131068 995438
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 133969 995407 134025 995887
rect 134613 995407 134669 995887
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 141421 995407 141477 995887
rect 142617 995407 142673 995887
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 181689 995466 181745 995887
rect 182333 995466 182389 995887
rect 181689 995407 181760 995466
rect 182333 995438 182496 995466
rect 182333 995407 182389 995438
rect 141436 990758 141464 995407
rect 141424 990752 141476 990758
rect 141424 990694 141476 990700
rect 181732 990690 181760 995407
rect 181720 990684 181772 990690
rect 181720 990626 181772 990632
rect 160192 990480 160244 990486
rect 121274 990448 121330 990457
rect 121274 990383 121330 990392
rect 131026 990448 131082 990457
rect 131026 990383 131082 990392
rect 160020 990428 160192 990434
rect 160020 990422 160244 990428
rect 160020 990406 160232 990422
rect 182468 990418 182496 995438
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 185369 995407 185425 995887
rect 186013 995407 186069 995887
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 192821 995466 192877 995887
rect 192821 995407 192892 995466
rect 194017 995407 194073 995887
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 233089 995466 233145 995887
rect 233733 995466 233789 995887
rect 233068 995407 233145 995466
rect 233712 995407 233789 995466
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 236769 995407 236825 995887
rect 237413 995407 237469 995887
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 244221 995466 244277 995887
rect 244200 995407 244277 995466
rect 245417 995407 245473 995887
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 284689 995452 284745 995887
rect 285333 995452 285389 995887
rect 284680 995407 284745 995452
rect 285324 995407 285389 995452
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 288369 995407 288425 995887
rect 289013 995407 289069 995887
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 295821 995452 295877 995887
rect 295812 995407 295877 995452
rect 297017 995407 297073 995887
rect 192864 990758 192892 995407
rect 192852 990752 192904 990758
rect 192852 990694 192904 990700
rect 192864 990486 192892 990694
rect 233068 990826 233096 995407
rect 233056 990820 233108 990826
rect 233056 990762 233108 990768
rect 194968 990752 195020 990758
rect 194968 990694 195020 990700
rect 194980 990486 195008 990694
rect 233712 990690 233740 995407
rect 244200 990758 244228 995407
rect 284680 990826 284708 995407
rect 284668 990820 284720 990826
rect 284668 990762 284720 990768
rect 244188 990752 244240 990758
rect 244188 990694 244240 990700
rect 285324 990690 285352 995407
rect 286968 990820 287020 990826
rect 286968 990762 287020 990768
rect 233700 990684 233752 990690
rect 233700 990626 233752 990632
rect 285312 990684 285364 990690
rect 285312 990626 285364 990632
rect 286980 990622 287008 990762
rect 295812 990758 295840 995407
rect 295800 990752 295852 990758
rect 295800 990694 295852 990700
rect 286968 990616 287020 990622
rect 286968 990558 287020 990564
rect 295812 990554 295840 990694
rect 342180 990690 342208 997405
rect 585044 997448 585104 997457
rect 585044 997379 585104 997388
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 386489 995452 386545 995887
rect 387133 995452 387189 995887
rect 386489 995407 386552 995452
rect 387133 995407 387196 995452
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 390169 995407 390225 995887
rect 390813 995407 390869 995887
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 397621 995452 397677 995887
rect 397621 995407 397684 995452
rect 398817 995407 398873 995887
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 475489 995452 475545 995887
rect 476133 995452 476189 995887
rect 475488 995407 475545 995452
rect 476132 995407 476189 995452
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 479169 995407 479225 995887
rect 479813 995407 479869 995887
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 486621 995452 486677 995887
rect 486620 995407 486677 995452
rect 487817 995407 487873 995887
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 526889 995407 526945 995887
rect 527533 995407 527589 995887
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 530569 995407 530625 995887
rect 531213 995407 531269 995887
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 538021 995407 538077 995887
rect 539217 995407 539273 995887
rect 372540 990826 372660 990842
rect 345112 990820 345164 990826
rect 345112 990762 345164 990768
rect 372528 990820 372672 990826
rect 372580 990814 372620 990820
rect 372528 990762 372580 990768
rect 372620 990762 372672 990768
rect 342168 990684 342220 990690
rect 342168 990626 342220 990632
rect 345020 990684 345072 990690
rect 345124 990672 345152 990762
rect 386524 990690 386552 995407
rect 345072 990644 345152 990672
rect 386420 990684 386472 990690
rect 345020 990626 345072 990632
rect 386420 990626 386472 990632
rect 386512 990684 386564 990690
rect 386512 990626 386564 990632
rect 295800 990548 295852 990554
rect 295800 990490 295852 990496
rect 386432 990486 386460 990626
rect 387168 990486 387196 995407
rect 397656 990826 397684 995407
rect 397460 990820 397512 990826
rect 397460 990762 397512 990768
rect 397644 990820 397696 990826
rect 397644 990762 397696 990768
rect 397472 990554 397500 990762
rect 400128 990752 400180 990758
rect 400128 990694 400180 990700
rect 419540 990752 419592 990758
rect 419540 990694 419592 990700
rect 438768 990752 438820 990758
rect 438768 990694 438820 990700
rect 458180 990752 458232 990758
rect 458180 990694 458232 990700
rect 397460 990548 397512 990554
rect 397460 990490 397512 990496
rect 400140 990486 400168 990694
rect 419552 990554 419580 990694
rect 438780 990554 438808 990694
rect 458192 990554 458220 990694
rect 475488 990690 475516 995407
rect 475476 990684 475528 990690
rect 475476 990626 475528 990632
rect 476132 990554 476160 995407
rect 486620 990826 486648 995407
rect 486608 990820 486660 990826
rect 486608 990762 486660 990768
rect 477408 990752 477460 990758
rect 477408 990694 477460 990700
rect 477420 990554 477448 990694
rect 526916 990690 526944 995407
rect 527560 990758 527588 995407
rect 538048 990826 538076 995407
rect 585060 992254 585088 997379
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 628689 995466 628745 995887
rect 629333 995466 629389 995887
rect 628668 995407 628745 995466
rect 629312 995407 629389 995466
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 632369 995407 632425 995887
rect 633013 995407 633069 995887
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 639821 995466 639877 995887
rect 639800 995407 639877 995466
rect 641017 995407 641073 995887
rect 585048 992248 585100 992254
rect 585048 992190 585100 992196
rect 538036 990820 538088 990826
rect 538036 990762 538088 990768
rect 527548 990752 527600 990758
rect 527548 990694 527600 990700
rect 526904 990684 526956 990690
rect 526904 990626 526956 990632
rect 626540 990684 626592 990690
rect 626540 990626 626592 990632
rect 419540 990548 419592 990554
rect 419540 990490 419592 990496
rect 438768 990548 438820 990554
rect 438768 990490 438820 990496
rect 458180 990548 458232 990554
rect 458180 990490 458232 990496
rect 476120 990548 476172 990554
rect 476120 990490 476172 990496
rect 477408 990548 477460 990554
rect 477408 990490 477460 990496
rect 192852 990480 192904 990486
rect 192852 990422 192904 990428
rect 194968 990480 195020 990486
rect 194968 990422 195020 990428
rect 386420 990480 386472 990486
rect 386420 990422 386472 990428
rect 387156 990480 387208 990486
rect 387156 990422 387208 990428
rect 400128 990480 400180 990486
rect 400128 990422 400180 990428
rect 173900 990412 173952 990418
rect 131040 990282 131068 990383
rect 160020 990350 160048 990406
rect 173900 990354 173952 990360
rect 182456 990412 182508 990418
rect 182456 990354 182508 990360
rect 140688 990344 140740 990350
rect 160008 990344 160060 990350
rect 140740 990292 140820 990298
rect 140688 990286 140820 990292
rect 160008 990286 160060 990292
rect 140700 990282 140820 990286
rect 173912 990282 173940 990354
rect 131028 990276 131080 990282
rect 140700 990276 140832 990282
rect 140700 990270 140780 990276
rect 131028 990218 131080 990224
rect 140780 990218 140832 990224
rect 173900 990276 173952 990282
rect 173900 990218 173952 990224
rect 89916 990146 90036 990162
rect 626552 990146 626580 990626
rect 628668 990146 628696 995407
rect 629312 990758 629340 995407
rect 639800 990826 639828 995407
rect 674748 992248 674800 992254
rect 674748 992190 674800 992196
rect 639788 990820 639840 990826
rect 639788 990762 639840 990768
rect 629300 990752 629352 990758
rect 629300 990694 629352 990700
rect 631232 990752 631284 990758
rect 631232 990694 631284 990700
rect 631244 990146 631272 990694
rect 639800 990214 639828 990762
rect 639788 990208 639840 990214
rect 639788 990150 639840 990156
rect 673644 990208 673696 990214
rect 673644 990150 673696 990156
rect 42340 990140 42392 990146
rect 42340 990082 42392 990088
rect 79508 990140 79560 990146
rect 79508 990082 79560 990088
rect 89904 990140 90036 990146
rect 89956 990134 90036 990140
rect 626540 990140 626592 990146
rect 89904 990082 89956 990088
rect 626540 990082 626592 990088
rect 628656 990140 628708 990146
rect 628656 990082 628708 990088
rect 631232 990140 631284 990146
rect 631232 990082 631284 990088
rect 673552 990140 673604 990146
rect 673552 990082 673604 990088
rect 42352 958118 42380 990082
rect 42524 990072 42576 990078
rect 42524 990014 42576 990020
rect 673460 990072 673512 990078
rect 673460 990014 673512 990020
rect 42536 968522 42564 990014
rect 42524 968516 42576 968522
rect 42524 968458 42576 968464
rect 42340 958112 42392 958118
rect 42340 958054 42392 958060
rect 42248 957772 42300 957778
rect 42248 957714 42300 957720
rect 41713 957533 42193 957589
rect 42248 957568 42300 957574
rect 42248 957510 42300 957516
rect 41713 956931 42193 956945
rect 42260 956931 42288 957510
rect 41713 956903 42288 956931
rect 41713 956889 42193 956903
rect 41713 956337 42193 956393
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 42246 870088 42302 870097
rect 42246 870023 42302 870032
rect 41713 799417 42193 799473
rect 41713 798221 42193 798277
rect 41800 797774 41828 798221
rect 41788 797768 41840 797774
rect 41788 797710 41840 797716
rect 41713 797577 42193 797633
rect 41713 796933 42193 796989
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41713 791413 42193 791469
rect 41713 790769 42193 790825
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 41713 787733 42193 787789
rect 41800 787302 41828 787733
rect 41788 787296 41840 787302
rect 41788 787238 41840 787244
rect 41713 787089 42193 787145
rect 41800 786690 41828 787089
rect 41788 786684 41840 786690
rect 41788 786626 41840 786632
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 41713 756217 42193 756273
rect 41713 755021 42193 755077
rect 41800 754526 41828 755021
rect 41788 754520 41840 754526
rect 41788 754462 41840 754468
rect 41713 754377 42193 754433
rect 41713 753733 42193 753789
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41713 748213 42193 748269
rect 41713 747569 42193 747625
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41713 744533 42193 744589
rect 41800 744190 41828 744533
rect 41788 744184 41840 744190
rect 41788 744126 41840 744132
rect 41788 744048 41840 744054
rect 41788 743990 41840 743996
rect 41800 743945 41828 743990
rect 41713 743889 42193 743945
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 41713 713017 42193 713073
rect 41713 711821 42193 711877
rect 41800 711346 41828 711821
rect 41788 711340 41840 711346
rect 41788 711282 41840 711288
rect 41713 711177 42193 711233
rect 41713 710533 42193 710589
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41713 705013 42193 705069
rect 41713 704369 42193 704425
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41713 701333 42193 701389
rect 41800 701010 41828 701333
rect 41788 701004 41840 701010
rect 41788 700946 41840 700952
rect 41788 700868 41840 700874
rect 41788 700810 41840 700816
rect 41800 700745 41828 700810
rect 41713 700689 42193 700745
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41713 669817 42193 669873
rect 41788 669112 41840 669118
rect 41788 669054 41840 669060
rect 41800 668677 41828 669054
rect 41713 668621 42193 668677
rect 41713 667977 42193 668033
rect 41713 667333 42193 667389
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 41713 661813 42193 661869
rect 41713 661169 42193 661225
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41788 658708 41840 658714
rect 41788 658650 41840 658656
rect 41800 658189 41828 658650
rect 41713 658133 42193 658189
rect 41788 658096 41840 658102
rect 41788 658038 41840 658044
rect 41800 657545 41828 658038
rect 41713 657489 42193 657545
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 41713 626617 42193 626673
rect 41713 625421 42193 625477
rect 41800 624986 41828 625421
rect 41788 624980 41840 624986
rect 41788 624922 41840 624928
rect 41713 624777 42193 624833
rect 41713 624133 42193 624189
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 41713 618613 42193 618669
rect 41713 617969 42193 618025
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41788 615528 41840 615534
rect 41788 615470 41840 615476
rect 41800 614989 41828 615470
rect 41713 614933 42193 614989
rect 41788 614848 41840 614854
rect 41788 614790 41840 614796
rect 41800 614345 41828 614790
rect 41713 614289 42193 614345
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 41713 583417 42193 583473
rect 41788 582684 41840 582690
rect 41788 582626 41840 582632
rect 41800 582277 41828 582626
rect 41713 582221 42193 582277
rect 41713 581577 42193 581633
rect 41713 580933 42193 580989
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 41713 575413 42193 575469
rect 41713 574769 42193 574825
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41713 571733 42193 571789
rect 41800 571266 41828 571733
rect 41788 571260 41840 571266
rect 41788 571202 41840 571208
rect 41713 571089 42193 571145
rect 41800 570722 41828 571089
rect 41788 570716 41840 570722
rect 41788 570658 41840 570664
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41713 540217 42193 540273
rect 41788 539504 41840 539510
rect 41788 539446 41840 539452
rect 41800 539077 41828 539446
rect 41713 539021 42193 539077
rect 41713 538377 42193 538433
rect 41713 537733 42193 537789
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41713 532213 42193 532269
rect 41713 531569 42193 531625
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 41713 528533 42193 528589
rect 41800 528086 41828 528533
rect 41788 528080 41840 528086
rect 41788 528022 41840 528028
rect 41713 527889 42193 527945
rect 41800 527542 41828 527889
rect 41788 527536 41840 527542
rect 41788 527478 41840 527484
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 41713 412617 42193 412673
rect 41713 411421 42193 411477
rect 41800 411262 41828 411421
rect 41788 411256 41840 411262
rect 41788 411198 41840 411204
rect 41713 410777 42193 410833
rect 41713 410133 42193 410189
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 41713 404613 42193 404669
rect 41713 403969 42193 404025
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41788 401396 41840 401402
rect 41788 401338 41840 401344
rect 41800 400989 41828 401338
rect 41713 400933 42193 400989
rect 41788 400852 41840 400858
rect 41788 400794 41840 400800
rect 41800 400345 41828 400794
rect 41713 400289 42193 400345
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41713 369417 42193 369473
rect 41788 368688 41840 368694
rect 41788 368630 41840 368636
rect 41800 368277 41828 368630
rect 41713 368221 42193 368277
rect 41713 367577 42193 367633
rect 41713 366933 42193 366989
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41713 361413 42193 361469
rect 41713 360769 42193 360825
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41788 358284 41840 358290
rect 41788 358226 41840 358232
rect 41800 357789 41828 358226
rect 41713 357733 42193 357789
rect 41788 357672 41840 357678
rect 41788 357614 41840 357620
rect 41800 357145 41828 357614
rect 41713 357089 42193 357145
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41713 326217 42193 326273
rect 41788 325508 41840 325514
rect 41788 325450 41840 325456
rect 41800 325077 41828 325450
rect 41713 325021 42193 325077
rect 41713 324377 42193 324433
rect 41713 323733 42193 323789
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41713 318213 42193 318269
rect 41713 317569 42193 317625
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41713 314533 42193 314589
rect 41800 314090 41828 314533
rect 41788 314084 41840 314090
rect 41788 314026 41840 314032
rect 41713 313889 42193 313945
rect 41800 313546 41828 313889
rect 41788 313540 41840 313546
rect 41788 313482 41840 313488
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 41713 283017 42193 283073
rect 41788 282328 41840 282334
rect 41788 282270 41840 282276
rect 41800 281877 41828 282270
rect 41713 281821 42193 281877
rect 41713 281177 42193 281233
rect 41713 280533 42193 280589
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41713 275013 42193 275069
rect 41713 274369 42193 274425
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41788 271924 41840 271930
rect 41788 271866 41840 271872
rect 41800 271389 41828 271866
rect 41713 271333 42193 271389
rect 41788 271244 41840 271250
rect 41788 271186 41840 271192
rect 41800 270745 41828 271186
rect 41713 270689 42193 270745
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 41713 239817 42193 239873
rect 41713 238621 42193 238677
rect 41800 238134 41828 238621
rect 41788 238128 41840 238134
rect 41788 238070 41840 238076
rect 41713 237977 42193 238033
rect 41713 237333 42193 237389
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 41713 231813 42193 231869
rect 41713 231169 42193 231225
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 41788 228676 41840 228682
rect 41788 228618 41840 228624
rect 41800 228189 41828 228618
rect 41713 228133 42193 228189
rect 41788 228064 41840 228070
rect 41788 228006 41840 228012
rect 41800 227545 41828 228006
rect 41713 227489 42193 227545
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41713 196617 42193 196673
rect 41713 195421 42193 195477
rect 41800 194954 41828 195421
rect 41788 194948 41840 194954
rect 41788 194890 41840 194896
rect 41713 194777 42193 194833
rect 41713 194133 42193 194189
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41713 188613 42193 188669
rect 41713 187969 42193 188025
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41788 185496 41840 185502
rect 41788 185438 41840 185444
rect 41800 184989 41828 185438
rect 41713 184933 42193 184989
rect 41788 184884 41840 184890
rect 41788 184826 41840 184832
rect 41800 184345 41828 184826
rect 41713 184289 42193 184345
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 42260 121514 42288 870023
rect 42536 797774 42564 968458
rect 673472 965326 673500 990014
rect 673460 965320 673512 965326
rect 673460 965262 673512 965268
rect 673472 875226 673500 965262
rect 673564 964782 673592 990082
rect 673552 964776 673604 964782
rect 673552 964718 673604 964724
rect 673460 875220 673512 875226
rect 673460 875162 673512 875168
rect 42524 797768 42576 797774
rect 42524 797710 42576 797716
rect 42708 797768 42760 797774
rect 42708 797710 42760 797716
rect 42616 787296 42668 787302
rect 42616 787238 42668 787244
rect 42524 786684 42576 786690
rect 42524 786626 42576 786632
rect 42432 767372 42484 767378
rect 42432 767314 42484 767320
rect 42444 754526 42472 767314
rect 42536 759014 42564 786626
rect 42524 759008 42576 759014
rect 42524 758950 42576 758956
rect 42432 754520 42484 754526
rect 42432 754462 42484 754468
rect 42340 744184 42392 744190
rect 42340 744126 42392 744132
rect 42352 739634 42380 744126
rect 42340 739628 42392 739634
rect 42340 739570 42392 739576
rect 42444 711346 42472 754462
rect 42524 753500 42576 753506
rect 42524 753442 42576 753448
rect 42536 744054 42564 753442
rect 42628 744190 42656 787238
rect 42720 767378 42748 797710
rect 673472 786622 673500 875162
rect 673564 874546 673592 964718
rect 673656 953358 673684 990150
rect 673644 953352 673696 953358
rect 673644 953294 673696 953300
rect 673552 874540 673604 874546
rect 673552 874482 673604 874488
rect 673460 786616 673512 786622
rect 673460 786558 673512 786564
rect 673564 786418 673592 874482
rect 673656 864482 673684 953294
rect 673644 864476 673696 864482
rect 673644 864418 673696 864424
rect 673552 786412 673604 786418
rect 673552 786354 673604 786360
rect 673460 774920 673512 774926
rect 673460 774862 673512 774868
rect 42708 767372 42760 767378
rect 42708 767314 42760 767320
rect 42800 759008 42852 759014
rect 42800 758950 42852 758956
rect 42812 753506 42840 758950
rect 42800 753500 42852 753506
rect 42800 753442 42852 753448
rect 42616 744184 42668 744190
rect 42616 744126 42668 744132
rect 42524 744048 42576 744054
rect 42524 743990 42576 743996
rect 42984 744048 43036 744054
rect 42984 743990 43036 743996
rect 42616 739628 42668 739634
rect 42616 739570 42668 739576
rect 42524 734188 42576 734194
rect 42524 734130 42576 734136
rect 42536 720390 42564 734130
rect 42524 720384 42576 720390
rect 42524 720326 42576 720332
rect 42432 711340 42484 711346
rect 42432 711282 42484 711288
rect 42628 701010 42656 739570
rect 42996 734194 43024 743990
rect 42984 734188 43036 734194
rect 42984 734130 43036 734136
rect 673472 730182 673500 774862
rect 673564 740722 673592 786354
rect 673656 774926 673684 864418
rect 674012 786616 674064 786622
rect 674012 786558 674064 786564
rect 673644 774920 673696 774926
rect 673644 774862 673696 774868
rect 674024 772818 674052 786558
rect 673736 772812 673788 772818
rect 673736 772754 673788 772760
rect 674012 772812 674064 772818
rect 674012 772754 674064 772760
rect 673748 753574 673776 772754
rect 673736 753568 673788 753574
rect 673736 753510 673788 753516
rect 673920 753568 673972 753574
rect 673920 753510 673972 753516
rect 673932 742014 673960 753510
rect 673644 742008 673696 742014
rect 673644 741950 673696 741956
rect 673920 742008 673972 742014
rect 673920 741950 673972 741956
rect 673552 740716 673604 740722
rect 673552 740658 673604 740664
rect 673460 730176 673512 730182
rect 673460 730118 673512 730124
rect 42892 720384 42944 720390
rect 42892 720326 42944 720332
rect 42708 711340 42760 711346
rect 42708 711282 42760 711288
rect 42616 701004 42668 701010
rect 42616 700946 42668 700952
rect 42432 695564 42484 695570
rect 42432 695506 42484 695512
rect 42444 681698 42472 695506
rect 42432 681692 42484 681698
rect 42432 681634 42484 681640
rect 42628 678570 42656 700946
rect 42616 678564 42668 678570
rect 42616 678506 42668 678512
rect 42720 678450 42748 711282
rect 42904 700874 42932 720326
rect 42892 700868 42944 700874
rect 42892 700810 42944 700816
rect 42904 695570 42932 700810
rect 42892 695564 42944 695570
rect 42892 695506 42944 695512
rect 673472 685234 673500 730118
rect 673564 695366 673592 740658
rect 673656 739838 673684 741950
rect 673644 739832 673696 739838
rect 673644 739774 673696 739780
rect 673644 739696 673696 739702
rect 673644 739638 673696 739644
rect 673656 720338 673684 739638
rect 673656 720310 673868 720338
rect 673840 701078 673868 720310
rect 673644 701072 673696 701078
rect 673644 701014 673696 701020
rect 673828 701072 673880 701078
rect 673828 701014 673880 701020
rect 673656 695910 673684 701014
rect 673644 695904 673696 695910
rect 673644 695846 673696 695852
rect 673552 695360 673604 695366
rect 673552 695302 673604 695308
rect 673460 685228 673512 685234
rect 673460 685170 673512 685176
rect 42800 681624 42852 681630
rect 42800 681566 42852 681572
rect 42628 678422 42748 678450
rect 42432 676184 42484 676190
rect 42432 676126 42484 676132
rect 42444 658714 42472 676126
rect 42628 672194 42656 678422
rect 42536 672166 42656 672194
rect 42536 669118 42564 672166
rect 42524 669112 42576 669118
rect 42524 669054 42576 669060
rect 42432 658708 42484 658714
rect 42432 658650 42484 658656
rect 42432 651432 42484 651438
rect 42432 651374 42484 651380
rect 42444 631938 42472 651374
rect 42536 632058 42564 669054
rect 42708 658708 42760 658714
rect 42708 658650 42760 658656
rect 42720 632058 42748 658650
rect 42812 658102 42840 681566
rect 42984 678564 43036 678570
rect 42984 678506 43036 678512
rect 42996 676190 43024 678506
rect 42984 676184 43036 676190
rect 42984 676126 43036 676132
rect 42800 658096 42852 658102
rect 42800 658038 42852 658044
rect 42812 651438 42840 658038
rect 42800 651432 42852 651438
rect 42800 651374 42852 651380
rect 673472 639742 673500 685170
rect 673564 651166 673592 695302
rect 673656 651778 673684 695846
rect 673644 651772 673696 651778
rect 673644 651714 673696 651720
rect 673552 651160 673604 651166
rect 673552 651102 673604 651108
rect 673460 639736 673512 639742
rect 673460 639678 673512 639684
rect 42524 632052 42576 632058
rect 42524 631994 42576 632000
rect 42708 632052 42760 632058
rect 42708 631994 42760 632000
rect 42984 632052 43036 632058
rect 42984 631994 43036 632000
rect 42444 631910 42564 631938
rect 42536 614854 42564 631910
rect 42800 631916 42852 631922
rect 42800 631858 42852 631864
rect 42812 624986 42840 631858
rect 42800 624980 42852 624986
rect 42800 624922 42852 624928
rect 42524 614848 42576 614854
rect 42524 614790 42576 614796
rect 42340 574116 42392 574122
rect 42340 574058 42392 574064
rect 42352 540546 42380 574058
rect 42536 570722 42564 614790
rect 42812 612882 42840 624922
rect 42996 615534 43024 631994
rect 42984 615528 43036 615534
rect 42984 615470 43036 615476
rect 42800 612876 42852 612882
rect 42800 612818 42852 612824
rect 42616 612808 42668 612814
rect 42996 612762 43024 615470
rect 42616 612750 42668 612756
rect 42628 612678 42656 612750
rect 42720 612734 43024 612762
rect 42616 612672 42668 612678
rect 42616 612614 42668 612620
rect 42720 571282 42748 612734
rect 42800 612672 42852 612678
rect 42800 612614 42852 612620
rect 42812 582690 42840 612614
rect 673564 606218 673592 651102
rect 673656 606762 673684 651714
rect 673920 639736 673972 639742
rect 673920 639678 673972 639684
rect 673644 606756 673696 606762
rect 673644 606698 673696 606704
rect 673552 606212 673604 606218
rect 673552 606154 673604 606160
rect 673656 595082 673684 606698
rect 673564 595054 673684 595082
rect 673564 585206 673592 595054
rect 673932 594930 673960 639678
rect 673644 594924 673696 594930
rect 673644 594866 673696 594872
rect 673920 594924 673972 594930
rect 673920 594866 673972 594872
rect 673552 585200 673604 585206
rect 673552 585142 673604 585148
rect 42800 582684 42852 582690
rect 42800 582626 42852 582632
rect 42812 574122 42840 582626
rect 42800 574116 42852 574122
rect 42800 574058 42852 574064
rect 42720 571266 42840 571282
rect 42720 571260 42852 571266
rect 42720 571254 42800 571260
rect 42800 571202 42852 571208
rect 42524 570716 42576 570722
rect 42524 570658 42576 570664
rect 42708 570716 42760 570722
rect 42708 570658 42760 570664
rect 42616 554804 42668 554810
rect 42616 554746 42668 554752
rect 42352 540518 42564 540546
rect 42536 539510 42564 540518
rect 42524 539504 42576 539510
rect 42524 539446 42576 539452
rect 42432 527536 42484 527542
rect 42432 527478 42484 527484
rect 42444 400858 42472 527478
rect 42536 411262 42564 539446
rect 42628 528086 42656 554746
rect 42616 528080 42668 528086
rect 42616 528022 42668 528028
rect 42628 444378 42656 528022
rect 42720 527542 42748 570658
rect 42812 554810 42840 571202
rect 673552 560584 673604 560590
rect 673552 560526 673604 560532
rect 42800 554804 42852 554810
rect 42800 554746 42852 554752
rect 673564 546446 673592 560526
rect 673656 550526 673684 594866
rect 673736 594788 673788 594794
rect 673736 594730 673788 594736
rect 673748 575482 673776 594730
rect 673828 585200 673880 585206
rect 673828 585142 673880 585148
rect 673736 575476 673788 575482
rect 673736 575418 673788 575424
rect 673840 560590 673868 585142
rect 674380 575476 674432 575482
rect 674380 575418 674432 575424
rect 673828 560584 673880 560590
rect 673828 560526 673880 560532
rect 674392 559978 674420 575418
rect 674012 559972 674064 559978
rect 674012 559914 674064 559920
rect 674380 559972 674432 559978
rect 674380 559914 674432 559920
rect 673644 550520 673696 550526
rect 673644 550462 673696 550468
rect 673552 546440 673604 546446
rect 673552 546382 673604 546388
rect 673828 546372 673880 546378
rect 673828 546314 673880 546320
rect 42708 527536 42760 527542
rect 42708 527478 42760 527484
rect 673734 521656 673790 521665
rect 673734 521591 673790 521600
rect 673748 502382 673776 521591
rect 673736 502376 673788 502382
rect 673736 502318 673788 502324
rect 673840 498234 673868 546314
rect 674024 521665 674052 559914
rect 674010 521656 674066 521665
rect 674010 521591 674066 521600
rect 673920 502376 673972 502382
rect 673920 502318 673972 502324
rect 673552 498228 673604 498234
rect 673552 498170 673604 498176
rect 673828 498228 673880 498234
rect 673828 498170 673880 498176
rect 673564 449614 673592 498170
rect 673932 488458 673960 502318
rect 673840 488430 673960 488458
rect 673840 469334 673868 488430
rect 673828 469328 673880 469334
rect 673828 469270 673880 469276
rect 673736 469192 673788 469198
rect 673736 469134 673788 469140
rect 673748 463690 673776 469134
rect 673736 463684 673788 463690
rect 673736 463626 673788 463632
rect 674012 463684 674064 463690
rect 674012 463626 674064 463632
rect 673552 449608 673604 449614
rect 673552 449550 673604 449556
rect 673828 449608 673880 449614
rect 673828 449550 673880 449556
rect 42616 444372 42668 444378
rect 42616 444314 42668 444320
rect 42800 444372 42852 444378
rect 42800 444314 42852 444320
rect 673736 444372 673788 444378
rect 673736 444314 673788 444320
rect 42812 441590 42840 444314
rect 42708 441584 42760 441590
rect 42708 441526 42760 441532
rect 42800 441584 42852 441590
rect 42800 441526 42852 441532
rect 42720 422346 42748 441526
rect 42616 422340 42668 422346
rect 42616 422282 42668 422288
rect 42708 422340 42760 422346
rect 42708 422282 42760 422288
rect 42524 411256 42576 411262
rect 42524 411198 42576 411204
rect 42432 400852 42484 400858
rect 42432 400794 42484 400800
rect 42444 357678 42472 400794
rect 42536 391898 42564 411198
rect 42628 405754 42656 422282
rect 673748 421002 673776 444314
rect 673656 420974 673776 421002
rect 673656 420782 673684 420974
rect 673840 420866 673868 449550
rect 674024 444378 674052 463626
rect 674012 444372 674064 444378
rect 674012 444314 674064 444320
rect 674760 427854 674788 992190
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 675407 965407 675887 965463
rect 675392 965320 675444 965326
rect 675392 965262 675444 965268
rect 675404 964911 675432 965262
rect 675404 964883 675887 964911
rect 675407 964855 675887 964883
rect 675392 964776 675444 964782
rect 675392 964718 675444 964724
rect 675404 964267 675432 964718
rect 675404 964239 675887 964267
rect 675407 964211 675887 964239
rect 675407 963567 675887 963623
rect 675407 963015 675887 963071
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 675407 961175 675887 961231
rect 675407 960531 675887 960587
rect 675407 959243 675887 959299
rect 675407 958691 675887 958747
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 675407 956207 675887 956263
rect 675407 955011 675887 955067
rect 675407 954367 675887 954423
rect 675407 953751 675887 953779
rect 675404 953723 675887 953751
rect 675404 953358 675432 953723
rect 675392 953352 675444 953358
rect 675392 953294 675444 953300
rect 675407 952527 675887 952583
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675407 875683 675887 875711
rect 675404 875655 675887 875683
rect 675404 875226 675432 875655
rect 675392 875220 675444 875226
rect 675392 875162 675444 875168
rect 675407 875039 675887 875067
rect 675404 875011 675887 875039
rect 675404 874546 675432 875011
rect 675392 874540 675444 874546
rect 675392 874482 675444 874488
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675887 872031
rect 675407 871331 675887 871387
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865811 675887 865867
rect 675407 865167 675887 865223
rect 675407 864551 675887 864579
rect 675404 864523 675887 864551
rect 675404 864482 675432 864523
rect 675392 864476 675444 864482
rect 675392 864418 675444 864424
rect 675407 863327 675887 863383
rect 677506 818408 677562 818417
rect 675300 818372 675352 818378
rect 677506 818343 677508 818352
rect 675300 818314 675352 818320
rect 677560 818343 677562 818352
rect 677508 818314 677560 818320
rect 675312 781658 675340 818314
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675392 786616 675444 786622
rect 675392 786558 675444 786564
rect 675404 786511 675432 786558
rect 675404 786483 675887 786511
rect 675407 786455 675887 786483
rect 675392 786412 675444 786418
rect 675392 786354 675444 786360
rect 675404 785867 675432 786354
rect 675404 785839 675887 785867
rect 675407 785811 675887 785839
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675887 782831
rect 675407 782131 675887 782187
rect 675300 781652 675352 781658
rect 675300 781594 675352 781600
rect 675300 781448 675352 781454
rect 675300 781390 675352 781396
rect 675312 736658 675340 781390
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 776611 675887 776667
rect 675407 775967 675887 776023
rect 675407 775351 675887 775379
rect 675404 775323 675887 775351
rect 675404 774926 675432 775323
rect 675392 774920 675444 774926
rect 675392 774862 675444 774868
rect 675407 774127 675887 774183
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 675392 741940 675444 741946
rect 675392 741882 675444 741888
rect 675404 741511 675432 741882
rect 675404 741483 675887 741511
rect 675407 741455 675887 741483
rect 675407 740860 675887 740867
rect 675404 740811 675887 740860
rect 675404 740722 675432 740811
rect 675392 740716 675444 740722
rect 675392 740658 675444 740664
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675887 737831
rect 675407 737131 675887 737187
rect 675220 736630 675340 736658
rect 675220 728362 675248 736630
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 731611 675887 731667
rect 675407 730967 675887 731023
rect 675407 730351 675887 730379
rect 675404 730323 675887 730351
rect 675404 730182 675432 730323
rect 675392 730176 675444 730182
rect 675392 730118 675444 730124
rect 675407 729127 675887 729183
rect 675220 728334 675340 728362
rect 675312 691642 675340 728334
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675407 696483 675887 696511
rect 675404 696455 675887 696483
rect 675404 695978 675432 696455
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675407 695844 675887 695867
rect 675404 695811 675887 695844
rect 675404 695366 675432 695811
rect 675392 695360 675444 695366
rect 675392 695302 675444 695308
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675887 692831
rect 675407 692131 675887 692187
rect 675220 691614 675340 691642
rect 675220 683346 675248 691614
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 686611 675887 686667
rect 675407 685967 675887 686023
rect 675407 685372 675887 685379
rect 675404 685323 675887 685372
rect 675404 685234 675432 685323
rect 675392 685228 675444 685234
rect 675392 685170 675444 685176
rect 675407 684127 675887 684183
rect 675220 683318 675340 683346
rect 675312 646898 675340 683318
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 675392 651772 675444 651778
rect 675392 651714 675444 651720
rect 675404 651311 675432 651714
rect 675404 651283 675887 651311
rect 675407 651255 675887 651283
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675404 650667 675432 651102
rect 675404 650639 675887 650667
rect 675407 650611 675887 650639
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675887 647631
rect 675407 646931 675887 646987
rect 675220 646870 675340 646898
rect 675220 646066 675248 646870
rect 675208 646060 675260 646066
rect 675208 646002 675260 646008
rect 675300 645788 675352 645794
rect 675300 645730 675352 645736
rect 675024 606212 675076 606218
rect 675024 606154 675076 606160
rect 675036 594794 675064 606154
rect 675024 594788 675076 594794
rect 675024 594730 675076 594736
rect 675312 593434 675340 645730
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 641411 675887 641467
rect 675407 640767 675887 640823
rect 675407 640151 675887 640179
rect 675404 640123 675887 640151
rect 675404 639742 675432 640123
rect 675392 639736 675444 639742
rect 675392 639678 675444 639684
rect 675407 638927 675887 638983
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 675392 606756 675444 606762
rect 675392 606698 675444 606704
rect 675404 606311 675432 606698
rect 675404 606283 675887 606311
rect 675407 606255 675887 606283
rect 675392 606212 675444 606218
rect 675392 606154 675444 606160
rect 675404 605667 675432 606154
rect 675404 605639 675887 605667
rect 675407 605611 675887 605639
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675887 602631
rect 675407 601931 675887 601987
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 596411 675887 596467
rect 675407 595767 675887 595823
rect 675407 595151 675887 595179
rect 675404 595123 675887 595151
rect 675404 594930 675432 595123
rect 675392 594924 675444 594930
rect 675392 594866 675444 594872
rect 675407 593927 675887 593983
rect 675300 593428 675352 593434
rect 675300 593370 675352 593376
rect 675300 593224 675352 593230
rect 675300 593166 675352 593172
rect 675312 556186 675340 593166
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 675407 561068 675887 561111
rect 675404 561055 675887 561068
rect 675404 560590 675432 561055
rect 675392 560584 675444 560590
rect 675392 560526 675444 560532
rect 675407 560439 675887 560467
rect 675404 560411 675887 560439
rect 675404 559978 675432 560411
rect 675392 559972 675444 559978
rect 675392 559914 675444 559920
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675887 557431
rect 675407 556731 675887 556787
rect 675220 556158 675340 556186
rect 675220 548298 675248 556158
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 551211 675887 551267
rect 675407 550567 675887 550623
rect 675392 550520 675444 550526
rect 675392 550462 675444 550468
rect 675404 549979 675432 550462
rect 675404 549951 675887 549979
rect 675407 549923 675887 549951
rect 675407 548727 675887 548783
rect 675220 548270 675340 548298
rect 675312 513806 675340 548270
rect 675300 513800 675352 513806
rect 677692 513800 677744 513806
rect 675300 513742 675352 513748
rect 677690 513768 677692 513777
rect 677744 513768 677746 513777
rect 677690 513703 677746 513712
rect 674748 427848 674800 427854
rect 674748 427790 674800 427796
rect 677124 427848 677176 427854
rect 677311 427836 677320 427852
rect 677176 427808 677320 427836
rect 677124 427790 677176 427796
rect 677311 427792 677320 427808
rect 677380 427792 677389 427852
rect 673748 420838 673868 420866
rect 673644 420776 673696 420782
rect 673644 420718 673696 420724
rect 42616 405748 42668 405754
rect 42616 405690 42668 405696
rect 42892 405748 42944 405754
rect 42892 405690 42944 405696
rect 42904 401402 42932 405690
rect 42892 401396 42944 401402
rect 42892 401338 42944 401344
rect 42904 401282 42932 401338
rect 42904 401254 43024 401282
rect 42536 391870 42656 391898
rect 42628 386374 42656 391870
rect 42616 386368 42668 386374
rect 42616 386310 42668 386316
rect 42892 386368 42944 386374
rect 42892 386310 42944 386316
rect 42800 372632 42852 372638
rect 42800 372574 42852 372580
rect 42812 367878 42840 372574
rect 42904 368694 42932 386310
rect 42996 372638 43024 401254
rect 673748 384334 673776 420838
rect 673828 420776 673880 420782
rect 673828 420718 673880 420724
rect 673840 401606 673868 420718
rect 673828 401600 673880 401606
rect 673828 401542 673880 401548
rect 675300 401600 675352 401606
rect 675300 401542 675352 401548
rect 673736 384328 673788 384334
rect 673736 384270 673788 384276
rect 673644 383240 673696 383246
rect 673644 383182 673696 383188
rect 673552 380928 673604 380934
rect 673552 380870 673604 380876
rect 42984 372632 43036 372638
rect 42984 372574 43036 372580
rect 42892 368688 42944 368694
rect 42892 368630 42944 368636
rect 42524 367872 42576 367878
rect 42524 367814 42576 367820
rect 42800 367872 42852 367878
rect 42800 367814 42852 367820
rect 42536 358290 42564 367814
rect 42904 367724 42932 368630
rect 42812 367696 42932 367724
rect 42524 358284 42576 358290
rect 42524 358226 42576 358232
rect 42432 357672 42484 357678
rect 42432 357614 42484 357620
rect 42432 325508 42484 325514
rect 42432 325450 42484 325456
rect 42444 322930 42472 325450
rect 42432 322924 42484 322930
rect 42432 322866 42484 322872
rect 42340 314220 42392 314226
rect 42340 314162 42392 314168
rect 42352 283703 42380 314162
rect 42536 314090 42564 358226
rect 42616 357672 42668 357678
rect 42616 357614 42668 357620
rect 42628 322862 42656 357614
rect 42812 342258 42840 367696
rect 42720 342230 42840 342258
rect 42720 325514 42748 342230
rect 673564 338162 673592 380870
rect 673552 338156 673604 338162
rect 673552 338098 673604 338104
rect 42708 325508 42760 325514
rect 42708 325450 42760 325456
rect 42616 322856 42668 322862
rect 42616 322798 42668 322804
rect 42708 322856 42760 322862
rect 42708 322798 42760 322804
rect 42720 314226 42748 322798
rect 42892 322788 42944 322794
rect 42892 322730 42944 322736
rect 42708 314220 42760 314226
rect 42708 314162 42760 314168
rect 42524 314084 42576 314090
rect 42524 314026 42576 314032
rect 42708 314084 42760 314090
rect 42708 314026 42760 314032
rect 42352 283675 42564 283703
rect 42536 282334 42564 283675
rect 42524 282328 42576 282334
rect 42524 282270 42576 282276
rect 42536 276026 42564 282270
rect 42352 275998 42564 276026
rect 42352 245614 42380 275998
rect 42720 271930 42748 314026
rect 42800 313472 42852 313478
rect 42904 313426 42932 322730
rect 42852 313420 42932 313426
rect 42800 313414 42932 313420
rect 42812 313398 42932 313414
rect 42708 271924 42760 271930
rect 42708 271866 42760 271872
rect 42524 271244 42576 271250
rect 42524 271186 42576 271192
rect 42340 245608 42392 245614
rect 42340 245550 42392 245556
rect 42536 245546 42564 271186
rect 42524 245540 42576 245546
rect 42524 245482 42576 245488
rect 42616 238128 42668 238134
rect 42616 238070 42668 238076
rect 42628 232898 42656 238070
rect 42340 232892 42392 232898
rect 42340 232834 42392 232840
rect 42616 232892 42668 232898
rect 42616 232834 42668 232840
rect 42352 208418 42380 232834
rect 42720 228682 42748 271866
rect 42812 271250 42840 313398
rect 673564 303618 673592 338098
rect 673656 337550 673684 383182
rect 673748 380934 673776 384270
rect 675312 383253 675340 401542
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675392 384328 675444 384334
rect 675392 384270 675444 384276
rect 675404 383911 675432 384270
rect 675404 383860 675887 383911
rect 675407 383855 675887 383860
rect 675407 383253 675887 383267
rect 675312 383246 675887 383253
rect 675300 383240 675887 383246
rect 675352 383225 675887 383240
rect 675407 383211 675887 383225
rect 675300 383182 675352 383188
rect 675312 383142 675340 383182
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 673736 380928 673788 380934
rect 673736 380870 673788 380876
rect 675407 380727 675887 380783
rect 675407 380175 675887 380231
rect 675407 379531 675887 379587
rect 673736 372360 673788 372366
rect 673736 372302 673788 372308
rect 673644 337544 673696 337550
rect 673644 337486 673696 337492
rect 673552 303612 673604 303618
rect 673552 303554 673604 303560
rect 673656 293622 673684 337486
rect 673748 328098 673776 372302
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 372751 675887 372779
rect 675404 372723 675887 372751
rect 675404 372366 675432 372723
rect 675392 372360 675444 372366
rect 675392 372302 675444 372308
rect 675407 371527 675887 371583
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675407 338708 675887 338711
rect 675404 338655 675887 338708
rect 675404 338162 675432 338655
rect 675392 338156 675444 338162
rect 675392 338098 675444 338104
rect 675407 338028 675887 338067
rect 675404 338011 675887 338028
rect 675404 337550 675432 338011
rect 675392 337544 675444 337550
rect 675392 337486 675444 337492
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675887 335031
rect 675407 334331 675887 334387
rect 673736 328092 673788 328098
rect 673736 328034 673788 328040
rect 673644 293616 673696 293622
rect 673644 293558 673696 293564
rect 673644 293480 673696 293486
rect 673644 293422 673696 293428
rect 42800 271244 42852 271250
rect 42800 271186 42852 271192
rect 673656 264994 673684 293422
rect 673748 282130 673776 328034
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675392 328092 675444 328098
rect 675392 328034 675444 328040
rect 675404 327579 675432 328034
rect 675404 327556 675887 327579
rect 675407 327523 675887 327556
rect 675407 326327 675887 326383
rect 675300 303612 675352 303618
rect 675300 303554 675352 303560
rect 675312 293706 675340 303554
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675407 293706 675887 293711
rect 675312 293678 675887 293706
rect 673920 293616 673972 293622
rect 673920 293558 673972 293564
rect 673736 282124 673788 282130
rect 673736 282066 673788 282072
rect 673460 264988 673512 264994
rect 673460 264930 673512 264936
rect 673644 264988 673696 264994
rect 673644 264930 673696 264936
rect 673472 248742 673500 264930
rect 673460 248736 673512 248742
rect 673460 248678 673512 248684
rect 673644 247512 673696 247518
rect 673644 247454 673696 247460
rect 42892 245608 42944 245614
rect 42892 245550 42944 245556
rect 42800 245540 42852 245546
rect 42800 245482 42852 245488
rect 42708 228676 42760 228682
rect 42708 228618 42760 228624
rect 42616 228064 42668 228070
rect 42616 228006 42668 228012
rect 42340 208412 42392 208418
rect 42340 208354 42392 208360
rect 42432 194948 42484 194954
rect 42432 194890 42484 194896
rect 42340 185496 42392 185502
rect 42340 185438 42392 185444
rect 42248 121508 42300 121514
rect 42248 121450 42300 121456
rect 41418 80608 41474 80617
rect 41418 80543 41474 80552
rect 41432 78305 41460 80543
rect 41418 78296 41474 78305
rect 41418 78231 41474 78240
rect 42352 45762 42380 185438
rect 42444 185366 42472 194890
rect 42432 185360 42484 185366
rect 42432 185302 42484 185308
rect 42628 184890 42656 228006
rect 42720 185502 42748 228618
rect 42812 228070 42840 245482
rect 42904 238134 42932 245550
rect 42892 238128 42944 238134
rect 42892 238070 42944 238076
rect 42800 228064 42852 228070
rect 42800 228006 42852 228012
rect 42892 208412 42944 208418
rect 42892 208354 42944 208360
rect 42904 194954 42932 208354
rect 673656 203386 673684 247454
rect 673748 244066 673776 282066
rect 673932 247518 673960 293558
rect 675312 293486 675340 293678
rect 675407 293655 675887 293678
rect 675392 293616 675444 293622
rect 675392 293558 675444 293564
rect 675300 293480 675352 293486
rect 675300 293422 675352 293428
rect 675404 293067 675432 293558
rect 675404 293012 675887 293067
rect 675407 293011 675887 293012
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675887 290031
rect 675407 289331 675887 289387
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675407 282540 675887 282579
rect 675404 282523 675887 282540
rect 675404 282130 675432 282523
rect 675392 282124 675444 282130
rect 675392 282066 675444 282072
rect 675407 281327 675887 281383
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675312 248742 675340 248773
rect 675300 248736 675352 248742
rect 675407 248690 675887 248711
rect 675352 248684 675887 248690
rect 675300 248678 675887 248684
rect 675312 248662 675887 248678
rect 673920 247512 673972 247518
rect 673920 247454 673972 247460
rect 673748 244038 673960 244066
rect 673828 243840 673880 243846
rect 673828 243782 673880 243788
rect 673840 218142 673868 243782
rect 673932 237726 673960 244038
rect 675312 243846 675340 248662
rect 675407 248655 675887 248662
rect 675407 248039 675887 248067
rect 675404 248011 675887 248039
rect 675404 247518 675432 248011
rect 675392 247512 675444 247518
rect 675392 247454 675444 247460
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675887 245031
rect 675407 244331 675887 244387
rect 675300 243840 675352 243846
rect 675300 243782 675352 243788
rect 673920 237720 673972 237726
rect 673920 237662 673972 237668
rect 673932 237386 673960 237662
rect 673920 237380 673972 237386
rect 673920 237322 673972 237328
rect 674104 237380 674156 237386
rect 674104 237322 674156 237328
rect 674116 231810 674144 237322
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675392 237720 675444 237726
rect 675392 237662 675444 237668
rect 675404 237579 675432 237662
rect 675404 237524 675887 237579
rect 675407 237523 675887 237524
rect 675407 236327 675887 236383
rect 674104 231804 674156 231810
rect 674104 231746 674156 231752
rect 674288 231804 674340 231810
rect 674288 231746 674340 231752
rect 673828 218136 673880 218142
rect 673828 218078 673880 218084
rect 673828 218000 673880 218006
rect 673828 217942 673880 217948
rect 673840 212566 673868 217942
rect 674300 212566 674328 231746
rect 673736 212560 673788 212566
rect 673736 212502 673788 212508
rect 673828 212560 673880 212566
rect 673828 212502 673880 212508
rect 674012 212560 674064 212566
rect 674012 212502 674064 212508
rect 674288 212560 674340 212566
rect 674288 212502 674340 212508
rect 673748 203930 673776 212502
rect 673736 203924 673788 203930
rect 673736 203866 673788 203872
rect 673644 203380 673696 203386
rect 673644 203322 673696 203328
rect 673656 203266 673684 203322
rect 673472 203238 673684 203266
rect 42892 194948 42944 194954
rect 42892 194890 42944 194896
rect 42708 185496 42760 185502
rect 42708 185438 42760 185444
rect 42708 185360 42760 185366
rect 42708 185302 42760 185308
rect 42432 184884 42484 184890
rect 42432 184826 42484 184832
rect 42616 184884 42668 184890
rect 42616 184826 42668 184832
rect 42340 45756 42392 45762
rect 42340 45698 42392 45704
rect 42444 45694 42472 184826
rect 42720 149122 42748 185302
rect 673472 157350 673500 203238
rect 673748 203130 673776 203866
rect 673564 203102 673776 203130
rect 673564 158370 673592 203102
rect 674024 198762 674052 212502
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 675392 203924 675444 203930
rect 675392 203866 675444 203872
rect 675404 203511 675432 203866
rect 675404 203483 675887 203511
rect 675407 203455 675887 203483
rect 675392 203380 675444 203386
rect 675392 203322 675444 203328
rect 675404 202867 675432 203322
rect 675404 202844 675887 202867
rect 675407 202811 675887 202844
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675887 199831
rect 675407 199131 675887 199187
rect 674012 198756 674064 198762
rect 674012 198698 674064 198704
rect 675208 198756 675260 198762
rect 675208 198698 675260 198704
rect 675220 192166 675248 198698
rect 674748 192160 674800 192166
rect 674748 192102 674800 192108
rect 675208 192160 675260 192166
rect 675208 192102 675260 192108
rect 674760 173942 674788 192102
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675407 192372 675887 192379
rect 675404 192323 675887 192372
rect 675404 192166 675432 192323
rect 675392 192160 675444 192166
rect 675392 192102 675444 192108
rect 675407 191127 675887 191183
rect 673828 173936 673880 173942
rect 673828 173878 673880 173884
rect 674748 173936 674800 173942
rect 674748 173878 674800 173884
rect 673552 158364 673604 158370
rect 673552 158306 673604 158312
rect 673460 157344 673512 157350
rect 673460 157286 673512 157292
rect 42524 149116 42576 149122
rect 42524 149058 42576 149064
rect 42708 149116 42760 149122
rect 42708 149058 42760 149064
rect 42536 129690 42564 149058
rect 42536 129662 42748 129690
rect 42720 110498 42748 129662
rect 44732 121508 44784 121514
rect 44732 121450 44784 121456
rect 44744 115938 44772 121450
rect 42984 115932 43036 115938
rect 42984 115874 43036 115880
rect 44732 115932 44784 115938
rect 44732 115874 44784 115880
rect 42524 110492 42576 110498
rect 42524 110434 42576 110440
rect 42708 110492 42760 110498
rect 42708 110434 42760 110440
rect 42536 91066 42564 110434
rect 42996 110401 43024 115874
rect 673472 112130 673500 157286
rect 673564 112810 673592 158306
rect 673840 154601 673868 173878
rect 675407 160295 675887 160351
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675407 158508 675887 158511
rect 675404 158455 675887 158508
rect 675404 158370 675432 158455
rect 675392 158364 675444 158370
rect 675392 158306 675444 158312
rect 675407 157828 675887 157867
rect 675404 157811 675887 157828
rect 675404 157350 675432 157811
rect 675392 157344 675444 157350
rect 675392 157286 675444 157292
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675887 154831
rect 673642 154592 673698 154601
rect 673642 154527 673698 154536
rect 673826 154592 673882 154601
rect 673826 154527 673882 154536
rect 673656 147150 673684 154527
rect 675407 154131 675887 154187
rect 673644 147144 673696 147150
rect 673644 147086 673696 147092
rect 675024 147144 675076 147150
rect 675024 147086 675076 147092
rect 675036 140690 675064 147086
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 147356 675887 147379
rect 675404 147323 675887 147356
rect 675404 147150 675432 147323
rect 675392 147144 675444 147150
rect 675392 147086 675444 147092
rect 675407 146127 675887 146183
rect 674012 140684 674064 140690
rect 674012 140626 674064 140632
rect 675024 140684 675076 140690
rect 675024 140626 675076 140632
rect 674024 116006 674052 140626
rect 673828 116000 673880 116006
rect 673828 115942 673880 115948
rect 674012 116000 674064 116006
rect 674012 115942 674064 115948
rect 673840 115870 673868 115942
rect 673828 115864 673880 115870
rect 673828 115806 673880 115812
rect 675024 115864 675076 115870
rect 675024 115806 675076 115812
rect 673552 112804 673604 112810
rect 673552 112746 673604 112752
rect 673460 112124 673512 112130
rect 673460 112066 673512 112072
rect 42982 110392 43038 110401
rect 42982 110327 43038 110336
rect 42996 96665 43024 110327
rect 42982 96656 43038 96665
rect 42982 96591 43038 96600
rect 44638 96656 44694 96665
rect 44638 96591 44694 96600
rect 42536 91038 42748 91066
rect 42720 80617 42748 91038
rect 44652 82890 44680 96591
rect 44640 82884 44692 82890
rect 44640 82826 44692 82832
rect 44824 82816 44876 82822
rect 44824 82758 44876 82764
rect 44836 82634 44864 82758
rect 44836 82606 44956 82634
rect 42706 80608 42762 80617
rect 42706 80543 42762 80552
rect 42432 45688 42484 45694
rect 42432 45630 42484 45636
rect 42720 45626 42748 80543
rect 42708 45620 42760 45626
rect 42708 45562 42760 45568
rect 44928 45558 44956 82606
rect 140964 45756 141016 45762
rect 140964 45698 141016 45704
rect 44916 45552 44968 45558
rect 44916 45494 44968 45500
rect 93768 41608 93820 41614
rect 121552 41608 121604 41614
rect 93768 41550 93820 41556
rect 121288 41556 121552 41562
rect 140872 41608 140924 41614
rect 121288 41550 121604 41556
rect 140700 41556 140872 41562
rect 140700 41550 140924 41556
rect 93780 40225 93808 41550
rect 121288 41546 121592 41550
rect 140700 41546 140912 41550
rect 121276 41540 121592 41546
rect 121328 41534 121592 41540
rect 140688 41540 140912 41546
rect 121276 41482 121328 41488
rect 140740 41534 140912 41540
rect 140688 41482 140740 41488
rect 93766 40216 93822 40225
rect 93766 40151 93822 40160
rect 140976 40202 141004 45698
rect 143632 45688 143684 45694
rect 143632 45630 143684 45636
rect 143540 45620 143592 45626
rect 143540 45562 143592 45568
rect 143552 40497 143580 45562
rect 143644 44402 143672 45630
rect 527456 45620 527508 45626
rect 527456 45562 527508 45568
rect 195980 45552 196032 45558
rect 195980 45494 196032 45500
rect 516324 45552 516376 45558
rect 516324 45494 516376 45500
rect 195992 44470 196020 45494
rect 405648 44804 405700 44810
rect 405648 44746 405700 44752
rect 411260 44804 411312 44810
rect 411260 44746 411312 44752
rect 359372 44736 359424 44742
rect 359372 44678 359424 44684
rect 354404 44532 354456 44538
rect 354404 44474 354456 44480
rect 195980 44464 196032 44470
rect 195980 44406 196032 44412
rect 304540 44464 304592 44470
rect 304540 44406 304592 44412
rect 143632 44396 143684 44402
rect 143632 44338 143684 44344
rect 145104 44396 145156 44402
rect 145104 44338 145156 44344
rect 195336 44396 195388 44402
rect 195336 44338 195388 44344
rect 144644 40792 144696 40798
rect 144644 40734 144696 40740
rect 143538 40488 143594 40497
rect 143538 40423 143594 40432
rect 143078 40216 143134 40225
rect 140976 40174 141036 40202
rect 141008 40118 141036 40174
rect 143078 40151 143134 40160
rect 143092 40118 143120 40151
rect 144656 40118 144684 40734
rect 145116 40202 145144 44338
rect 188528 44328 188580 44334
rect 188528 44270 188580 44276
rect 192852 44328 192904 44334
rect 192852 44270 192904 44276
rect 188540 42193 188568 44270
rect 192864 42193 192892 44270
rect 195348 42193 195376 44338
rect 195992 42193 196020 44406
rect 199660 44396 199712 44402
rect 199660 44338 199712 44344
rect 200856 44396 200908 44402
rect 200856 44338 200908 44344
rect 241336 44396 241388 44402
rect 241336 44338 241388 44344
rect 251088 44396 251140 44402
rect 251088 44338 251140 44344
rect 199672 44266 199700 44338
rect 199660 44260 199712 44266
rect 199660 44202 199712 44208
rect 199672 42193 199700 44202
rect 200868 42193 200896 44338
rect 201500 44328 201552 44334
rect 201500 44270 201552 44276
rect 201512 42193 201540 44270
rect 146300 42016 146352 42022
rect 146300 41958 146352 41964
rect 146312 40798 146340 41958
rect 149612 41812 149664 41818
rect 149612 41754 149664 41760
rect 146300 40792 146352 40798
rect 146300 40734 146352 40740
rect 149624 40361 149652 41754
rect 168288 41744 168340 41750
rect 187327 41713 187383 42193
rect 187700 41948 187752 41954
rect 187700 41890 187752 41896
rect 187712 41818 187740 41890
rect 187700 41812 187752 41818
rect 187700 41754 187752 41760
rect 188523 41970 188579 42193
rect 188448 41954 188579 41970
rect 188436 41948 188579 41954
rect 188488 41942 188579 41948
rect 188436 41890 188488 41896
rect 188523 41713 188579 41942
rect 189167 41834 189223 42193
rect 189167 41818 189304 41834
rect 189167 41812 189316 41818
rect 189167 41806 189264 41812
rect 189167 41713 189223 41806
rect 189264 41754 189316 41760
rect 191007 41834 191063 42193
rect 191007 41818 191144 41834
rect 191007 41812 191156 41818
rect 191007 41806 191104 41812
rect 191007 41713 191063 41806
rect 191104 41754 191156 41760
rect 192203 41834 192259 42193
rect 192203 41818 192340 41834
rect 192203 41812 192352 41818
rect 192203 41806 192300 41812
rect 192203 41713 192259 41806
rect 192300 41754 192352 41760
rect 192847 41713 192903 42193
rect 193491 41834 193547 42193
rect 193491 41818 193628 41834
rect 193491 41812 193640 41818
rect 193491 41806 193588 41812
rect 193491 41713 193547 41806
rect 193588 41754 193640 41760
rect 194043 41713 194099 42193
rect 195331 41713 195387 42193
rect 195975 41713 196031 42193
rect 196527 41834 196583 42193
rect 197171 41834 197227 42193
rect 197815 41834 197871 42193
rect 198367 41834 198423 42193
rect 198924 41948 198976 41954
rect 198924 41890 198976 41896
rect 198464 41880 198516 41886
rect 196452 41828 198464 41834
rect 198936 41834 198964 41890
rect 199011 41834 199067 42193
rect 196452 41822 198516 41828
rect 196452 41818 198504 41822
rect 198844 41818 199067 41834
rect 196440 41812 198504 41818
rect 196492 41806 198504 41812
rect 198832 41812 199067 41818
rect 196440 41754 196492 41760
rect 196527 41713 196583 41806
rect 197171 41713 197227 41806
rect 197815 41713 197871 41806
rect 198367 41713 198423 41806
rect 198884 41806 199067 41812
rect 198832 41754 198884 41760
rect 199011 41713 199067 41806
rect 199655 41713 199711 42193
rect 200120 41880 200172 41886
rect 200207 41834 200263 42193
rect 200851 41834 200907 42193
rect 200172 41828 200907 41834
rect 200120 41822 200907 41828
rect 200132 41806 200907 41822
rect 200207 41713 200263 41806
rect 200851 41713 200907 41806
rect 201495 41713 201551 42193
rect 168288 41686 168340 41692
rect 168300 41546 168328 41686
rect 168288 41540 168340 41546
rect 168288 41482 168340 41488
rect 149610 40352 149666 40361
rect 149610 40287 149666 40296
rect 145103 40174 145144 40202
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143080 40112 143132 40118
rect 143080 40054 143132 40060
rect 144644 40112 144696 40118
rect 144644 40054 144696 40060
rect 141008 40000 141036 40054
rect 143092 40000 143120 40054
rect 144656 40000 144684 40054
rect 145103 40000 145131 40174
rect 140996 39872 141048 40000
rect 141667 39934 141813 40000
rect 143068 39450 143128 40000
rect 144573 39803 144689 40000
rect 145091 39706 145143 40000
rect 241348 39953 241376 44338
rect 251100 42090 251128 44338
rect 297088 44328 297140 44334
rect 297088 44270 297140 44276
rect 299572 44328 299624 44334
rect 299572 44270 299624 44276
rect 297100 42193 297128 44270
rect 299584 42193 299612 44270
rect 303896 44260 303948 44266
rect 303896 44202 303948 44208
rect 303908 42193 303936 44202
rect 304552 42193 304580 44406
rect 306380 44396 306432 44402
rect 306380 44338 306432 44344
rect 309416 44396 309468 44402
rect 309416 44338 309468 44344
rect 352564 44396 352616 44402
rect 352564 44338 352616 44344
rect 305736 44328 305788 44334
rect 305736 44270 305788 44276
rect 305748 42193 305776 44270
rect 306392 42193 306420 44338
rect 308220 44260 308272 44266
rect 308220 44202 308272 44208
rect 308232 42193 308260 44202
rect 309428 42193 309456 44338
rect 351920 44328 351972 44334
rect 351920 44270 351972 44276
rect 351932 42193 351960 44270
rect 352576 42193 352604 44338
rect 354416 44334 354444 44474
rect 359384 44402 359412 44678
rect 405660 44577 405688 44746
rect 406752 44736 406804 44742
rect 406752 44678 406804 44684
rect 386418 44568 386474 44577
rect 360568 44532 360620 44538
rect 360568 44474 360620 44480
rect 360660 44532 360712 44538
rect 405646 44568 405702 44577
rect 386418 44503 386420 44512
rect 360660 44474 360712 44480
rect 386472 44503 386474 44512
rect 399668 44532 399720 44538
rect 386420 44474 386472 44480
rect 406764 44538 406792 44678
rect 411272 44538 411300 44746
rect 425060 44736 425112 44742
rect 425060 44678 425112 44684
rect 444196 44736 444248 44742
rect 444196 44678 444248 44684
rect 483018 44704 483074 44713
rect 425072 44606 425100 44678
rect 425060 44600 425112 44606
rect 425060 44542 425112 44548
rect 405646 44503 405702 44512
rect 406752 44532 406804 44538
rect 399668 44474 399720 44480
rect 406752 44474 406804 44480
rect 411260 44532 411312 44538
rect 411260 44474 411312 44480
rect 355416 44396 355468 44402
rect 355416 44338 355468 44344
rect 359372 44396 359424 44402
rect 359372 44338 359424 44344
rect 354404 44328 354456 44334
rect 354404 44270 354456 44276
rect 355428 44282 355456 44338
rect 358728 44328 358780 44334
rect 354416 42193 354444 44270
rect 355428 44266 355640 44282
rect 358728 44270 358780 44276
rect 355428 44260 355652 44266
rect 355428 44254 355600 44260
rect 355600 44202 355652 44208
rect 355612 42193 355640 44202
rect 358740 44198 358768 44270
rect 358728 44192 358780 44198
rect 358728 44134 358780 44140
rect 358740 42193 358768 44134
rect 359384 42193 359412 44338
rect 360580 44334 360608 44474
rect 360672 44402 360700 44474
rect 360660 44396 360712 44402
rect 360660 44338 360712 44344
rect 364248 44396 364300 44402
rect 364248 44338 364300 44344
rect 360568 44328 360620 44334
rect 360568 44270 360620 44276
rect 359924 44260 359976 44266
rect 359924 44202 359976 44208
rect 359936 42193 359964 44202
rect 360580 42193 360608 44270
rect 363052 44260 363104 44266
rect 363052 44202 363104 44208
rect 363064 42193 363092 44202
rect 364260 42193 364288 44338
rect 399680 44334 399708 44474
rect 399668 44328 399720 44334
rect 399668 44270 399720 44276
rect 406764 42193 406792 44474
rect 414204 44464 414256 44470
rect 414204 44406 414256 44412
rect 419816 44464 419868 44470
rect 419816 44406 419868 44412
rect 444208 44418 444236 44678
rect 483018 44639 483020 44648
rect 483072 44639 483074 44648
rect 502062 44704 502118 44713
rect 502062 44639 502118 44648
rect 483020 44610 483072 44616
rect 461492 44600 461544 44606
rect 461492 44542 461544 44548
rect 469128 44600 469180 44606
rect 469220 44600 469272 44606
rect 469180 44548 469220 44554
rect 469128 44542 469272 44548
rect 444288 44532 444340 44538
rect 444288 44474 444340 44480
rect 444300 44418 444328 44474
rect 407396 44396 407448 44402
rect 407396 44338 407448 44344
rect 410432 44396 410484 44402
rect 410432 44338 410484 44344
rect 407408 42193 407436 44338
rect 410444 42193 410472 44338
rect 413560 44328 413612 44334
rect 413560 44270 413612 44276
rect 411076 44260 411128 44266
rect 411076 44202 411128 44208
rect 411088 42193 411116 44202
rect 413572 42193 413600 44270
rect 414216 42193 414244 44406
rect 419080 44396 419132 44402
rect 419080 44338 419132 44344
rect 417884 44328 417936 44334
rect 417884 44270 417936 44276
rect 417896 42193 417924 44270
rect 419092 42193 419120 44338
rect 419828 44266 419856 44406
rect 444208 44390 444328 44418
rect 419724 44260 419776 44266
rect 419724 44202 419776 44208
rect 419816 44260 419868 44266
rect 419816 44202 419868 44208
rect 419736 42193 419764 44202
rect 461504 42193 461532 44542
rect 469140 44526 469260 44542
rect 502076 44418 502104 44639
rect 516336 44538 516364 45494
rect 502248 44532 502300 44538
rect 502248 44474 502300 44480
rect 516324 44532 516376 44538
rect 516324 44474 516376 44480
rect 502260 44418 502288 44474
rect 462136 44396 462188 44402
rect 462136 44338 462188 44344
rect 465172 44396 465224 44402
rect 465172 44338 465224 44344
rect 473820 44396 473872 44402
rect 502076 44390 502288 44418
rect 473820 44338 473872 44344
rect 462148 42193 462176 44338
rect 465184 42193 465212 44338
rect 468300 44328 468352 44334
rect 465814 44296 465870 44305
rect 468300 44270 468352 44276
rect 472624 44328 472676 44334
rect 472624 44270 472676 44276
rect 465814 44231 465870 44240
rect 465828 42193 465856 44231
rect 468312 42193 468340 44270
rect 468944 44260 468996 44266
rect 468944 44202 468996 44208
rect 468956 42193 468984 44202
rect 472636 42193 472664 44270
rect 473832 42193 473860 44338
rect 474462 44296 474518 44305
rect 474462 44231 474518 44240
rect 474476 42193 474504 44231
rect 516336 42193 516364 44474
rect 516968 44396 517020 44402
rect 516968 44338 517020 44344
rect 520004 44396 520056 44402
rect 520004 44338 520056 44344
rect 516980 42193 517008 44338
rect 518806 44296 518862 44305
rect 518806 44231 518862 44240
rect 518820 42193 518848 44231
rect 520016 42193 520044 44338
rect 523132 44328 523184 44334
rect 523132 44270 523184 44276
rect 524970 44296 525026 44305
rect 523144 44198 523172 44270
rect 523776 44260 523828 44266
rect 524970 44231 525026 44240
rect 523776 44202 523828 44208
rect 523132 44192 523184 44198
rect 523132 44134 523184 44140
rect 523144 42193 523172 44134
rect 523788 42193 523816 44202
rect 524984 42193 525012 44231
rect 527468 44198 527496 45562
rect 527456 44192 527508 44198
rect 527456 44134 527508 44140
rect 527468 42193 527496 44134
rect 673472 42770 673500 112066
rect 673564 45626 673592 112746
rect 675036 102338 675064 115806
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675407 113283 675887 113311
rect 675404 113255 675887 113283
rect 675404 112810 675432 113255
rect 675392 112804 675444 112810
rect 675392 112746 675444 112752
rect 675407 112639 675887 112667
rect 675404 112611 675887 112639
rect 675404 112130 675432 112611
rect 675392 112124 675444 112130
rect 675392 112066 675444 112072
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 109575 675887 109631
rect 675407 108931 675887 108987
rect 673644 102332 673696 102338
rect 673644 102274 673696 102280
rect 675024 102332 675076 102338
rect 675024 102274 675076 102280
rect 673552 45620 673604 45626
rect 673552 45562 673604 45568
rect 673656 45558 673684 102274
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675392 102332 675444 102338
rect 675392 102274 675444 102280
rect 675404 102179 675432 102274
rect 675404 102151 675887 102179
rect 675407 102123 675887 102151
rect 675407 100927 675887 100983
rect 673644 45552 673696 45558
rect 673644 45494 673696 45500
rect 576768 42764 576820 42770
rect 576768 42706 576820 42712
rect 673460 42764 673512 42770
rect 673460 42706 673512 42712
rect 251088 42084 251140 42090
rect 251088 42026 251140 42032
rect 255228 42084 255280 42090
rect 255228 42026 255280 42032
rect 255240 41886 255268 42026
rect 255228 41880 255280 41886
rect 255228 41822 255280 41828
rect 297100 41806 297179 42193
rect 297640 41880 297692 41886
rect 297767 41834 297823 42193
rect 297692 41828 297823 41834
rect 297640 41822 297823 41828
rect 297652 41806 297823 41822
rect 297123 41713 297179 41806
rect 297767 41713 297823 41806
rect 299584 41806 299663 42193
rect 299607 41713 299663 41806
rect 300676 41880 300728 41886
rect 300803 41834 300859 42193
rect 301447 41834 301503 42193
rect 302091 41834 302147 42193
rect 300728 41828 302280 41834
rect 300676 41822 302280 41828
rect 300688 41818 302280 41822
rect 300688 41812 302292 41818
rect 300688 41806 302240 41812
rect 300803 41713 300859 41806
rect 301447 41713 301503 41806
rect 302091 41713 302147 41806
rect 302240 41754 302292 41760
rect 302643 41713 302699 42193
rect 303908 41806 303987 42193
rect 304552 41806 304631 42193
rect 305127 41834 305183 42193
rect 305012 41818 305183 41834
rect 303931 41713 303987 41806
rect 304575 41713 304631 41806
rect 305000 41812 305183 41818
rect 305052 41806 305183 41812
rect 305748 41806 305827 42193
rect 306392 41834 306471 42193
rect 306300 41818 306471 41834
rect 305000 41754 305052 41760
rect 305127 41713 305183 41806
rect 305771 41713 305827 41806
rect 306288 41812 306471 41818
rect 306340 41806 306471 41812
rect 306288 41754 306340 41760
rect 306415 41713 306471 41806
rect 306967 41713 307023 42193
rect 307484 41948 307536 41954
rect 307484 41890 307536 41896
rect 307496 41834 307524 41890
rect 307611 41834 307667 42193
rect 307496 41806 307667 41834
rect 308232 41806 308311 42193
rect 307611 41713 307667 41806
rect 308255 41713 308311 41806
rect 308807 41834 308863 42193
rect 309428 41834 309507 42193
rect 308807 41806 309507 41834
rect 308807 41713 308863 41806
rect 309451 41713 309507 41806
rect 310095 41713 310151 42193
rect 349618 41848 349674 41857
rect 349618 41783 349674 41792
rect 314580 41682 314700 41698
rect 241334 39944 241390 39953
rect 241334 39879 241390 39888
rect 314568 41676 314712 41682
rect 314620 41670 314660 41676
rect 314568 41618 314620 41624
rect 314660 41618 314712 41624
rect 349632 41614 349660 41783
rect 351923 41713 351979 42193
rect 352567 41713 352623 42193
rect 354407 41713 354463 42193
rect 355603 41834 355659 42193
rect 356247 41834 356303 42193
rect 356891 41834 356947 42193
rect 355603 41806 356947 41834
rect 355603 41713 355659 41806
rect 356247 41713 356303 41806
rect 356891 41713 356947 41806
rect 357443 41713 357499 42193
rect 358731 41713 358787 42193
rect 359375 41713 359431 42193
rect 359927 41834 359983 42193
rect 360016 41880 360068 41886
rect 359927 41828 360016 41834
rect 359927 41822 360068 41828
rect 359927 41806 360056 41822
rect 359927 41713 359983 41806
rect 360571 41713 360627 42193
rect 361120 41880 361172 41886
rect 361215 41834 361271 42193
rect 361172 41828 361271 41834
rect 361120 41822 361271 41828
rect 361132 41806 361271 41822
rect 361215 41713 361271 41806
rect 361767 41713 361823 42193
rect 362411 41936 362467 42193
rect 362500 41948 362552 41954
rect 362411 41908 362500 41936
rect 362411 41857 362467 41908
rect 362500 41890 362552 41896
rect 362406 41848 362467 41857
rect 362462 41792 362467 41848
rect 362406 41783 362467 41792
rect 362411 41713 362467 41783
rect 363055 41713 363111 42193
rect 363512 41880 363564 41886
rect 363607 41834 363663 42193
rect 364251 41834 364307 42193
rect 363564 41828 364307 41834
rect 363512 41822 364307 41828
rect 363524 41806 364307 41822
rect 363607 41713 363663 41806
rect 364251 41713 364307 41806
rect 364895 41713 364951 42193
rect 367098 41984 367154 41993
rect 367098 41919 367100 41928
rect 367152 41919 367154 41928
rect 386142 41984 386198 41993
rect 386142 41919 386198 41928
rect 367100 41890 367152 41896
rect 349620 41608 349672 41614
rect 349620 41550 349672 41556
rect 386156 41562 386184 41919
rect 405527 41713 405583 42193
rect 406723 41820 406792 42193
rect 407367 41820 407436 42193
rect 406723 41713 406779 41820
rect 407367 41713 407423 41820
rect 409207 41834 409263 42193
rect 409207 41818 409368 41834
rect 409207 41812 409380 41818
rect 409207 41806 409328 41812
rect 409207 41713 409263 41806
rect 409328 41754 409380 41760
rect 410403 41834 410472 42193
rect 410524 41880 410576 41886
rect 410403 41828 410524 41834
rect 410403 41822 410576 41828
rect 410403 41806 410564 41822
rect 411047 41820 411116 42193
rect 411691 41834 411747 42193
rect 411812 41880 411864 41886
rect 411691 41828 411812 41834
rect 411691 41822 411864 41828
rect 412243 41834 412299 42193
rect 410403 41713 410459 41806
rect 411047 41713 411103 41820
rect 411691 41806 411852 41822
rect 412243 41818 412404 41834
rect 413531 41820 413600 42193
rect 414175 41820 414244 42193
rect 414727 41834 414783 42193
rect 414848 41880 414900 41886
rect 414727 41828 414848 41834
rect 415371 41834 415427 42193
rect 414727 41822 414900 41828
rect 412243 41812 412416 41818
rect 412243 41806 412364 41812
rect 411691 41713 411747 41806
rect 412243 41713 412299 41806
rect 412364 41754 412416 41760
rect 413531 41713 413587 41820
rect 414175 41713 414231 41820
rect 414727 41806 414888 41822
rect 415228 41818 415427 41834
rect 415216 41812 415427 41818
rect 414727 41713 414783 41806
rect 415268 41806 415427 41812
rect 415216 41754 415268 41760
rect 415371 41713 415427 41806
rect 416015 41834 416071 42193
rect 416136 41880 416188 41886
rect 416015 41828 416136 41834
rect 416015 41822 416188 41828
rect 416015 41806 416176 41822
rect 416015 41713 416071 41806
rect 416567 41713 416623 42193
rect 417211 41834 417267 42193
rect 417068 41818 417267 41834
rect 417056 41812 417267 41818
rect 417108 41806 417267 41812
rect 417056 41754 417108 41760
rect 417211 41713 417267 41806
rect 417855 41820 417924 42193
rect 418407 41834 418463 42193
rect 418540 41886 418568 41917
rect 418528 41880 418580 41886
rect 418407 41828 418528 41834
rect 419051 41834 419120 42193
rect 418580 41828 419120 41834
rect 418407 41820 419120 41828
rect 419695 41820 419764 42193
rect 417855 41713 417911 41820
rect 418407 41806 419107 41820
rect 418407 41713 418463 41806
rect 419051 41713 419107 41806
rect 419695 41713 419751 41820
rect 460327 41713 460383 42193
rect 461504 41806 461579 42193
rect 462148 41806 462223 42193
rect 461523 41713 461579 41806
rect 462167 41713 462223 41806
rect 464007 41834 464063 42193
rect 464160 41880 464212 41886
rect 464007 41828 464160 41834
rect 464007 41822 464212 41828
rect 464007 41806 464200 41822
rect 464007 41713 464063 41806
rect 465184 41834 465259 42193
rect 465184 41818 465396 41834
rect 465184 41812 465408 41818
rect 465184 41806 465356 41812
rect 465203 41713 465259 41806
rect 465828 41806 465903 42193
rect 466491 41834 466547 42193
rect 466380 41818 466547 41834
rect 465356 41754 465408 41760
rect 465847 41713 465903 41806
rect 466368 41812 466547 41818
rect 466420 41806 466547 41812
rect 466368 41754 466420 41760
rect 466491 41713 466547 41806
rect 467043 41834 467099 42193
rect 467196 41880 467248 41886
rect 467043 41828 467196 41834
rect 467043 41822 467248 41828
rect 467043 41806 467236 41822
rect 468312 41806 468387 42193
rect 468956 41806 469031 42193
rect 467043 41713 467099 41806
rect 468331 41713 468387 41806
rect 468975 41713 469031 41806
rect 469527 41834 469583 42193
rect 470048 41880 470100 41886
rect 469527 41818 469720 41834
rect 470171 41834 470227 42193
rect 470100 41828 470227 41834
rect 470048 41822 470227 41828
rect 469527 41812 469732 41818
rect 469527 41806 469680 41812
rect 469527 41713 469583 41806
rect 470060 41806 470227 41822
rect 469680 41754 469732 41760
rect 470171 41713 470227 41806
rect 470815 41834 470871 42193
rect 470968 41880 471020 41886
rect 470815 41828 470968 41834
rect 470815 41822 471020 41828
rect 470815 41806 471008 41822
rect 470815 41713 470871 41806
rect 471367 41713 471423 42193
rect 472011 41834 472067 42193
rect 471900 41818 472067 41834
rect 471888 41812 472067 41818
rect 471940 41806 472067 41812
rect 472636 41806 472711 42193
rect 473084 41880 473136 41886
rect 473207 41834 473263 42193
rect 473832 41834 473907 42193
rect 473136 41828 473907 41834
rect 473084 41822 473907 41828
rect 473096 41806 473907 41822
rect 474476 41806 474551 42193
rect 471888 41754 471940 41760
rect 472011 41713 472067 41806
rect 472655 41713 472711 41806
rect 473207 41713 473263 41806
rect 473851 41713 473907 41806
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516323 41713 516379 42193
rect 516967 41713 517023 42193
rect 518807 41713 518863 42193
rect 520003 41834 520059 42193
rect 520096 41880 520148 41886
rect 520003 41828 520096 41834
rect 520003 41822 520148 41828
rect 520003 41806 520136 41822
rect 520003 41713 520059 41806
rect 520647 41713 520703 42193
rect 521200 41880 521252 41886
rect 521291 41834 521347 42193
rect 521252 41828 521347 41834
rect 521200 41822 521347 41828
rect 521212 41806 521347 41822
rect 521291 41713 521347 41806
rect 521843 41713 521899 42193
rect 523131 41713 523187 42193
rect 523775 41713 523831 42193
rect 524236 41880 524288 41886
rect 524327 41834 524383 42193
rect 524288 41828 524383 41834
rect 524236 41822 524383 41828
rect 524248 41806 524383 41822
rect 524327 41713 524383 41806
rect 524971 41713 525027 42193
rect 525524 41880 525576 41886
rect 525615 41834 525671 42193
rect 525576 41828 525671 41834
rect 525524 41822 525671 41828
rect 525536 41806 525671 41822
rect 525615 41713 525671 41806
rect 526167 41713 526223 42193
rect 526811 41834 526867 42193
rect 526732 41818 526867 41834
rect 526720 41812 526867 41818
rect 526772 41806 526867 41812
rect 526720 41754 526772 41760
rect 526811 41713 526867 41806
rect 527455 41713 527511 42193
rect 527916 41880 527968 41886
rect 528007 41834 528063 42193
rect 528651 41834 528707 42193
rect 527968 41828 528707 41834
rect 527916 41822 528707 41828
rect 527928 41806 528707 41822
rect 528007 41713 528063 41806
rect 528651 41713 528707 41806
rect 529295 41713 529351 42193
rect 576780 42022 576808 42706
rect 569132 42016 569184 42022
rect 569132 41958 569184 41964
rect 576768 42016 576820 42022
rect 576768 41958 576820 41964
rect 386328 41676 386380 41682
rect 386328 41618 386380 41624
rect 386340 41562 386368 41618
rect 386156 41534 386368 41562
rect 507860 41608 507912 41614
rect 507780 41556 507860 41562
rect 507780 41550 507912 41556
rect 507780 41546 507900 41550
rect 507768 41540 507900 41546
rect 507820 41534 507900 41540
rect 507768 41482 507820 41488
rect 569144 40225 569172 41958
rect 569130 40216 569186 40225
rect 569130 40151 569186 40160
<< via2 >>
rect 342164 997414 342224 997474
rect 121274 990392 121330 990448
rect 131026 990392 131082 990448
rect 585044 997388 585104 997448
rect 42246 870032 42302 870088
rect 673734 521600 673790 521656
rect 674010 521600 674066 521656
rect 677506 818372 677562 818408
rect 677506 818352 677508 818372
rect 677508 818352 677560 818372
rect 677560 818352 677562 818372
rect 677690 513748 677692 513768
rect 677692 513748 677744 513768
rect 677744 513748 677746 513768
rect 677690 513712 677746 513748
rect 677320 427792 677380 427852
rect 41418 80552 41474 80608
rect 41418 78240 41474 78296
rect 673642 154536 673698 154592
rect 673826 154536 673882 154592
rect 42982 110336 43038 110392
rect 42982 96600 43038 96656
rect 44638 96600 44694 96656
rect 42706 80552 42762 80608
rect 93766 40160 93822 40216
rect 143538 40432 143594 40488
rect 143078 40160 143134 40216
rect 149610 40296 149666 40352
rect 386418 44532 386474 44568
rect 386418 44512 386420 44532
rect 386420 44512 386472 44532
rect 386472 44512 386474 44532
rect 405646 44512 405702 44568
rect 483018 44668 483074 44704
rect 483018 44648 483020 44668
rect 483020 44648 483072 44668
rect 483072 44648 483074 44668
rect 502062 44648 502118 44704
rect 465814 44240 465870 44296
rect 474462 44240 474518 44296
rect 518806 44240 518862 44296
rect 524970 44240 525026 44296
rect 349618 41792 349674 41848
rect 241334 39888 241390 39944
rect 362406 41792 362462 41848
rect 367098 41948 367154 41984
rect 367098 41928 367100 41948
rect 367100 41928 367152 41948
rect 367152 41928 367154 41948
rect 386142 41928 386198 41984
rect 569130 40160 569186 40216
<< obsm2 >>
rect 76242 995943 92183 1037600
rect 76242 995887 76441 995943
rect 76609 995887 76993 995943
rect 77161 995887 77637 995943
rect 77805 995887 78281 995943
rect 78449 995887 78833 995943
rect 79001 995887 79477 995943
rect 79645 995887 80121 995943
rect 80289 995887 80673 995943
rect 80841 995887 81317 995943
rect 81485 995887 81961 995943
rect 82129 995887 82513 995943
rect 82681 995887 83157 995943
rect 83325 995887 83801 995943
rect 83969 995887 84445 995943
rect 84613 995887 84997 995943
rect 85165 995887 85641 995943
rect 85809 995887 86285 995943
rect 86453 995887 86837 995943
rect 87005 995887 87481 995943
rect 87649 995887 88125 995943
rect 88293 995887 88677 995943
rect 88845 995887 89321 995943
rect 89489 995887 89965 995943
rect 90133 995887 90517 995943
rect 90685 995887 91161 995943
rect 91329 995887 91805 995943
rect 91973 995887 92183 995943
rect 127642 995943 143583 1037600
rect 127642 995887 127841 995943
rect 128009 995887 128393 995943
rect 128561 995887 129037 995943
rect 129205 995887 129681 995943
rect 129849 995887 130233 995943
rect 130401 995887 130877 995943
rect 131045 995887 131521 995943
rect 131689 995887 132073 995943
rect 132241 995887 132717 995943
rect 132885 995887 133361 995943
rect 133529 995887 133913 995943
rect 134081 995887 134557 995943
rect 134725 995887 135201 995943
rect 135369 995887 135845 995943
rect 136013 995887 136397 995943
rect 136565 995887 137041 995943
rect 137209 995887 137685 995943
rect 137853 995887 138237 995943
rect 138405 995887 138881 995943
rect 139049 995887 139525 995943
rect 139693 995887 140077 995943
rect 140245 995887 140721 995943
rect 140889 995887 141365 995943
rect 141533 995887 141917 995943
rect 142085 995887 142561 995943
rect 142729 995887 143205 995943
rect 143373 995887 143583 995943
rect 179042 995943 194983 1037600
rect 179042 995887 179241 995943
rect 179409 995887 179793 995943
rect 179961 995887 180437 995943
rect 180605 995887 181081 995943
rect 181249 995887 181633 995943
rect 181801 995887 182277 995943
rect 182445 995887 182921 995943
rect 183089 995887 183473 995943
rect 183641 995887 184117 995943
rect 184285 995887 184761 995943
rect 184929 995887 185313 995943
rect 185481 995887 185957 995943
rect 186125 995887 186601 995943
rect 186769 995887 187245 995943
rect 187413 995887 187797 995943
rect 187965 995887 188441 995943
rect 188609 995887 189085 995943
rect 189253 995887 189637 995943
rect 189805 995887 190281 995943
rect 190449 995887 190925 995943
rect 191093 995887 191477 995943
rect 191645 995887 192121 995943
rect 192289 995887 192765 995943
rect 192933 995887 193317 995943
rect 193485 995887 193961 995943
rect 194129 995887 194605 995943
rect 194773 995887 194983 995943
rect 230442 995943 246383 1037600
rect 230442 995887 230641 995943
rect 230809 995887 231193 995943
rect 231361 995887 231837 995943
rect 232005 995887 232481 995943
rect 232649 995887 233033 995943
rect 233201 995887 233677 995943
rect 233845 995887 234321 995943
rect 234489 995887 234873 995943
rect 235041 995887 235517 995943
rect 235685 995887 236161 995943
rect 236329 995887 236713 995943
rect 236881 995887 237357 995943
rect 237525 995887 238001 995943
rect 238169 995887 238645 995943
rect 238813 995887 239197 995943
rect 239365 995887 239841 995943
rect 240009 995887 240485 995943
rect 240653 995887 241037 995943
rect 241205 995887 241681 995943
rect 241849 995887 242325 995943
rect 242493 995887 242877 995943
rect 243045 995887 243521 995943
rect 243689 995887 244165 995943
rect 244333 995887 244717 995943
rect 244885 995887 245361 995943
rect 245529 995887 246005 995943
rect 246173 995887 246383 995943
rect 282042 995943 297983 1037600
rect 333453 998007 348258 1036615
rect 333499 997600 338279 998007
rect 338579 997600 338979 997984
rect 343478 997600 348258 998007
rect 282042 995887 282241 995943
rect 282409 995887 282793 995943
rect 282961 995887 283437 995943
rect 283605 995887 284081 995943
rect 284249 995887 284633 995943
rect 284801 995887 285277 995943
rect 285445 995887 285921 995943
rect 286089 995887 286473 995943
rect 286641 995887 287117 995943
rect 287285 995887 287761 995943
rect 287929 995887 288313 995943
rect 288481 995887 288957 995943
rect 289125 995887 289601 995943
rect 289769 995887 290245 995943
rect 290413 995887 290797 995943
rect 290965 995887 291441 995943
rect 291609 995887 292085 995943
rect 292253 995887 292637 995943
rect 292805 995887 293281 995943
rect 293449 995887 293925 995943
rect 294093 995887 294477 995943
rect 294645 995887 295121 995943
rect 295289 995887 295765 995943
rect 295933 995887 296317 995943
rect 296485 995887 296961 995943
rect 297129 995887 297605 995943
rect 297773 995887 297983 995943
rect 76497 995407 76553 995887
rect 83857 995466 83913 995887
rect 84016 995590 84068 995654
rect 84028 995466 84056 995590
rect 83857 995438 84056 995466
rect 83857 995407 83913 995438
rect 86893 995407 86949 995887
rect 88181 995407 88237 995887
rect 90573 995407 90629 995887
rect 91744 995590 91796 995654
rect 91756 995466 91784 995590
rect 91861 995466 91917 995887
rect 91756 995438 91917 995466
rect 91861 995407 91917 995438
rect 127897 995407 127953 995887
rect 0 969973 41713 970183
rect 0 969805 41657 969973
rect 41713 969861 42193 969917
rect 0 969329 41713 969805
rect 41800 969406 41828 969861
rect 41788 969342 41840 969406
rect 0 969161 41657 969329
rect 0 968685 41713 969161
rect 0 968517 41657 968685
rect 41713 968573 42193 968629
rect 0 968133 41713 968517
rect 0 967965 41657 968133
rect 0 967489 41713 967965
rect 0 967321 41657 967489
rect 0 966845 41713 967321
rect 0 966677 41657 966845
rect 0 966293 41713 966677
rect 0 966125 41657 966293
rect 41713 966181 42193 966237
rect 0 965649 41713 966125
rect 0 965481 41657 965649
rect 0 965005 41713 965481
rect 0 964837 41657 965005
rect 41713 964893 42193 964949
rect 0 964453 41713 964837
rect 0 964285 41657 964453
rect 0 963809 41713 964285
rect 0 963641 41657 963809
rect 0 963165 41713 963641
rect 0 962997 41657 963165
rect 0 962613 41713 962997
rect 0 962445 41657 962613
rect 0 961969 41713 962445
rect 41788 962406 41840 962470
rect 0 961801 41657 961969
rect 41800 961913 41828 962406
rect 41713 961857 42193 961913
rect 0 961325 41713 961801
rect 0 961157 41657 961325
rect 0 960681 41713 961157
rect 0 960513 41657 960681
rect 0 960129 41713 960513
rect 0 959961 41657 960129
rect 0 959485 41713 959961
rect 0 959317 41657 959485
rect 0 958841 41713 959317
rect 0 958673 41657 958841
rect 0 958289 41713 958673
rect 0 958121 41657 958289
rect 0 957645 41713 958121
rect 0 957477 41657 957645
rect 135257 995466 135313 995887
rect 135352 995466 135404 995518
rect 135257 995454 135404 995466
rect 135257 995438 135392 995454
rect 135257 995407 135313 995438
rect 138293 995407 138349 995887
rect 139581 995407 139637 995887
rect 141973 995407 142029 995887
rect 143172 995466 143224 995518
rect 143261 995466 143317 995887
rect 143172 995454 143317 995466
rect 143184 995438 143317 995454
rect 143261 995407 143317 995438
rect 179297 995407 179353 995887
rect 186657 995466 186713 995887
rect 186657 995407 186728 995466
rect 189693 995407 189749 995887
rect 190981 995407 191037 995887
rect 193373 995407 193429 995887
rect 194661 995466 194717 995887
rect 194661 995407 194732 995466
rect 230697 995407 230753 995887
rect 238057 995466 238113 995887
rect 238208 995590 238260 995654
rect 238220 995466 238248 995590
rect 238057 995438 238248 995466
rect 238057 995407 238113 995438
rect 241093 995407 241149 995887
rect 242381 995407 242437 995887
rect 244773 995407 244829 995887
rect 245936 995590 245988 995654
rect 245948 995466 245976 995590
rect 246061 995466 246117 995887
rect 245948 995438 246117 995466
rect 246061 995407 246117 995438
rect 282297 995407 282353 995887
rect 289657 995452 289713 995887
rect 289648 995407 289713 995452
rect 292693 995407 292749 995887
rect 293981 995407 294037 995887
rect 296373 995407 296429 995887
rect 297661 995452 297717 995887
rect 297652 995407 297717 995452
rect 186700 990622 186728 995407
rect 186688 990558 186740 990622
rect 194704 990622 194732 995407
rect 194692 990558 194744 990622
rect 289648 995314 289676 995407
rect 289636 995250 289688 995314
rect 297652 995314 297680 995407
rect 297640 995250 297692 995314
rect 383842 995943 399783 1037600
rect 383842 995887 384041 995943
rect 384209 995887 384593 995943
rect 384761 995887 385237 995943
rect 385405 995887 385881 995943
rect 386049 995887 386433 995943
rect 386601 995887 387077 995943
rect 387245 995887 387721 995943
rect 387889 995887 388273 995943
rect 388441 995887 388917 995943
rect 389085 995887 389561 995943
rect 389729 995887 390113 995943
rect 390281 995887 390757 995943
rect 390925 995887 391401 995943
rect 391569 995887 392045 995943
rect 392213 995887 392597 995943
rect 392765 995887 393241 995943
rect 393409 995887 393885 995943
rect 394053 995887 394437 995943
rect 394605 995887 395081 995943
rect 395249 995887 395725 995943
rect 395893 995887 396277 995943
rect 396445 995887 396921 995943
rect 397089 995887 397565 995943
rect 397733 995887 398117 995943
rect 398285 995887 398761 995943
rect 398929 995887 399405 995943
rect 399573 995887 399783 995943
rect 472842 995943 488783 1037600
rect 472842 995887 473041 995943
rect 473209 995887 473593 995943
rect 473761 995887 474237 995943
rect 474405 995887 474881 995943
rect 475049 995887 475433 995943
rect 475601 995887 476077 995943
rect 476245 995887 476721 995943
rect 476889 995887 477273 995943
rect 477441 995887 477917 995943
rect 478085 995887 478561 995943
rect 478729 995887 479113 995943
rect 479281 995887 479757 995943
rect 479925 995887 480401 995943
rect 480569 995887 481045 995943
rect 481213 995887 481597 995943
rect 481765 995887 482241 995943
rect 482409 995887 482885 995943
rect 483053 995887 483437 995943
rect 483605 995887 484081 995943
rect 484249 995887 484725 995943
rect 484893 995887 485277 995943
rect 485445 995887 485921 995943
rect 486089 995887 486565 995943
rect 486733 995887 487117 995943
rect 487285 995887 487761 995943
rect 487929 995887 488405 995943
rect 488573 995887 488783 995943
rect 524242 995943 540183 1037600
rect 575653 998007 590458 1036615
rect 575699 997600 580479 998007
rect 580779 997600 581179 997984
rect 585678 997600 590458 998007
rect 524242 995887 524441 995943
rect 524609 995887 524993 995943
rect 525161 995887 525637 995943
rect 525805 995887 526281 995943
rect 526449 995887 526833 995943
rect 527001 995887 527477 995943
rect 527645 995887 528121 995943
rect 528289 995887 528673 995943
rect 528841 995887 529317 995943
rect 529485 995887 529961 995943
rect 530129 995887 530513 995943
rect 530681 995887 531157 995943
rect 531325 995887 531801 995943
rect 531969 995887 532445 995943
rect 532613 995887 532997 995943
rect 533165 995887 533641 995943
rect 533809 995887 534285 995943
rect 534453 995887 534837 995943
rect 535005 995887 535481 995943
rect 535649 995887 536125 995943
rect 536293 995887 536677 995943
rect 536845 995887 537321 995943
rect 537489 995887 537965 995943
rect 538133 995887 538517 995943
rect 538685 995887 539161 995943
rect 539329 995887 539805 995943
rect 539973 995887 540183 995943
rect 384097 995407 384153 995887
rect 391457 995452 391513 995887
rect 391457 995407 391520 995452
rect 394493 995407 394549 995887
rect 395781 995407 395837 995887
rect 398173 995407 398229 995887
rect 399461 995452 399517 995887
rect 399461 995407 399524 995452
rect 473097 995407 473153 995887
rect 480457 995452 480513 995887
rect 480456 995407 480513 995452
rect 483493 995407 483549 995887
rect 484781 995407 484837 995887
rect 487173 995407 487229 995887
rect 488461 995452 488517 995887
rect 488460 995407 488517 995452
rect 524497 995407 524553 995887
rect 531857 995466 531913 995887
rect 531964 995590 532016 995654
rect 531976 995466 532004 995590
rect 531857 995438 532004 995466
rect 531857 995407 531913 995438
rect 534893 995407 534949 995887
rect 536181 995407 536237 995887
rect 538573 995407 538629 995887
rect 539692 995590 539744 995654
rect 539704 995466 539732 995590
rect 539861 995466 539917 995887
rect 539704 995438 539917 995466
rect 539861 995407 539917 995438
rect 391492 995314 391520 995407
rect 391480 995250 391532 995314
rect 399496 995314 399524 995407
rect 399484 995250 399536 995314
rect 480456 995314 480484 995407
rect 480444 995250 480496 995314
rect 488460 995314 488488 995407
rect 488448 995250 488500 995314
rect 626042 995943 641983 1037600
rect 626042 995887 626241 995943
rect 626409 995887 626793 995943
rect 626961 995887 627437 995943
rect 627605 995887 628081 995943
rect 628249 995887 628633 995943
rect 628801 995887 629277 995943
rect 629445 995887 629921 995943
rect 630089 995887 630473 995943
rect 630641 995887 631117 995943
rect 631285 995887 631761 995943
rect 631929 995887 632313 995943
rect 632481 995887 632957 995943
rect 633125 995887 633601 995943
rect 633769 995887 634245 995943
rect 634413 995887 634797 995943
rect 634965 995887 635441 995943
rect 635609 995887 636085 995943
rect 636253 995887 636637 995943
rect 636805 995887 637281 995943
rect 637449 995887 637925 995943
rect 638093 995887 638477 995943
rect 638645 995887 639121 995943
rect 639289 995887 639765 995943
rect 639933 995887 640317 995943
rect 640485 995887 640961 995943
rect 641129 995887 641605 995943
rect 641773 995887 641983 995943
rect 626297 995407 626353 995887
rect 633657 995466 633713 995887
rect 633808 995466 633860 995518
rect 633657 995454 633860 995466
rect 633657 995438 633848 995454
rect 633657 995407 633713 995438
rect 636693 995407 636749 995887
rect 637981 995407 638037 995887
rect 640373 995407 640429 995887
rect 641536 995466 641588 995518
rect 641661 995466 641717 995887
rect 641536 995454 641717 995466
rect 641548 995438 641717 995454
rect 641661 995407 641717 995438
rect 42432 969342 42484 969406
rect 42444 962470 42472 969342
rect 42432 962406 42484 962470
rect 0 957001 41713 957477
rect 0 956833 41657 957001
rect 0 956449 41713 956833
rect 0 956281 41657 956449
rect 0 955805 41713 956281
rect 0 955637 41657 955805
rect 0 955161 41713 955637
rect 0 954993 41657 955161
rect 0 954609 41713 954993
rect 0 954441 41657 954609
rect 41713 954497 42193 954553
rect 0 954242 41713 954441
rect 30753 927000 31683 929228
rect 31928 927049 32702 929239
rect 714 926940 39593 927000
rect 714 922819 39600 926940
rect 714 922707 39593 922819
rect 714 916185 39600 922707
rect 714 916099 39593 916185
rect 714 912100 39600 916099
rect 714 912098 39593 912100
rect 985 879878 40000 884658
rect 985 874679 39593 879878
rect 39616 874979 40000 875379
rect 985 869899 40000 874679
rect 985 869853 39593 869899
rect 985 837678 40000 842458
rect 985 832479 39593 837678
rect 39616 832779 40000 833179
rect 985 827699 40000 832479
rect 985 827653 39593 827699
rect 0 800173 41713 800383
rect 0 800005 41657 800173
rect 41713 800061 42193 800117
rect 0 799529 41713 800005
rect 41800 799610 41828 800061
rect 41788 799546 41840 799610
rect 0 799361 41657 799529
rect 0 798885 41713 799361
rect 0 798717 41657 798885
rect 41713 798773 42193 798829
rect 0 798333 41713 798717
rect 0 798165 41657 798333
rect 0 797689 41713 798165
rect 0 797521 41657 797689
rect 0 797045 41713 797521
rect 0 796877 41657 797045
rect 0 796493 41713 796877
rect 0 796325 41657 796493
rect 41713 796381 42193 796437
rect 0 795849 41713 796325
rect 0 795681 41657 795849
rect 0 795205 41713 795681
rect 0 795037 41657 795205
rect 41713 795093 42193 795149
rect 0 794653 41713 795037
rect 0 794485 41657 794653
rect 0 794009 41713 794485
rect 0 793841 41657 794009
rect 0 793365 41713 793841
rect 0 793197 41657 793365
rect 0 792813 41713 793197
rect 0 792645 41657 792813
rect 0 792169 41713 792645
rect 41788 792542 41840 792606
rect 0 792001 41657 792169
rect 41800 792113 41828 792542
rect 41713 792057 42193 792113
rect 0 791525 41713 792001
rect 0 791357 41657 791525
rect 0 790881 41713 791357
rect 0 790713 41657 790881
rect 0 790329 41713 790713
rect 0 790161 41657 790329
rect 0 789685 41713 790161
rect 0 789517 41657 789685
rect 0 789041 41713 789517
rect 0 788873 41657 789041
rect 0 788489 41713 788873
rect 0 788321 41657 788489
rect 0 787845 41713 788321
rect 0 787677 41657 787845
rect 0 787201 41713 787677
rect 0 787033 41657 787201
rect 0 786649 41713 787033
rect 0 786481 41657 786649
rect 0 786005 41713 786481
rect 0 785837 41657 786005
rect 0 785361 41713 785837
rect 0 785193 41657 785361
rect 0 784809 41713 785193
rect 0 784641 41657 784809
rect 41713 784697 42193 784753
rect 0 784442 41713 784641
rect 0 756973 41713 757183
rect 0 756805 41657 756973
rect 41722 756917 41828 756922
rect 41713 756861 42193 756917
rect 0 756329 41713 756805
rect 41800 756430 41828 756861
rect 41788 756366 41840 756430
rect 0 756161 41657 756329
rect 0 755685 41713 756161
rect 0 755517 41657 755685
rect 41713 755573 42193 755629
rect 0 755133 41713 755517
rect 0 754965 41657 755133
rect 0 754489 41713 754965
rect 0 754321 41657 754489
rect 0 753845 41713 754321
rect 0 753677 41657 753845
rect 0 753293 41713 753677
rect 0 753125 41657 753293
rect 41713 753181 42193 753237
rect 0 752649 41713 753125
rect 0 752481 41657 752649
rect 0 752005 41713 752481
rect 0 751837 41657 752005
rect 41713 751893 42193 751949
rect 0 751453 41713 751837
rect 0 751285 41657 751453
rect 0 750809 41713 751285
rect 0 750641 41657 750809
rect 0 750165 41713 750641
rect 0 749997 41657 750165
rect 0 749613 41713 749997
rect 0 749445 41657 749613
rect 0 748969 41713 749445
rect 41788 749362 41840 749426
rect 0 748801 41657 748969
rect 41800 748913 41828 749362
rect 41713 748857 42193 748913
rect 0 748325 41713 748801
rect 0 748157 41657 748325
rect 0 747681 41713 748157
rect 0 747513 41657 747681
rect 0 747129 41713 747513
rect 0 746961 41657 747129
rect 0 746485 41713 746961
rect 0 746317 41657 746485
rect 0 745841 41713 746317
rect 0 745673 41657 745841
rect 0 745289 41713 745673
rect 0 745121 41657 745289
rect 0 744645 41713 745121
rect 0 744477 41657 744645
rect 0 744001 41713 744477
rect 0 743833 41657 744001
rect 0 743449 41713 743833
rect 0 743281 41657 743449
rect 0 742805 41713 743281
rect 0 742637 41657 742805
rect 0 742161 41713 742637
rect 0 741993 41657 742161
rect 0 741609 41713 741993
rect 0 741441 41657 741609
rect 41713 741497 42193 741553
rect 0 741242 41713 741441
rect 0 713773 41713 713983
rect 0 713605 41657 713773
rect 41713 713661 42193 713717
rect 0 713129 41713 713605
rect 41800 713182 41828 713661
rect 0 712961 41657 713129
rect 41788 713118 41840 713182
rect 0 712485 41713 712961
rect 0 712317 41657 712485
rect 41713 712373 42193 712429
rect 0 711933 41713 712317
rect 0 711765 41657 711933
rect 0 711289 41713 711765
rect 0 711121 41657 711289
rect 0 710645 41713 711121
rect 0 710477 41657 710645
rect 0 710093 41713 710477
rect 0 709925 41657 710093
rect 41713 709981 42193 710037
rect 0 709449 41713 709925
rect 0 709281 41657 709449
rect 0 708805 41713 709281
rect 0 708637 41657 708805
rect 41713 708693 42193 708749
rect 0 708253 41713 708637
rect 0 708085 41657 708253
rect 0 707609 41713 708085
rect 0 707441 41657 707609
rect 0 706965 41713 707441
rect 0 706797 41657 706965
rect 0 706413 41713 706797
rect 0 706245 41657 706413
rect 0 705769 41713 706245
rect 41788 706182 41840 706246
rect 0 705601 41657 705769
rect 41800 705713 41828 706182
rect 41713 705657 42193 705713
rect 0 705125 41713 705601
rect 0 704957 41657 705125
rect 0 704481 41713 704957
rect 0 704313 41657 704481
rect 0 703929 41713 704313
rect 0 703761 41657 703929
rect 0 703285 41713 703761
rect 0 703117 41657 703285
rect 0 702641 41713 703117
rect 0 702473 41657 702641
rect 0 702089 41713 702473
rect 0 701921 41657 702089
rect 0 701445 41713 701921
rect 0 701277 41657 701445
rect 0 700801 41713 701277
rect 0 700633 41657 700801
rect 0 700249 41713 700633
rect 0 700081 41657 700249
rect 0 699605 41713 700081
rect 0 699437 41657 699605
rect 0 698961 41713 699437
rect 0 698793 41657 698961
rect 0 698409 41713 698793
rect 0 698241 41657 698409
rect 41713 698297 42193 698353
rect 0 698042 41713 698241
rect 0 670573 41713 670783
rect 0 670405 41657 670573
rect 41713 670461 42193 670517
rect 0 669929 41713 670405
rect 41800 670002 41828 670461
rect 41788 669938 41840 670002
rect 0 669761 41657 669929
rect 0 669285 41713 669761
rect 0 669117 41657 669285
rect 41713 669173 42193 669229
rect 0 668733 41713 669117
rect 0 668565 41657 668733
rect 0 668089 41713 668565
rect 0 667921 41657 668089
rect 0 667445 41713 667921
rect 0 667277 41657 667445
rect 0 666893 41713 667277
rect 0 666725 41657 666893
rect 41713 666781 42193 666837
rect 0 666249 41713 666725
rect 0 666081 41657 666249
rect 0 665605 41713 666081
rect 0 665437 41657 665605
rect 41713 665493 42193 665549
rect 0 665053 41713 665437
rect 0 664885 41657 665053
rect 0 664409 41713 664885
rect 0 664241 41657 664409
rect 0 663765 41713 664241
rect 0 663597 41657 663765
rect 0 663213 41713 663597
rect 0 663045 41657 663213
rect 0 662569 41713 663045
rect 41788 663002 41840 663066
rect 0 662401 41657 662569
rect 41800 662513 41828 663002
rect 41713 662457 42193 662513
rect 0 661925 41713 662401
rect 0 661757 41657 661925
rect 0 661281 41713 661757
rect 0 661113 41657 661281
rect 0 660729 41713 661113
rect 0 660561 41657 660729
rect 0 660085 41713 660561
rect 0 659917 41657 660085
rect 0 659441 41713 659917
rect 0 659273 41657 659441
rect 0 658889 41713 659273
rect 0 658721 41657 658889
rect 0 658245 41713 658721
rect 0 658077 41657 658245
rect 0 657601 41713 658077
rect 0 657433 41657 657601
rect 0 657049 41713 657433
rect 0 656881 41657 657049
rect 0 656405 41713 656881
rect 0 656237 41657 656405
rect 0 655761 41713 656237
rect 0 655593 41657 655761
rect 0 655209 41713 655593
rect 0 655041 41657 655209
rect 41713 655097 42193 655153
rect 0 654842 41713 655041
rect 0 627373 41713 627583
rect 0 627205 41657 627373
rect 41713 627261 42193 627317
rect 0 626729 41713 627205
rect 41800 626822 41828 627261
rect 41788 626758 41840 626822
rect 0 626561 41657 626729
rect 0 626085 41713 626561
rect 0 625917 41657 626085
rect 41713 625973 42193 626029
rect 0 625533 41713 625917
rect 0 625365 41657 625533
rect 0 624889 41713 625365
rect 0 624721 41657 624889
rect 0 624245 41713 624721
rect 0 624077 41657 624245
rect 0 623693 41713 624077
rect 0 623525 41657 623693
rect 41713 623581 42193 623637
rect 0 623049 41713 623525
rect 0 622881 41657 623049
rect 0 622405 41713 622881
rect 0 622237 41657 622405
rect 41713 622293 42193 622349
rect 0 621853 41713 622237
rect 0 621685 41657 621853
rect 0 621209 41713 621685
rect 0 621041 41657 621209
rect 0 620565 41713 621041
rect 0 620397 41657 620565
rect 0 620013 41713 620397
rect 0 619845 41657 620013
rect 0 619369 41713 619845
rect 41788 619754 41840 619818
rect 0 619201 41657 619369
rect 41800 619313 41828 619754
rect 41713 619257 42193 619313
rect 0 618725 41713 619201
rect 0 618557 41657 618725
rect 0 618081 41713 618557
rect 0 617913 41657 618081
rect 0 617529 41713 617913
rect 0 617361 41657 617529
rect 0 616885 41713 617361
rect 0 616717 41657 616885
rect 0 616241 41713 616717
rect 0 616073 41657 616241
rect 0 615689 41713 616073
rect 0 615521 41657 615689
rect 0 615045 41713 615521
rect 0 614877 41657 615045
rect 0 614401 41713 614877
rect 0 614233 41657 614401
rect 0 613849 41713 614233
rect 0 613681 41657 613849
rect 0 613205 41713 613681
rect 0 613037 41657 613205
rect 0 612561 41713 613037
rect 0 612393 41657 612561
rect 0 612009 41713 612393
rect 0 611841 41657 612009
rect 41713 611897 42193 611953
rect 0 611642 41713 611841
rect 0 584173 41713 584383
rect 0 584005 41657 584173
rect 41713 584061 42193 584117
rect 0 583529 41713 584005
rect 41800 583574 41828 584061
rect 0 583361 41657 583529
rect 41788 583510 41840 583574
rect 0 582885 41713 583361
rect 0 582717 41657 582885
rect 41713 582773 42193 582829
rect 0 582333 41713 582717
rect 0 582165 41657 582333
rect 0 581689 41713 582165
rect 0 581521 41657 581689
rect 0 581045 41713 581521
rect 0 580877 41657 581045
rect 0 580493 41713 580877
rect 0 580325 41657 580493
rect 41713 580381 42193 580437
rect 0 579849 41713 580325
rect 0 579681 41657 579849
rect 0 579205 41713 579681
rect 0 579037 41657 579205
rect 41713 579093 42193 579149
rect 0 578653 41713 579037
rect 0 578485 41657 578653
rect 0 578009 41713 578485
rect 0 577841 41657 578009
rect 0 577365 41713 577841
rect 0 577197 41657 577365
rect 0 576813 41713 577197
rect 0 576645 41657 576813
rect 0 576169 41713 576645
rect 41788 576574 41840 576638
rect 0 576001 41657 576169
rect 41800 576113 41828 576574
rect 41713 576057 42193 576113
rect 0 575525 41713 576001
rect 0 575357 41657 575525
rect 0 574881 41713 575357
rect 0 574713 41657 574881
rect 0 574329 41713 574713
rect 0 574161 41657 574329
rect 0 573685 41713 574161
rect 0 573517 41657 573685
rect 0 573041 41713 573517
rect 0 572873 41657 573041
rect 0 572489 41713 572873
rect 0 572321 41657 572489
rect 0 571845 41713 572321
rect 0 571677 41657 571845
rect 0 571201 41713 571677
rect 0 571033 41657 571201
rect 0 570649 41713 571033
rect 0 570481 41657 570649
rect 0 570005 41713 570481
rect 0 569837 41657 570005
rect 0 569361 41713 569837
rect 0 569193 41657 569361
rect 0 568809 41713 569193
rect 0 568641 41657 568809
rect 41713 568697 42193 568753
rect 0 568442 41713 568641
rect 0 540973 41713 541183
rect 0 540805 41657 540973
rect 41713 540861 42193 540917
rect 0 540329 41713 540805
rect 41800 540394 41828 540861
rect 41788 540330 41840 540394
rect 0 540161 41657 540329
rect 0 539685 41713 540161
rect 0 539517 41657 539685
rect 41713 539573 42193 539629
rect 0 539133 41713 539517
rect 0 538965 41657 539133
rect 0 538489 41713 538965
rect 0 538321 41657 538489
rect 0 537845 41713 538321
rect 0 537677 41657 537845
rect 0 537293 41713 537677
rect 0 537125 41657 537293
rect 41713 537181 42193 537237
rect 0 536649 41713 537125
rect 0 536481 41657 536649
rect 0 536005 41713 536481
rect 0 535837 41657 536005
rect 41713 535893 42193 535949
rect 0 535453 41713 535837
rect 0 535285 41657 535453
rect 0 534809 41713 535285
rect 0 534641 41657 534809
rect 0 534165 41713 534641
rect 0 533997 41657 534165
rect 0 533613 41713 533997
rect 0 533445 41657 533613
rect 0 532969 41713 533445
rect 41788 533394 41840 533458
rect 0 532801 41657 532969
rect 41800 532913 41828 533394
rect 41713 532857 42193 532913
rect 0 532325 41713 532801
rect 0 532157 41657 532325
rect 0 531681 41713 532157
rect 0 531513 41657 531681
rect 0 531129 41713 531513
rect 0 530961 41657 531129
rect 0 530485 41713 530961
rect 0 530317 41657 530485
rect 0 529841 41713 530317
rect 0 529673 41657 529841
rect 0 529289 41713 529673
rect 0 529121 41657 529289
rect 0 528645 41713 529121
rect 0 528477 41657 528645
rect 0 528001 41713 528477
rect 0 527833 41657 528001
rect 0 527449 41713 527833
rect 0 527281 41657 527449
rect 0 526805 41713 527281
rect 0 526637 41657 526805
rect 0 526161 41713 526637
rect 0 525993 41657 526161
rect 0 525609 41713 525993
rect 0 525441 41657 525609
rect 41713 525497 42193 525553
rect 0 525242 41713 525441
rect 985 493078 40000 497858
rect 985 487879 39593 493078
rect 39616 488179 40000 488579
rect 985 483099 40000 487879
rect 985 483053 39593 483099
rect 30753 455800 31683 458028
rect 31928 455849 32702 458039
rect 714 455740 39593 455800
rect 714 451619 39600 455740
rect 714 451507 39593 451619
rect 714 444985 39600 451507
rect 714 444899 39593 444985
rect 714 440900 39600 444899
rect 0 413373 41713 413583
rect 0 413205 41657 413373
rect 41713 413261 42193 413317
rect 0 412729 41713 413205
rect 41800 412826 41828 413261
rect 41788 412762 41840 412826
rect 0 412561 41657 412729
rect 0 412085 41713 412561
rect 0 411917 41657 412085
rect 41713 411973 42193 412029
rect 0 411533 41713 411917
rect 0 411365 41657 411533
rect 0 410889 41713 411365
rect 0 410721 41657 410889
rect 0 410245 41713 410721
rect 0 410077 41657 410245
rect 0 409693 41713 410077
rect 0 409525 41657 409693
rect 41713 409581 42193 409637
rect 0 409049 41713 409525
rect 0 408881 41657 409049
rect 0 408405 41713 408881
rect 0 408237 41657 408405
rect 41713 408293 42193 408349
rect 0 407853 41713 408237
rect 0 407685 41657 407853
rect 0 407209 41713 407685
rect 0 407041 41657 407209
rect 0 406565 41713 407041
rect 0 406397 41657 406565
rect 0 406013 41713 406397
rect 0 405845 41657 406013
rect 0 405369 41713 405845
rect 41788 405758 41840 405822
rect 0 405201 41657 405369
rect 41800 405313 41828 405758
rect 41713 405257 42193 405313
rect 0 404725 41713 405201
rect 0 404557 41657 404725
rect 0 404081 41713 404557
rect 0 403913 41657 404081
rect 0 403529 41713 403913
rect 0 403361 41657 403529
rect 0 402885 41713 403361
rect 0 402717 41657 402885
rect 0 402241 41713 402717
rect 0 402073 41657 402241
rect 0 401689 41713 402073
rect 0 401521 41657 401689
rect 0 401045 41713 401521
rect 0 400877 41657 401045
rect 0 400401 41713 400877
rect 0 400233 41657 400401
rect 0 399849 41713 400233
rect 0 399681 41657 399849
rect 0 399205 41713 399681
rect 0 399037 41657 399205
rect 0 398561 41713 399037
rect 0 398393 41657 398561
rect 0 398009 41713 398393
rect 0 397841 41657 398009
rect 41713 397897 42193 397953
rect 0 397642 41713 397841
rect 0 370173 41713 370383
rect 0 370005 41657 370173
rect 41713 370061 42193 370117
rect 0 369529 41713 370005
rect 41800 369578 41828 370061
rect 0 369361 41657 369529
rect 41788 369514 41840 369578
rect 0 368885 41713 369361
rect 0 368717 41657 368885
rect 41713 368773 42193 368829
rect 0 368333 41713 368717
rect 0 368165 41657 368333
rect 0 367689 41713 368165
rect 0 367521 41657 367689
rect 0 367045 41713 367521
rect 0 366877 41657 367045
rect 0 366493 41713 366877
rect 0 366325 41657 366493
rect 41713 366381 42193 366437
rect 0 365849 41713 366325
rect 0 365681 41657 365849
rect 0 365205 41713 365681
rect 0 365037 41657 365205
rect 41713 365093 42193 365149
rect 0 364653 41713 365037
rect 0 364485 41657 364653
rect 0 364009 41713 364485
rect 0 363841 41657 364009
rect 0 363365 41713 363841
rect 0 363197 41657 363365
rect 0 362813 41713 363197
rect 0 362645 41657 362813
rect 0 362169 41713 362645
rect 41788 362578 41840 362642
rect 0 362001 41657 362169
rect 41800 362113 41828 362578
rect 41713 362057 42193 362113
rect 0 361525 41713 362001
rect 0 361357 41657 361525
rect 0 360881 41713 361357
rect 0 360713 41657 360881
rect 0 360329 41713 360713
rect 0 360161 41657 360329
rect 0 359685 41713 360161
rect 0 359517 41657 359685
rect 0 359041 41713 359517
rect 0 358873 41657 359041
rect 0 358489 41713 358873
rect 0 358321 41657 358489
rect 0 357845 41713 358321
rect 0 357677 41657 357845
rect 0 357201 41713 357677
rect 0 357033 41657 357201
rect 0 356649 41713 357033
rect 0 356481 41657 356649
rect 0 356005 41713 356481
rect 0 355837 41657 356005
rect 0 355361 41713 355837
rect 0 355193 41657 355361
rect 0 354809 41713 355193
rect 0 354641 41657 354809
rect 41713 354697 42193 354753
rect 0 354442 41713 354641
rect 0 326973 41713 327183
rect 0 326805 41657 326973
rect 41713 326861 42193 326917
rect 0 326329 41713 326805
rect 41800 326398 41828 326861
rect 41788 326334 41840 326398
rect 0 326161 41657 326329
rect 0 325685 41713 326161
rect 0 325517 41657 325685
rect 41713 325573 42193 325629
rect 0 325133 41713 325517
rect 0 324965 41657 325133
rect 0 324489 41713 324965
rect 0 324321 41657 324489
rect 0 323845 41713 324321
rect 0 323677 41657 323845
rect 0 323293 41713 323677
rect 0 323125 41657 323293
rect 41713 323181 42193 323237
rect 0 322649 41713 323125
rect 0 322481 41657 322649
rect 0 322005 41713 322481
rect 0 321837 41657 322005
rect 41713 321893 42193 321949
rect 0 321453 41713 321837
rect 0 321285 41657 321453
rect 0 320809 41713 321285
rect 0 320641 41657 320809
rect 0 320165 41713 320641
rect 0 319997 41657 320165
rect 0 319613 41713 319997
rect 0 319445 41657 319613
rect 0 318969 41713 319445
rect 41788 319398 41840 319462
rect 0 318801 41657 318969
rect 41800 318913 41828 319398
rect 41713 318857 42193 318913
rect 0 318325 41713 318801
rect 0 318157 41657 318325
rect 0 317681 41713 318157
rect 0 317513 41657 317681
rect 0 317129 41713 317513
rect 0 316961 41657 317129
rect 0 316485 41713 316961
rect 0 316317 41657 316485
rect 0 315841 41713 316317
rect 0 315673 41657 315841
rect 0 315289 41713 315673
rect 0 315121 41657 315289
rect 0 314645 41713 315121
rect 0 314477 41657 314645
rect 0 314001 41713 314477
rect 0 313833 41657 314001
rect 0 313449 41713 313833
rect 0 313281 41657 313449
rect 0 312805 41713 313281
rect 0 312637 41657 312805
rect 0 312161 41713 312637
rect 0 311993 41657 312161
rect 0 311609 41713 311993
rect 0 311441 41657 311609
rect 41713 311497 42193 311553
rect 0 311242 41713 311441
rect 0 283773 41713 283983
rect 0 283605 41657 283773
rect 41713 283661 42193 283717
rect 0 283129 41713 283605
rect 41800 283218 41828 283661
rect 41788 283154 41840 283218
rect 0 282961 41657 283129
rect 0 282485 41713 282961
rect 0 282317 41657 282485
rect 41713 282373 42193 282429
rect 0 281933 41713 282317
rect 0 281765 41657 281933
rect 0 281289 41713 281765
rect 0 281121 41657 281289
rect 0 280645 41713 281121
rect 0 280477 41657 280645
rect 0 280093 41713 280477
rect 0 279925 41657 280093
rect 41713 279981 42193 280037
rect 0 279449 41713 279925
rect 0 279281 41657 279449
rect 0 278805 41713 279281
rect 0 278637 41657 278805
rect 41713 278693 42193 278749
rect 0 278253 41713 278637
rect 0 278085 41657 278253
rect 0 277609 41713 278085
rect 0 277441 41657 277609
rect 0 276965 41713 277441
rect 0 276797 41657 276965
rect 0 276413 41713 276797
rect 0 276245 41657 276413
rect 0 275769 41713 276245
rect 41788 276150 41840 276214
rect 0 275601 41657 275769
rect 41800 275713 41828 276150
rect 41713 275657 42193 275713
rect 0 275125 41713 275601
rect 0 274957 41657 275125
rect 0 274481 41713 274957
rect 0 274313 41657 274481
rect 0 273929 41713 274313
rect 0 273761 41657 273929
rect 0 273285 41713 273761
rect 0 273117 41657 273285
rect 0 272641 41713 273117
rect 0 272473 41657 272641
rect 0 272089 41713 272473
rect 0 271921 41657 272089
rect 0 271445 41713 271921
rect 0 271277 41657 271445
rect 0 270801 41713 271277
rect 0 270633 41657 270801
rect 0 270249 41713 270633
rect 0 270081 41657 270249
rect 0 269605 41713 270081
rect 0 269437 41657 269605
rect 0 268961 41713 269437
rect 0 268793 41657 268961
rect 0 268409 41713 268793
rect 0 268241 41657 268409
rect 41713 268297 42193 268353
rect 0 268042 41713 268241
rect 0 240573 41713 240783
rect 0 240405 41657 240573
rect 41722 240517 41828 240530
rect 41713 240461 42193 240517
rect 0 239929 41713 240405
rect 41800 239970 41828 240461
rect 0 239761 41657 239929
rect 41788 239906 41840 239970
rect 0 239285 41713 239761
rect 0 239117 41657 239285
rect 41713 239173 42193 239229
rect 0 238733 41713 239117
rect 0 238565 41657 238733
rect 0 238089 41713 238565
rect 0 237921 41657 238089
rect 0 237445 41713 237921
rect 0 237277 41657 237445
rect 0 236893 41713 237277
rect 0 236725 41657 236893
rect 41713 236781 42193 236837
rect 0 236249 41713 236725
rect 0 236081 41657 236249
rect 0 235605 41713 236081
rect 0 235437 41657 235605
rect 41713 235493 42193 235549
rect 0 235053 41713 235437
rect 0 234885 41657 235053
rect 0 234409 41713 234885
rect 0 234241 41657 234409
rect 0 233765 41713 234241
rect 0 233597 41657 233765
rect 0 233213 41713 233597
rect 0 233045 41657 233213
rect 0 232569 41713 233045
rect 41788 232970 41840 233034
rect 0 232401 41657 232569
rect 41800 232513 41828 232970
rect 41713 232457 42193 232513
rect 0 231925 41713 232401
rect 0 231757 41657 231925
rect 0 231281 41713 231757
rect 0 231113 41657 231281
rect 0 230729 41713 231113
rect 0 230561 41657 230729
rect 0 230085 41713 230561
rect 0 229917 41657 230085
rect 0 229441 41713 229917
rect 0 229273 41657 229441
rect 0 228889 41713 229273
rect 0 228721 41657 228889
rect 0 228245 41713 228721
rect 0 228077 41657 228245
rect 0 227601 41713 228077
rect 0 227433 41657 227601
rect 0 227049 41713 227433
rect 0 226881 41657 227049
rect 0 226405 41713 226881
rect 0 226237 41657 226405
rect 0 225761 41713 226237
rect 0 225593 41657 225761
rect 0 225209 41713 225593
rect 0 225041 41657 225209
rect 41713 225097 42193 225153
rect 0 224842 41713 225041
rect 0 197373 41713 197583
rect 0 197205 41657 197373
rect 41713 197261 42193 197317
rect 0 196729 41713 197205
rect 41800 196790 41828 197261
rect 0 196561 41657 196729
rect 41788 196726 41840 196790
rect 0 196085 41713 196561
rect 0 195917 41657 196085
rect 41713 195973 42193 196029
rect 0 195533 41713 195917
rect 0 195365 41657 195533
rect 0 194889 41713 195365
rect 0 194721 41657 194889
rect 0 194245 41713 194721
rect 0 194077 41657 194245
rect 0 193693 41713 194077
rect 0 193525 41657 193693
rect 41713 193581 42193 193637
rect 0 193049 41713 193525
rect 0 192881 41657 193049
rect 0 192405 41713 192881
rect 0 192237 41657 192405
rect 41713 192293 42193 192349
rect 0 191853 41713 192237
rect 0 191685 41657 191853
rect 0 191209 41713 191685
rect 0 191041 41657 191209
rect 0 190565 41713 191041
rect 0 190397 41657 190565
rect 0 190013 41713 190397
rect 0 189845 41657 190013
rect 0 189369 41713 189845
rect 41788 189790 41840 189854
rect 0 189201 41657 189369
rect 41800 189313 41828 189790
rect 41713 189257 42193 189313
rect 0 188725 41713 189201
rect 0 188557 41657 188725
rect 0 188081 41713 188557
rect 0 187913 41657 188081
rect 0 187529 41713 187913
rect 0 187361 41657 187529
rect 0 186885 41713 187361
rect 0 186717 41657 186885
rect 0 186241 41713 186717
rect 0 186073 41657 186241
rect 0 185689 41713 186073
rect 0 185521 41657 185689
rect 0 185045 41713 185521
rect 0 184877 41657 185045
rect 0 184401 41713 184877
rect 0 184233 41657 184401
rect 0 183849 41713 184233
rect 0 183681 41657 183849
rect 0 183205 41713 183681
rect 0 183037 41657 183205
rect 0 182561 41713 183037
rect 0 182393 41657 182561
rect 0 182009 41713 182393
rect 0 181841 41657 182009
rect 41713 181897 42193 181953
rect 0 181642 41713 181841
rect 985 120278 40000 125058
rect 42340 799546 42392 799610
rect 42352 792606 42380 799546
rect 42340 792542 42392 792606
rect 42340 756366 42392 756430
rect 42352 749426 42380 756366
rect 42340 749362 42392 749426
rect 42340 713118 42392 713182
rect 42352 706246 42380 713118
rect 673736 870130 673788 870194
rect 42340 706182 42392 706246
rect 673748 863258 673776 870130
rect 673736 863194 673788 863258
rect 42340 669938 42392 670002
rect 42352 663066 42380 669938
rect 42340 663002 42392 663066
rect 42340 626758 42392 626822
rect 42352 619818 42380 626758
rect 42340 619754 42392 619818
rect 42340 583510 42392 583574
rect 42352 576638 42380 583510
rect 42340 576574 42392 576638
rect 42340 540330 42392 540394
rect 42352 533458 42380 540330
rect 42340 533394 42392 533458
rect 42340 412762 42392 412826
rect 42352 405822 42380 412762
rect 42340 405758 42392 405822
rect 42340 369514 42392 369578
rect 42352 362642 42380 369514
rect 42340 362578 42392 362642
rect 675887 967359 717600 967558
rect 675407 967247 675887 967303
rect 675943 967191 717600 967359
rect 675887 966807 717600 967191
rect 675943 966639 717600 966807
rect 675887 966163 717600 966639
rect 675943 965995 717600 966163
rect 675887 965519 717600 965995
rect 675943 965351 717600 965519
rect 675887 964967 717600 965351
rect 675943 964799 717600 964967
rect 675887 964323 717600 964799
rect 675943 964155 717600 964323
rect 675887 963679 717600 964155
rect 675943 963511 717600 963679
rect 675887 963127 717600 963511
rect 675943 962959 717600 963127
rect 675887 962483 717600 962959
rect 675943 962315 717600 962483
rect 675887 961839 717600 962315
rect 675943 961671 717600 961839
rect 675887 961287 717600 961671
rect 675943 961119 717600 961287
rect 675887 960643 717600 961119
rect 675943 960475 717600 960643
rect 675887 959999 717600 960475
rect 675407 959929 675887 959943
rect 675312 959901 675887 959929
rect 675312 951810 675340 959901
rect 675407 959887 675887 959901
rect 675943 959831 717600 959999
rect 675887 959355 717600 959831
rect 675943 959187 717600 959355
rect 675887 958803 717600 959187
rect 675943 958635 717600 958803
rect 675887 958159 717600 958635
rect 675943 957991 717600 958159
rect 675887 957515 717600 957991
rect 675943 957347 717600 957515
rect 675887 956963 717600 957347
rect 675407 956851 675887 956907
rect 675943 956795 717600 956963
rect 675887 956319 717600 956795
rect 675943 956151 717600 956319
rect 675887 955675 717600 956151
rect 675407 955563 675887 955619
rect 675943 955507 717600 955675
rect 675887 955123 717600 955507
rect 675943 954955 717600 955123
rect 675887 954479 717600 954955
rect 675943 954311 717600 954479
rect 675887 953835 717600 954311
rect 675943 953667 717600 953835
rect 675887 953283 717600 953667
rect 675407 953171 675887 953227
rect 675943 953115 717600 953283
rect 675887 952639 717600 953115
rect 675943 952471 717600 952639
rect 675887 951995 717600 952471
rect 675407 951932 675887 951939
rect 675404 951883 675887 951932
rect 675404 951810 675432 951883
rect 675943 951827 717600 951995
rect 675312 951782 675432 951810
rect 675887 951617 717600 951827
rect 678007 922500 716886 922502
rect 678000 918501 716886 922500
rect 678007 918415 716886 918501
rect 678000 911893 716886 918415
rect 678007 911781 716886 911893
rect 678000 907660 716886 911781
rect 678007 907600 716886 907660
rect 684898 905361 685672 907551
rect 685917 905372 686847 907600
rect 675887 878159 717600 878358
rect 675407 878047 675887 878103
rect 675943 877991 717600 878159
rect 675887 877607 717600 877991
rect 675943 877439 717600 877607
rect 675887 876963 717600 877439
rect 675943 876795 717600 876963
rect 675887 876319 717600 876795
rect 675943 876151 717600 876319
rect 675887 875767 717600 876151
rect 675943 875599 717600 875767
rect 675887 875123 717600 875599
rect 675943 874955 717600 875123
rect 675887 874479 717600 874955
rect 675943 874311 717600 874479
rect 675887 873927 717600 874311
rect 675943 873759 717600 873927
rect 675887 873283 717600 873759
rect 675943 873115 717600 873283
rect 675887 872639 717600 873115
rect 675943 872471 717600 872639
rect 675887 872087 717600 872471
rect 675943 871919 717600 872087
rect 675887 871443 717600 871919
rect 675943 871275 717600 871443
rect 675887 870799 717600 871275
rect 675407 870740 675887 870743
rect 675404 870687 675887 870740
rect 675404 870194 675432 870687
rect 675943 870631 717600 870799
rect 675392 870130 675444 870194
rect 675887 870155 717600 870631
rect 675943 869987 717600 870155
rect 675887 869603 717600 869987
rect 675943 869435 717600 869603
rect 675887 868959 717600 869435
rect 675943 868791 717600 868959
rect 675887 868315 717600 868791
rect 675943 868147 717600 868315
rect 675887 867763 717600 868147
rect 675407 867651 675887 867707
rect 675943 867595 717600 867763
rect 675887 867119 717600 867595
rect 675943 866951 717600 867119
rect 675887 866475 717600 866951
rect 675407 866363 675887 866419
rect 675943 866307 717600 866475
rect 675887 865923 717600 866307
rect 675943 865755 717600 865923
rect 675887 865279 717600 865755
rect 675943 865111 717600 865279
rect 675887 864635 717600 865111
rect 675943 864467 717600 864635
rect 675887 864083 717600 864467
rect 675407 863971 675887 864027
rect 675943 863915 717600 864083
rect 675887 863439 717600 863915
rect 675943 863271 717600 863439
rect 675392 863194 675444 863258
rect 675404 862739 675432 863194
rect 675887 862795 717600 863271
rect 675404 862716 675887 862739
rect 675407 862683 675887 862716
rect 675943 862627 717600 862795
rect 675887 862417 717600 862627
rect 678007 833301 716615 833347
rect 677600 828521 716615 833301
rect 677600 827821 677984 828221
rect 678007 823322 716615 828521
rect 677600 818542 716615 823322
rect 675887 788959 717600 789158
rect 675407 788847 675887 788903
rect 675943 788791 717600 788959
rect 675887 788407 717600 788791
rect 675943 788239 717600 788407
rect 675887 787763 717600 788239
rect 675943 787595 717600 787763
rect 675887 787119 717600 787595
rect 675943 786951 717600 787119
rect 675887 786567 717600 786951
rect 675943 786399 717600 786567
rect 675887 785923 717600 786399
rect 675943 785755 717600 785923
rect 675887 785279 717600 785755
rect 675943 785111 717600 785279
rect 675887 784727 717600 785111
rect 675943 784559 717600 784727
rect 675887 784083 717600 784559
rect 675943 783915 717600 784083
rect 675887 783439 717600 783915
rect 675943 783271 717600 783439
rect 675887 782887 717600 783271
rect 675943 782719 717600 782887
rect 675887 782243 717600 782719
rect 675943 782075 717600 782243
rect 675887 781599 717600 782075
rect 675407 781538 675887 781543
rect 675220 781510 675887 781538
rect 675220 774042 675248 781510
rect 675407 781487 675887 781510
rect 675943 781431 717600 781599
rect 675208 773978 675260 774042
rect 675887 780955 717600 781431
rect 675943 780787 717600 780955
rect 675887 780403 717600 780787
rect 675943 780235 717600 780403
rect 675887 779759 717600 780235
rect 675943 779591 717600 779759
rect 675887 779115 717600 779591
rect 675943 778947 717600 779115
rect 675887 778563 717600 778947
rect 675407 778451 675887 778507
rect 675943 778395 717600 778563
rect 675887 777919 717600 778395
rect 675943 777751 717600 777919
rect 675887 777275 717600 777751
rect 675407 777163 675887 777219
rect 675943 777107 717600 777275
rect 675887 776723 717600 777107
rect 675943 776555 717600 776723
rect 675887 776079 717600 776555
rect 675943 775911 717600 776079
rect 675887 775435 717600 775911
rect 675943 775267 717600 775435
rect 675887 774883 717600 775267
rect 675407 774771 675887 774827
rect 675943 774715 717600 774883
rect 675887 774239 717600 774715
rect 675943 774071 717600 774239
rect 675392 773978 675444 774042
rect 675404 773539 675432 773978
rect 675887 773595 717600 774071
rect 675404 773500 675887 773539
rect 675407 773483 675887 773500
rect 675943 773427 717600 773595
rect 675887 773217 717600 773427
rect 675887 743959 717600 744158
rect 675407 743847 675887 743903
rect 675943 743791 717600 743959
rect 675887 743407 717600 743791
rect 675943 743239 717600 743407
rect 675887 742763 717600 743239
rect 675943 742595 717600 742763
rect 675887 742119 717600 742595
rect 675943 741951 717600 742119
rect 675887 741567 717600 741951
rect 675943 741399 717600 741567
rect 675887 740923 717600 741399
rect 675943 740755 717600 740923
rect 675887 740279 717600 740755
rect 675943 740111 717600 740279
rect 675887 739727 717600 740111
rect 675943 739559 717600 739727
rect 675887 739083 717600 739559
rect 675943 738915 717600 739083
rect 675887 738439 717600 738915
rect 675943 738271 717600 738439
rect 675887 737887 717600 738271
rect 675943 737719 717600 737887
rect 675887 737243 717600 737719
rect 675943 737075 717600 737243
rect 675887 736599 717600 737075
rect 675407 736522 675887 736543
rect 675312 736494 675887 736522
rect 675312 729042 675340 736494
rect 675407 736487 675887 736494
rect 675943 736431 717600 736599
rect 675887 735955 717600 736431
rect 675943 735787 717600 735955
rect 675887 735403 717600 735787
rect 675943 735235 717600 735403
rect 675887 734759 717600 735235
rect 675943 734591 717600 734759
rect 675887 734115 717600 734591
rect 675943 733947 717600 734115
rect 675887 733563 717600 733947
rect 675407 733451 675887 733507
rect 675943 733395 717600 733563
rect 675887 732919 717600 733395
rect 675943 732751 717600 732919
rect 675887 732275 717600 732751
rect 675407 732163 675887 732219
rect 675943 732107 717600 732275
rect 675887 731723 717600 732107
rect 675943 731555 717600 731723
rect 675887 731079 717600 731555
rect 675943 730911 717600 731079
rect 675887 730435 717600 730911
rect 675943 730267 717600 730435
rect 675887 729883 717600 730267
rect 675407 729771 675887 729827
rect 675943 729715 717600 729883
rect 675887 729239 717600 729715
rect 675943 729071 717600 729239
rect 675312 729014 675432 729042
rect 675404 728539 675432 729014
rect 675887 728595 717600 729071
rect 675404 728484 675887 728539
rect 675407 728483 675887 728484
rect 675943 728427 717600 728595
rect 675887 728217 717600 728427
rect 675887 698959 717600 699158
rect 675407 698847 675887 698903
rect 675943 698791 717600 698959
rect 675887 698407 717600 698791
rect 675943 698239 717600 698407
rect 675887 697763 717600 698239
rect 675943 697595 717600 697763
rect 675887 697119 717600 697595
rect 675943 696951 717600 697119
rect 675887 696567 717600 696951
rect 675943 696399 717600 696567
rect 675887 695923 717600 696399
rect 675943 695755 717600 695923
rect 675887 695279 717600 695755
rect 675943 695111 717600 695279
rect 675887 694727 717600 695111
rect 675943 694559 717600 694727
rect 675887 694083 717600 694559
rect 675943 693915 717600 694083
rect 675887 693439 717600 693915
rect 675943 693271 717600 693439
rect 675887 692887 717600 693271
rect 675943 692719 717600 692887
rect 675887 692243 717600 692719
rect 675943 692075 717600 692243
rect 675887 691599 717600 692075
rect 675407 691487 675887 691543
rect 675418 691478 675524 691487
rect 675496 690962 675524 691478
rect 675943 691431 717600 691599
rect 675312 690934 675524 690962
rect 675887 690955 717600 691431
rect 675312 683525 675340 690934
rect 675943 690787 717600 690955
rect 675887 690403 717600 690787
rect 675943 690235 717600 690403
rect 675887 689759 717600 690235
rect 675943 689591 717600 689759
rect 675887 689115 717600 689591
rect 675943 688947 717600 689115
rect 675887 688563 717600 688947
rect 675407 688451 675887 688507
rect 675943 688395 717600 688563
rect 675887 687919 717600 688395
rect 675943 687751 717600 687919
rect 675887 687275 717600 687751
rect 675407 687163 675887 687219
rect 675943 687107 717600 687275
rect 675887 686723 717600 687107
rect 675943 686555 717600 686723
rect 675887 686079 717600 686555
rect 675943 685911 717600 686079
rect 675887 685435 717600 685911
rect 675943 685267 717600 685435
rect 675887 684883 717600 685267
rect 675407 684771 675887 684827
rect 675943 684715 717600 684883
rect 675887 684239 717600 684715
rect 675943 684071 717600 684239
rect 675887 683595 717600 684071
rect 675407 683525 675887 683539
rect 675312 683497 675887 683525
rect 675407 683483 675887 683497
rect 675943 683427 717600 683595
rect 675887 683217 717600 683427
rect 675887 653759 717600 653958
rect 675407 653647 675887 653703
rect 675943 653591 717600 653759
rect 675887 653207 717600 653591
rect 675943 653039 717600 653207
rect 675887 652563 717600 653039
rect 675943 652395 717600 652563
rect 675887 651919 717600 652395
rect 675943 651751 717600 651919
rect 675887 651367 717600 651751
rect 675943 651199 717600 651367
rect 675887 650723 717600 651199
rect 675943 650555 717600 650723
rect 675887 650079 717600 650555
rect 675943 649911 717600 650079
rect 675887 649527 717600 649911
rect 675943 649359 717600 649527
rect 675887 648883 717600 649359
rect 675943 648715 717600 648883
rect 675887 648239 717600 648715
rect 675943 648071 717600 648239
rect 675887 647687 717600 648071
rect 675943 647519 717600 647687
rect 675887 647043 717600 647519
rect 675943 646875 717600 647043
rect 675887 646399 717600 646875
rect 675407 646340 675887 646343
rect 675404 646287 675887 646340
rect 675404 645946 675432 646287
rect 675943 646231 717600 646399
rect 675220 645918 675432 645946
rect 675220 638858 675248 645918
rect 675887 645755 717600 646231
rect 675208 638794 675260 638858
rect 675208 600782 675260 600846
rect 675220 593314 675248 600782
rect 675943 645587 717600 645755
rect 675887 645203 717600 645587
rect 675943 645035 717600 645203
rect 675887 644559 717600 645035
rect 675943 644391 717600 644559
rect 675887 643915 717600 644391
rect 675943 643747 717600 643915
rect 675887 643363 717600 643747
rect 675407 643251 675887 643307
rect 675943 643195 717600 643363
rect 675887 642719 717600 643195
rect 675943 642551 717600 642719
rect 675887 642075 717600 642551
rect 675407 641963 675887 642019
rect 675943 641907 717600 642075
rect 675887 641523 717600 641907
rect 675943 641355 717600 641523
rect 675887 640879 717600 641355
rect 675943 640711 717600 640879
rect 675887 640235 717600 640711
rect 675943 640067 717600 640235
rect 675887 639683 717600 640067
rect 675407 639571 675887 639627
rect 675943 639515 717600 639683
rect 675887 639039 717600 639515
rect 675943 638871 717600 639039
rect 675392 638794 675444 638858
rect 675404 638339 675432 638794
rect 675887 638395 717600 638871
rect 675404 638316 675887 638339
rect 675407 638283 675887 638316
rect 675943 638227 717600 638395
rect 675887 638017 717600 638227
rect 675887 608759 717600 608958
rect 675407 608647 675887 608703
rect 675943 608591 717600 608759
rect 675887 608207 717600 608591
rect 675943 608039 717600 608207
rect 675887 607563 717600 608039
rect 675943 607395 717600 607563
rect 675887 606919 717600 607395
rect 675943 606751 717600 606919
rect 675887 606367 717600 606751
rect 675943 606199 717600 606367
rect 675887 605723 717600 606199
rect 675943 605555 717600 605723
rect 675887 605079 717600 605555
rect 675943 604911 717600 605079
rect 675887 604527 717600 604911
rect 675943 604359 717600 604527
rect 675887 603883 717600 604359
rect 675943 603715 717600 603883
rect 675887 603239 717600 603715
rect 675943 603071 717600 603239
rect 675887 602687 717600 603071
rect 675943 602519 717600 602687
rect 675887 602043 717600 602519
rect 675943 601875 717600 602043
rect 675887 601399 717600 601875
rect 675407 601324 675887 601343
rect 675404 601287 675887 601324
rect 675404 600846 675432 601287
rect 675943 601231 717600 601399
rect 675392 600782 675444 600846
rect 675887 600755 717600 601231
rect 675943 600587 717600 600755
rect 675887 600203 717600 600587
rect 675943 600035 717600 600203
rect 675887 599559 717600 600035
rect 675943 599391 717600 599559
rect 675887 598915 717600 599391
rect 675943 598747 717600 598915
rect 675887 598363 717600 598747
rect 675407 598251 675887 598307
rect 675943 598195 717600 598363
rect 675887 597719 717600 598195
rect 675943 597551 717600 597719
rect 675887 597075 717600 597551
rect 675407 596963 675887 597019
rect 675943 596907 717600 597075
rect 675887 596523 717600 596907
rect 675943 596355 717600 596523
rect 675887 595879 717600 596355
rect 675943 595711 717600 595879
rect 675887 595235 717600 595711
rect 675943 595067 717600 595235
rect 675887 594683 717600 595067
rect 675407 594571 675887 594627
rect 675943 594515 717600 594683
rect 675887 594039 717600 594515
rect 675943 593871 717600 594039
rect 675887 593395 717600 593871
rect 675407 593314 675887 593339
rect 675220 593286 675887 593314
rect 675407 593283 675887 593286
rect 675943 593227 717600 593395
rect 675887 593017 717600 593227
rect 675887 563559 717600 563758
rect 675407 563447 675887 563503
rect 675943 563391 717600 563559
rect 675887 563007 717600 563391
rect 675943 562839 717600 563007
rect 675887 562363 717600 562839
rect 675943 562195 717600 562363
rect 675887 561719 717600 562195
rect 675943 561551 717600 561719
rect 675887 561167 717600 561551
rect 675943 560999 717600 561167
rect 675887 560523 717600 560999
rect 675943 560355 717600 560523
rect 675887 559879 717600 560355
rect 675943 559711 717600 559879
rect 675887 559327 717600 559711
rect 675943 559159 717600 559327
rect 675887 558683 717600 559159
rect 675943 558515 717600 558683
rect 675887 558039 717600 558515
rect 675943 557871 717600 558039
rect 675887 557487 717600 557871
rect 675943 557319 717600 557487
rect 675887 556843 717600 557319
rect 675943 556675 717600 556843
rect 675887 556199 717600 556675
rect 675407 556129 675887 556143
rect 675312 556101 675887 556129
rect 675312 548570 675340 556101
rect 675407 556087 675887 556101
rect 675943 556031 717600 556199
rect 675887 555555 717600 556031
rect 675943 555387 717600 555555
rect 675887 555003 717600 555387
rect 675943 554835 717600 555003
rect 675887 554359 717600 554835
rect 675943 554191 717600 554359
rect 675887 553715 717600 554191
rect 675943 553547 717600 553715
rect 675887 553163 717600 553547
rect 675407 553051 675887 553107
rect 675943 552995 717600 553163
rect 675887 552519 717600 552995
rect 675943 552351 717600 552519
rect 675887 551875 717600 552351
rect 675407 551763 675887 551819
rect 675943 551707 717600 551875
rect 675887 551323 717600 551707
rect 675943 551155 717600 551323
rect 675887 550679 717600 551155
rect 675943 550511 717600 550679
rect 675887 550035 717600 550511
rect 675943 549867 717600 550035
rect 675887 549483 717600 549867
rect 675407 549371 675887 549427
rect 675943 549315 717600 549483
rect 675887 548839 717600 549315
rect 675943 548671 717600 548839
rect 675312 548542 675432 548570
rect 675404 548139 675432 548542
rect 675887 548195 717600 548671
rect 675404 548111 675887 548139
rect 675407 548083 675887 548111
rect 675943 548027 717600 548195
rect 675887 547817 717600 548027
rect 678007 518701 716615 518747
rect 677600 513921 716615 518701
rect 677600 513221 677984 513621
rect 678007 508722 716615 513921
rect 677600 503942 716615 508722
rect 678000 470701 716886 474700
rect 678007 470615 716886 470701
rect 678000 464093 716886 470615
rect 678007 463981 716886 464093
rect 678000 459860 716886 463981
rect 678007 459800 716886 459860
rect 684898 457561 685672 459751
rect 685917 457572 686847 459800
rect 678007 430501 716615 430547
rect 677600 425721 716615 430501
rect 677600 425021 677984 425421
rect 678007 420522 716615 425721
rect 677600 415742 716615 420522
rect 42340 326334 42392 326398
rect 42352 319462 42380 326334
rect 42340 319398 42392 319462
rect 42340 283154 42392 283218
rect 42352 276214 42380 283154
rect 42340 276150 42392 276214
rect 42340 239906 42392 239970
rect 42352 233034 42380 239906
rect 42340 232970 42392 233034
rect 675887 386359 717600 386558
rect 675407 386247 675887 386303
rect 675943 386191 717600 386359
rect 675887 385807 717600 386191
rect 675943 385639 717600 385807
rect 675887 385163 717600 385639
rect 675943 384995 717600 385163
rect 675887 384519 717600 384995
rect 675943 384351 717600 384519
rect 675887 383967 717600 384351
rect 675943 383799 717600 383967
rect 675887 383323 717600 383799
rect 675943 383155 717600 383323
rect 675887 382679 717600 383155
rect 675943 382511 717600 382679
rect 675887 382127 717600 382511
rect 675943 381959 717600 382127
rect 675887 381483 717600 381959
rect 675943 381315 717600 381483
rect 675887 380839 717600 381315
rect 675943 380671 717600 380839
rect 675887 380287 717600 380671
rect 675943 380119 717600 380287
rect 675887 379643 717600 380119
rect 675943 379475 717600 379643
rect 675887 378999 717600 379475
rect 675407 378929 675887 378943
rect 675312 378901 675887 378929
rect 675312 370925 675340 378901
rect 675407 378887 675887 378901
rect 675943 378831 717600 378999
rect 675887 378355 717600 378831
rect 675943 378187 717600 378355
rect 675887 377803 717600 378187
rect 675943 377635 717600 377803
rect 675887 377159 717600 377635
rect 675943 376991 717600 377159
rect 675887 376515 717600 376991
rect 675943 376347 717600 376515
rect 675887 375963 717600 376347
rect 675407 375851 675887 375907
rect 675943 375795 717600 375963
rect 675887 375319 717600 375795
rect 675943 375151 717600 375319
rect 675887 374675 717600 375151
rect 675407 374563 675887 374619
rect 675943 374507 717600 374675
rect 675887 374123 717600 374507
rect 675407 374011 675887 374067
rect 675943 373955 717600 374123
rect 675887 373479 717600 373955
rect 675943 373311 717600 373479
rect 675887 372835 717600 373311
rect 675943 372667 717600 372835
rect 675887 372283 717600 372667
rect 675407 372171 675887 372227
rect 675943 372115 717600 372283
rect 675887 371639 717600 372115
rect 675943 371471 717600 371639
rect 675887 370995 717600 371471
rect 675407 370925 675887 370939
rect 675312 370897 675887 370925
rect 675407 370883 675887 370897
rect 675943 370827 717600 370995
rect 675887 370617 717600 370827
rect 675887 341159 717600 341358
rect 675407 341047 675887 341103
rect 675943 340991 717600 341159
rect 675887 340607 717600 340991
rect 675943 340439 717600 340607
rect 675887 339963 717600 340439
rect 675943 339795 717600 339963
rect 675887 339319 717600 339795
rect 675943 339151 717600 339319
rect 675887 338767 717600 339151
rect 675943 338599 717600 338767
rect 675887 338123 717600 338599
rect 675943 337955 717600 338123
rect 675887 337479 717600 337955
rect 675943 337311 717600 337479
rect 675887 336927 717600 337311
rect 675943 336759 717600 336927
rect 675887 336283 717600 336759
rect 675943 336115 717600 336283
rect 675887 335639 717600 336115
rect 675943 335471 717600 335639
rect 675887 335087 717600 335471
rect 675943 334919 717600 335087
rect 675887 334443 717600 334919
rect 675943 334275 717600 334443
rect 675887 333799 717600 334275
rect 675407 333729 675887 333743
rect 675312 333701 675887 333729
rect 675312 325725 675340 333701
rect 675407 333687 675887 333701
rect 675943 333631 717600 333799
rect 675887 333155 717600 333631
rect 675943 332987 717600 333155
rect 675887 332603 717600 332987
rect 675943 332435 717600 332603
rect 675887 331959 717600 332435
rect 675943 331791 717600 331959
rect 675887 331315 717600 331791
rect 675943 331147 717600 331315
rect 675887 330763 717600 331147
rect 675407 330651 675887 330707
rect 675943 330595 717600 330763
rect 675887 330119 717600 330595
rect 675943 329951 717600 330119
rect 675887 329475 717600 329951
rect 675407 329363 675887 329419
rect 675943 329307 717600 329475
rect 675887 328923 717600 329307
rect 675407 328811 675887 328867
rect 675943 328755 717600 328923
rect 675887 328279 717600 328755
rect 675943 328111 717600 328279
rect 675887 327635 717600 328111
rect 675943 327467 717600 327635
rect 675887 327083 717600 327467
rect 675407 326971 675887 327027
rect 675943 326915 717600 327083
rect 675887 326439 717600 326915
rect 675943 326271 717600 326439
rect 675887 325795 717600 326271
rect 675407 325725 675887 325739
rect 675312 325697 675887 325725
rect 675407 325683 675887 325697
rect 675943 325627 717600 325795
rect 675887 325417 717600 325627
rect 675887 296159 717600 296358
rect 675407 296047 675887 296103
rect 675943 295991 717600 296159
rect 675887 295607 717600 295991
rect 675943 295439 717600 295607
rect 675887 294963 717600 295439
rect 675943 294795 717600 294963
rect 675887 294319 717600 294795
rect 675943 294151 717600 294319
rect 675887 293767 717600 294151
rect 42340 196726 42392 196790
rect 42352 189854 42380 196726
rect 42340 189790 42392 189854
rect 985 115079 39593 120278
rect 39616 115379 40000 115779
rect 985 110299 40000 115079
rect 985 110253 39593 110299
rect 7 83240 30281 85187
rect 30753 83000 31683 85228
rect 32033 83240 34915 85187
rect 7 82940 39593 83000
rect 7 78819 39600 82940
rect 7 78707 39593 78819
rect 7 72185 39600 78707
rect 7 72099 39593 72185
rect 7 68100 39600 72099
rect 7 68000 39593 68100
rect 30760 65805 31690 68000
rect 675943 293599 717600 293767
rect 675887 293123 717600 293599
rect 675943 292955 717600 293123
rect 675887 292479 717600 292955
rect 675943 292311 717600 292479
rect 675887 291927 717600 292311
rect 675943 291759 717600 291927
rect 675887 291283 717600 291759
rect 675943 291115 717600 291283
rect 675887 290639 717600 291115
rect 675943 290471 717600 290639
rect 675887 290087 717600 290471
rect 675943 289919 717600 290087
rect 675887 289443 717600 289919
rect 675943 289275 717600 289443
rect 675887 288799 717600 289275
rect 675407 288729 675887 288743
rect 675312 288701 675887 288729
rect 675312 280725 675340 288701
rect 675407 288687 675887 288701
rect 675943 288631 717600 288799
rect 675887 288155 717600 288631
rect 675943 287987 717600 288155
rect 675887 287603 717600 287987
rect 675943 287435 717600 287603
rect 675887 286959 717600 287435
rect 675943 286791 717600 286959
rect 675887 286315 717600 286791
rect 675943 286147 717600 286315
rect 675887 285763 717600 286147
rect 675407 285651 675887 285707
rect 675943 285595 717600 285763
rect 675887 285119 717600 285595
rect 675943 284951 717600 285119
rect 675887 284475 717600 284951
rect 675407 284363 675887 284419
rect 675943 284307 717600 284475
rect 675887 283923 717600 284307
rect 675407 283811 675887 283867
rect 675943 283755 717600 283923
rect 675887 283279 717600 283755
rect 675943 283111 717600 283279
rect 675887 282635 717600 283111
rect 675943 282467 717600 282635
rect 675887 282083 717600 282467
rect 675407 281971 675887 282027
rect 675943 281915 717600 282083
rect 675887 281439 717600 281915
rect 675943 281271 717600 281439
rect 675887 280795 717600 281271
rect 675407 280725 675887 280739
rect 675312 280697 675887 280725
rect 675407 280683 675887 280697
rect 675943 280627 717600 280795
rect 675887 280417 717600 280627
rect 675887 251159 717600 251358
rect 675407 251047 675887 251103
rect 675943 250991 717600 251159
rect 675887 250607 717600 250991
rect 675943 250439 717600 250607
rect 675887 249963 717600 250439
rect 675943 249795 717600 249963
rect 675887 249319 717600 249795
rect 675943 249151 717600 249319
rect 675887 248767 717600 249151
rect 675943 248599 717600 248767
rect 675887 248123 717600 248599
rect 675943 247955 717600 248123
rect 675887 247479 717600 247955
rect 675943 247311 717600 247479
rect 675887 246927 717600 247311
rect 675943 246759 717600 246927
rect 675887 246283 717600 246759
rect 675943 246115 717600 246283
rect 675887 245639 717600 246115
rect 675943 245471 717600 245639
rect 675887 245087 717600 245471
rect 675943 244919 717600 245087
rect 675887 244443 717600 244919
rect 675943 244275 717600 244443
rect 675887 243799 717600 244275
rect 675407 243729 675887 243743
rect 675312 243701 675887 243729
rect 675312 235725 675340 243701
rect 675407 243687 675887 243701
rect 675943 243631 717600 243799
rect 675887 243155 717600 243631
rect 675943 242987 717600 243155
rect 675887 242603 717600 242987
rect 675943 242435 717600 242603
rect 675887 241959 717600 242435
rect 675943 241791 717600 241959
rect 675887 241315 717600 241791
rect 675943 241147 717600 241315
rect 675887 240763 717600 241147
rect 675407 240651 675887 240707
rect 675943 240595 717600 240763
rect 675887 240119 717600 240595
rect 675943 239951 717600 240119
rect 675887 239475 717600 239951
rect 675407 239363 675887 239419
rect 675943 239307 717600 239475
rect 675887 238923 717600 239307
rect 675407 238811 675887 238867
rect 675943 238755 717600 238923
rect 675887 238279 717600 238755
rect 675943 238111 717600 238279
rect 675887 237635 717600 238111
rect 675943 237467 717600 237635
rect 675887 237083 717600 237467
rect 675407 236971 675887 237027
rect 675943 236915 717600 237083
rect 675887 236439 717600 236915
rect 675943 236271 717600 236439
rect 675887 235795 717600 236271
rect 675407 235725 675887 235739
rect 675312 235697 675887 235725
rect 675407 235683 675887 235697
rect 675943 235627 717600 235795
rect 675887 235417 717600 235627
rect 675887 205959 717600 206158
rect 675407 205847 675887 205903
rect 675943 205791 717600 205959
rect 675887 205407 717600 205791
rect 675943 205239 717600 205407
rect 675887 204763 717600 205239
rect 675943 204595 717600 204763
rect 675887 204119 717600 204595
rect 675943 203951 717600 204119
rect 675887 203567 717600 203951
rect 675943 203399 717600 203567
rect 675887 202923 717600 203399
rect 675943 202755 717600 202923
rect 675887 202279 717600 202755
rect 675943 202111 717600 202279
rect 675887 201727 717600 202111
rect 675943 201559 717600 201727
rect 675887 201083 717600 201559
rect 675943 200915 717600 201083
rect 675887 200439 717600 200915
rect 675943 200271 717600 200439
rect 675887 199887 717600 200271
rect 675943 199719 717600 199887
rect 675887 199243 717600 199719
rect 675943 199075 717600 199243
rect 675312 198614 675432 198642
rect 675312 190525 675340 198614
rect 675404 198543 675432 198614
rect 675887 198599 717600 199075
rect 675404 198492 675887 198543
rect 675407 198487 675887 198492
rect 675943 198431 717600 198599
rect 675887 197955 717600 198431
rect 675943 197787 717600 197955
rect 675887 197403 717600 197787
rect 675943 197235 717600 197403
rect 675887 196759 717600 197235
rect 675943 196591 717600 196759
rect 675887 196115 717600 196591
rect 675943 195947 717600 196115
rect 675887 195563 717600 195947
rect 675407 195451 675887 195507
rect 675943 195395 717600 195563
rect 675887 194919 717600 195395
rect 675943 194751 717600 194919
rect 675887 194275 717600 194751
rect 675407 194163 675887 194219
rect 675943 194107 717600 194275
rect 675887 193723 717600 194107
rect 675407 193611 675887 193667
rect 675943 193555 717600 193723
rect 675887 193079 717600 193555
rect 675943 192911 717600 193079
rect 675887 192435 717600 192911
rect 675943 192267 717600 192435
rect 675887 191883 717600 192267
rect 675407 191771 675887 191827
rect 675943 191715 717600 191883
rect 675887 191239 717600 191715
rect 675943 191071 717600 191239
rect 675887 190595 717600 191071
rect 675407 190525 675887 190539
rect 675312 190497 675887 190525
rect 675407 190483 675887 190497
rect 675943 190427 717600 190595
rect 675887 190217 717600 190427
rect 675887 160959 717600 161158
rect 675407 160847 675887 160903
rect 675943 160791 717600 160959
rect 675887 160407 717600 160791
rect 675943 160239 717600 160407
rect 675887 159763 717600 160239
rect 675943 159595 717600 159763
rect 675887 159119 717600 159595
rect 675943 158951 717600 159119
rect 675887 158567 717600 158951
rect 675943 158399 717600 158567
rect 675887 157923 717600 158399
rect 675943 157755 717600 157923
rect 675887 157279 717600 157755
rect 675943 157111 717600 157279
rect 675887 156727 717600 157111
rect 675943 156559 717600 156727
rect 675887 156083 717600 156559
rect 675943 155915 717600 156083
rect 675887 155439 717600 155915
rect 675943 155271 717600 155439
rect 675887 154887 717600 155271
rect 675943 154719 717600 154887
rect 675887 154243 717600 154719
rect 675943 154075 717600 154243
rect 675887 153599 717600 154075
rect 675407 153529 675887 153543
rect 675312 153501 675887 153529
rect 675312 145525 675340 153501
rect 675407 153487 675887 153501
rect 675943 153431 717600 153599
rect 675887 152955 717600 153431
rect 675943 152787 717600 152955
rect 675887 152403 717600 152787
rect 675943 152235 717600 152403
rect 675887 151759 717600 152235
rect 675943 151591 717600 151759
rect 675887 151115 717600 151591
rect 675943 150947 717600 151115
rect 675887 150563 717600 150947
rect 675407 150451 675887 150507
rect 675943 150395 717600 150563
rect 675887 149919 717600 150395
rect 675943 149751 717600 149919
rect 675887 149275 717600 149751
rect 675407 149163 675887 149219
rect 675943 149107 717600 149275
rect 675887 148723 717600 149107
rect 675407 148611 675887 148667
rect 675943 148555 717600 148723
rect 675887 148079 717600 148555
rect 675943 147911 717600 148079
rect 675887 147435 717600 147911
rect 675943 147267 717600 147435
rect 675887 146883 717600 147267
rect 675407 146771 675887 146827
rect 675943 146715 717600 146883
rect 675887 146239 717600 146715
rect 675943 146071 717600 146239
rect 675887 145595 717600 146071
rect 675407 145525 675887 145539
rect 675312 145497 675887 145525
rect 675407 145483 675887 145497
rect 675943 145427 717600 145595
rect 675887 145217 717600 145427
rect 135168 40225 135220 40254
rect 135166 40151 135222 40225
rect 143540 40225 143592 40254
rect 143538 40151 143594 40225
rect 186688 44202 186740 44266
rect 186700 42193 186728 44202
rect 194692 44202 194744 44266
rect 194704 42193 194732 44202
rect 186683 41713 186739 42193
rect 187971 41713 188027 42193
rect 189811 41713 189867 42193
rect 190363 41713 190419 42193
rect 191651 41713 191707 42193
rect 194687 41713 194743 42193
rect 202047 41713 202103 42193
rect 186417 41657 186627 41713
rect 186795 41657 187271 41713
rect 187439 41657 187915 41713
rect 188083 41657 188467 41713
rect 188635 41657 189111 41713
rect 189279 41657 189755 41713
rect 189923 41657 190307 41713
rect 190475 41657 190951 41713
rect 191119 41657 191595 41713
rect 191763 41657 192147 41713
rect 192315 41657 192791 41713
rect 192959 41657 193435 41713
rect 193603 41657 193987 41713
rect 194155 41657 194631 41713
rect 194799 41657 195275 41713
rect 195443 41657 195919 41713
rect 196087 41657 196471 41713
rect 196639 41657 197115 41713
rect 197283 41657 197759 41713
rect 197927 41657 198311 41713
rect 198479 41657 198955 41713
rect 199123 41657 199599 41713
rect 199767 41657 200151 41713
rect 200319 41657 200795 41713
rect 200963 41657 201439 41713
rect 201607 41657 201991 41713
rect 202159 41657 202358 41713
rect 78942 39593 83722 40000
rect 88221 39616 88621 40000
rect 88921 39593 93701 40000
rect 132617 39878 132897 40000
rect 132953 39934 133157 40000
rect 133213 39878 140940 40000
rect 132617 39816 140940 39878
rect 141104 39878 141313 40000
rect 141369 39934 141499 40000
rect 141555 39878 141611 40000
rect 141869 39878 141898 40000
rect 141954 39934 142084 40000
rect 142140 39878 143012 40000
rect 141104 39816 143012 39878
rect 78942 985 93747 39593
rect 132617 39450 143012 39816
rect 143184 39662 143299 40000
rect 143355 39718 143585 40000
rect 143641 39831 143762 40000
rect 143818 39887 144151 40000
rect 144207 39831 144517 40000
rect 143641 39747 144517 39831
rect 144745 39747 145035 40000
rect 143641 39662 145035 39747
rect 145199 39878 145765 40000
rect 145821 39934 145915 40000
rect 145971 39878 147532 40000
rect 143184 39650 145035 39662
rect 145199 39650 147532 39878
rect 143184 39450 147532 39650
rect 132617 158 147532 39450
rect 186417 0 202358 41657
rect 295248 44134 295300 44198
rect 295260 42193 295288 44134
rect 303252 44134 303304 44198
rect 303264 42193 303292 44134
rect 350080 44134 350132 44198
rect 350092 42193 350120 44134
rect 358084 44134 358136 44198
rect 358096 42193 358124 44134
rect 404912 44134 404964 44198
rect 404924 42193 404952 44134
rect 412916 44134 412968 44198
rect 412928 42193 412956 44134
rect 459652 44134 459704 44198
rect 459664 42193 459692 44134
rect 467656 44134 467708 44198
rect 467668 42193 467696 44134
rect 514484 44134 514536 44198
rect 514496 42193 514524 44134
rect 522488 44134 522540 44198
rect 522500 42193 522528 44134
rect 675887 115759 717600 115958
rect 675407 115647 675887 115703
rect 675943 115591 717600 115759
rect 675887 115207 717600 115591
rect 675943 115039 717600 115207
rect 675887 114563 717600 115039
rect 675943 114395 717600 114563
rect 675887 113919 717600 114395
rect 675943 113751 717600 113919
rect 675887 113367 717600 113751
rect 675943 113199 717600 113367
rect 675887 112723 717600 113199
rect 675943 112555 717600 112723
rect 675887 112079 717600 112555
rect 675943 111911 717600 112079
rect 675887 111527 717600 111911
rect 675943 111359 717600 111527
rect 675887 110883 717600 111359
rect 675943 110715 717600 110883
rect 675887 110239 717600 110715
rect 675943 110071 717600 110239
rect 675887 109687 717600 110071
rect 675943 109519 717600 109687
rect 675887 109043 717600 109519
rect 675943 108875 717600 109043
rect 675887 108399 717600 108875
rect 675407 108338 675887 108343
rect 675312 108310 675887 108338
rect 675312 100314 675340 108310
rect 675407 108287 675887 108310
rect 675943 108231 717600 108399
rect 675887 107755 717600 108231
rect 675943 107587 717600 107755
rect 675887 107203 717600 107587
rect 675943 107035 717600 107203
rect 675887 106559 717600 107035
rect 675943 106391 717600 106559
rect 675887 105915 717600 106391
rect 675943 105747 717600 105915
rect 675887 105363 717600 105747
rect 675407 105251 675887 105307
rect 675943 105195 717600 105363
rect 675887 104719 717600 105195
rect 675943 104551 717600 104719
rect 675887 104075 717600 104551
rect 675407 103963 675887 104019
rect 675943 103907 717600 104075
rect 675887 103523 717600 103907
rect 675407 103411 675887 103467
rect 675943 103355 717600 103523
rect 675887 102879 717600 103355
rect 675943 102711 717600 102879
rect 675887 102235 717600 102711
rect 675943 102067 717600 102235
rect 675887 101683 717600 102067
rect 675407 101571 675887 101627
rect 675943 101515 717600 101683
rect 675887 101039 717600 101515
rect 675943 100871 717600 101039
rect 675887 100395 717600 100871
rect 675407 100314 675887 100339
rect 675312 100286 675887 100314
rect 675407 100283 675887 100286
rect 675943 100227 717600 100395
rect 675887 100017 717600 100227
rect 295260 41806 295339 42193
rect 295283 41713 295339 41806
rect 295927 41713 295983 42193
rect 296571 41713 296627 42193
rect 298411 41713 298467 42193
rect 298963 41713 299019 42193
rect 300251 41713 300307 42193
rect 303264 41806 303343 42193
rect 303287 41713 303343 41806
rect 310647 41713 310703 42193
rect 295017 41657 295227 41713
rect 295395 41657 295871 41713
rect 296039 41657 296515 41713
rect 296683 41657 297067 41713
rect 297235 41657 297711 41713
rect 297879 41657 298355 41713
rect 298523 41657 298907 41713
rect 299075 41657 299551 41713
rect 299719 41657 300195 41713
rect 300363 41657 300747 41713
rect 300915 41657 301391 41713
rect 301559 41657 302035 41713
rect 302203 41657 302587 41713
rect 302755 41657 303231 41713
rect 303399 41657 303875 41713
rect 304043 41657 304519 41713
rect 304687 41657 305071 41713
rect 305239 41657 305715 41713
rect 305883 41657 306359 41713
rect 306527 41657 306911 41713
rect 307079 41657 307555 41713
rect 307723 41657 308199 41713
rect 308367 41657 308751 41713
rect 308919 41657 309395 41713
rect 309563 41657 310039 41713
rect 310207 41657 310591 41713
rect 310759 41657 310958 41713
rect 241260 39593 245381 39600
rect 245493 39593 252015 39600
rect 252101 39593 256100 39600
rect 239013 32033 240960 34915
rect 241200 31690 256200 39593
rect 241200 31683 258395 31690
rect 238972 30760 258395 31683
rect 238972 30753 256200 30760
rect 239013 7 240960 30281
rect 241200 7 256200 30753
rect 295017 0 310958 41657
rect 350083 41713 350139 42193
rect 350727 41713 350783 42193
rect 351371 41713 351427 42193
rect 353211 41713 353267 42193
rect 353763 41713 353819 42193
rect 355051 41713 355107 42193
rect 358087 41713 358143 42193
rect 365447 41713 365503 42193
rect 349817 41657 350027 41713
rect 350195 41657 350671 41713
rect 350839 41657 351315 41713
rect 351483 41657 351867 41713
rect 352035 41657 352511 41713
rect 352679 41657 353155 41713
rect 353323 41657 353707 41713
rect 353875 41657 354351 41713
rect 354519 41657 354995 41713
rect 355163 41657 355547 41713
rect 355715 41657 356191 41713
rect 356359 41657 356835 41713
rect 357003 41657 357387 41713
rect 357555 41657 358031 41713
rect 358199 41657 358675 41713
rect 358843 41657 359319 41713
rect 359487 41657 359871 41713
rect 360039 41657 360515 41713
rect 360683 41657 361159 41713
rect 361327 41657 361711 41713
rect 361879 41657 362355 41713
rect 362523 41657 362999 41713
rect 363167 41657 363551 41713
rect 363719 41657 364195 41713
rect 364363 41657 364839 41713
rect 365007 41657 365391 41713
rect 365559 41657 365758 41713
rect 349817 0 365758 41657
rect 404883 41820 404952 42193
rect 404883 41713 404939 41820
rect 406171 41713 406227 42193
rect 408011 41713 408067 42193
rect 408563 41713 408619 42193
rect 409851 41713 409907 42193
rect 412887 41820 412956 42193
rect 412887 41713 412943 41820
rect 420247 41713 420303 42193
rect 459664 41806 459739 42193
rect 459683 41713 459739 41806
rect 460971 41713 461027 42193
rect 462811 41713 462867 42193
rect 463363 41713 463419 42193
rect 464651 41713 464707 42193
rect 467668 41806 467743 42193
rect 467687 41713 467743 41806
rect 475047 41713 475103 42193
rect 514483 41713 514539 42193
rect 515771 41713 515827 42193
rect 517611 41713 517667 42193
rect 518163 41713 518219 42193
rect 519451 41713 519507 42193
rect 522487 41713 522543 42193
rect 529847 41713 529903 42193
rect 404617 41657 404827 41713
rect 404995 41657 405471 41713
rect 405639 41657 406115 41713
rect 406283 41657 406667 41713
rect 406835 41657 407311 41713
rect 407479 41657 407955 41713
rect 408123 41657 408507 41713
rect 408675 41657 409151 41713
rect 409319 41657 409795 41713
rect 409963 41657 410347 41713
rect 410515 41657 410991 41713
rect 411159 41657 411635 41713
rect 411803 41657 412187 41713
rect 412355 41657 412831 41713
rect 412999 41657 413475 41713
rect 413643 41657 414119 41713
rect 414287 41657 414671 41713
rect 414839 41657 415315 41713
rect 415483 41657 415959 41713
rect 416127 41657 416511 41713
rect 416679 41657 417155 41713
rect 417323 41657 417799 41713
rect 417967 41657 418351 41713
rect 418519 41657 418995 41713
rect 419163 41657 419639 41713
rect 419807 41657 420191 41713
rect 420359 41657 420558 41713
rect 404617 0 420558 41657
rect 459417 41657 459627 41713
rect 459795 41657 460271 41713
rect 460439 41657 460915 41713
rect 461083 41657 461467 41713
rect 461635 41657 462111 41713
rect 462279 41657 462755 41713
rect 462923 41657 463307 41713
rect 463475 41657 463951 41713
rect 464119 41657 464595 41713
rect 464763 41657 465147 41713
rect 465315 41657 465791 41713
rect 465959 41657 466435 41713
rect 466603 41657 466987 41713
rect 467155 41657 467631 41713
rect 467799 41657 468275 41713
rect 468443 41657 468919 41713
rect 469087 41657 469471 41713
rect 469639 41657 470115 41713
rect 470283 41657 470759 41713
rect 470927 41657 471311 41713
rect 471479 41657 471955 41713
rect 472123 41657 472599 41713
rect 472767 41657 473151 41713
rect 473319 41657 473795 41713
rect 473963 41657 474439 41713
rect 474607 41657 474991 41713
rect 475159 41657 475358 41713
rect 459417 0 475358 41657
rect 514217 41657 514427 41713
rect 514595 41657 515071 41713
rect 515239 41657 515715 41713
rect 515883 41657 516267 41713
rect 516435 41657 516911 41713
rect 517079 41657 517555 41713
rect 517723 41657 518107 41713
rect 518275 41657 518751 41713
rect 518919 41657 519395 41713
rect 519563 41657 519947 41713
rect 520115 41657 520591 41713
rect 520759 41657 521235 41713
rect 521403 41657 521787 41713
rect 521955 41657 522431 41713
rect 522599 41657 523075 41713
rect 523243 41657 523719 41713
rect 523887 41657 524271 41713
rect 524439 41657 524915 41713
rect 525083 41657 525559 41713
rect 525727 41657 526111 41713
rect 526279 41657 526755 41713
rect 526923 41657 527399 41713
rect 527567 41657 527951 41713
rect 528119 41657 528595 41713
rect 528763 41657 529239 41713
rect 529407 41657 529791 41713
rect 529959 41657 530158 41713
rect 514217 0 530158 41657
rect 569142 39593 573922 40000
rect 578421 39616 578821 40000
rect 579121 39593 583901 40000
rect 622942 39593 627722 40000
rect 632221 39616 632621 40000
rect 632921 39593 637701 40000
rect 569142 985 583947 39593
rect 622942 985 637747 39593
<< metal3 >>
rect 333499 997600 338279 1002770
rect 343478 997600 348258 1002770
rect 342159 997478 342229 997479
rect 343590 997478 343650 997600
rect 342159 997474 343650 997478
rect 342159 997414 342164 997474
rect 342224 997418 343650 997474
rect 342224 997414 342229 997418
rect 342159 997409 342229 997414
rect 575699 997600 580479 1004103
rect 585678 997600 590458 1004952
rect 585039 997448 585109 997453
rect 585039 997388 585044 997448
rect 585104 997446 585109 997448
rect 585734 997446 585794 997600
rect 585104 997388 585794 997446
rect 585039 997386 585794 997388
rect 585039 997383 585109 997386
rect 121269 990450 121335 990453
rect 131021 990450 131087 990453
rect 121269 990448 131087 990450
rect 121269 990392 121274 990448
rect 121330 990392 131026 990448
rect 131082 990392 131087 990448
rect 121269 990390 131087 990392
rect 121269 990387 121335 990390
rect 131021 990387 131087 990390
rect 38220 922151 39600 926940
rect 678000 917700 679380 922500
rect 38220 912100 39600 916900
rect 678000 907660 679380 912449
rect 36040 870090 40000 874679
rect 42241 870090 42307 870093
rect 36040 870088 42307 870090
rect 36040 870032 42246 870088
rect 42302 870032 42307 870088
rect 36040 870030 42307 870032
rect 36040 869899 40000 870030
rect 42241 870027 42307 870030
rect 32648 837678 40000 842458
rect 33497 827699 40000 832479
rect 677600 828521 680592 833301
rect 677600 818542 680592 823322
rect 677501 818410 677567 818413
rect 677734 818410 677794 818542
rect 677501 818408 677794 818410
rect 677501 818352 677506 818408
rect 677562 818352 677794 818408
rect 677501 818350 677794 818352
rect 677501 818347 677567 818350
rect 673729 521658 673795 521661
rect 674005 521658 674071 521661
rect 673729 521656 674071 521658
rect 673729 521600 673734 521656
rect 673790 521600 674010 521656
rect 674066 521600 674071 521656
rect 673729 521598 674071 521600
rect 673729 521595 673795 521598
rect 674005 521595 674071 521598
rect 677600 513921 680592 518701
rect 677734 513773 677794 513921
rect 677685 513768 677794 513773
rect 677685 513712 677690 513768
rect 677746 513712 677794 513768
rect 677685 513710 677794 513712
rect 677685 513707 677751 513710
rect 37008 493078 40000 497858
rect 37008 483099 40000 487879
rect 678000 469900 685920 474700
rect 678000 459860 685920 464649
rect 31680 450951 39600 455740
rect 31680 440900 39600 445700
rect 677315 427852 677385 427857
rect 677600 427852 684103 430501
rect 677315 427792 677320 427852
rect 677380 427792 684103 427852
rect 677315 427787 677385 427792
rect 677600 425721 684103 427792
rect 673637 154594 673703 154597
rect 673821 154594 673887 154597
rect 673637 154592 673887 154594
rect 673637 154536 673642 154592
rect 673698 154536 673826 154592
rect 673882 154536 673887 154592
rect 673637 154534 673887 154536
rect 673637 154531 673703 154534
rect 673821 154531 673887 154534
rect 36040 120278 40000 125058
rect 36040 110394 40000 115079
rect 42977 110394 43043 110397
rect 36040 110392 43043 110394
rect 36040 110336 42982 110392
rect 43038 110336 43043 110392
rect 36040 110334 43043 110336
rect 36040 110299 40000 110334
rect 42977 110331 43043 110334
rect 42977 96658 43043 96661
rect 44633 96658 44699 96661
rect 42977 96656 44699 96658
rect 42977 96600 42982 96656
rect 43038 96600 44638 96656
rect 44694 96600 44699 96656
rect 42977 96598 44699 96600
rect 42977 96595 43043 96598
rect 44633 96595 44699 96598
rect 38220 78298 39600 82940
rect 41413 80610 41479 80613
rect 42701 80610 42767 80613
rect 41413 80608 42767 80610
rect 41413 80552 41418 80608
rect 41474 80552 42706 80608
rect 42762 80552 42767 80608
rect 41413 80550 42767 80552
rect 41413 80547 41479 80550
rect 42701 80547 42767 80550
rect 41413 78298 41479 78301
rect 38220 78296 41479 78298
rect 38220 78240 41418 78296
rect 41474 78240 41479 78296
rect 38220 78238 41479 78240
rect 38220 78151 39600 78238
rect 41413 78235 41479 78238
rect 38220 68100 39600 72900
rect 483013 44706 483079 44709
rect 502057 44706 502123 44709
rect 483013 44704 502123 44706
rect 483013 44648 483018 44704
rect 483074 44648 502062 44704
rect 502118 44648 502123 44704
rect 483013 44646 502123 44648
rect 483013 44643 483079 44646
rect 502057 44643 502123 44646
rect 386413 44570 386479 44573
rect 405641 44570 405707 44573
rect 386413 44568 405707 44570
rect 386413 44512 386418 44568
rect 386474 44512 405646 44568
rect 405702 44512 405707 44568
rect 386413 44510 405707 44512
rect 386413 44507 386479 44510
rect 405641 44507 405707 44510
rect 465809 44298 465875 44301
rect 474457 44298 474523 44301
rect 465809 44296 474523 44298
rect 465809 44240 465814 44296
rect 465870 44240 474462 44296
rect 474518 44240 474523 44296
rect 465809 44238 474523 44240
rect 465809 44235 465875 44238
rect 474457 44235 474523 44238
rect 518801 44298 518867 44301
rect 524965 44298 525031 44301
rect 518801 44296 525031 44298
rect 518801 44240 518806 44296
rect 518862 44240 524970 44296
rect 525026 44240 525031 44296
rect 518801 44238 525031 44240
rect 518801 44235 518867 44238
rect 524965 44235 525031 44238
rect 367093 41986 367159 41989
rect 386137 41986 386203 41989
rect 367093 41984 386203 41986
rect 367093 41928 367098 41984
rect 367154 41928 386142 41984
rect 386198 41928 386203 41984
rect 367093 41926 386203 41928
rect 367093 41923 367159 41926
rect 386137 41923 386203 41926
rect 349613 41850 349679 41853
rect 362401 41850 362467 41853
rect 349613 41848 362467 41850
rect 349613 41792 349618 41848
rect 349674 41792 362406 41848
rect 362462 41792 362467 41848
rect 349613 41790 362467 41792
rect 349613 41787 349679 41790
rect 362401 41787 362467 41790
rect 143533 40490 143599 40493
rect 143533 40488 145850 40490
rect 143533 40432 143538 40488
rect 143594 40432 145850 40488
rect 143533 40430 145850 40432
rect 143533 40427 143599 40430
rect 145790 40354 145850 40430
rect 149605 40354 149671 40357
rect 145790 40352 149671 40354
rect 145790 40296 149610 40352
rect 149666 40296 149671 40352
rect 145790 40294 149671 40296
rect 93761 40218 93827 40221
rect 91142 40216 93827 40218
rect 91142 40160 93766 40216
rect 93822 40160 93827 40216
rect 91142 40158 93827 40160
rect 91142 40000 91202 40158
rect 93761 40155 93827 40158
rect 143073 40218 143139 40221
rect 143073 40216 143458 40218
rect 143073 40160 143078 40216
rect 143134 40160 143458 40216
rect 143073 40158 143458 40160
rect 143073 40155 143139 40158
rect 143398 40000 143458 40158
rect 145838 40014 145898 40294
rect 149605 40291 149671 40294
rect 145820 40000 145898 40014
rect 78942 32648 83722 40000
rect 88921 33497 93701 40000
rect 141667 39450 141813 40000
rect 143355 39450 143585 40000
rect 145816 39450 145920 40000
rect 241329 39946 241395 39949
rect 241286 39944 241395 39946
rect 241286 39888 241334 39944
rect 241390 39888 241395 39944
rect 241286 39883 241395 39888
rect 241286 39600 241346 39883
rect 241260 31680 246049 39600
rect 251300 31680 256100 39600
rect 569125 40218 569191 40221
rect 569125 40216 569234 40218
rect 569125 40160 569130 40216
rect 569186 40160 569234 40216
rect 569125 40155 569234 40160
rect 569174 40000 569234 40155
rect 569142 34830 573922 40000
rect 579121 34830 583901 40000
rect 622942 37008 627722 40000
rect 632921 37008 637701 40000
<< obsm3 >>
rect 76262 997338 92114 1037600
rect 127662 997338 143514 1037600
rect 179062 997338 194914 1037600
rect 230462 997338 246314 1037600
rect 282062 997338 297914 1037600
rect 333448 1002850 348258 1037600
rect 338359 998007 343398 1002850
rect 338579 997600 340779 998007
rect 340978 997600 343178 998007
rect 383862 997338 399714 1037600
rect 472862 997338 488714 1037600
rect 524262 997338 540114 1037600
rect 575648 1005032 590458 1036620
rect 575648 1004183 585598 1005032
rect 580559 998007 585598 1004183
rect 580779 997600 582979 998007
rect 583178 997600 585378 998007
rect 626062 997338 641914 1037600
rect 0 954262 40262 970114
rect 677338 951686 717600 967538
rect 30753 927121 31683 929228
rect 31961 927088 32654 929228
rect 879 922071 38140 927000
rect 879 921851 39593 922071
rect 879 919676 39600 921851
rect 879 919376 39593 919676
rect 879 917200 39600 919376
rect 679460 917620 716721 922502
rect 678007 917400 716721 917620
rect 879 916980 39593 917200
rect 879 912098 38140 916980
rect 678000 915224 716721 917400
rect 678007 914924 716721 915224
rect 678000 912749 716721 914924
rect 678007 912529 716721 912749
rect 679460 907600 716721 912529
rect 684946 905372 685639 907512
rect 685917 905372 686847 907479
rect 0 879798 35960 884658
rect 36040 879878 40000 884658
rect 0 879578 39593 879798
rect 0 877378 40000 879578
rect 0 877179 39593 877378
rect 0 874979 40000 877179
rect 0 874759 39593 874979
rect 0 869848 35960 874759
rect 677338 862486 717600 878338
rect 980 837598 32568 842458
rect 980 837378 39593 837598
rect 980 835178 40000 837378
rect 980 834979 39593 835178
rect 980 832779 40000 834979
rect 980 832559 39593 832779
rect 980 827648 33417 832559
rect 680672 828441 717600 833352
rect 678007 828221 717600 828441
rect 677600 826021 717600 828221
rect 678007 825822 717600 826021
rect 677600 823622 717600 825822
rect 678007 823402 717600 823622
rect 680672 818469 717600 823402
rect 0 784462 40262 800314
rect 677338 773286 717600 789138
rect 0 741262 40262 757114
rect 677338 728286 717600 744138
rect 0 698062 40262 713914
rect 677338 683286 717600 699138
rect 0 654862 40262 670714
rect 677338 638086 717600 653938
rect 0 611662 40262 627514
rect 677338 593086 717600 608938
rect 0 568462 40262 584314
rect 677338 547886 717600 563738
rect 0 525262 40262 541114
rect 680672 513841 717600 518752
rect 678007 513621 717600 513841
rect 677600 511421 717600 513621
rect 678007 511222 717600 511421
rect 677600 509022 717600 511222
rect 678007 508802 717600 509022
rect 677600 503942 680592 508722
rect 680672 503869 717600 508802
rect 0 492998 36928 497931
rect 0 492778 39593 492998
rect 0 490578 40000 492778
rect 0 490379 39593 490578
rect 0 488179 40000 490379
rect 0 487959 39593 488179
rect 0 483048 36928 487959
rect 686000 469820 716721 474700
rect 678007 469600 716721 469820
rect 678000 467424 716721 469600
rect 678007 467124 716721 467424
rect 678000 464949 716721 467124
rect 678007 464729 716721 464949
rect 686000 459800 716721 464729
rect 30753 455921 31683 458028
rect 31961 455888 32654 458028
rect 684946 457572 685639 459712
rect 685917 457572 686847 459679
rect 879 450871 31600 455800
rect 879 450651 39593 450871
rect 879 448476 39600 450651
rect 879 448176 39593 448476
rect 879 446000 39600 448176
rect 879 445780 39593 446000
rect 879 440900 31600 445780
rect 684183 425641 716620 430552
rect 678007 425421 716620 425641
rect 677600 423221 716620 425421
rect 678007 423022 716620 423221
rect 677600 420822 716620 423022
rect 678007 420602 716620 420822
rect 677600 415742 684952 420522
rect 685032 415742 716620 420602
rect 0 397662 40262 413514
rect 677338 370686 717600 386538
rect 0 354462 40262 370314
rect 0 311262 40262 327114
rect 677338 325486 717600 341338
rect 0 268062 40262 283914
rect 677338 280486 717600 296338
rect 0 224862 40262 240714
rect 677338 235486 717600 251338
rect 0 181662 40262 197514
rect 677338 190286 717600 206138
rect 677338 145286 717600 161138
rect 0 120198 35960 125058
rect 0 119978 39593 120198
rect 0 117778 40000 119978
rect 0 117579 39593 117778
rect 0 115379 40000 117579
rect 0 115159 39593 115379
rect 0 110248 35960 115159
rect 677338 100086 717600 115938
rect 7 83240 4850 85187
rect 30753 83121 31683 85228
rect 33910 83240 34840 85187
rect 7 78071 38140 83000
rect 7 77851 39593 78071
rect 7 75676 39600 77851
rect 7 75376 39593 75676
rect 7 73200 39600 75376
rect 7 72980 39593 73200
rect 7 68020 38140 72980
rect 7 68000 39593 68020
rect 30760 65805 31690 67821
rect 135161 40218 135227 40221
rect 133094 40158 135227 40218
rect 133094 40000 133154 40158
rect 135161 40155 135227 40158
rect 143533 40218 143599 40221
rect 143533 40158 144010 40218
rect 143533 40155 143599 40158
rect 143950 40000 144010 40158
rect 47600 32953 51202 36017
rect 51600 32953 55202 36017
rect 55600 32953 59202 36017
rect 59600 32953 63202 36017
rect 63600 32953 67202 36017
rect 67600 32953 71202 36017
rect 84022 39593 86222 40000
rect 86421 39593 88621 40000
rect 83802 33417 88841 39593
rect 83802 32568 93752 33417
rect 101400 32953 105002 36017
rect 105400 32953 109002 36017
rect 109400 32953 113002 36017
rect 113400 32953 117002 36017
rect 117400 32953 121002 36017
rect 121400 32953 125002 36017
rect 78942 980 93752 32568
rect 132660 30216 132868 39875
rect 132660 26680 132735 30216
rect 132948 30136 133162 40000
rect 132815 30016 133162 30136
rect 133242 39450 141587 39875
rect 141893 39450 143275 39875
rect 143665 39450 143738 39875
rect 143818 39450 144151 40000
rect 144231 39450 145736 39875
rect 146000 39450 147407 39875
rect 132815 30003 132948 30016
rect 132815 27080 133162 30003
rect 133242 27160 147407 39450
rect 155200 32953 158802 36017
rect 159200 32953 162802 36017
rect 163200 32953 166802 36017
rect 167200 32953 170802 36017
rect 171200 32953 174802 36017
rect 175200 32953 178802 36017
rect 132815 26760 133482 27080
rect 133562 26840 147407 27160
rect 132660 26360 133082 26680
rect 133162 26480 133762 26760
rect 133842 26560 147407 26840
rect 133162 26450 133949 26480
rect 133162 26440 133482 26450
rect 133482 26390 133739 26440
rect 133762 26390 133949 26450
rect 132660 26103 133402 26360
rect 133482 26293 133949 26390
rect 134029 26373 147407 26560
rect 133482 26270 133942 26293
rect 133482 26240 133739 26270
rect 133949 26240 134122 26293
rect 133482 26210 134122 26240
rect 133482 26183 133739 26210
rect 133739 26180 133929 26183
rect 133949 26180 134122 26210
rect 134202 26200 147407 26373
rect 133739 26120 134122 26180
rect 132660 25913 133659 26103
rect 133739 26090 134392 26120
rect 133739 26060 133929 26090
rect 134122 26060 134392 26090
rect 133739 26000 134392 26060
rect 133739 25993 133929 26000
rect 134122 25993 134392 26000
rect 132660 25720 133849 25913
rect 133929 25850 134392 25993
rect 134472 25930 147407 26200
rect 133929 25820 134628 25850
rect 133929 25800 134122 25820
rect 134122 25760 134364 25800
rect 134392 25760 134628 25820
rect 132660 25478 134042 25720
rect 134122 25584 134628 25760
rect 134122 25558 134364 25584
rect 134368 25558 134628 25584
rect 134364 25520 134628 25558
rect 132660 25440 134284 25478
rect 132660 20991 134322 25440
rect 134402 21071 134628 25520
rect 134708 20991 147407 25930
rect 132660 0 147407 20991
rect 186486 0 202338 40262
rect 210000 32953 213602 36017
rect 214000 32953 217602 36017
rect 218000 32953 221602 36017
rect 222000 32953 225602 36017
rect 226000 32953 229602 36017
rect 230000 32953 233602 36017
rect 239013 33910 240960 34840
rect 238972 30753 241079 31683
rect 246349 39593 248524 39600
rect 248824 39593 251000 39600
rect 246129 31600 251220 39593
rect 256180 31600 256200 39593
rect 263800 32953 267402 36017
rect 267800 32953 271402 36017
rect 271800 32953 275402 36017
rect 275800 32953 279402 36017
rect 279800 32953 283402 36017
rect 283800 32953 287402 36017
rect 239013 7 240960 4850
rect 241200 7 256200 31600
rect 256379 30760 258395 31690
rect 295086 0 310938 40262
rect 318600 32953 322202 36017
rect 322600 32953 326202 36017
rect 326600 32953 330202 36017
rect 330600 32953 334202 36017
rect 334600 32953 338202 36017
rect 338600 32953 342202 36017
rect 349886 0 365738 40262
rect 373400 32953 377002 36017
rect 377400 32953 381002 36017
rect 381400 32953 385002 36017
rect 385400 32953 389002 36017
rect 389400 32953 393002 36017
rect 393400 32953 397002 36017
rect 404686 0 420538 40262
rect 428200 32953 431802 36017
rect 432200 32953 435802 36017
rect 436200 32953 439802 36017
rect 440200 32953 443802 36017
rect 444200 32953 447802 36017
rect 448200 32953 451802 36017
rect 459486 0 475338 40262
rect 483000 32953 486602 36017
rect 487000 32953 490602 36017
rect 491000 32953 494602 36017
rect 495000 32953 498602 36017
rect 499000 32953 502602 36017
rect 503000 32953 506602 36017
rect 514286 0 530138 40262
rect 537800 32953 541402 36017
rect 541800 32953 545402 36017
rect 545800 32953 549402 36017
rect 549800 32953 553402 36017
rect 553800 32953 557402 36017
rect 557800 32953 561402 36017
rect 574222 39593 576422 40000
rect 576621 39593 578821 40000
rect 574002 34750 579041 39593
rect 628022 39593 630222 40000
rect 630421 39593 632621 40000
rect 627802 36928 632841 39593
rect 569142 0 583952 34750
rect 591600 32953 595202 36017
rect 595600 32953 599202 36017
rect 599600 32953 603202 36017
rect 603600 32953 607202 36017
rect 607600 32953 611202 36017
rect 611600 32953 615202 36017
rect 622869 0 637752 36928
rect 645400 32953 649002 36017
rect 649400 32953 653002 36017
rect 653400 32953 657002 36017
rect 657400 32953 661002 36017
rect 661400 32953 665002 36017
rect 665400 32953 669002 36017
<< metal4 >>
rect 333400 1032757 333654 1037600
rect 348146 1032757 348400 1037600
rect 533618 1008881 575854 1008947
rect 590346 1008881 626522 1008947
rect 575600 1007929 575854 1008165
rect 590346 1007929 590600 1008165
rect 533618 1007147 575854 1007213
rect 590346 1007147 626522 1007213
rect 539946 1004947 575854 1005637
rect 590346 1004947 626254 1005637
rect 297746 1002767 333654 1003697
rect 348146 1002767 384054 1003697
rect 28653 842346 28719 954722
rect 28653 793818 28719 827854
rect 29435 842346 29671 842600
rect 29435 827600 29671 827854
rect 30387 842346 30453 954722
rect 37293 926746 38223 954454
rect 679377 922346 680307 951854
rect 37293 884546 38223 912254
rect 679377 878146 680307 907854
rect 31963 842346 32653 870054
rect 680587 833207 681277 862606
rect 30387 793818 30453 827854
rect 31963 800146 32653 827854
rect 680587 789007 681277 818593
rect 36323 497807 37013 525393
rect 30753 455546 31683 483254
rect 36323 455607 37013 483193
rect 685917 474546 686847 504054
rect 30753 413346 31683 441054
rect 685917 430346 686847 460054
rect 21000 124946 25993 125400
rect 21000 109800 25993 110454
rect 35113 124946 36043 181854
rect 35113 82746 36043 110454
rect 37293 82746 38223 110454
rect 37293 40546 38223 68254
rect 583807 36323 622993 37013
rect 637607 36323 677051 37013
rect 39733 31963 79054 32653
rect 93546 31963 132854 32653
rect 202146 30753 241454 31683
rect 255946 30753 295254 31683
rect 36085 30387 79054 30453
rect 93546 30387 192982 30453
rect 78800 29435 79054 29671
rect 93546 29435 93800 29671
rect 35365 28653 79054 28719
rect 93546 28653 192982 28719
<< obsm4 >>
rect 0 1032677 40466 1037600
rect 40546 1032757 76454 1037600
rect 0 1016680 40549 1032677
rect 40800 1032407 76200 1032757
rect 76534 1032677 91866 1037600
rect 91946 1032757 127854 1037600
rect 0 1011527 40349 1016680
rect 40800 1016600 76200 1017007
rect 76393 1016680 91994 1032677
rect 92200 1032407 127600 1032757
rect 127934 1032677 143266 1037600
rect 143346 1032757 179254 1037600
rect 40429 1011607 76454 1016600
rect 0 1011387 40549 1011527
rect 40800 1011387 76200 1011607
rect 76534 1011527 91866 1016680
rect 92200 1016600 127600 1017007
rect 127793 1016680 143394 1032677
rect 143600 1032407 179000 1032757
rect 179334 1032677 194666 1037600
rect 194746 1032757 230654 1037600
rect 91946 1011607 127854 1016600
rect 76393 1011387 91994 1011527
rect 92200 1011387 127600 1011607
rect 127934 1011527 143266 1016680
rect 143600 1016600 179000 1017007
rect 179193 1016680 194794 1032677
rect 195000 1032407 230400 1032757
rect 230734 1032677 246066 1037600
rect 246146 1032757 282254 1037600
rect 143346 1011607 179254 1016600
rect 127793 1011387 143394 1011527
rect 143600 1011387 179000 1011607
rect 179334 1011527 194666 1016680
rect 195000 1016600 230400 1017007
rect 230593 1016680 246194 1032677
rect 246400 1032407 282000 1032757
rect 282334 1032677 297666 1037600
rect 297746 1032757 333400 1037600
rect 194746 1011607 230654 1016600
rect 179193 1011387 194794 1011527
rect 195000 1011387 230400 1011607
rect 230734 1011527 246066 1016680
rect 246400 1016600 282000 1017007
rect 282193 1016680 297794 1032677
rect 298000 1032407 333400 1032757
rect 333734 1032677 348066 1037600
rect 348400 1032757 384054 1037600
rect 246146 1011607 282254 1016600
rect 230593 1011387 246194 1011527
rect 246400 1011387 282000 1011607
rect 282334 1011527 297666 1016680
rect 298000 1016600 333400 1017007
rect 333593 1016680 348207 1032677
rect 348400 1032407 383800 1032757
rect 384134 1032677 399466 1037600
rect 399546 1032757 473054 1037600
rect 297746 1011607 333654 1016600
rect 282193 1011387 297794 1011527
rect 298000 1011387 333400 1011607
rect 333734 1011527 348066 1016680
rect 348400 1016600 383800 1017007
rect 383993 1016680 399594 1032677
rect 399800 1032407 435200 1032757
rect 437200 1032407 472800 1032757
rect 473134 1032677 488466 1037600
rect 488546 1032757 524454 1037600
rect 348146 1011607 384054 1016600
rect 333593 1011387 348207 1011527
rect 348400 1011387 383800 1011607
rect 384134 1011527 399466 1016680
rect 399800 1016600 435200 1017007
rect 437200 1016600 472800 1017007
rect 472993 1016680 488594 1032677
rect 488800 1032407 524200 1032757
rect 524534 1032677 539866 1037600
rect 539946 1032757 575854 1037600
rect 399546 1011607 473054 1016600
rect 383993 1011387 399594 1011527
rect 399800 1011387 435200 1011607
rect 437200 1011387 472800 1011607
rect 473134 1011527 488466 1016680
rect 488800 1016600 524200 1017007
rect 524393 1016680 539994 1032677
rect 540200 1032407 575600 1032757
rect 575934 1032677 590266 1037600
rect 590346 1032757 626254 1037600
rect 488546 1011607 524454 1016600
rect 472993 1011387 488594 1011527
rect 488800 1011387 524200 1011607
rect 524534 1011527 539866 1016680
rect 540200 1016600 575600 1017007
rect 575793 1016680 590407 1032677
rect 590600 1032407 626000 1032757
rect 626334 1032677 641666 1037600
rect 641746 1032757 677887 1037600
rect 642000 1032677 677600 1032757
rect 677967 1032677 717600 1037600
rect 539946 1011607 575854 1016600
rect 524393 1011387 539994 1011527
rect 540200 1011387 575600 1011607
rect 575934 1011527 590266 1016680
rect 590600 1016600 626000 1017007
rect 626193 1016680 641794 1032677
rect 642000 1032407 717600 1032677
rect 677600 1017007 717600 1032407
rect 642000 1016680 717600 1017007
rect 590346 1011607 626254 1016600
rect 575793 1011387 590407 1011527
rect 590600 1011387 626000 1011607
rect 626334 1011527 641666 1016680
rect 642000 1016600 677600 1016680
rect 641746 1011607 678129 1016600
rect 642000 1011527 677600 1011607
rect 678209 1011527 717600 1016680
rect 626193 1011387 641794 1011527
rect 642000 1011387 717600 1011527
rect 0 1010337 40466 1011387
rect 40546 1010417 76454 1011307
rect 76534 1010337 91866 1011387
rect 91946 1010417 127854 1011307
rect 127934 1010337 143266 1011387
rect 143346 1010417 179254 1011307
rect 179334 1010337 194666 1011387
rect 194746 1010417 230654 1011307
rect 230734 1010337 246066 1011387
rect 246146 1010417 282254 1011307
rect 282334 1010337 297666 1011387
rect 297746 1010417 333654 1011307
rect 333734 1010337 348066 1011387
rect 348146 1010417 384054 1011307
rect 384134 1010337 399466 1011387
rect 399546 1010417 473054 1011307
rect 473134 1010337 488466 1011387
rect 488546 1010417 524454 1011307
rect 524534 1010337 539866 1011387
rect 539946 1010417 575854 1011307
rect 575934 1010337 590266 1011387
rect 590346 1010417 626254 1011307
rect 626334 1010337 641666 1011387
rect 641746 1010417 677896 1011307
rect 677976 1010337 717600 1011387
rect 0 1010217 40549 1010337
rect 40800 1010217 75800 1010337
rect 76393 1010217 91994 1010337
rect 92200 1010217 127200 1010337
rect 127793 1010217 143394 1010337
rect 143600 1010217 178600 1010337
rect 179193 1010217 194794 1010337
rect 195000 1010217 230000 1010337
rect 230593 1010217 246194 1010337
rect 246400 1010217 281400 1010337
rect 282193 1010217 297794 1010337
rect 298000 1010217 333000 1010337
rect 333593 1010217 348207 1010337
rect 348400 1010217 383400 1010337
rect 383993 1010217 399594 1010337
rect 399800 1010217 434800 1010337
rect 437200 1010217 472200 1010337
rect 472993 1010217 488594 1010337
rect 488800 1010217 523800 1010337
rect 524393 1010217 539994 1010337
rect 540200 1010217 575200 1010337
rect 575793 1010217 590407 1010337
rect 590600 1010217 625600 1010337
rect 626193 1010217 641794 1010337
rect 642000 1010217 677000 1010337
rect 677600 1010217 717600 1010337
rect 0 1009167 40466 1010217
rect 40546 1009247 76454 1010137
rect 76534 1009167 91866 1010217
rect 91946 1009247 127854 1010137
rect 127934 1009167 143266 1010217
rect 143346 1009247 179254 1010137
rect 179334 1009167 194666 1010217
rect 194746 1009247 230654 1010137
rect 230734 1009167 246066 1010217
rect 246146 1009247 282254 1010137
rect 282334 1009167 297666 1010217
rect 297746 1009247 333654 1010137
rect 333734 1009167 348066 1010217
rect 348146 1009247 384054 1010137
rect 384134 1009167 399466 1010217
rect 399546 1009247 473054 1010137
rect 473134 1009167 488466 1010217
rect 488546 1009247 524454 1010137
rect 524534 1009167 539866 1010217
rect 539946 1009247 575854 1010137
rect 575934 1009167 590266 1010217
rect 590346 1009247 626254 1010137
rect 626334 1009167 641666 1010217
rect 641746 1009247 677925 1010137
rect 678005 1009167 717600 1010217
rect 0 1009027 40549 1009167
rect 40800 1009027 76200 1009167
rect 76393 1009027 91994 1009167
rect 92200 1009027 127600 1009167
rect 127793 1009027 143394 1009167
rect 143600 1009027 179000 1009167
rect 179193 1009027 194794 1009167
rect 195000 1009027 230400 1009167
rect 230593 1009027 246194 1009167
rect 246400 1009027 282000 1009167
rect 282193 1009027 297794 1009167
rect 298000 1009027 333400 1009167
rect 333593 1009027 348207 1009167
rect 348400 1009027 383800 1009167
rect 383993 1009027 399594 1009167
rect 399800 1009027 435200 1009167
rect 437200 1009027 472800 1009167
rect 472993 1009027 488594 1009167
rect 488800 1009027 524200 1009167
rect 524393 1009027 539994 1009167
rect 540200 1009027 575600 1009167
rect 575793 1009027 590407 1009167
rect 590600 1009027 626000 1009167
rect 626193 1009027 641794 1009167
rect 642000 1009027 717600 1009167
rect 0 1008801 35285 1009027
rect 35365 1008881 76722 1008947
rect 76802 1008901 85538 1009027
rect 0 1008145 35338 1008801
rect 35418 1008225 83488 1008821
rect 36489 1008145 40800 1008165
rect 76200 1008145 76454 1008165
rect 83568 1008145 83872 1008901
rect 85618 1008881 128122 1008947
rect 128202 1008901 136938 1009027
rect 83952 1008225 134888 1008821
rect 91946 1008145 92200 1008165
rect 127600 1008145 127854 1008165
rect 134968 1008145 135272 1008901
rect 137018 1008881 179522 1008947
rect 179602 1008901 188338 1009027
rect 135352 1008225 186288 1008821
rect 143346 1008145 143600 1008165
rect 179000 1008145 179254 1008165
rect 186368 1008145 186672 1008901
rect 188418 1008881 230922 1008947
rect 231002 1008901 239738 1009027
rect 186752 1008225 237688 1008821
rect 194746 1008145 195000 1008165
rect 230400 1008145 230654 1008165
rect 237768 1008145 238072 1008901
rect 239818 1008881 282522 1008947
rect 282602 1008901 291338 1009027
rect 238152 1008225 289288 1008821
rect 246146 1008145 246400 1008165
rect 282000 1008145 282254 1008165
rect 289368 1008145 289672 1008901
rect 291418 1008881 384322 1008947
rect 384402 1008901 393138 1009027
rect 289752 1008225 391088 1008821
rect 297746 1008145 298000 1008165
rect 333400 1008145 333654 1008165
rect 348146 1008145 348400 1008165
rect 383800 1008145 384054 1008165
rect 391168 1008145 391472 1008901
rect 393218 1008881 435200 1008947
rect 436200 1008881 473322 1008947
rect 473402 1008901 482138 1009027
rect 391552 1008225 480088 1008821
rect 399546 1008145 399800 1008165
rect 436200 1008145 437200 1008165
rect 472800 1008145 473054 1008165
rect 480168 1008145 480472 1008901
rect 482218 1008881 524722 1008947
rect 524802 1008901 533538 1009027
rect 480552 1008225 531488 1008821
rect 488546 1008145 488800 1008165
rect 524200 1008145 524454 1008165
rect 531568 1008145 531872 1008901
rect 575934 1008901 590266 1009027
rect 626602 1008901 635338 1009027
rect 531952 1008225 633288 1008821
rect 539946 1008145 540200 1008165
rect 0 1007849 36409 1008145
rect 36489 1007949 76454 1008145
rect 76534 1007949 91866 1008145
rect 91946 1007949 127854 1008145
rect 127934 1007949 143266 1008145
rect 143346 1007949 179254 1008145
rect 179334 1007949 194666 1008145
rect 194746 1007949 230654 1008145
rect 230734 1007949 246066 1008145
rect 246146 1007949 282254 1008145
rect 282334 1007949 297666 1008145
rect 297746 1007949 333654 1008145
rect 333734 1007949 348066 1008145
rect 348146 1007949 384054 1008145
rect 384134 1007949 399466 1008145
rect 399546 1007949 435200 1008145
rect 436200 1007949 473054 1008145
rect 473134 1007949 488466 1008145
rect 488546 1007949 524454 1008145
rect 524534 1007949 539866 1008145
rect 539946 1007949 575600 1008145
rect 36489 1007929 40800 1007949
rect 76200 1007929 76454 1007949
rect 0 1007293 36545 1007849
rect 0 1007067 36005 1007293
rect 36625 1007273 86629 1007869
rect 86709 1007293 87013 1007949
rect 91946 1007929 92200 1007949
rect 127600 1007929 127854 1007949
rect 87093 1007273 138029 1007869
rect 138109 1007293 138413 1007949
rect 143346 1007929 143600 1007949
rect 179000 1007929 179254 1007949
rect 138493 1007273 189429 1007869
rect 189509 1007293 189813 1007949
rect 194746 1007929 195000 1007949
rect 230400 1007929 230654 1007949
rect 189893 1007273 240829 1007869
rect 240909 1007293 241213 1007949
rect 246146 1007929 246400 1007949
rect 282000 1007929 282254 1007949
rect 241293 1007273 292429 1007869
rect 292509 1007293 292813 1007949
rect 297746 1007929 298000 1007949
rect 333400 1007929 333654 1007949
rect 348146 1007929 348400 1007949
rect 383800 1007929 384054 1007949
rect 292893 1007273 394229 1007869
rect 394309 1007293 394613 1007949
rect 399546 1007929 399800 1007949
rect 436200 1007929 437200 1007949
rect 472800 1007929 473054 1007949
rect 394693 1007273 483229 1007869
rect 483309 1007293 483613 1007949
rect 488546 1007929 488800 1007949
rect 524200 1007929 524454 1007949
rect 483693 1007273 534629 1007869
rect 534709 1007293 535013 1007949
rect 539946 1007929 540200 1007949
rect 575934 1007949 590266 1008145
rect 626000 1008145 626254 1008165
rect 633368 1008145 633672 1008901
rect 635418 1008881 682235 1008947
rect 633752 1008225 682182 1008821
rect 682315 1008801 717600 1009027
rect 641746 1008145 642000 1008165
rect 677600 1008145 681910 1008165
rect 682262 1008145 717600 1008801
rect 590600 1007949 626254 1008145
rect 626334 1007949 641666 1008145
rect 641746 1007949 681910 1008145
rect 626000 1007929 626254 1007949
rect 535093 1007273 636429 1007869
rect 636509 1007293 636813 1007949
rect 641746 1007929 642000 1007949
rect 677600 1007929 681910 1007949
rect 636893 1007273 681787 1007869
rect 681990 1007849 717600 1008145
rect 36085 1007147 76722 1007213
rect 76802 1007067 85538 1007193
rect 85618 1007147 128122 1007213
rect 128202 1007067 136938 1007193
rect 137018 1007147 179522 1007213
rect 179602 1007067 188338 1007193
rect 188418 1007147 230922 1007213
rect 231002 1007067 239738 1007193
rect 239818 1007147 282522 1007213
rect 282602 1007067 291338 1007193
rect 291418 1007147 384322 1007213
rect 384402 1007067 393138 1007193
rect 393218 1007147 435200 1007213
rect 436200 1007147 473322 1007213
rect 473402 1007067 482138 1007193
rect 482218 1007147 524722 1007213
rect 524802 1007067 533538 1007193
rect 575934 1007067 590266 1007193
rect 626602 1007067 635338 1007193
rect 635418 1007147 681515 1007213
rect 681867 1007193 717600 1007849
rect 681595 1007067 717600 1007193
rect 0 1006927 40549 1007067
rect 76393 1006927 91994 1007067
rect 127793 1006927 143394 1007067
rect 179193 1006927 194794 1007067
rect 230593 1006927 246194 1007067
rect 282193 1006927 297794 1007067
rect 333593 1006927 348207 1007067
rect 383993 1006927 399594 1007067
rect 472993 1006927 488594 1007067
rect 524393 1006927 539994 1007067
rect 575793 1006927 590407 1007067
rect 626193 1006927 641794 1007067
rect 677600 1006927 717600 1007067
rect 0 1005837 40466 1006927
rect 40546 1005917 76454 1006847
rect 76534 1005837 91866 1006927
rect 91946 1005917 127854 1006847
rect 127934 1005837 143266 1006927
rect 143346 1005917 179254 1006847
rect 179334 1005837 194666 1006927
rect 194746 1005917 230654 1006847
rect 230734 1005837 246066 1006927
rect 246146 1005917 282254 1006847
rect 282334 1005837 297666 1006927
rect 297746 1005917 333654 1006847
rect 333734 1005837 348066 1006927
rect 348146 1005917 384054 1006847
rect 384134 1005837 399466 1006927
rect 399546 1005917 436200 1006847
rect 437200 1005917 473054 1006847
rect 473134 1005837 488466 1006927
rect 488546 1005917 524454 1006847
rect 524534 1005837 539866 1006927
rect 539946 1005917 575854 1006847
rect 575934 1005837 590266 1006927
rect 590346 1005917 626254 1006847
rect 626334 1005837 641666 1006927
rect 641746 1005917 677895 1006847
rect 677975 1005837 717600 1006927
rect 0 1005717 40549 1005837
rect 76393 1005717 91994 1005837
rect 127793 1005717 143394 1005837
rect 179193 1005717 194794 1005837
rect 230593 1005717 246194 1005837
rect 282193 1005717 297794 1005837
rect 333593 1005717 348207 1005837
rect 383993 1005717 399594 1005837
rect 472993 1005717 488594 1005837
rect 524393 1005717 539994 1005837
rect 575793 1005717 590407 1005837
rect 626193 1005717 641794 1005837
rect 677600 1005717 717600 1005837
rect 0 1004867 40466 1005717
rect 40546 1004947 76454 1005637
rect 76534 1004867 91866 1005717
rect 91946 1004947 127854 1005637
rect 127934 1004867 143266 1005717
rect 143346 1004947 179254 1005637
rect 179334 1004867 194666 1005717
rect 194746 1004947 230654 1005637
rect 230734 1004867 246066 1005717
rect 246146 1004947 282254 1005637
rect 282334 1004867 297666 1005717
rect 297746 1004947 333654 1005637
rect 333734 1004867 348066 1005717
rect 348146 1004947 384054 1005637
rect 384134 1004867 399466 1005717
rect 399546 1004947 435200 1005637
rect 436200 1004947 473054 1005637
rect 473134 1004867 488466 1005717
rect 488546 1004947 524454 1005637
rect 524534 1004867 539866 1005717
rect 575934 1004867 590266 1005717
rect 626334 1004867 641666 1005717
rect 641746 1004947 677867 1005637
rect 677947 1004867 717600 1005717
rect 0 1004747 40549 1004867
rect 76393 1004747 91994 1004867
rect 127793 1004747 143394 1004867
rect 179193 1004747 194794 1004867
rect 230593 1004747 246194 1004867
rect 282193 1004747 297794 1004867
rect 333593 1004747 348207 1004867
rect 383993 1004747 399594 1004867
rect 472993 1004747 488594 1004867
rect 524393 1004747 539994 1004867
rect 575793 1004747 590407 1004867
rect 626193 1004747 641794 1004867
rect 677600 1004747 717600 1004867
rect 0 1003897 40466 1004747
rect 40546 1003977 76454 1004667
rect 76534 1003897 91866 1004747
rect 91946 1003977 127854 1004667
rect 127934 1003897 143266 1004747
rect 143346 1003977 179254 1004667
rect 179334 1003897 194666 1004747
rect 194746 1003977 230654 1004667
rect 230734 1003897 246066 1004747
rect 246146 1003977 282254 1004667
rect 282334 1003897 297666 1004747
rect 297746 1003977 333654 1004667
rect 333734 1003897 348066 1004747
rect 348146 1003977 384054 1004667
rect 384134 1003897 399466 1004747
rect 399546 1003977 473054 1004667
rect 473134 1003897 488466 1004747
rect 488546 1003977 524454 1004667
rect 524534 1003897 539866 1004747
rect 539946 1003977 575854 1004667
rect 575934 1003897 590266 1004747
rect 590346 1003977 626254 1004667
rect 626334 1003897 641666 1004747
rect 641746 1003977 677877 1004667
rect 677957 1003897 717600 1004747
rect 0 1003777 40549 1003897
rect 76393 1003777 91994 1003897
rect 127793 1003777 143394 1003897
rect 179193 1003777 194794 1003897
rect 230593 1003777 246194 1003897
rect 282193 1003777 297794 1003897
rect 333593 1003777 348207 1003897
rect 383993 1003777 399594 1003897
rect 472993 1003777 488594 1003897
rect 524393 1003777 539994 1003897
rect 575793 1003777 590407 1003897
rect 626193 1003777 641794 1003897
rect 677600 1003777 717600 1003897
rect 0 1002687 40466 1003777
rect 40546 1002767 76454 1003697
rect 76534 1002687 91866 1003777
rect 91946 1002767 127854 1003697
rect 127934 1002687 143266 1003777
rect 143346 1002767 179254 1003697
rect 179334 1002687 194666 1003777
rect 194746 1002767 230654 1003697
rect 230734 1002687 246066 1003777
rect 246146 1002767 282254 1003697
rect 282334 1002687 297666 1003777
rect 333734 1002687 348066 1003777
rect 384134 1002687 399466 1003777
rect 399546 1002767 473054 1003697
rect 473134 1002687 488466 1003777
rect 488546 1002767 524454 1003697
rect 524534 1002687 539866 1003777
rect 539946 1002767 575854 1003697
rect 575934 1002687 590266 1003777
rect 590346 1002767 626254 1003697
rect 626334 1002687 641666 1003777
rect 641746 1002767 677920 1003697
rect 678000 1002687 717600 1003777
rect 0 1002567 40549 1002687
rect 76393 1002567 91994 1002687
rect 127793 1002567 143394 1002687
rect 179193 1002567 194794 1002687
rect 230593 1002567 246194 1002687
rect 282193 1002567 297794 1002687
rect 333593 1002567 348207 1002687
rect 383993 1002567 399594 1002687
rect 472993 1002567 488594 1002687
rect 524393 1002567 539994 1002687
rect 575793 1002567 590407 1002687
rect 626193 1002567 641794 1002687
rect 677600 1002567 717600 1002687
rect 0 1002315 40466 1002567
rect 0 998209 28573 1002315
rect 28799 1002262 40466 1002315
rect 0 997967 20920 998209
rect 0 997600 4843 997887
rect 4923 997600 20920 997967
rect 21000 997600 25993 998129
rect 26073 998005 28573 998209
rect 26073 997976 27383 998005
rect 26073 997600 26213 997976
rect 0 970200 5193 997600
rect 20593 970200 26213 997600
rect 0 969946 4843 970200
rect 4923 969866 20920 969994
rect 21000 969946 25993 970200
rect 26073 969866 26213 969994
rect 26293 969946 27183 997896
rect 27263 997600 27383 997976
rect 27263 970200 27383 997200
rect 27263 969866 27383 969994
rect 27463 969946 28353 997925
rect 28433 970200 28573 998005
rect 28433 969866 28573 969994
rect 0 963538 28573 969866
rect 28653 963618 28719 1002235
rect 0 961872 28699 963538
rect 28779 961952 29375 1002182
rect 29455 1001990 40466 1002262
rect 29435 997600 29671 1001910
rect 29751 1001867 40466 1001990
rect 29455 970200 29651 997600
rect 29435 969946 29671 970200
rect 29455 965013 29651 969866
rect 29731 965093 30327 1001787
rect 30407 1001595 40466 1001867
rect 29455 964709 30307 965013
rect 29455 961872 29651 964709
rect 0 961568 29651 961872
rect 0 954802 28699 961568
rect 0 954534 28573 954802
rect 0 954200 4843 954454
rect 4923 954393 20920 954534
rect 21000 954200 25993 954454
rect 26073 954393 26213 954534
rect 0 927000 5193 954200
rect 20593 927000 26213 954200
rect 0 926746 4843 927000
rect 4923 926666 20920 927000
rect 21000 926746 25993 927000
rect 26073 926666 26213 927000
rect 26293 926746 27183 954454
rect 27263 954393 27383 954534
rect 27263 926666 27383 954000
rect 27463 926746 28353 954454
rect 28433 954393 28573 954534
rect 28433 926666 28573 954200
rect 0 912334 28573 926666
rect 0 912000 4843 912254
rect 4923 912193 20920 912334
rect 21000 912000 25993 912254
rect 26073 912193 26213 912334
rect 0 884800 5193 912000
rect 20593 884800 26213 912000
rect 0 884546 4843 884800
rect 4923 884466 20920 884607
rect 21000 884546 25993 884800
rect 26073 884466 26213 884607
rect 26293 884546 27183 912254
rect 27263 912193 27383 912334
rect 27263 884800 27383 911800
rect 27263 884466 27383 884607
rect 27463 884546 28353 912254
rect 28433 912193 28573 912334
rect 28433 884800 28573 912000
rect 28433 884466 28573 884607
rect 0 870134 28573 884466
rect 0 869800 4843 870054
rect 4923 869993 20920 870134
rect 21000 869800 25993 870054
rect 26073 869993 26213 870134
rect 0 842600 5193 869800
rect 20593 842600 26213 869800
rect 0 842346 4843 842600
rect 4923 842266 20920 842407
rect 21000 842346 25993 842600
rect 26073 842266 26213 842407
rect 26293 842346 27183 870054
rect 27263 869993 27383 870134
rect 27263 842600 27383 869600
rect 27263 842266 27383 842407
rect 27463 842346 28353 870054
rect 28433 869993 28573 870134
rect 28433 842600 28573 869800
rect 28433 842266 28573 842407
rect 0 827934 28699 842266
rect 0 827600 4843 827854
rect 4923 827793 20920 827934
rect 21000 827600 25993 827854
rect 26073 827793 26213 827934
rect 0 800400 5193 827600
rect 20593 800400 26213 827600
rect 0 800146 4843 800400
rect 4923 800066 20920 800194
rect 21000 800146 25993 800400
rect 26073 800066 26213 800194
rect 26293 800146 27183 827854
rect 27263 827793 27383 827934
rect 27263 800400 27383 827400
rect 27263 800066 27383 800194
rect 27463 800146 28353 827854
rect 28433 827793 28573 827934
rect 28433 800400 28573 827600
rect 28433 800066 28573 800194
rect 0 793738 28573 800066
rect 0 792072 28699 793738
rect 28779 792152 29375 961488
rect 29455 954534 29651 961568
rect 29435 954200 29671 954454
rect 29455 927000 29651 954200
rect 29435 926746 29671 927000
rect 29455 912334 29651 926666
rect 29435 912000 29671 912254
rect 29455 884800 29651 912000
rect 29435 884546 29671 884800
rect 29455 870134 29651 884466
rect 29435 869800 29671 870054
rect 29455 842600 29651 869800
rect 29455 827934 29651 842266
rect 29455 800400 29651 827600
rect 29435 800146 29671 800400
rect 29455 795213 29651 800066
rect 29731 795293 30327 964629
rect 30387 963618 30453 1001515
rect 30533 1001477 40466 1001595
rect 40546 1001557 76454 1002487
rect 76534 1001477 91866 1002567
rect 91946 1001557 127854 1002487
rect 127934 1001477 143266 1002567
rect 143346 1001557 179254 1002487
rect 179334 1001477 194666 1002567
rect 194746 1001557 230654 1002487
rect 230734 1001477 246066 1002567
rect 246146 1001557 282254 1002487
rect 282334 1001477 297666 1002567
rect 297746 1001557 333654 1002487
rect 333734 1001477 348066 1002567
rect 348146 1001557 384054 1002487
rect 384134 1001477 399466 1002567
rect 399546 1001557 473054 1002487
rect 473134 1001477 488466 1002567
rect 488546 1001557 524454 1002487
rect 524534 1001477 539866 1002567
rect 539946 1001557 575854 1002487
rect 575934 1001477 590266 1002567
rect 590346 1001557 626254 1002487
rect 626334 1001477 641666 1002567
rect 641746 1001557 677905 1002487
rect 677985 1002315 717600 1002567
rect 677985 1002262 688801 1002315
rect 677985 1001595 688145 1002262
rect 677985 1001477 687067 1001595
rect 30533 1001357 40549 1001477
rect 76393 1001357 91994 1001477
rect 127793 1001357 143394 1001477
rect 179193 1001357 194794 1001477
rect 230593 1001357 246194 1001477
rect 282193 1001357 297794 1001477
rect 333593 1001357 348207 1001477
rect 383993 1001357 399594 1001477
rect 472993 1001357 488594 1001477
rect 524393 1001357 539994 1001477
rect 575793 1001357 590407 1001477
rect 626193 1001357 641794 1001477
rect 677600 1001357 687067 1001477
rect 30533 1000507 40469 1001357
rect 40549 1000587 76393 1001277
rect 76473 1000507 91914 1001357
rect 91994 1000587 127793 1001277
rect 127873 1000507 143314 1001357
rect 143394 1000587 179193 1001277
rect 179273 1000507 194714 1001357
rect 194794 1000587 230593 1001277
rect 230673 1000507 246114 1001357
rect 246194 1000587 282193 1001277
rect 282273 1000507 297714 1001357
rect 297794 1000587 333593 1001277
rect 333673 1000507 348127 1001357
rect 348207 1000587 383993 1001277
rect 384073 1000507 399514 1001357
rect 399594 1000587 435200 1001277
rect 436200 1000587 472993 1001277
rect 473073 1000507 488514 1001357
rect 488594 1000587 524393 1001277
rect 524473 1000507 539914 1001357
rect 539994 1000587 575793 1001277
rect 575873 1000507 590327 1001357
rect 590407 1000587 626193 1001277
rect 626273 1000507 641714 1001357
rect 641794 1000587 677894 1001277
rect 677974 1000507 687067 1001357
rect 30533 1000387 40549 1000507
rect 76393 1000387 91994 1000507
rect 127793 1000387 143394 1000507
rect 179193 1000387 194794 1000507
rect 230593 1000387 246194 1000507
rect 282193 1000387 297794 1000507
rect 333593 1000387 348207 1000507
rect 383993 1000387 399594 1000507
rect 472993 1000387 488594 1000507
rect 524393 1000387 539994 1000507
rect 575793 1000387 590407 1000507
rect 626193 1000387 641794 1000507
rect 677600 1000387 687067 1000507
rect 30533 999297 40466 1000387
rect 40546 999377 76454 1000307
rect 76534 999297 91866 1000387
rect 91946 999377 127854 1000307
rect 127934 999297 143266 1000387
rect 143346 999377 179254 1000307
rect 179334 999297 194666 1000387
rect 194746 999377 230654 1000307
rect 230734 999297 246066 1000387
rect 246146 999377 282254 1000307
rect 282334 999297 297666 1000387
rect 297746 999377 333654 1000307
rect 333734 999297 348066 1000387
rect 348146 999377 384054 1000307
rect 384134 999297 399466 1000387
rect 399546 999377 436200 1000307
rect 437200 999377 473054 1000307
rect 473134 999297 488466 1000387
rect 488546 999377 524454 1000307
rect 524534 999297 539866 1000387
rect 539946 999377 575854 1000307
rect 575934 999297 590266 1000387
rect 590346 999377 626254 1000307
rect 626334 999297 641666 1000387
rect 641746 999377 678357 1000307
rect 678437 999297 687067 1000387
rect 30533 999177 40549 999297
rect 76393 999177 91994 999297
rect 127793 999177 143394 999297
rect 179193 999177 194794 999297
rect 230593 999177 246194 999297
rect 282193 999177 297794 999297
rect 333593 999177 348207 999297
rect 383993 999177 399594 999297
rect 472993 999177 488594 999297
rect 524393 999177 539994 999297
rect 575793 999177 590407 999297
rect 626193 999177 641794 999297
rect 677600 999177 687067 999297
rect 30533 998437 40466 999177
rect 30533 998000 37213 998437
rect 30533 997975 33823 998000
rect 30533 997600 30673 997975
rect 31763 997957 33823 997975
rect 31763 997947 32853 997957
rect 30533 969866 30673 969994
rect 30753 969946 31683 997895
rect 31763 997600 31883 997947
rect 31763 969866 31883 969994
rect 31963 969946 32653 997867
rect 32733 997600 32853 997947
rect 32733 969866 32853 969994
rect 32933 969946 33623 997877
rect 33703 997600 33823 997957
rect 34913 997985 37213 998000
rect 33703 969866 33823 969994
rect 33903 969946 34833 997920
rect 34913 997600 35033 997985
rect 36123 997974 37213 997985
rect 34913 969866 35033 969994
rect 35113 969946 36043 997905
rect 36123 997600 36243 997974
rect 36323 969994 37013 997894
rect 37093 997600 37213 997974
rect 36123 969914 36243 969994
rect 37093 969914 37213 969994
rect 37293 969946 38223 998357
rect 38303 998150 40466 998437
rect 38303 997600 38423 998150
rect 38503 998007 39593 998070
rect 39673 998007 40466 998150
rect 40546 998007 76454 999097
rect 38503 997927 40466 998007
rect 76534 997927 91866 999177
rect 91946 998007 127854 999097
rect 127934 997927 143266 999177
rect 143346 998007 179254 999097
rect 179334 997927 194666 999177
rect 194746 998007 230654 999097
rect 230734 997927 246066 999177
rect 246146 998007 282254 999097
rect 282334 997927 297666 999177
rect 297746 998007 333654 999097
rect 333734 998007 348066 999177
rect 348146 998007 384054 999097
rect 384134 997927 399466 999177
rect 399546 998007 473054 999097
rect 473134 997927 488466 999177
rect 488546 998007 524454 999097
rect 524534 997927 539866 999177
rect 539946 998007 575854 999097
rect 575934 998007 590266 999177
rect 590346 998007 626254 999097
rect 626334 997927 641666 999177
rect 641746 998007 678070 999097
tri 677600 997927 677680 998007 ne
rect 677680 997927 678007 998007
rect 678150 997927 687067 999177
rect 38503 997680 40549 997927
rect 76393 997707 91994 997927
rect 127793 997707 143394 997927
rect 179193 997707 194794 997927
rect 230593 997707 246194 997927
rect 282193 997707 297794 997927
rect 383993 997707 399594 997927
rect 472993 997707 488594 997927
rect 524393 997707 539994 997927
rect 626193 997707 641794 997927
rect 36123 969866 37213 969914
rect 38303 969866 38423 969994
rect 38503 969946 39593 997680
tri 39593 997600 39673 997680 nw
rect 39673 997600 40549 997680
rect 677600 997134 687067 997927
rect 677600 997051 677927 997134
rect 39673 969866 39893 969994
rect 30533 963538 39893 969866
rect 30407 954802 39893 963538
rect 30533 954534 39893 954802
rect 30533 954393 30673 954534
rect 30533 926666 30673 927000
rect 30753 926746 31683 954454
rect 31763 954393 31883 954534
rect 31763 926666 31883 927000
rect 31963 926746 32653 954454
rect 32733 954393 32853 954534
rect 32733 926666 32853 927000
rect 32933 926746 33623 954454
rect 33703 954393 33823 954534
rect 33703 926666 33823 927000
rect 33903 926746 34833 954454
rect 34913 954393 35033 954534
rect 36123 954473 37213 954534
rect 34913 926666 35033 927000
rect 35113 926746 36043 954454
rect 36123 954393 36243 954473
rect 37093 954393 37213 954473
rect 36123 926727 36243 927000
rect 36323 926807 37013 954393
rect 37093 926727 37213 927000
rect 38303 954393 38423 954534
rect 36123 926666 37213 926727
rect 38303 926666 38423 927000
rect 38503 926746 39593 954454
rect 39673 954393 39893 954534
rect 677707 967266 677927 967407
rect 678007 967346 679097 997054
rect 679177 997051 679297 997134
rect 680387 997131 681477 997134
rect 679177 967266 679297 967407
rect 679377 967346 680307 997054
rect 680387 997051 680507 997131
rect 681357 997051 681477 997131
rect 680587 967407 681277 997051
rect 680387 967327 680507 967407
rect 681357 967327 681477 967407
rect 681557 967346 682487 997054
rect 682567 997051 682687 997134
rect 680387 967266 681477 967327
rect 682567 967266 682687 967407
rect 682767 967346 683697 997054
rect 683777 997051 683897 997134
rect 683777 967266 683897 967407
rect 683977 967346 684667 997054
rect 684747 997051 684867 997134
rect 684747 967266 684867 967407
rect 684947 967346 685637 997054
rect 685717 997051 685837 997134
rect 685717 967266 685837 967407
rect 685917 967346 686847 997054
rect 686927 997051 687067 997134
rect 686927 967266 687067 967407
rect 677707 966998 687067 967266
rect 687147 967078 687213 1001515
rect 687293 1001191 688145 1001595
rect 687293 1001055 687849 1001191
rect 677707 958262 687193 966998
rect 677707 951934 687067 958262
rect 677707 951806 677927 951934
rect 30533 912334 39593 926666
rect 678007 922346 679097 951854
rect 679177 951806 679297 951934
rect 680387 951886 681477 951934
rect 679177 922266 679297 922407
rect 680387 951806 680507 951886
rect 681357 951806 681477 951886
rect 680587 922407 681277 951806
rect 680387 922327 680507 922407
rect 681357 922327 681477 922407
rect 681557 922346 682487 951854
rect 682567 951806 682687 951934
rect 680387 922266 681477 922327
rect 682567 922266 682687 922407
rect 682767 922346 683697 951854
rect 683777 951806 683897 951934
rect 683777 922266 683897 922407
rect 683977 922346 684667 951854
rect 684747 951806 684867 951934
rect 684747 922266 684867 922407
rect 684947 922346 685637 951854
rect 685717 951806 685837 951934
rect 685717 922266 685837 922407
rect 685917 922346 686847 951854
rect 686927 951806 687067 951934
rect 686927 922266 687067 922407
rect 30533 912193 30673 912334
rect 30533 884466 30673 884607
rect 30753 884546 31683 912254
rect 31763 912193 31883 912334
rect 31763 884466 31883 884607
rect 31963 884546 32653 912254
rect 32733 912193 32853 912334
rect 32733 884466 32853 884607
rect 32933 884546 33623 912254
rect 33703 912193 33823 912334
rect 33703 884466 33823 884607
rect 33903 884546 34833 912254
rect 34913 912193 35033 912334
rect 36123 912273 37213 912334
rect 34913 884466 35033 884607
rect 35113 884546 36043 912254
rect 36123 912193 36243 912273
rect 37093 912193 37213 912273
rect 36323 884607 37013 912193
rect 36123 884527 36243 884607
rect 37093 884527 37213 884607
rect 38303 912193 38423 912334
rect 36123 884466 37213 884527
rect 38303 884466 38423 884607
rect 38503 884546 39593 912254
rect 678007 907934 687067 922266
rect 30533 870134 39593 884466
rect 677707 878066 677927 878207
rect 678007 878146 679097 907854
rect 679177 907600 679297 907934
rect 680387 907873 681477 907934
rect 679177 878066 679297 878207
rect 680387 907600 680507 907873
rect 680587 878207 681277 907793
rect 681357 907600 681477 907873
rect 680387 878127 680507 878207
rect 681357 878127 681477 878207
rect 681557 878146 682487 907854
rect 682567 907600 682687 907934
rect 680387 878066 681477 878127
rect 682567 878066 682687 878207
rect 682767 878146 683697 907854
rect 683777 907600 683897 907934
rect 683777 878066 683897 878207
rect 683977 878146 684667 907854
rect 684747 907600 684867 907934
rect 684747 878066 684867 878207
rect 684947 878146 685637 907854
rect 685717 907600 685837 907934
rect 685717 878066 685837 878207
rect 685917 878146 686847 907854
rect 686927 907600 687067 907934
rect 686927 878066 687067 878207
rect 677707 877798 687067 878066
rect 687147 877878 687213 958182
rect 687273 957171 687869 1000975
rect 687929 996800 688165 1001111
rect 687949 967600 688145 996800
rect 687929 967346 688165 967600
rect 687949 960232 688145 967266
rect 688225 960312 688821 1002182
rect 688881 967078 688947 1002235
rect 689027 997251 717600 1002315
rect 689027 997134 691527 997251
rect 689027 997051 689167 997134
rect 689027 967600 689167 996800
rect 689027 967266 689167 967407
rect 689247 967346 690137 997054
rect 690217 997051 690337 997134
rect 690217 967600 690337 996600
rect 690217 967266 690337 967407
rect 690417 967346 691307 997054
rect 691387 997051 691527 997134
rect 691607 996800 696600 997171
rect 696680 997134 717600 997251
rect 696680 997051 712677 997134
rect 712757 996800 717600 997054
rect 691387 967600 697007 996800
rect 712407 967600 717600 996800
rect 691387 967266 691527 967407
rect 691607 967346 696600 967600
rect 696680 967266 712677 967407
rect 712757 967346 717600 967600
rect 689027 966998 717600 967266
rect 688901 960232 717600 966998
rect 687949 959928 717600 960232
rect 687949 957091 688145 959928
rect 687293 956787 688145 957091
rect 30533 869993 30673 870134
rect 30533 842266 30673 842407
rect 30753 842346 31683 870054
rect 31763 869993 31883 870134
rect 31763 842266 31883 842407
rect 32733 869993 32853 870134
rect 32733 842266 32853 842407
rect 32933 842346 33623 870054
rect 33703 869993 33823 870134
rect 33703 842266 33823 842407
rect 33903 842346 34833 870054
rect 34913 869993 35033 870134
rect 36123 870073 37213 870134
rect 34913 842266 35033 842407
rect 35113 842346 36043 870054
rect 36123 869993 36243 870073
rect 37093 869993 37213 870073
rect 36323 842407 37013 869993
rect 36123 842327 36243 842407
rect 37093 842327 37213 842407
rect 37293 842346 38223 870054
rect 38303 869993 38423 870134
rect 36123 842266 37213 842327
rect 38303 842266 38423 842407
rect 38503 842346 39593 870054
rect 677707 869062 687193 877798
rect 677707 862734 687067 869062
rect 677707 862606 677927 862734
rect 30407 827934 39593 842266
rect 678007 833146 679097 862654
rect 679177 862606 679297 862734
rect 680387 862686 681477 862734
rect 679177 833066 679297 833207
rect 679377 833146 680307 862654
rect 680387 862606 680507 862686
rect 681357 862606 681477 862686
rect 680387 833127 680507 833207
rect 681357 833127 681477 833207
rect 681557 833146 682487 862654
rect 682567 862606 682687 862734
rect 680387 833066 681477 833127
rect 682567 833066 682687 833207
rect 682767 833146 683697 862654
rect 683777 862606 683897 862734
rect 683777 833066 683897 833207
rect 683977 833146 684667 862654
rect 684747 862606 684867 862734
rect 684747 833066 684867 833207
rect 684947 833146 685637 862654
rect 685717 862606 685837 862734
rect 685717 833066 685837 833207
rect 685917 833146 686847 862654
rect 686927 862606 687067 862734
rect 686927 833066 687067 833207
rect 29455 794909 30307 795213
rect 29455 792072 29651 794909
rect 0 791768 29651 792072
rect 0 785002 28699 791768
rect 0 784734 28573 785002
rect 0 784400 4843 784654
rect 4923 784593 20920 784734
rect 21000 784400 25993 784654
rect 26073 784593 26213 784734
rect 0 757200 5193 784400
rect 20593 757200 26213 784400
rect 0 756946 4843 757200
rect 4923 756866 20920 756994
rect 21000 756946 25993 757200
rect 26073 756866 26213 756994
rect 26293 756946 27183 784654
rect 27263 784593 27383 784734
rect 27263 757200 27383 784200
rect 27263 756866 27383 756994
rect 27463 756946 28353 784654
rect 28433 784593 28573 784734
rect 28433 757200 28573 784400
rect 28433 756866 28573 756994
rect 0 750538 28573 756866
rect 28653 750618 28719 784922
rect 0 748872 28699 750538
rect 28779 748952 29375 791688
rect 29455 784734 29651 791768
rect 29435 784400 29671 784654
rect 29455 757200 29651 784400
rect 29435 756946 29671 757200
rect 29455 752013 29651 756866
rect 29731 752093 30327 794829
rect 30533 827793 30673 827934
rect 30533 800066 30673 800194
rect 30753 800146 31683 827854
rect 31763 827793 31883 827934
rect 31763 800066 31883 800194
rect 32733 827793 32853 827934
rect 32733 800066 32853 800194
rect 32933 800146 33623 827854
rect 33703 827793 33823 827934
rect 33703 800066 33823 800194
rect 33903 800146 34833 827854
rect 34913 827793 35033 827934
rect 36123 827873 37213 827934
rect 34913 800066 35033 800194
rect 35113 800146 36043 827854
rect 36123 827793 36243 827873
rect 37093 827793 37213 827873
rect 36323 800194 37013 827793
rect 36123 800114 36243 800194
rect 37093 800114 37213 800194
rect 37293 800146 38223 827854
rect 38303 827793 38423 827934
rect 36123 800066 37213 800114
rect 38303 800066 38423 800194
rect 38503 800146 39593 827854
rect 678007 818734 687067 833066
rect 39673 800066 39893 800194
rect 30533 793738 39893 800066
rect 30407 785002 39893 793738
rect 29455 751709 30307 752013
rect 29455 748872 29651 751709
rect 0 748568 29651 748872
rect 0 741802 28699 748568
rect 0 741534 28573 741802
rect 0 741200 4843 741454
rect 4923 741393 20920 741534
rect 21000 741200 25993 741454
rect 26073 741393 26213 741534
rect 0 714000 5193 741200
rect 20593 714000 26213 741200
rect 0 713746 4843 714000
rect 4923 713666 20920 713794
rect 21000 713746 25993 714000
rect 26073 713666 26213 713794
rect 26293 713746 27183 741454
rect 27263 741393 27383 741534
rect 27263 714000 27383 741000
rect 27263 713666 27383 713794
rect 27463 713746 28353 741454
rect 28433 741393 28573 741534
rect 28433 714000 28573 741200
rect 28433 713666 28573 713794
rect 0 707338 28573 713666
rect 28653 707418 28719 741722
rect 0 705672 28699 707338
rect 28779 705752 29375 748488
rect 29455 741534 29651 748568
rect 29435 741200 29671 741454
rect 29455 714000 29651 741200
rect 29435 713746 29671 714000
rect 29455 708813 29651 713666
rect 29731 708893 30327 751629
rect 30387 750618 30453 784922
rect 30533 784734 39893 785002
rect 30533 784593 30673 784734
rect 30533 756866 30673 756994
rect 30753 756946 31683 784654
rect 31763 784593 31883 784734
rect 31763 756866 31883 756994
rect 31963 756946 32653 784654
rect 32733 784593 32853 784734
rect 32733 756866 32853 756994
rect 32933 756946 33623 784654
rect 33703 784593 33823 784734
rect 33703 756866 33823 756994
rect 33903 756946 34833 784654
rect 34913 784593 35033 784734
rect 36123 784673 37213 784734
rect 34913 756866 35033 756994
rect 35113 756946 36043 784654
rect 36123 784593 36243 784673
rect 37093 784593 37213 784673
rect 36323 756994 37013 784593
rect 36123 756914 36243 756994
rect 37093 756914 37213 756994
rect 37293 756946 38223 784654
rect 38303 784593 38423 784734
rect 36123 756866 37213 756914
rect 38303 756866 38423 756994
rect 38503 756946 39593 784654
rect 39673 784593 39893 784734
rect 677707 788866 677927 789007
rect 678007 788946 679097 818654
rect 679177 818593 679297 818734
rect 680387 818673 681477 818734
rect 679177 788866 679297 789007
rect 679377 788946 680307 818654
rect 680387 818593 680507 818673
rect 681357 818593 681477 818673
rect 680387 788927 680507 789007
rect 681357 788927 681477 789007
rect 681557 788946 682487 818654
rect 682567 818593 682687 818734
rect 680387 788866 681477 788927
rect 682567 788866 682687 789007
rect 682767 788946 683697 818654
rect 683777 818593 683897 818734
rect 683777 788866 683897 789007
rect 683977 788946 684667 818654
rect 684747 818593 684867 818734
rect 684747 788866 684867 789007
rect 684947 788946 685637 818654
rect 685717 818593 685837 818734
rect 685717 788866 685837 789007
rect 685917 788946 686847 818654
rect 686927 818593 687067 818734
rect 686927 788866 687067 789007
rect 677707 788598 687067 788866
rect 687147 788678 687213 868982
rect 687273 867971 687869 956707
rect 687949 951934 688145 956787
rect 687929 951600 688165 951854
rect 687949 922600 688145 951600
rect 687929 922346 688165 922600
rect 687949 907934 688145 922266
rect 687929 907600 688165 907854
rect 687949 878400 688145 907600
rect 687929 878146 688165 878400
rect 687949 871032 688145 878066
rect 688225 871112 688821 959848
rect 688901 958262 717600 959928
rect 688881 877878 688947 958182
rect 689027 951934 717600 958262
rect 689027 951806 689167 951934
rect 689027 922600 689167 951600
rect 689027 922266 689167 922407
rect 689247 922346 690137 951854
rect 690217 951806 690337 951934
rect 690217 922600 690337 951600
rect 690217 922266 690337 922407
rect 690417 922346 691307 951854
rect 691387 951806 691527 951934
rect 691607 951600 696600 951854
rect 696680 951806 712677 951934
rect 712757 951600 717600 951854
rect 691387 922600 697007 951600
rect 712407 922600 717600 951600
rect 691387 922266 691527 922407
rect 691607 922346 696600 922600
rect 696680 922266 712677 922407
rect 712757 922346 717600 922600
rect 689027 907934 717600 922266
rect 689027 878400 689167 907934
rect 689027 878066 689167 878207
rect 689247 878146 690137 907854
rect 690217 907600 690337 907934
rect 690217 878400 690337 907400
rect 690217 878066 690337 878207
rect 690417 878146 691307 907854
rect 691387 907600 691527 907934
rect 691607 907600 696600 907854
rect 696680 907600 712677 907934
rect 712757 907600 717600 907854
rect 691387 878400 697007 907600
rect 712407 878400 717600 907600
rect 691387 878066 691527 878207
rect 691607 878146 696600 878400
rect 696680 878066 712677 878207
rect 712757 878146 717600 878400
rect 689027 877798 717600 878066
rect 688901 871032 717600 877798
rect 687949 870728 717600 871032
rect 687949 867891 688145 870728
rect 687293 867587 688145 867891
rect 677707 779862 687193 788598
rect 677707 773534 687067 779862
rect 677707 773406 677927 773534
rect 39673 756866 39893 756994
rect 30533 750538 39893 756866
rect 30407 741802 39893 750538
rect 29455 708509 30307 708813
rect 29455 705672 29651 708509
rect 0 705368 29651 705672
rect 0 698602 28699 705368
rect 0 698334 28573 698602
rect 0 698000 4843 698254
rect 4923 698193 20920 698334
rect 21000 698000 25993 698254
rect 26073 698193 26213 698334
rect 0 670800 5193 698000
rect 20593 670800 26213 698000
rect 0 670546 4843 670800
rect 4923 670466 20920 670594
rect 21000 670546 25993 670800
rect 26073 670466 26213 670594
rect 26293 670546 27183 698254
rect 27263 698193 27383 698334
rect 27263 670800 27383 697800
rect 27263 670466 27383 670594
rect 27463 670546 28353 698254
rect 28433 698193 28573 698334
rect 28433 670800 28573 698000
rect 28433 670466 28573 670594
rect 0 664138 28573 670466
rect 28653 664218 28719 698522
rect 0 662472 28699 664138
rect 28779 662552 29375 705288
rect 29455 698334 29651 705368
rect 29435 698000 29671 698254
rect 29455 670800 29651 698000
rect 29435 670546 29671 670800
rect 29455 665613 29651 670466
rect 29731 665693 30327 708429
rect 30387 707418 30453 741722
rect 30533 741534 39893 741802
rect 30533 741393 30673 741534
rect 30533 713666 30673 713794
rect 30753 713746 31683 741454
rect 31763 741393 31883 741534
rect 31763 713666 31883 713794
rect 31963 713746 32653 741454
rect 32733 741393 32853 741534
rect 32733 713666 32853 713794
rect 32933 713746 33623 741454
rect 33703 741393 33823 741534
rect 33703 713666 33823 713794
rect 33903 713746 34833 741454
rect 34913 741393 35033 741534
rect 36123 741473 37213 741534
rect 34913 713666 35033 713794
rect 35113 713746 36043 741454
rect 36123 741393 36243 741473
rect 37093 741393 37213 741473
rect 36323 713794 37013 741393
rect 36123 713714 36243 713794
rect 37093 713714 37213 713794
rect 37293 713746 38223 741454
rect 38303 741393 38423 741534
rect 36123 713666 37213 713714
rect 38303 713666 38423 713794
rect 38503 713746 39593 741454
rect 39673 741393 39893 741534
rect 677707 743866 677927 744007
rect 678007 743946 679097 773454
rect 679177 773406 679297 773534
rect 680387 773486 681477 773534
rect 679177 743866 679297 744007
rect 679377 743946 680307 773454
rect 680387 773406 680507 773486
rect 681357 773406 681477 773486
rect 680587 744007 681277 773406
rect 680387 743927 680507 744007
rect 681357 743927 681477 744007
rect 681557 743946 682487 773454
rect 682567 773406 682687 773534
rect 680387 743866 681477 743927
rect 682567 743866 682687 744007
rect 682767 743946 683697 773454
rect 683777 773406 683897 773534
rect 683777 743866 683897 744007
rect 683977 743946 684667 773454
rect 684747 773406 684867 773534
rect 684747 743866 684867 744007
rect 684947 743946 685637 773454
rect 685717 773406 685837 773534
rect 685717 743866 685837 744007
rect 685917 743946 686847 773454
rect 686927 773406 687067 773534
rect 686927 743866 687067 744007
rect 677707 743598 687067 743866
rect 687147 743678 687213 779782
rect 687273 778771 687869 867507
rect 687949 862734 688145 867587
rect 687929 862400 688165 862654
rect 687949 833400 688145 862400
rect 687929 833146 688165 833400
rect 687949 818734 688145 833066
rect 687929 818400 688165 818654
rect 687949 789200 688145 818400
rect 687929 788946 688165 789200
rect 687949 781832 688145 788866
rect 688225 781912 688821 870648
rect 688901 869062 717600 870728
rect 688881 788678 688947 868982
rect 689027 862734 717600 869062
rect 689027 862606 689167 862734
rect 689027 833400 689167 862400
rect 689027 833066 689167 833207
rect 689247 833146 690137 862654
rect 690217 862606 690337 862734
rect 690217 833400 690337 862400
rect 690217 833066 690337 833207
rect 690417 833146 691307 862654
rect 691387 862606 691527 862734
rect 691607 862400 696600 862654
rect 696680 862606 712677 862734
rect 712757 862400 717600 862654
rect 691387 833400 697007 862400
rect 712407 833400 717600 862400
rect 691387 833066 691527 833207
rect 691607 833146 696600 833400
rect 696680 833066 712677 833207
rect 712757 833146 717600 833400
rect 689027 818734 717600 833066
rect 689027 818593 689167 818734
rect 689027 789200 689167 818400
rect 689027 788866 689167 789007
rect 689247 788946 690137 818654
rect 690217 818593 690337 818734
rect 690217 789200 690337 818200
rect 690217 788866 690337 789007
rect 690417 788946 691307 818654
rect 691387 818593 691527 818734
rect 691607 818400 696600 818654
rect 696680 818593 712677 818734
rect 712757 818400 717600 818654
rect 691387 789200 697007 818400
rect 712407 789200 717600 818400
rect 691387 788866 691527 789007
rect 691607 788946 696600 789200
rect 696680 788866 712677 789007
rect 712757 788946 717600 789200
rect 689027 788598 717600 788866
rect 688901 781832 717600 788598
rect 687949 781528 717600 781832
rect 687949 778691 688145 781528
rect 687293 778387 688145 778691
rect 677707 734862 687193 743598
rect 677707 728534 687067 734862
rect 677707 728406 677927 728534
rect 39673 713666 39893 713794
rect 30533 707338 39893 713666
rect 30407 698602 39893 707338
rect 29455 665309 30307 665613
rect 29455 662472 29651 665309
rect 0 662168 29651 662472
rect 0 655402 28699 662168
rect 0 655134 28573 655402
rect 0 654800 4843 655054
rect 4923 654993 20920 655134
rect 21000 654800 25993 655054
rect 26073 654993 26213 655134
rect 0 627600 5193 654800
rect 20593 627600 26213 654800
rect 0 627346 4843 627600
rect 4923 627266 20920 627394
rect 21000 627346 25993 627600
rect 26073 627266 26213 627394
rect 26293 627346 27183 655054
rect 27263 654993 27383 655134
rect 27263 627600 27383 654600
rect 27263 627266 27383 627394
rect 27463 627346 28353 655054
rect 28433 654993 28573 655134
rect 28433 627600 28573 654800
rect 28433 627266 28573 627394
rect 0 620938 28573 627266
rect 28653 621018 28719 655322
rect 0 619272 28699 620938
rect 28779 619352 29375 662088
rect 29455 655134 29651 662168
rect 29435 654800 29671 655054
rect 29455 627600 29651 654800
rect 29435 627346 29671 627600
rect 29455 622413 29651 627266
rect 29731 622493 30327 665229
rect 30387 664218 30453 698522
rect 30533 698334 39893 698602
rect 30533 698193 30673 698334
rect 30533 670466 30673 670594
rect 30753 670546 31683 698254
rect 31763 698193 31883 698334
rect 31763 670466 31883 670594
rect 31963 670546 32653 698254
rect 32733 698193 32853 698334
rect 32733 670466 32853 670594
rect 32933 670546 33623 698254
rect 33703 698193 33823 698334
rect 33703 670466 33823 670594
rect 33903 670546 34833 698254
rect 34913 698193 35033 698334
rect 36123 698273 37213 698334
rect 34913 670466 35033 670594
rect 35113 670546 36043 698254
rect 36123 698193 36243 698273
rect 37093 698193 37213 698273
rect 36323 670594 37013 698193
rect 36123 670514 36243 670594
rect 37093 670514 37213 670594
rect 37293 670546 38223 698254
rect 38303 698193 38423 698334
rect 36123 670466 37213 670514
rect 38303 670466 38423 670594
rect 38503 670546 39593 698254
rect 39673 698193 39893 698334
rect 677707 698866 677927 699007
rect 678007 698946 679097 728454
rect 679177 728406 679297 728534
rect 680387 728486 681477 728534
rect 679177 698866 679297 699007
rect 679377 698946 680307 728454
rect 680387 728406 680507 728486
rect 681357 728406 681477 728486
rect 680587 699007 681277 728406
rect 680387 698927 680507 699007
rect 681357 698927 681477 699007
rect 681557 698946 682487 728454
rect 682567 728406 682687 728534
rect 680387 698866 681477 698927
rect 682567 698866 682687 699007
rect 682767 698946 683697 728454
rect 683777 728406 683897 728534
rect 683777 698866 683897 699007
rect 683977 698946 684667 728454
rect 684747 728406 684867 728534
rect 684747 698866 684867 699007
rect 684947 698946 685637 728454
rect 685717 728406 685837 728534
rect 685717 698866 685837 699007
rect 685917 698946 686847 728454
rect 686927 728406 687067 728534
rect 686927 698866 687067 699007
rect 677707 698598 687067 698866
rect 687147 698678 687213 734782
rect 687273 733771 687869 778307
rect 687949 773534 688145 778387
rect 687929 773200 688165 773454
rect 687949 744200 688145 773200
rect 687929 743946 688165 744200
rect 687949 736832 688145 743866
rect 688225 736912 688821 781448
rect 688901 779862 717600 781528
rect 688881 743678 688947 779782
rect 689027 773534 717600 779862
rect 689027 773406 689167 773534
rect 689027 744200 689167 773200
rect 689027 743866 689167 744007
rect 689247 743946 690137 773454
rect 690217 773406 690337 773534
rect 690217 744200 690337 773200
rect 690217 743866 690337 744007
rect 690417 743946 691307 773454
rect 691387 773406 691527 773534
rect 691607 773200 696600 773454
rect 696680 773406 712677 773534
rect 712757 773200 717600 773454
rect 691387 744200 697007 773200
rect 712407 744200 717600 773200
rect 691387 743866 691527 744007
rect 691607 743946 696600 744200
rect 696680 743866 712677 744007
rect 712757 743946 717600 744200
rect 689027 743598 717600 743866
rect 688901 736832 717600 743598
rect 687949 736528 717600 736832
rect 687949 733691 688145 736528
rect 687293 733387 688145 733691
rect 677707 689862 687193 698598
rect 677707 683534 687067 689862
rect 677707 683406 677927 683534
rect 39673 670466 39893 670594
rect 30533 664138 39893 670466
rect 30407 655402 39893 664138
rect 29455 622109 30307 622413
rect 29455 619272 29651 622109
rect 0 618968 29651 619272
rect 0 612202 28699 618968
rect 0 611934 28573 612202
rect 0 611600 4843 611854
rect 4923 611793 20920 611934
rect 21000 611600 25993 611854
rect 26073 611793 26213 611934
rect 0 584400 5193 611600
rect 20593 584400 26213 611600
rect 0 584146 4843 584400
rect 4923 584066 20920 584194
rect 21000 584146 25993 584400
rect 26073 584066 26213 584194
rect 26293 584146 27183 611854
rect 27263 611793 27383 611934
rect 27263 584400 27383 611400
rect 27263 584066 27383 584194
rect 27463 584146 28353 611854
rect 28433 611793 28573 611934
rect 28433 584400 28573 611600
rect 28433 584066 28573 584194
rect 0 577738 28573 584066
rect 28653 577818 28719 612122
rect 0 576072 28699 577738
rect 28779 576152 29375 618888
rect 29455 611934 29651 618968
rect 29435 611600 29671 611854
rect 29455 584400 29651 611600
rect 29435 584146 29671 584400
rect 29455 579213 29651 584066
rect 29731 579293 30327 622029
rect 30387 621018 30453 655322
rect 30533 655134 39893 655402
rect 30533 654993 30673 655134
rect 30533 627266 30673 627394
rect 30753 627346 31683 655054
rect 31763 654993 31883 655134
rect 31763 627266 31883 627394
rect 31963 627346 32653 655054
rect 32733 654993 32853 655134
rect 32733 627266 32853 627394
rect 32933 627346 33623 655054
rect 33703 654993 33823 655134
rect 33703 627266 33823 627394
rect 33903 627346 34833 655054
rect 34913 654993 35033 655134
rect 36123 655073 37213 655134
rect 34913 627266 35033 627394
rect 35113 627346 36043 655054
rect 36123 654993 36243 655073
rect 37093 654993 37213 655073
rect 36323 627394 37013 654993
rect 36123 627314 36243 627394
rect 37093 627314 37213 627394
rect 37293 627346 38223 655054
rect 38303 654993 38423 655134
rect 36123 627266 37213 627314
rect 38303 627266 38423 627394
rect 38503 627346 39593 655054
rect 39673 654993 39893 655134
rect 677707 653666 677927 653807
rect 678007 653746 679097 683454
rect 679177 683406 679297 683534
rect 680387 683486 681477 683534
rect 679177 653666 679297 653807
rect 679377 653746 680307 683454
rect 680387 683406 680507 683486
rect 681357 683406 681477 683486
rect 680587 653807 681277 683406
rect 680387 653727 680507 653807
rect 681357 653727 681477 653807
rect 681557 653746 682487 683454
rect 682567 683406 682687 683534
rect 680387 653666 681477 653727
rect 682567 653666 682687 653807
rect 682767 653746 683697 683454
rect 683777 683406 683897 683534
rect 683777 653666 683897 653807
rect 683977 653746 684667 683454
rect 684747 683406 684867 683534
rect 684747 653666 684867 653807
rect 684947 653746 685637 683454
rect 685717 683406 685837 683534
rect 685717 653666 685837 653807
rect 685917 653746 686847 683454
rect 686927 683406 687067 683534
rect 686927 653666 687067 653807
rect 677707 653398 687067 653666
rect 687147 653478 687213 689782
rect 687273 688771 687869 733307
rect 687949 728534 688145 733387
rect 687929 728200 688165 728454
rect 687949 699200 688145 728200
rect 687929 698946 688165 699200
rect 687949 691832 688145 698866
rect 688225 691912 688821 736448
rect 688901 734862 717600 736528
rect 688881 698678 688947 734782
rect 689027 728534 717600 734862
rect 689027 728406 689167 728534
rect 689027 699200 689167 728200
rect 689027 698866 689167 699007
rect 689247 698946 690137 728454
rect 690217 728406 690337 728534
rect 690217 699200 690337 728200
rect 690217 698866 690337 699007
rect 690417 698946 691307 728454
rect 691387 728406 691527 728534
rect 691607 728200 696600 728454
rect 696680 728406 712677 728534
rect 712757 728200 717600 728454
rect 691387 699200 697007 728200
rect 712407 699200 717600 728200
rect 691387 698866 691527 699007
rect 691607 698946 696600 699200
rect 696680 698866 712677 699007
rect 712757 698946 717600 699200
rect 689027 698598 717600 698866
rect 688901 691832 717600 698598
rect 687949 691528 717600 691832
rect 687949 688691 688145 691528
rect 687293 688387 688145 688691
rect 677707 644662 687193 653398
rect 677707 638334 687067 644662
rect 677707 638206 677927 638334
rect 39673 627266 39893 627394
rect 30533 620938 39893 627266
rect 30407 612202 39893 620938
rect 29455 578909 30307 579213
rect 29455 576072 29651 578909
rect 0 575768 29651 576072
rect 0 569002 28699 575768
rect 0 568734 28573 569002
rect 0 568400 4843 568654
rect 4923 568593 20920 568734
rect 21000 568400 25993 568654
rect 26073 568593 26213 568734
rect 0 541200 5193 568400
rect 20593 541200 26213 568400
rect 0 540946 4843 541200
rect 4923 540866 20920 540994
rect 21000 540946 25993 541200
rect 26073 540866 26213 540994
rect 26293 540946 27183 568654
rect 27263 568593 27383 568734
rect 27263 541200 27383 568200
rect 27263 540866 27383 540994
rect 27463 540946 28353 568654
rect 28433 568593 28573 568734
rect 28433 541200 28573 568400
rect 28433 540866 28573 540994
rect 0 534538 28573 540866
rect 28653 534618 28719 568922
rect 0 532872 28699 534538
rect 28779 532952 29375 575688
rect 29455 568734 29651 575768
rect 29435 568400 29671 568654
rect 29455 541200 29651 568400
rect 29435 540946 29671 541200
rect 29455 536013 29651 540866
rect 29731 536093 30327 578829
rect 30387 577818 30453 612122
rect 30533 611934 39893 612202
rect 30533 611793 30673 611934
rect 30533 584066 30673 584194
rect 30753 584146 31683 611854
rect 31763 611793 31883 611934
rect 31763 584066 31883 584194
rect 31963 584146 32653 611854
rect 32733 611793 32853 611934
rect 32733 584066 32853 584194
rect 32933 584146 33623 611854
rect 33703 611793 33823 611934
rect 33703 584066 33823 584194
rect 33903 584146 34833 611854
rect 34913 611793 35033 611934
rect 36123 611873 37213 611934
rect 34913 584066 35033 584194
rect 35113 584146 36043 611854
rect 36123 611793 36243 611873
rect 37093 611793 37213 611873
rect 36323 584194 37013 611793
rect 36123 584114 36243 584194
rect 37093 584114 37213 584194
rect 37293 584146 38223 611854
rect 38303 611793 38423 611934
rect 36123 584066 37213 584114
rect 38303 584066 38423 584194
rect 38503 584146 39593 611854
rect 39673 611793 39893 611934
rect 677707 608666 677927 608807
rect 678007 608746 679097 638254
rect 679177 638206 679297 638334
rect 680387 638286 681477 638334
rect 679177 608666 679297 608807
rect 679377 608746 680307 638254
rect 680387 638206 680507 638286
rect 681357 638206 681477 638286
rect 680587 608807 681277 638206
rect 680387 608727 680507 608807
rect 681357 608727 681477 608807
rect 681557 608746 682487 638254
rect 682567 638206 682687 638334
rect 680387 608666 681477 608727
rect 682567 608666 682687 608807
rect 682767 608746 683697 638254
rect 683777 638206 683897 638334
rect 683777 608666 683897 608807
rect 683977 608746 684667 638254
rect 684747 638206 684867 638334
rect 684747 608666 684867 608807
rect 684947 608746 685637 638254
rect 685717 638206 685837 638334
rect 685717 608666 685837 608807
rect 685917 608746 686847 638254
rect 686927 638206 687067 638334
rect 686927 608666 687067 608807
rect 677707 608398 687067 608666
rect 687147 608478 687213 644582
rect 687273 643571 687869 688307
rect 687949 683534 688145 688387
rect 687929 683200 688165 683454
rect 687949 654000 688145 683200
rect 687929 653746 688165 654000
rect 687949 646632 688145 653666
rect 688225 646712 688821 691448
rect 688901 689862 717600 691528
rect 688881 653478 688947 689782
rect 689027 683534 717600 689862
rect 689027 683406 689167 683534
rect 689027 654000 689167 683200
rect 689027 653666 689167 653807
rect 689247 653746 690137 683454
rect 690217 683406 690337 683534
rect 690217 654000 690337 683000
rect 690217 653666 690337 653807
rect 690417 653746 691307 683454
rect 691387 683406 691527 683534
rect 691607 683200 696600 683454
rect 696680 683406 712677 683534
rect 712757 683200 717600 683454
rect 691387 654000 697007 683200
rect 712407 654000 717600 683200
rect 691387 653666 691527 653807
rect 691607 653746 696600 654000
rect 696680 653666 712677 653807
rect 712757 653746 717600 654000
rect 689027 653398 717600 653666
rect 688901 646632 717600 653398
rect 687949 646328 717600 646632
rect 687949 643491 688145 646328
rect 687293 643187 688145 643491
rect 677707 599662 687193 608398
rect 677707 593334 687067 599662
rect 677707 593206 677927 593334
rect 39673 584066 39893 584194
rect 30533 577738 39893 584066
rect 30407 569002 39893 577738
rect 29455 535709 30307 536013
rect 29455 532872 29651 535709
rect 0 532568 29651 532872
rect 0 525802 28699 532568
rect 0 525534 28573 525802
rect 0 525200 4843 525454
rect 4923 525393 20920 525534
rect 21000 525200 25993 525454
rect 26073 525393 26213 525534
rect 0 498000 5193 525200
rect 20593 498000 26213 525200
rect 0 497746 4843 498000
rect 4923 497666 20920 497807
rect 21000 497746 25993 498000
rect 26073 497666 26213 497807
rect 26293 497746 27183 525454
rect 27263 525393 27383 525534
rect 27263 498000 27383 525000
rect 27263 497666 27383 497807
rect 27463 497746 28353 525454
rect 28433 525393 28573 525534
rect 28433 498000 28573 525200
rect 28433 497666 28573 497807
rect 0 483334 28573 497666
rect 0 483000 4843 483254
rect 4923 483193 20920 483334
rect 21000 483000 25993 483254
rect 26073 483193 26213 483334
rect 0 455800 5193 483000
rect 20593 455800 26213 483000
rect 0 455546 4843 455800
rect 4923 455466 20920 455800
rect 21000 455546 25993 455800
rect 26073 455466 26213 455800
rect 26293 455546 27183 483254
rect 27263 483193 27383 483334
rect 27263 455466 27383 482800
rect 27463 455546 28353 483254
rect 28433 483193 28573 483334
rect 28433 455466 28573 483000
rect 0 441134 28573 455466
rect 0 440800 4843 441054
rect 4923 440993 20920 441134
rect 21000 440800 25993 441054
rect 26073 440993 26213 441134
rect 0 413600 5193 440800
rect 20593 413600 26213 440800
rect 0 413346 4843 413600
rect 4923 413266 20920 413394
rect 21000 413346 25993 413600
rect 26073 413266 26213 413394
rect 26293 413346 27183 441054
rect 27263 440993 27383 441134
rect 27263 413600 27383 440600
rect 27263 413266 27383 413394
rect 27463 413346 28353 441054
rect 28433 440993 28573 441134
rect 28433 413600 28573 440800
rect 28433 413266 28573 413394
rect 0 406938 28573 413266
rect 28653 407018 28719 525722
rect 0 405272 28699 406938
rect 28779 405352 29375 532488
rect 29455 525534 29651 532568
rect 29435 525200 29671 525454
rect 29455 498000 29651 525200
rect 29435 497746 29671 498000
rect 29455 483334 29651 497666
rect 29435 483000 29671 483254
rect 29455 455800 29651 483000
rect 29435 455546 29671 455800
rect 29455 441134 29651 455466
rect 29435 440800 29671 441054
rect 29455 413600 29651 440800
rect 29435 413346 29671 413600
rect 29455 408413 29651 413266
rect 29731 408493 30327 535629
rect 30387 534618 30453 568922
rect 30533 568734 39893 569002
rect 30533 568593 30673 568734
rect 30533 540866 30673 540994
rect 30753 540946 31683 568654
rect 31763 568593 31883 568734
rect 31763 540866 31883 540994
rect 31963 540946 32653 568654
rect 32733 568593 32853 568734
rect 32733 540866 32853 540994
rect 32933 540946 33623 568654
rect 33703 568593 33823 568734
rect 33703 540866 33823 540994
rect 33903 540946 34833 568654
rect 34913 568593 35033 568734
rect 36123 568673 37213 568734
rect 34913 540866 35033 540994
rect 35113 540946 36043 568654
rect 36123 568593 36243 568673
rect 37093 568593 37213 568673
rect 36323 540994 37013 568593
rect 36123 540914 36243 540994
rect 37093 540914 37213 540994
rect 37293 540946 38223 568654
rect 38303 568593 38423 568734
rect 36123 540866 37213 540914
rect 38303 540866 38423 540994
rect 38503 540946 39593 568654
rect 39673 568593 39893 568734
rect 677707 563466 677927 563607
rect 678007 563546 679097 593254
rect 679177 593206 679297 593334
rect 680387 593286 681477 593334
rect 679177 563466 679297 563607
rect 679377 563546 680307 593254
rect 680387 593206 680507 593286
rect 681357 593206 681477 593286
rect 680587 563607 681277 593206
rect 680387 563527 680507 563607
rect 681357 563527 681477 563607
rect 681557 563546 682487 593254
rect 682567 593206 682687 593334
rect 680387 563466 681477 563527
rect 682567 563466 682687 563607
rect 682767 563546 683697 593254
rect 683777 593206 683897 593334
rect 683777 563466 683897 563607
rect 683977 563546 684667 593254
rect 684747 593206 684867 593334
rect 684747 563466 684867 563607
rect 684947 563546 685637 593254
rect 685717 593206 685837 593334
rect 685717 563466 685837 563607
rect 685917 563546 686847 593254
rect 686927 593206 687067 593334
rect 686927 563466 687067 563607
rect 677707 563198 687067 563466
rect 687147 563278 687213 599582
rect 687273 598571 687869 643107
rect 687949 638334 688145 643187
rect 687929 638000 688165 638254
rect 687949 609000 688145 638000
rect 687929 608746 688165 609000
rect 687949 601632 688145 608666
rect 688225 601712 688821 646248
rect 688901 644662 717600 646328
rect 688881 608478 688947 644582
rect 689027 638334 717600 644662
rect 689027 638206 689167 638334
rect 689027 609000 689167 638000
rect 689027 608666 689167 608807
rect 689247 608746 690137 638254
rect 690217 638206 690337 638334
rect 690217 609000 690337 638000
rect 690217 608666 690337 608807
rect 690417 608746 691307 638254
rect 691387 638206 691527 638334
rect 691607 638000 696600 638254
rect 696680 638206 712677 638334
rect 712757 638000 717600 638254
rect 691387 609000 697007 638000
rect 712407 609000 717600 638000
rect 691387 608666 691527 608807
rect 691607 608746 696600 609000
rect 696680 608666 712677 608807
rect 712757 608746 717600 609000
rect 689027 608398 717600 608666
rect 688901 601632 717600 608398
rect 687949 601328 717600 601632
rect 687949 598491 688145 601328
rect 687293 598187 688145 598491
rect 677707 554462 687193 563198
rect 677707 548134 687067 554462
rect 677707 548006 677927 548134
rect 39673 540866 39893 540994
rect 30533 534538 39893 540866
rect 30407 525802 39893 534538
rect 29455 408109 30307 408413
rect 29455 405272 29651 408109
rect 0 404968 29651 405272
rect 0 398202 28699 404968
rect 0 397934 28573 398202
rect 0 397600 4843 397854
rect 4923 397793 20920 397934
rect 21000 397600 25993 397854
rect 26073 397793 26213 397934
rect 0 370400 5193 397600
rect 20593 370400 26213 397600
rect 0 370146 4843 370400
rect 4923 370066 20920 370194
rect 21000 370146 25993 370400
rect 26073 370066 26213 370194
rect 26293 370146 27183 397854
rect 27263 397793 27383 397934
rect 27263 370400 27383 397400
rect 27263 370066 27383 370194
rect 27463 370146 28353 397854
rect 28433 397793 28573 397934
rect 28433 370400 28573 397600
rect 28433 370066 28573 370194
rect 0 363738 28573 370066
rect 28653 363818 28719 398122
rect 0 362072 28699 363738
rect 28779 362152 29375 404888
rect 29455 397934 29651 404968
rect 29435 397600 29671 397854
rect 29455 370400 29651 397600
rect 29435 370146 29671 370400
rect 29455 365213 29651 370066
rect 29731 365293 30327 408029
rect 30387 407018 30453 525722
rect 30533 525534 39893 525802
rect 30533 525393 30673 525534
rect 30533 497666 30673 497807
rect 30753 497746 31683 525454
rect 31763 525393 31883 525534
rect 31763 497666 31883 497807
rect 31963 497746 32653 525454
rect 32733 525393 32853 525534
rect 32733 497666 32853 497807
rect 32933 497746 33623 525454
rect 33703 525393 33823 525534
rect 33703 497666 33823 497807
rect 33903 497746 34833 525454
rect 34913 525393 35033 525534
rect 36123 525473 37213 525534
rect 34913 497666 35033 497807
rect 35113 497746 36043 525454
rect 36123 525393 36243 525473
rect 37093 525393 37213 525473
rect 36123 497727 36243 497807
rect 37093 497727 37213 497807
rect 37293 497746 38223 525454
rect 38303 525393 38423 525534
rect 36123 497666 37213 497727
rect 38303 497666 38423 497807
rect 38503 497746 39593 525454
rect 39673 525393 39893 525534
rect 678007 518546 679097 548054
rect 679177 548006 679297 548134
rect 680387 548086 681477 548134
rect 679177 518466 679297 518607
rect 679377 518546 680307 548054
rect 680387 548006 680507 548086
rect 681357 548006 681477 548086
rect 680587 518607 681277 548006
rect 680387 518527 680507 518607
rect 681357 518527 681477 518607
rect 681557 518546 682487 548054
rect 682567 548006 682687 548134
rect 680387 518466 681477 518527
rect 682567 518466 682687 518607
rect 682767 518546 683697 548054
rect 683777 548006 683897 548134
rect 683777 518466 683897 518607
rect 683977 518546 684667 548054
rect 684747 548006 684867 548134
rect 684747 518466 684867 518607
rect 684947 518546 685637 548054
rect 685717 548006 685837 548134
rect 685717 518466 685837 518607
rect 685917 518546 686847 548054
rect 686927 548006 687067 548134
rect 686927 518466 687067 518607
rect 678007 504134 687067 518466
rect 30533 483334 39593 497666
rect 30533 483193 30673 483334
rect 30533 455466 30673 455800
rect 31763 483193 31883 483334
rect 31763 455466 31883 455800
rect 31963 455546 32653 483254
rect 32733 483193 32853 483334
rect 32733 455466 32853 455800
rect 32933 455546 33623 483254
rect 33703 483193 33823 483334
rect 33703 455466 33823 455800
rect 33903 455546 34833 483254
rect 34913 483193 35033 483334
rect 36123 483273 37213 483334
rect 34913 455466 35033 455800
rect 35113 455546 36043 483254
rect 36123 483193 36243 483273
rect 37093 483193 37213 483273
rect 36123 455527 36243 455800
rect 37093 455527 37213 455800
rect 37293 455546 38223 483254
rect 38303 483193 38423 483334
rect 36123 455466 37213 455527
rect 38303 455466 38423 455800
rect 38503 455546 39593 483254
rect 678007 474546 679097 504054
rect 679177 503993 679297 504134
rect 680387 504073 681477 504134
rect 679177 474466 679297 474607
rect 679377 474546 680307 504054
rect 680387 503993 680507 504073
rect 681357 503993 681477 504073
rect 680587 474607 681277 503993
rect 680387 474527 680507 474607
rect 681357 474527 681477 474607
rect 681557 474546 682487 504054
rect 682567 503993 682687 504134
rect 680387 474466 681477 474527
rect 682567 474466 682687 474607
rect 682767 474546 683697 504054
rect 683777 503993 683897 504134
rect 683777 474466 683897 474607
rect 683977 474546 684667 504054
rect 684747 503993 684867 504134
rect 684747 474466 684867 474607
rect 684947 474546 685637 504054
rect 685717 503993 685837 504134
rect 685717 474466 685837 474607
rect 686927 503993 687067 504134
rect 686927 474466 687067 474607
rect 678007 460134 687067 474466
rect 30533 441134 39593 455466
rect 30533 440993 30673 441134
rect 30533 413266 30673 413394
rect 31763 440993 31883 441134
rect 31763 413266 31883 413394
rect 31963 413346 32653 441054
rect 32733 440993 32853 441134
rect 32733 413266 32853 413394
rect 32933 413346 33623 441054
rect 33703 440993 33823 441134
rect 33703 413266 33823 413394
rect 33903 413346 34833 441054
rect 34913 440993 35033 441134
rect 36123 441073 37213 441134
rect 34913 413266 35033 413394
rect 35113 413346 36043 441054
rect 36123 440993 36243 441073
rect 37093 440993 37213 441073
rect 36323 413394 37013 440993
rect 36123 413314 36243 413394
rect 37093 413314 37213 413394
rect 37293 413346 38223 441054
rect 38303 440993 38423 441134
rect 36123 413266 37213 413314
rect 38303 413266 38423 413394
rect 38503 413346 39593 441054
rect 678007 430346 679097 460054
rect 679177 459800 679297 460134
rect 680387 460073 681477 460134
rect 679177 430266 679297 430407
rect 679377 430346 680307 460054
rect 680387 459800 680507 460073
rect 680587 430407 681277 459993
rect 681357 459800 681477 460073
rect 680387 430327 680507 430407
rect 681357 430327 681477 430407
rect 681557 430346 682487 460054
rect 682567 459800 682687 460134
rect 680387 430266 681477 430327
rect 682567 430266 682687 430407
rect 682767 430346 683697 460054
rect 683777 459800 683897 460134
rect 683777 430266 683897 430407
rect 683977 430346 684667 460054
rect 684747 459800 684867 460134
rect 684747 430266 684867 430407
rect 684947 430346 685637 460054
rect 685717 459800 685837 460134
rect 685717 430266 685837 430407
rect 686927 459800 687067 460134
rect 686927 430266 687067 430407
rect 687147 430346 687213 554382
rect 687273 553371 687869 598107
rect 687949 593334 688145 598187
rect 687929 593000 688165 593254
rect 687949 563800 688145 593000
rect 687929 563546 688165 563800
rect 687949 556432 688145 563466
rect 688225 556512 688821 601248
rect 688901 599662 717600 601328
rect 688881 563278 688947 599582
rect 689027 593334 717600 599662
rect 689027 593206 689167 593334
rect 689027 563800 689167 593000
rect 689027 563466 689167 563607
rect 689247 563546 690137 593254
rect 690217 593206 690337 593334
rect 690217 563800 690337 592800
rect 690217 563466 690337 563607
rect 690417 563546 691307 593254
rect 691387 593206 691527 593334
rect 691607 593000 696600 593254
rect 696680 593206 712677 593334
rect 712757 593000 717600 593254
rect 691387 563800 697007 593000
rect 712407 563800 717600 593000
rect 691387 563466 691527 563607
rect 691607 563546 696600 563800
rect 696680 563466 712677 563607
rect 712757 563546 717600 563800
rect 689027 563198 717600 563466
rect 688901 556432 717600 563198
rect 687949 556128 717600 556432
rect 687949 553291 688145 556128
rect 687293 552987 688145 553291
rect 678007 415934 687193 430266
rect 39673 413266 39893 413394
rect 30533 406938 39893 413266
rect 30407 398202 39893 406938
rect 29455 364909 30307 365213
rect 29455 362072 29651 364909
rect 0 361768 29651 362072
rect 0 355002 28699 361768
rect 0 354734 28573 355002
rect 0 354400 4843 354654
rect 4923 354593 20920 354734
rect 21000 354400 25993 354654
rect 26073 354593 26213 354734
rect 0 327200 5193 354400
rect 20593 327200 26213 354400
rect 0 326946 4843 327200
rect 4923 326866 20920 326994
rect 21000 326946 25993 327200
rect 26073 326866 26213 326994
rect 26293 326946 27183 354654
rect 27263 354593 27383 354734
rect 27263 327200 27383 354200
rect 27263 326866 27383 326994
rect 27463 326946 28353 354654
rect 28433 354593 28573 354734
rect 28433 327200 28573 354400
rect 28433 326866 28573 326994
rect 0 320538 28573 326866
rect 28653 320618 28719 354922
rect 0 318872 28699 320538
rect 28779 318952 29375 361688
rect 29455 354734 29651 361768
rect 29435 354400 29671 354654
rect 29455 327200 29651 354400
rect 29435 326946 29671 327200
rect 29455 322013 29651 326866
rect 29731 322093 30327 364829
rect 30387 363818 30453 398122
rect 30533 397934 39893 398202
rect 30533 397793 30673 397934
rect 30533 370066 30673 370194
rect 30753 370146 31683 397854
rect 31763 397793 31883 397934
rect 31763 370066 31883 370194
rect 31963 370146 32653 397854
rect 32733 397793 32853 397934
rect 32733 370066 32853 370194
rect 32933 370146 33623 397854
rect 33703 397793 33823 397934
rect 33703 370066 33823 370194
rect 33903 370146 34833 397854
rect 34913 397793 35033 397934
rect 36123 397873 37213 397934
rect 34913 370066 35033 370194
rect 35113 370146 36043 397854
rect 36123 397793 36243 397873
rect 37093 397793 37213 397873
rect 36323 370194 37013 397793
rect 36123 370114 36243 370194
rect 37093 370114 37213 370194
rect 37293 370146 38223 397854
rect 38303 397793 38423 397934
rect 36123 370066 37213 370114
rect 38303 370066 38423 370194
rect 38503 370146 39593 397854
rect 39673 397793 39893 397934
rect 677707 386266 677927 386407
rect 678007 386346 679097 415854
rect 679177 415793 679297 415934
rect 680387 415873 681477 415934
rect 679177 386266 679297 386407
rect 679377 386346 680307 415854
rect 680387 415793 680507 415873
rect 681357 415793 681477 415873
rect 680587 386407 681277 415793
rect 680387 386327 680507 386407
rect 681357 386327 681477 386407
rect 681557 386346 682487 415854
rect 682567 415793 682687 415934
rect 680387 386266 681477 386327
rect 682567 386266 682687 386407
rect 682767 386346 683697 415854
rect 683777 415793 683897 415934
rect 683777 386266 683897 386407
rect 683977 386346 684667 415854
rect 684747 415793 684867 415934
rect 684747 386266 684867 386407
rect 684947 386346 685637 415854
rect 685717 415793 685837 415934
rect 685717 386266 685837 386407
rect 685917 386346 686847 415854
rect 686927 415793 687067 415934
rect 686927 386266 687067 386407
rect 677707 385998 687067 386266
rect 687147 386078 687213 415854
rect 677707 377262 687193 385998
rect 677707 370934 687067 377262
rect 677707 370806 677927 370934
rect 39673 370066 39893 370194
rect 30533 363738 39893 370066
rect 30407 355002 39893 363738
rect 29455 321709 30307 322013
rect 29455 318872 29651 321709
rect 0 318568 29651 318872
rect 0 311802 28699 318568
rect 0 311534 28573 311802
rect 0 311200 4843 311454
rect 4923 311393 20920 311534
rect 21000 311200 25993 311454
rect 26073 311393 26213 311534
rect 0 284000 5193 311200
rect 20593 284000 26213 311200
rect 0 283746 4843 284000
rect 4923 283666 20920 283794
rect 21000 283746 25993 284000
rect 26073 283666 26213 283794
rect 26293 283746 27183 311454
rect 27263 311393 27383 311534
rect 27263 284000 27383 311000
rect 27263 283666 27383 283794
rect 27463 283746 28353 311454
rect 28433 311393 28573 311534
rect 28433 284000 28573 311200
rect 28433 283666 28573 283794
rect 0 277338 28573 283666
rect 28653 277418 28719 311722
rect 0 275672 28699 277338
rect 28779 275752 29375 318488
rect 29455 311534 29651 318568
rect 29435 311200 29671 311454
rect 29455 284000 29651 311200
rect 29435 283746 29671 284000
rect 29455 278813 29651 283666
rect 29731 278893 30327 321629
rect 30387 320618 30453 354922
rect 30533 354734 39893 355002
rect 30533 354593 30673 354734
rect 30533 326866 30673 326994
rect 30753 326946 31683 354654
rect 31763 354593 31883 354734
rect 31763 326866 31883 326994
rect 31963 326946 32653 354654
rect 32733 354593 32853 354734
rect 32733 326866 32853 326994
rect 32933 326946 33623 354654
rect 33703 354593 33823 354734
rect 33703 326866 33823 326994
rect 33903 326946 34833 354654
rect 34913 354593 35033 354734
rect 36123 354673 37213 354734
rect 34913 326866 35033 326994
rect 35113 326946 36043 354654
rect 36123 354593 36243 354673
rect 37093 354593 37213 354673
rect 36323 326994 37013 354593
rect 36123 326914 36243 326994
rect 37093 326914 37213 326994
rect 37293 326946 38223 354654
rect 38303 354593 38423 354734
rect 36123 326866 37213 326914
rect 38303 326866 38423 326994
rect 38503 326946 39593 354654
rect 39673 354593 39893 354734
rect 677707 341066 677927 341207
rect 678007 341146 679097 370854
rect 679177 370806 679297 370934
rect 680387 370886 681477 370934
rect 679177 341066 679297 341207
rect 679377 341146 680307 370854
rect 680387 370806 680507 370886
rect 681357 370806 681477 370886
rect 680587 341207 681277 370806
rect 680387 341127 680507 341207
rect 681357 341127 681477 341207
rect 681557 341146 682487 370854
rect 682567 370806 682687 370934
rect 680387 341066 681477 341127
rect 682567 341066 682687 341207
rect 682767 341146 683697 370854
rect 683777 370806 683897 370934
rect 683777 341066 683897 341207
rect 683977 341146 684667 370854
rect 684747 370806 684867 370934
rect 684747 341066 684867 341207
rect 684947 341146 685637 370854
rect 685717 370806 685837 370934
rect 685717 341066 685837 341207
rect 685917 341146 686847 370854
rect 686927 370806 687067 370934
rect 686927 341066 687067 341207
rect 677707 340798 687067 341066
rect 687147 340878 687213 377182
rect 687273 376171 687869 552907
rect 687949 548134 688145 552987
rect 687929 547800 688165 548054
rect 687949 518800 688145 547800
rect 687929 518546 688165 518800
rect 687949 504134 688145 518466
rect 687929 503800 688165 504054
rect 687949 474800 688145 503800
rect 687929 474546 688165 474800
rect 687949 460134 688145 474466
rect 687929 459800 688165 460054
rect 687949 430600 688145 459800
rect 687929 430346 688165 430600
rect 687949 415934 688145 430266
rect 687929 415600 688165 415854
rect 687949 386600 688145 415600
rect 687929 386346 688165 386600
rect 687949 379232 688145 386266
rect 688225 379312 688821 556048
rect 688901 554462 717600 556128
rect 688881 430346 688947 554382
rect 689027 548134 717600 554462
rect 689027 548006 689167 548134
rect 689027 518800 689167 547800
rect 689027 518466 689167 518607
rect 689247 518546 690137 548054
rect 690217 548006 690337 548134
rect 690217 518800 690337 547800
rect 690217 518466 690337 518607
rect 690417 518546 691307 548054
rect 691387 548006 691527 548134
rect 691607 547800 696600 548054
rect 696680 548006 712677 548134
rect 712757 547800 717600 548054
rect 691387 518800 697007 547800
rect 712407 518800 717600 547800
rect 691387 518466 691527 518607
rect 691607 518546 696600 518800
rect 696680 518466 712677 518607
rect 712757 518546 717600 518800
rect 689027 504134 717600 518466
rect 689027 503993 689167 504134
rect 689027 474800 689167 503800
rect 689027 474466 689167 474607
rect 689247 474546 690137 504054
rect 690217 503993 690337 504134
rect 690217 474800 690337 503800
rect 690217 474466 690337 474607
rect 690417 474546 691307 504054
rect 691387 503993 691527 504134
rect 691607 503800 696600 504054
rect 696680 503993 712677 504134
rect 712757 503800 717600 504054
rect 691387 474800 697007 503800
rect 712407 474800 717600 503800
rect 691387 474466 691527 474607
rect 691607 474546 696600 474800
rect 696680 474466 712677 474607
rect 712757 474546 717600 474800
rect 689027 460134 717600 474466
rect 689027 430600 689167 460134
rect 689027 430266 689167 430407
rect 689247 430346 690137 460054
rect 690217 459800 690337 460134
rect 690217 430600 690337 459600
rect 690217 430266 690337 430407
rect 690417 430346 691307 460054
rect 691387 459800 691527 460134
rect 691607 459800 696600 460054
rect 696680 459800 712677 460134
rect 712757 459800 717600 460054
rect 691387 430600 697007 459800
rect 712407 430600 717600 459800
rect 691387 430266 691527 430407
rect 691607 430346 696600 430600
rect 696680 430266 712677 430407
rect 712757 430346 717600 430600
rect 688901 415934 717600 430266
rect 688881 386078 688947 415854
rect 689027 415793 689167 415934
rect 689027 386600 689167 415600
rect 689027 386266 689167 386407
rect 689247 386346 690137 415854
rect 690217 415793 690337 415934
rect 690217 386600 690337 415600
rect 690217 386266 690337 386407
rect 690417 386346 691307 415854
rect 691387 415793 691527 415934
rect 691607 415600 696600 415854
rect 696680 415793 712677 415934
rect 712757 415600 717600 415854
rect 691387 386600 697007 415600
rect 712407 386600 717600 415600
rect 691387 386266 691527 386407
rect 691607 386346 696600 386600
rect 696680 386266 712677 386407
rect 712757 386346 717600 386600
rect 689027 385998 717600 386266
rect 688901 379232 717600 385998
rect 687949 378928 717600 379232
rect 687949 376091 688145 378928
rect 687293 375787 688145 376091
rect 677707 332062 687193 340798
rect 39673 326866 39893 326994
rect 30533 320538 39893 326866
rect 677707 325734 687067 332062
rect 677707 325606 677927 325734
rect 30407 311802 39893 320538
rect 29455 278509 30307 278813
rect 29455 275672 29651 278509
rect 0 275368 29651 275672
rect 0 268602 28699 275368
rect 0 268334 28573 268602
rect 0 268000 4843 268254
rect 4923 268193 20920 268334
rect 21000 268000 25993 268254
rect 26073 268193 26213 268334
rect 0 240800 5193 268000
rect 20593 240800 26213 268000
rect 0 240546 4843 240800
rect 4923 240466 20920 240594
rect 21000 240546 25993 240800
rect 26073 240466 26213 240594
rect 26293 240546 27183 268254
rect 27263 268193 27383 268334
rect 27263 240800 27383 267800
rect 27263 240466 27383 240594
rect 27463 240546 28353 268254
rect 28433 268193 28573 268334
rect 28433 240800 28573 268000
rect 28433 240466 28573 240594
rect 0 234138 28573 240466
rect 28653 234218 28719 268522
rect 0 232472 28699 234138
rect 28779 232552 29375 275288
rect 29455 268334 29651 275368
rect 29435 268000 29671 268254
rect 29455 240800 29651 268000
rect 29435 240546 29671 240800
rect 29455 235613 29651 240466
rect 29731 235693 30327 278429
rect 30387 277418 30453 311722
rect 30533 311534 39893 311802
rect 30533 311393 30673 311534
rect 30533 283666 30673 283794
rect 30753 283746 31683 311454
rect 31763 311393 31883 311534
rect 31763 283666 31883 283794
rect 31963 283746 32653 311454
rect 32733 311393 32853 311534
rect 32733 283666 32853 283794
rect 32933 283746 33623 311454
rect 33703 311393 33823 311534
rect 33703 283666 33823 283794
rect 33903 283746 34833 311454
rect 34913 311393 35033 311534
rect 36123 311473 37213 311534
rect 34913 283666 35033 283794
rect 35113 283746 36043 311454
rect 36123 311393 36243 311473
rect 37093 311393 37213 311473
rect 36323 283794 37013 311393
rect 36123 283714 36243 283794
rect 37093 283714 37213 283794
rect 37293 283746 38223 311454
rect 38303 311393 38423 311534
rect 36123 283666 37213 283714
rect 38303 283666 38423 283794
rect 38503 283746 39593 311454
rect 39673 311393 39893 311534
rect 677707 296066 677927 296207
rect 678007 296146 679097 325654
rect 679177 325606 679297 325734
rect 680387 325686 681477 325734
rect 679177 296066 679297 296207
rect 679377 296146 680307 325654
rect 680387 325606 680507 325686
rect 681357 325606 681477 325686
rect 680587 296207 681277 325606
rect 680387 296127 680507 296207
rect 681357 296127 681477 296207
rect 681557 296146 682487 325654
rect 682567 325606 682687 325734
rect 680387 296066 681477 296127
rect 682567 296066 682687 296207
rect 682767 296146 683697 325654
rect 683777 325606 683897 325734
rect 683777 296066 683897 296207
rect 683977 296146 684667 325654
rect 684747 325606 684867 325734
rect 684747 296066 684867 296207
rect 684947 296146 685637 325654
rect 685717 325606 685837 325734
rect 685717 296066 685837 296207
rect 685917 296146 686847 325654
rect 686927 325606 687067 325734
rect 686927 296066 687067 296207
rect 677707 295798 687067 296066
rect 687147 295878 687213 331982
rect 687273 330971 687869 375707
rect 687949 370934 688145 375787
rect 687929 370600 688165 370854
rect 687949 341400 688145 370600
rect 687929 341146 688165 341400
rect 687949 334032 688145 341066
rect 688225 334112 688821 378848
rect 688901 377262 717600 378928
rect 688881 340878 688947 377182
rect 689027 370934 717600 377262
rect 689027 370806 689167 370934
rect 689027 341400 689167 370600
rect 689027 341066 689167 341207
rect 689247 341146 690137 370854
rect 690217 370806 690337 370934
rect 690217 341400 690337 370400
rect 690217 341066 690337 341207
rect 690417 341146 691307 370854
rect 691387 370806 691527 370934
rect 691607 370600 696600 370854
rect 696680 370806 712677 370934
rect 712757 370600 717600 370854
rect 691387 341400 697007 370600
rect 712407 341400 717600 370600
rect 691387 341066 691527 341207
rect 691607 341146 696600 341400
rect 696680 341066 712677 341207
rect 712757 341146 717600 341400
rect 689027 340798 717600 341066
rect 688901 334032 717600 340798
rect 687949 333728 717600 334032
rect 687949 330891 688145 333728
rect 687293 330587 688145 330891
rect 677707 287062 687193 295798
rect 39673 283666 39893 283794
rect 30533 277338 39893 283666
rect 677707 280734 687067 287062
rect 677707 280606 677927 280734
rect 30407 268602 39893 277338
rect 29455 235309 30307 235613
rect 29455 232472 29651 235309
rect 0 232168 29651 232472
rect 0 225402 28699 232168
rect 0 225134 28573 225402
rect 0 224800 4843 225054
rect 4923 224993 20920 225134
rect 21000 224800 25993 225054
rect 26073 224993 26213 225134
rect 0 197600 5193 224800
rect 20593 197600 26213 224800
rect 0 197346 4843 197600
rect 4923 197266 20920 197394
rect 21000 197346 25993 197600
rect 26073 197266 26213 197394
rect 26293 197346 27183 225054
rect 27263 224993 27383 225134
rect 27263 197600 27383 224600
rect 27263 197266 27383 197394
rect 27463 197346 28353 225054
rect 28433 224993 28573 225134
rect 28433 197600 28573 224800
rect 28433 197266 28573 197394
rect 0 190938 28573 197266
rect 28653 191018 28719 225322
rect 0 189272 28699 190938
rect 28779 189352 29375 232088
rect 29455 225134 29651 232168
rect 29435 224800 29671 225054
rect 29455 197600 29651 224800
rect 29435 197346 29671 197600
rect 29455 192413 29651 197266
rect 29731 192493 30327 235229
rect 30387 234218 30453 268522
rect 30533 268334 39893 268602
rect 30533 268193 30673 268334
rect 30533 240466 30673 240594
rect 30753 240546 31683 268254
rect 31763 268193 31883 268334
rect 31763 240466 31883 240594
rect 31963 240546 32653 268254
rect 32733 268193 32853 268334
rect 32733 240466 32853 240594
rect 32933 240546 33623 268254
rect 33703 268193 33823 268334
rect 33703 240466 33823 240594
rect 33903 240546 34833 268254
rect 34913 268193 35033 268334
rect 36123 268273 37213 268334
rect 34913 240466 35033 240594
rect 35113 240546 36043 268254
rect 36123 268193 36243 268273
rect 37093 268193 37213 268273
rect 36323 240594 37013 268193
rect 36123 240514 36243 240594
rect 37093 240514 37213 240594
rect 37293 240546 38223 268254
rect 38303 268193 38423 268334
rect 36123 240466 37213 240514
rect 38303 240466 38423 240594
rect 38503 240546 39593 268254
rect 39673 268193 39893 268334
rect 677707 251066 677927 251207
rect 678007 251146 679097 280654
rect 679177 280606 679297 280734
rect 680387 280686 681477 280734
rect 679177 251066 679297 251207
rect 679377 251146 680307 280654
rect 680387 280606 680507 280686
rect 681357 280606 681477 280686
rect 680587 251207 681277 280606
rect 680387 251127 680507 251207
rect 681357 251127 681477 251207
rect 681557 251146 682487 280654
rect 682567 280606 682687 280734
rect 680387 251066 681477 251127
rect 682567 251066 682687 251207
rect 682767 251146 683697 280654
rect 683777 280606 683897 280734
rect 683777 251066 683897 251207
rect 683977 251146 684667 280654
rect 684747 280606 684867 280734
rect 684747 251066 684867 251207
rect 684947 251146 685637 280654
rect 685717 280606 685837 280734
rect 685717 251066 685837 251207
rect 685917 251146 686847 280654
rect 686927 280606 687067 280734
rect 686927 251066 687067 251207
rect 677707 250798 687067 251066
rect 687147 250878 687213 286982
rect 687273 285971 687869 330507
rect 687949 325734 688145 330587
rect 687929 325400 688165 325654
rect 687949 296400 688145 325400
rect 687929 296146 688165 296400
rect 687949 289032 688145 296066
rect 688225 289112 688821 333648
rect 688901 332062 717600 333728
rect 688881 295878 688947 331982
rect 689027 325734 717600 332062
rect 689027 325606 689167 325734
rect 689027 296400 689167 325400
rect 689027 296066 689167 296207
rect 689247 296146 690137 325654
rect 690217 325606 690337 325734
rect 690217 296400 690337 325400
rect 690217 296066 690337 296207
rect 690417 296146 691307 325654
rect 691387 325606 691527 325734
rect 691607 325400 696600 325654
rect 696680 325606 712677 325734
rect 712757 325400 717600 325654
rect 691387 296400 697007 325400
rect 712407 296400 717600 325400
rect 691387 296066 691527 296207
rect 691607 296146 696600 296400
rect 696680 296066 712677 296207
rect 712757 296146 717600 296400
rect 689027 295798 717600 296066
rect 688901 289032 717600 295798
rect 687949 288728 717600 289032
rect 687949 285891 688145 288728
rect 687293 285587 688145 285891
rect 677707 242062 687193 250798
rect 39673 240466 39893 240594
rect 30533 234138 39893 240466
rect 677707 235734 687067 242062
rect 677707 235606 677927 235734
rect 30407 225402 39893 234138
rect 29455 192109 30307 192413
rect 29455 189272 29651 192109
rect 0 188968 29651 189272
rect 0 182202 28699 188968
rect 0 181934 28573 182202
rect 0 181600 4843 181854
rect 4923 181793 20920 181934
rect 21000 181600 25993 181854
rect 26073 181793 26213 181934
rect 0 154400 5193 181600
rect 20593 154400 26213 181600
rect 0 152400 4843 154400
rect 21000 152400 25993 154400
rect 0 125200 5193 152400
rect 20593 125400 26213 152400
rect 20593 125200 21000 125400
rect 0 124946 4843 125200
rect 4923 124866 20920 125007
rect 25993 125200 26213 125400
rect 26073 124866 26213 125007
rect 26293 124946 27183 181854
rect 27263 181793 27383 181934
rect 27263 154400 27383 181400
rect 27263 125200 27383 152200
rect 27263 124866 27383 125007
rect 27463 124946 28353 181854
rect 28433 181793 28573 181934
rect 28433 154400 28573 181600
rect 28653 153400 28719 182122
rect 28433 125200 28573 152400
rect 28433 124866 28573 125007
rect 0 110534 28573 124866
rect 0 110200 4843 110454
rect 4923 110393 20920 110534
rect 0 83000 5193 110200
rect 20593 109800 21000 110200
rect 26073 110393 26213 110534
rect 25993 109800 26213 110200
rect 20593 83000 26213 109800
rect 0 82957 4850 83000
rect 0 82746 4843 82957
rect 4923 82666 20920 83000
rect 21000 82746 25993 83000
rect 26073 82666 26213 83000
rect 26293 82746 27183 110454
rect 27263 110393 27383 110534
rect 27263 82666 27383 110000
rect 27463 82746 28353 110454
rect 28433 110393 28573 110534
rect 28433 82666 28573 110200
rect 0 68334 28573 82666
rect 0 68000 4843 68254
rect 4923 68000 20920 68334
rect 21000 68000 25993 68254
rect 26073 68000 26213 68334
rect 0 40800 5193 68000
rect 20593 40800 26213 68000
rect 0 40546 4843 40800
rect 4923 40466 20920 40549
rect 0 40349 20920 40466
rect 21000 40429 25993 40800
rect 26073 40466 26213 40549
rect 26293 40546 27183 68254
rect 27263 68000 27383 68334
rect 27263 40800 27383 67800
rect 27263 40466 27383 40549
rect 27463 40546 28353 68254
rect 28433 40800 28573 68334
rect 28433 40466 28573 40549
rect 26073 40349 28573 40466
rect 0 35285 28573 40349
rect 28653 35365 28719 152400
rect 28779 35418 29375 188888
rect 29455 181934 29651 188968
rect 29435 181600 29671 181854
rect 29455 154400 29651 181600
rect 29435 153400 29671 154400
rect 29455 125200 29651 152400
rect 29435 124946 29671 125200
rect 29455 110534 29651 124866
rect 29435 110200 29671 110454
rect 29455 83000 29651 110200
rect 29435 82746 29671 83000
rect 29455 68334 29651 82666
rect 29435 68000 29671 68254
rect 29455 40800 29651 68000
rect 29435 36489 29671 40800
rect 29731 36625 30327 192029
rect 30387 191018 30453 225322
rect 30533 225134 39893 225402
rect 30533 224993 30673 225134
rect 30533 197266 30673 197394
rect 30753 197346 31683 225054
rect 31763 224993 31883 225134
rect 31763 197266 31883 197394
rect 31963 197346 32653 225054
rect 32733 224993 32853 225134
rect 32733 197266 32853 197394
rect 32933 197346 33623 225054
rect 33703 224993 33823 225134
rect 33703 197266 33823 197394
rect 33903 197346 34833 225054
rect 34913 224993 35033 225134
rect 36123 225073 37213 225134
rect 34913 197266 35033 197394
rect 35113 197346 36043 225054
rect 36123 224993 36243 225073
rect 37093 224993 37213 225073
rect 36323 197394 37013 224993
rect 36123 197314 36243 197394
rect 37093 197314 37213 197394
rect 37293 197346 38223 225054
rect 38303 224993 38423 225134
rect 36123 197266 37213 197314
rect 38303 197266 38423 197394
rect 38503 197346 39593 225054
rect 39673 224993 39893 225134
rect 677707 205866 677927 206007
rect 678007 205946 679097 235654
rect 679177 235606 679297 235734
rect 680387 235686 681477 235734
rect 679177 205866 679297 206007
rect 679377 205946 680307 235654
rect 680387 235606 680507 235686
rect 681357 235606 681477 235686
rect 680587 206007 681277 235606
rect 680387 205927 680507 206007
rect 681357 205927 681477 206007
rect 681557 205946 682487 235654
rect 682567 235606 682687 235734
rect 680387 205866 681477 205927
rect 682567 205866 682687 206007
rect 682767 205946 683697 235654
rect 683777 235606 683897 235734
rect 683777 205866 683897 206007
rect 683977 205946 684667 235654
rect 684747 235606 684867 235734
rect 684747 205866 684867 206007
rect 684947 205946 685637 235654
rect 685717 235606 685837 235734
rect 685717 205866 685837 206007
rect 685917 205946 686847 235654
rect 686927 235606 687067 235734
rect 686927 205866 687067 206007
rect 677707 205598 687067 205866
rect 687147 205678 687213 241982
rect 687273 240971 687869 285507
rect 687949 280734 688145 285587
rect 687929 280400 688165 280654
rect 687949 251400 688145 280400
rect 687929 251146 688165 251400
rect 687949 244032 688145 251066
rect 688225 244112 688821 288648
rect 688901 287062 717600 288728
rect 688881 250878 688947 286982
rect 689027 280734 717600 287062
rect 689027 280606 689167 280734
rect 689027 251400 689167 280400
rect 689027 251066 689167 251207
rect 689247 251146 690137 280654
rect 690217 280606 690337 280734
rect 690217 251400 690337 280400
rect 690217 251066 690337 251207
rect 690417 251146 691307 280654
rect 691387 280606 691527 280734
rect 691607 280400 696600 280654
rect 696680 280606 712677 280734
rect 712757 280400 717600 280654
rect 691387 251400 697007 280400
rect 712407 251400 717600 280400
rect 691387 251066 691527 251207
rect 691607 251146 696600 251400
rect 696680 251066 712677 251207
rect 712757 251146 717600 251400
rect 689027 250798 717600 251066
rect 688901 244032 717600 250798
rect 687949 243728 717600 244032
rect 687949 240891 688145 243728
rect 687293 240587 688145 240891
rect 39673 197266 39893 197394
rect 30533 190938 39893 197266
rect 30407 182202 39893 190938
rect 677707 196862 687193 205598
rect 677707 190534 687067 196862
rect 677707 190406 677927 190534
rect 30387 153400 30453 182122
rect 30533 181934 39893 182202
rect 30533 181793 30673 181934
rect 30753 154400 31683 181854
rect 31763 181793 31883 181934
rect 31963 153400 32653 181854
rect 32733 181793 32853 181934
rect 29751 36409 30307 36545
rect 29455 36005 30307 36409
rect 30387 36085 30453 152400
rect 30533 124866 30673 125007
rect 30753 124946 31683 153400
rect 31763 124866 31883 125007
rect 31963 124946 32653 152400
rect 32733 124866 32853 125007
rect 32933 124946 33623 181854
rect 33703 181793 33823 181934
rect 33703 124866 33823 125007
rect 33903 124946 34833 181854
rect 34913 181793 35033 181934
rect 36123 181873 37213 181934
rect 34913 124866 35033 125007
rect 36123 181793 36243 181873
rect 37093 181793 37213 181873
rect 36323 153400 37013 181793
rect 37293 154400 38223 181854
rect 38303 181793 38423 181934
rect 36323 125007 37013 152400
rect 36123 124927 36243 125007
rect 37093 124927 37213 125007
rect 37293 124946 38223 153400
rect 36123 124866 37213 124927
rect 38303 124866 38423 125007
rect 38503 124946 39593 181854
rect 39673 181793 39893 181934
rect 677707 160866 677927 161007
rect 678007 160946 679097 190454
rect 679177 190406 679297 190534
rect 680387 190486 681477 190534
rect 679177 160866 679297 161007
rect 679377 160946 680307 190454
rect 680387 190406 680507 190486
rect 681357 190406 681477 190486
rect 680587 161007 681277 190406
rect 680387 160927 680507 161007
rect 681357 160927 681477 161007
rect 681557 160946 682487 190454
rect 682567 190406 682687 190534
rect 680387 160866 681477 160927
rect 682567 160866 682687 161007
rect 682767 160946 683697 190454
rect 683777 190406 683897 190534
rect 683777 160866 683897 161007
rect 683977 160946 684667 190454
rect 684747 190406 684867 190534
rect 684747 160866 684867 161007
rect 684947 160946 685637 190454
rect 685717 190406 685837 190534
rect 685717 160866 685837 161007
rect 685917 160946 686847 190454
rect 686927 190406 687067 190534
rect 686927 160866 687067 161007
rect 677707 160598 687067 160866
rect 687147 160678 687213 196782
rect 687273 195771 687869 240507
rect 687949 235734 688145 240587
rect 687929 235400 688165 235654
rect 687949 206200 688145 235400
rect 687929 205946 688165 206200
rect 687949 198832 688145 205866
rect 688225 198912 688821 243648
rect 688901 242062 717600 243728
rect 688881 205678 688947 241982
rect 689027 235734 717600 242062
rect 689027 235606 689167 235734
rect 689027 206200 689167 235400
rect 689027 205866 689167 206007
rect 689247 205946 690137 235654
rect 690217 235606 690337 235734
rect 690217 206200 690337 235200
rect 690217 205866 690337 206007
rect 690417 205946 691307 235654
rect 691387 235606 691527 235734
rect 691607 235400 696600 235654
rect 696680 235606 712677 235734
rect 712757 235400 717600 235654
rect 691387 206200 697007 235400
rect 712407 206200 717600 235400
rect 691387 205866 691527 206007
rect 691607 205946 696600 206200
rect 696680 205866 712677 206007
rect 712757 205946 717600 206200
rect 689027 205598 717600 205866
rect 688901 198832 717600 205598
rect 687949 198528 717600 198832
rect 687949 195691 688145 198528
rect 687293 195387 688145 195691
rect 677707 151862 687193 160598
rect 677707 145534 687067 151862
rect 677707 145406 677927 145534
rect 30533 110534 39593 124866
rect 677707 115666 677927 115807
rect 678007 115746 679097 145454
rect 679177 145406 679297 145534
rect 680387 145486 681477 145534
rect 679177 115666 679297 115807
rect 679377 115746 680307 145454
rect 680387 145406 680507 145486
rect 681357 145406 681477 145486
rect 680587 115807 681277 145406
rect 680387 115727 680507 115807
rect 681357 115727 681477 115807
rect 681557 115746 682487 145454
rect 682567 145406 682687 145534
rect 680387 115666 681477 115727
rect 682567 115666 682687 115807
rect 682767 115746 683697 145454
rect 683777 145406 683897 145534
rect 683777 115666 683897 115807
rect 683977 115746 684667 145454
rect 684747 145406 684867 145534
rect 684747 115666 684867 115807
rect 684947 115746 685637 145454
rect 685717 145406 685837 145534
rect 685717 115666 685837 115807
rect 685917 115746 686847 145454
rect 686927 145406 687067 145534
rect 686927 115666 687067 115807
rect 677707 115398 687067 115666
rect 687147 115478 687213 151782
rect 687273 150771 687869 195307
rect 687949 190534 688145 195387
rect 687929 190200 688165 190454
rect 687949 161200 688145 190200
rect 687929 160946 688165 161200
rect 687949 153832 688145 160866
rect 688225 153912 688821 198448
rect 688901 196862 717600 198528
rect 688881 160678 688947 196782
rect 689027 190534 717600 196862
rect 689027 190406 689167 190534
rect 689027 161200 689167 190200
rect 689027 160866 689167 161007
rect 689247 160946 690137 190454
rect 690217 190406 690337 190534
rect 690217 161200 690337 190200
rect 690217 160866 690337 161007
rect 690417 160946 691307 190454
rect 691387 190406 691527 190534
rect 691607 190200 696600 190454
rect 696680 190406 712677 190534
rect 712757 190200 717600 190454
rect 691387 161200 697007 190200
rect 712407 161200 717600 190200
rect 691387 160866 691527 161007
rect 691607 160946 696600 161200
rect 696680 160866 712677 161007
rect 712757 160946 717600 161200
rect 689027 160598 717600 160866
rect 688901 153832 717600 160598
rect 687949 153528 717600 153832
rect 687949 150691 688145 153528
rect 687293 150387 688145 150691
rect 30533 110393 30673 110534
rect 30533 82666 30673 83000
rect 30753 82746 31683 110454
rect 31763 110393 31883 110534
rect 31763 82666 31883 83000
rect 31963 82746 32653 110454
rect 32733 110393 32853 110534
rect 32733 82666 32853 83000
rect 32933 82746 33623 110454
rect 33703 110393 33823 110534
rect 33903 85187 34833 110454
rect 34913 110393 35033 110534
rect 36123 110473 37213 110534
rect 33703 82666 33823 83000
rect 33903 82987 34840 85187
rect 33903 82746 34833 82987
rect 34913 82666 35033 83000
rect 36123 110393 36243 110473
rect 37093 110393 37213 110473
rect 36123 82727 36243 83000
rect 36323 82807 37013 110393
rect 37093 82727 37213 83000
rect 38303 110393 38423 110534
rect 36123 82666 37213 82727
rect 38303 82666 38423 83000
rect 38503 82746 39593 110454
rect 677707 106662 687193 115398
rect 677707 100334 687067 106662
rect 677707 100206 677927 100334
rect 30533 68334 39593 82666
rect 30533 68000 30673 68334
rect 30753 68014 31683 68254
rect 30753 65805 31690 68014
rect 31763 68000 31883 68334
rect 30533 40466 30673 40549
rect 30753 40546 31683 65805
rect 31763 40466 31883 40549
rect 31963 40546 32653 68254
rect 32733 68000 32853 68334
rect 32733 40466 32853 40549
rect 32933 40546 33623 68254
rect 33703 68000 33823 68334
rect 33703 40466 33823 40549
rect 33903 40546 34833 68254
rect 34913 68000 35033 68334
rect 36123 68273 37213 68334
rect 34913 40466 35033 40549
rect 35113 40546 36043 68254
rect 36123 68000 36243 68273
rect 36323 40549 37013 68193
rect 37093 68000 37213 68273
rect 36123 40469 36243 40549
rect 37093 40469 37213 40549
rect 38303 68000 38423 68334
rect 36123 40466 37213 40469
rect 38303 40466 38423 40549
rect 38503 40546 39593 68254
rect 39673 40466 40000 40549
rect 30533 39673 40000 40466
rect 677051 39920 677927 40000
tri 677927 39920 678007 40000 se
rect 678007 39920 679097 100254
rect 679177 100206 679297 100334
rect 680387 100286 681477 100334
rect 679377 71000 680307 100254
rect 680387 100206 680507 100286
rect 681357 100206 681477 100286
rect 680587 70000 681277 100206
rect 186606 39673 202207 39893
rect 295206 39673 310807 39893
rect 350006 39673 365607 39893
rect 404806 39673 420407 39893
rect 459606 39673 475207 39893
rect 514406 39673 530007 39893
rect 677051 39673 679097 39920
rect 30533 38423 39450 39673
rect 39593 39593 39920 39673
tri 39920 39593 40000 39673 sw
rect 39530 38503 79054 39593
rect 79134 38423 93466 39593
rect 93546 38503 132854 39593
rect 132934 38423 147266 39593
rect 147346 38503 186654 39593
rect 186734 38423 202066 39673
rect 202146 38503 241454 39593
rect 241534 38423 255866 39593
rect 255946 38503 295254 39593
rect 295334 38423 310666 39673
rect 310746 38503 350054 39593
rect 350134 38423 365466 39673
rect 365546 38503 404854 39593
rect 404934 38423 420266 39673
rect 420346 38503 459654 39593
rect 459734 38423 475066 39673
rect 475146 38503 514454 39593
rect 514534 38423 529866 39673
rect 677134 39593 679097 39673
rect 529946 38503 569254 39593
rect 569334 38423 583666 39593
rect 583746 38503 623054 39593
rect 623134 38423 637466 39593
rect 637546 38503 677054 39593
rect 677134 39450 677927 39593
rect 678007 39530 679097 39593
rect 679177 39450 679297 40000
rect 677134 39163 679297 39450
rect 679377 39243 680307 70000
rect 680387 39626 680507 40000
rect 680587 39706 681277 69000
rect 681357 39626 681477 40000
rect 681557 39695 682487 100254
rect 682567 100206 682687 100334
rect 680387 39615 681477 39626
rect 682567 39615 682687 40000
rect 682767 39680 683697 100254
rect 683777 100206 683897 100334
rect 680387 39600 682687 39615
rect 683777 39643 683897 40000
rect 683977 39723 684667 100254
rect 684747 100206 684867 100334
rect 684947 70000 685637 100254
rect 685717 100206 685837 100334
rect 685917 71000 686847 100254
rect 686927 100206 687067 100334
rect 687147 70000 687213 106582
rect 687273 105571 687869 150307
rect 687949 145534 688145 150387
rect 687929 145200 688165 145454
rect 687949 116000 688145 145200
rect 687929 115746 688165 116000
rect 687949 108632 688145 115666
rect 688225 108712 688821 153448
rect 688901 151862 717600 153528
rect 688881 115478 688947 151782
rect 689027 145534 717600 151862
rect 689027 145406 689167 145534
rect 689027 116000 689167 145200
rect 689027 115666 689167 115807
rect 689247 115746 690137 145454
rect 690217 145406 690337 145534
rect 690217 116000 690337 145000
rect 690217 115666 690337 115807
rect 690417 115746 691307 145454
rect 691387 145406 691527 145534
rect 691607 145200 696600 145454
rect 696680 145406 712677 145534
rect 712757 145200 717600 145454
rect 691387 116000 697007 145200
rect 712407 116000 717600 145200
rect 691387 115666 691527 115807
rect 691607 115746 696600 116000
rect 696680 115666 712677 115807
rect 712757 115746 717600 116000
rect 689027 115398 717600 115666
rect 688901 108632 717600 115398
rect 687949 108328 717600 108632
rect 687949 105491 688145 108328
rect 687293 105187 688145 105491
rect 684747 39653 684867 40000
rect 684947 39733 685637 69000
rect 685717 39653 685837 40000
rect 685917 39705 686847 70000
rect 684747 39643 685837 39653
rect 683777 39625 685837 39643
rect 686927 39625 687067 40000
rect 683777 39600 687067 39625
rect 680387 39163 687067 39600
rect 677134 38423 687067 39163
rect 30533 38303 40000 38423
rect 78993 38303 93607 38423
rect 132793 38303 147407 38423
rect 186606 38303 202207 38423
rect 241200 38303 256200 38423
rect 295206 38303 310807 38423
rect 350006 38303 365607 38423
rect 404806 38303 420407 38423
rect 459606 38303 475207 38423
rect 514406 38303 530007 38423
rect 569193 38303 583807 38423
rect 622993 38303 637607 38423
rect 677051 38303 687067 38423
rect 30533 37213 39163 38303
rect 39243 37293 79054 38223
rect 79134 37213 93466 38303
rect 93546 37293 132854 38223
rect 132934 37213 147266 38303
rect 147346 37293 186654 38223
rect 186734 37213 202066 38303
rect 202146 37293 241454 38223
rect 241534 37213 255866 38303
rect 255946 37293 295254 38223
rect 295334 37213 310666 38303
rect 310746 37293 350054 38223
rect 350134 37213 365466 38303
rect 365546 37293 404854 38223
rect 404934 37213 420266 38303
rect 420346 37293 459654 38223
rect 459734 37213 475066 38303
rect 475146 37293 514454 38223
rect 514534 37213 529866 38303
rect 529946 37293 569254 38223
rect 569334 37213 583666 38303
rect 583746 37293 623054 38223
rect 623134 37213 637466 38303
rect 637546 37293 677054 38223
rect 677134 37213 687067 38303
rect 30533 37093 40000 37213
rect 78993 37093 93607 37213
rect 132793 37093 147407 37213
rect 186606 37093 202207 37213
rect 241200 37093 256200 37213
rect 295206 37093 310807 37213
rect 350006 37093 365607 37213
rect 404806 37093 420407 37213
rect 459606 37093 475207 37213
rect 514406 37093 530007 37213
rect 569193 37093 583807 37213
rect 622993 37093 637607 37213
rect 677051 37093 687067 37213
rect 30533 36243 39626 37093
rect 39706 36323 78993 37013
rect 79073 36243 93527 37093
rect 93607 36323 132793 37013
rect 132873 36243 147327 37093
rect 147407 36323 186606 37013
rect 186686 36243 202127 37093
rect 202207 36323 241393 37013
rect 241473 36243 255927 37093
rect 256007 36323 295206 37013
rect 295286 36243 310727 37093
rect 310807 36323 350006 37013
rect 350086 36243 365527 37093
rect 365607 36323 404806 37013
rect 404886 36243 420327 37093
rect 420407 36323 459606 37013
rect 459686 36243 475127 37093
rect 475207 36323 514406 37013
rect 514486 36243 529927 37093
rect 530007 36323 569193 37013
rect 569273 36243 583727 37093
rect 623073 36243 637527 37093
rect 677131 36243 687067 37093
rect 30533 36123 40000 36243
rect 78993 36123 93607 36243
rect 132793 36123 147407 36243
rect 186606 36123 202207 36243
rect 241200 36123 256200 36243
rect 295206 36123 310807 36243
rect 350006 36123 365607 36243
rect 404806 36123 420407 36243
rect 459606 36123 475207 36243
rect 514406 36123 530007 36243
rect 569193 36123 583807 36243
rect 622993 36123 637607 36243
rect 677051 36123 687067 36243
rect 30533 36005 39615 36123
rect 29455 35338 39615 36005
rect 28799 35285 39615 35338
rect 0 35033 39615 35285
rect 39695 35113 79054 36043
rect 79134 35033 93466 36123
rect 93546 35113 132854 36043
rect 132934 35033 147266 36123
rect 147346 35113 186654 36043
rect 186734 35033 202066 36123
rect 202146 35113 241454 36043
rect 241534 35033 255866 36123
rect 255946 35113 295254 36043
rect 295334 35033 310666 36123
rect 310746 35113 350054 36043
rect 350134 35033 365466 36123
rect 365546 35113 404854 36043
rect 404934 35033 420266 36123
rect 420346 35113 459654 36043
rect 459734 35033 475066 36123
rect 475146 35113 514454 36043
rect 514534 35033 529866 36123
rect 529946 35113 569254 36043
rect 569334 35033 583666 36123
rect 583746 35113 623054 36043
rect 623134 35033 637466 36123
rect 637546 35113 677054 36043
rect 677134 36005 687067 36123
rect 687147 36085 687213 69000
rect 677134 35733 687193 36005
rect 687273 35813 687869 105107
rect 687949 100334 688145 105187
rect 687929 100000 688165 100254
rect 687949 71000 688145 100000
rect 687929 70000 688165 71000
rect 687949 40000 688145 69000
rect 677134 35610 687849 35733
rect 687929 35690 688165 40000
rect 677134 35338 688145 35610
rect 688225 35418 688821 108248
rect 688901 106662 717600 108328
rect 688881 70000 688947 106582
rect 689027 100334 717600 106662
rect 689027 100206 689167 100334
rect 689027 71000 689167 100000
rect 688881 35365 688947 69000
rect 689027 39595 689167 69000
rect 689247 39675 690137 100254
rect 690217 100206 690337 100334
rect 690217 71000 690337 100000
rect 690217 39624 690337 69000
rect 690417 39704 691307 100254
rect 691387 100206 691527 100334
rect 691607 100000 696600 100254
rect 696680 100206 712677 100334
rect 712757 100000 717600 100254
rect 691387 71000 697007 100000
rect 712407 71000 717600 100000
rect 691607 69000 696600 71000
rect 712757 69000 717600 71000
rect 691387 40000 697007 69000
rect 712407 40000 717600 69000
rect 691387 39624 691527 40000
rect 690217 39595 691527 39624
rect 689027 39391 691527 39595
rect 691607 39471 696600 40000
rect 696680 39633 712677 40000
rect 712757 39713 717600 40000
rect 696680 39391 717600 39633
rect 677134 35285 688801 35338
rect 689027 35285 717600 39391
rect 677134 35033 717600 35285
rect 0 34913 40000 35033
rect 78993 34913 93607 35033
rect 132793 34913 147407 35033
rect 186606 34913 202207 35033
rect 241200 34913 256200 35033
rect 295206 34913 310807 35033
rect 350006 34913 365607 35033
rect 404806 34913 420407 35033
rect 459606 34913 475207 35033
rect 514406 34913 530007 35033
rect 569193 34913 583807 35033
rect 622993 34913 637607 35033
rect 677051 34913 717600 35033
rect 0 33823 39600 34913
rect 39680 33903 79054 34833
rect 79134 33823 93466 34913
rect 93546 33903 132854 34833
rect 132934 33823 147266 34913
rect 147346 33903 186654 34833
rect 186734 33823 202066 34913
rect 239013 34833 241213 34840
rect 202146 33903 241454 34833
rect 241534 33823 255866 34913
rect 255946 33903 295254 34833
rect 295334 33823 310666 34913
rect 310746 33903 350054 34833
rect 350134 33823 365466 34913
rect 365546 33903 404854 34833
rect 404934 33823 420266 34913
rect 420346 33903 459654 34833
rect 459734 33823 475066 34913
rect 475146 33903 514454 34833
rect 514534 33823 529866 34913
rect 529946 33903 569254 34833
rect 569334 33823 583666 34913
rect 583746 33903 623054 34833
rect 623134 33823 637466 34913
rect 637546 33903 677054 34833
rect 677134 33823 717600 34913
rect 0 33703 40000 33823
rect 78993 33703 93607 33823
rect 132793 33703 147407 33823
rect 186606 33703 202207 33823
rect 241200 33703 256200 33823
rect 295206 33703 310807 33823
rect 350006 33703 365607 33823
rect 404806 33703 420407 33823
rect 459606 33703 475207 33823
rect 514406 33703 530007 33823
rect 569193 33703 583807 33823
rect 622993 33703 637607 33823
rect 677051 33703 717600 33823
rect 0 32853 39643 33703
rect 39723 32933 79054 33623
rect 79134 32853 93466 33703
rect 93546 32933 132854 33623
rect 132934 32853 147266 33703
rect 147346 32933 186654 33623
rect 186734 32853 202066 33703
rect 202146 32933 241454 33623
rect 241534 32853 255866 33703
rect 255946 32933 295254 33623
rect 295334 32853 310666 33703
rect 310746 32933 350054 33623
rect 350134 32853 365466 33703
rect 365546 32933 404854 33623
rect 404934 32853 420266 33703
rect 420346 32933 459654 33623
rect 459734 32853 475066 33703
rect 475146 32933 514454 33623
rect 514534 32853 529866 33703
rect 529946 32933 569254 33623
rect 569334 32853 583666 33703
rect 583746 32933 623054 33623
rect 623134 32853 637466 33703
rect 637546 32933 677054 33623
rect 677134 32853 717600 33703
rect 0 32733 40000 32853
rect 78993 32733 93607 32853
rect 132793 32733 147407 32853
rect 186606 32733 202207 32853
rect 241200 32733 256200 32853
rect 295206 32733 310807 32853
rect 350006 32733 365607 32853
rect 404806 32733 420407 32853
rect 459606 32733 475207 32853
rect 514406 32733 530007 32853
rect 569193 32733 583807 32853
rect 622993 32733 637607 32853
rect 677051 32733 717600 32853
rect 0 31883 39653 32733
rect 79134 31883 93466 32733
rect 132934 31883 147266 32733
rect 147346 31963 186654 32653
rect 186734 31883 202066 32733
rect 202146 31963 241454 32653
rect 241534 31883 255866 32733
rect 255946 31963 295254 32653
rect 295334 31883 310666 32733
rect 310746 31963 350054 32653
rect 350134 31883 365466 32733
rect 365546 31963 404854 32653
rect 404934 31883 420266 32733
rect 420346 31963 459654 32653
rect 459734 31883 475066 32733
rect 475146 31963 514454 32653
rect 514534 31883 529866 32733
rect 529946 31963 569254 32653
rect 569334 31883 583666 32733
rect 583746 31963 623054 32653
rect 623134 31883 637466 32733
rect 637546 31963 677054 32653
rect 677134 31883 717600 32733
rect 0 31763 40000 31883
rect 78993 31763 93607 31883
rect 132793 31763 147407 31883
rect 186606 31763 202207 31883
rect 241200 31763 256200 31883
rect 295206 31763 310807 31883
rect 350006 31763 365607 31883
rect 404806 31763 420407 31883
rect 459606 31763 475207 31883
rect 514406 31763 530007 31883
rect 569193 31763 583807 31883
rect 622993 31763 637607 31883
rect 677051 31763 717600 31883
rect 0 30673 39625 31763
rect 39705 30753 79054 31683
rect 79134 30673 93466 31763
rect 132934 31754 147266 31763
rect 93546 31674 132854 31683
rect 93546 30762 132869 31674
rect 93546 30753 132854 30762
rect 132949 30682 147266 31754
rect 147346 30753 186654 31683
rect 132934 30673 147266 30682
rect 186734 30673 202066 31763
rect 241534 30673 255866 31763
rect 256186 31683 258395 31690
rect 295334 30673 310666 31763
rect 310746 30753 350054 31683
rect 350134 30673 365466 31763
rect 365546 30753 404854 31683
rect 404934 30673 420266 31763
rect 420346 30753 459654 31683
rect 459734 30673 475066 31763
rect 475146 30753 514454 31683
rect 514534 30673 529866 31763
rect 529946 30753 569254 31683
rect 569334 30673 583666 31763
rect 583746 30753 623054 31683
rect 623134 30673 637466 31763
rect 637546 30753 677054 31683
rect 677134 30673 717600 31763
rect 0 30533 40000 30673
rect 78993 30533 93607 30673
rect 132793 30533 147407 30673
rect 186606 30533 202207 30673
rect 241200 30533 256200 30673
rect 295206 30533 310807 30673
rect 350006 30533 365607 30673
rect 404806 30533 420407 30673
rect 459606 30533 475207 30673
rect 514406 30533 530007 30673
rect 569193 30533 583807 30673
rect 622993 30533 637607 30673
rect 677051 30533 717600 30673
rect 0 30407 36005 30533
rect 0 29751 35733 30407
rect 79134 30407 93466 30533
rect 193062 30407 201798 30533
rect 201878 30387 301582 30453
rect 301662 30407 310398 30533
rect 310478 30387 356382 30453
rect 356462 30407 365198 30533
rect 365278 30387 411182 30453
rect 411262 30407 419998 30533
rect 420078 30387 465982 30453
rect 466062 30407 474798 30533
rect 474878 30387 520782 30453
rect 520862 30407 529598 30533
rect 529678 30387 681515 30453
rect 0 29455 35610 29751
rect 35813 29731 191507 30327
rect 35690 29651 40000 29671
rect 47400 29651 71400 29671
rect 35690 29455 78800 29651
rect 0 28799 35338 29455
rect 35690 29435 40000 29455
rect 47400 29435 71400 29455
rect 79134 29455 93466 29651
rect 101200 29651 125200 29671
rect 132600 29651 132854 29671
rect 147346 29651 147600 29671
rect 155000 29651 179000 29671
rect 186400 29651 186654 29671
rect 191587 29651 191891 30307
rect 191971 29731 300107 30327
rect 202146 29651 202400 29671
rect 209800 29651 233800 29671
rect 241200 29651 241454 29671
rect 255946 29651 256200 29671
rect 263600 29651 287600 29671
rect 295000 29651 295254 29671
rect 300187 29651 300491 30307
rect 300571 29731 354907 30327
rect 310746 29651 311000 29671
rect 318400 29651 342400 29671
rect 349800 29651 350054 29671
rect 354987 29651 355291 30307
rect 355371 29731 409707 30327
rect 365546 29651 365800 29671
rect 373200 29651 397200 29671
rect 404600 29651 404854 29671
rect 409787 29651 410091 30307
rect 410171 29731 464507 30327
rect 420346 29651 420600 29671
rect 428000 29651 452000 29671
rect 459400 29651 459654 29671
rect 464587 29651 464891 30307
rect 464971 29731 519307 30327
rect 475146 29651 475400 29671
rect 482800 29651 506800 29671
rect 514200 29651 514454 29671
rect 519387 29651 519691 30307
rect 519771 29731 680975 30327
rect 681595 30307 717600 30533
rect 681055 29751 717600 30307
rect 529946 29651 530200 29671
rect 537600 29651 561600 29671
rect 569000 29651 569254 29671
rect 583746 29651 584000 29671
rect 591400 29651 615400 29671
rect 622800 29651 623054 29671
rect 637546 29651 637800 29671
rect 645200 29651 669200 29671
rect 676800 29651 681111 29671
rect 93800 29455 132854 29651
rect 132934 29455 147266 29651
rect 147346 29455 186654 29651
rect 186734 29455 202066 29651
rect 202146 29455 241454 29651
rect 241534 29455 255866 29651
rect 255946 29455 295254 29651
rect 295334 29455 310666 29651
rect 310746 29455 350054 29651
rect 350134 29455 365466 29651
rect 365546 29455 404854 29651
rect 404934 29455 420266 29651
rect 420346 29455 459654 29651
rect 459734 29455 475066 29651
rect 475146 29455 514454 29651
rect 514534 29455 529866 29651
rect 529946 29455 569254 29651
rect 569334 29455 583666 29651
rect 583746 29455 623054 29651
rect 623134 29455 637466 29651
rect 637546 29455 681111 29651
rect 681191 29455 717600 29751
rect 101200 29435 125200 29455
rect 132600 29435 132854 29455
rect 147346 29435 147600 29455
rect 155000 29435 179000 29455
rect 186400 29435 186654 29455
rect 0 28573 35285 28799
rect 35418 28779 194648 29375
rect 79134 28573 93466 28699
rect 194728 28699 195032 29455
rect 202146 29435 202400 29455
rect 209800 29435 233800 29455
rect 241200 29435 241454 29455
rect 255946 29435 256200 29455
rect 263600 29435 287600 29455
rect 295000 29435 295254 29455
rect 195112 28779 303248 29375
rect 193062 28573 201798 28699
rect 201878 28653 301582 28719
rect 303328 28699 303632 29455
rect 310746 29435 311000 29455
rect 318400 29435 342400 29455
rect 349800 29435 350054 29455
rect 303712 28779 358048 29375
rect 301662 28573 310398 28699
rect 310478 28653 356382 28719
rect 358128 28699 358432 29455
rect 365546 29435 365800 29455
rect 373200 29435 397200 29455
rect 404600 29435 404854 29455
rect 358512 28779 412848 29375
rect 356462 28573 365198 28699
rect 365278 28653 411182 28719
rect 412928 28699 413232 29455
rect 420346 29435 420600 29455
rect 428000 29435 452000 29455
rect 459400 29435 459654 29455
rect 413312 28779 467648 29375
rect 411262 28573 419998 28699
rect 420078 28653 465982 28719
rect 467728 28699 468032 29455
rect 475146 29435 475400 29455
rect 482800 29435 506800 29455
rect 514200 29435 514454 29455
rect 468112 28779 522448 29375
rect 466062 28573 474798 28699
rect 474878 28653 520782 28719
rect 522528 28699 522832 29455
rect 529946 29435 530200 29455
rect 537600 29435 561600 29455
rect 569000 29435 569254 29455
rect 583746 29435 584000 29455
rect 591400 29435 615400 29455
rect 622800 29435 623054 29455
rect 637546 29435 637800 29455
rect 645200 29435 669200 29455
rect 676800 29435 681111 29455
rect 522912 28779 682182 29375
rect 682262 28799 717600 29455
rect 520862 28573 529598 28699
rect 529678 28653 682235 28719
rect 682315 28573 717600 28799
rect 0 28433 47400 28573
rect 71400 28433 78800 28573
rect 78993 28433 93607 28573
rect 93800 28433 101200 28573
rect 125200 28433 132600 28573
rect 132793 28433 147407 28573
rect 147600 28433 155000 28573
rect 179000 28433 186400 28573
rect 186606 28433 202207 28573
rect 202400 28433 209800 28573
rect 233800 28433 263600 28573
rect 287600 28433 295000 28573
rect 295206 28433 310807 28573
rect 311000 28433 318400 28573
rect 342400 28433 349800 28573
rect 350006 28433 365607 28573
rect 365800 28433 373200 28573
rect 397200 28433 404600 28573
rect 404806 28433 420407 28573
rect 420600 28433 428000 28573
rect 452000 28433 459400 28573
rect 459606 28433 475207 28573
rect 475400 28433 482800 28573
rect 506800 28433 514200 28573
rect 514406 28433 530007 28573
rect 530200 28433 537600 28573
rect 561600 28433 569000 28573
rect 569193 28433 583807 28573
rect 584000 28433 591400 28573
rect 615400 28433 622800 28573
rect 622993 28433 637607 28573
rect 637800 28433 645200 28573
rect 669200 28433 676800 28573
rect 677051 28433 717600 28573
rect 0 27383 39595 28433
rect 39675 27463 79054 28353
rect 79134 27383 93466 28433
rect 93546 27463 132854 28353
rect 132934 27383 147266 28433
rect 147346 27463 186654 28353
rect 186734 27383 202066 28433
rect 202146 27463 241454 28353
rect 241534 27383 255866 28433
rect 255946 27463 295254 28353
rect 295334 27383 310666 28433
rect 310746 27463 350054 28353
rect 350134 27383 365466 28433
rect 365546 27463 404854 28353
rect 404934 27383 420266 28433
rect 420346 27463 459654 28353
rect 459734 27383 475066 28433
rect 475146 27463 514454 28353
rect 514534 27383 529866 28433
rect 529946 27463 569254 28353
rect 569334 27383 583666 28433
rect 583746 27463 623054 28353
rect 623134 27383 637466 28433
rect 637546 27463 677054 28353
rect 677134 27383 717600 28433
rect 0 27263 47000 27383
rect 71400 27263 78400 27383
rect 78993 27263 93607 27383
rect 93800 27263 100800 27383
rect 125200 27263 132200 27383
rect 132793 27263 147407 27383
rect 147600 27263 154600 27383
rect 179000 27263 186000 27383
rect 186606 27263 202207 27383
rect 202400 27263 209400 27383
rect 233800 27263 240800 27383
rect 241200 27263 263200 27383
rect 287600 27263 294600 27383
rect 295206 27263 310807 27383
rect 311000 27263 318000 27383
rect 342400 27263 349400 27383
rect 350006 27263 365607 27383
rect 365800 27263 372800 27383
rect 397200 27263 404200 27383
rect 404806 27263 420407 27383
rect 420600 27263 427600 27383
rect 452000 27263 459000 27383
rect 459606 27263 475207 27383
rect 475400 27263 482400 27383
rect 506800 27263 513800 27383
rect 514406 27263 530007 27383
rect 530200 27263 537200 27383
rect 561600 27263 568600 27383
rect 569193 27263 583807 27383
rect 584000 27263 591000 27383
rect 615400 27263 622400 27383
rect 622993 27263 637607 27383
rect 637800 27263 644800 27383
rect 669200 27263 676200 27383
rect 677051 27263 717600 27383
rect 0 26213 39624 27263
rect 39704 26293 79054 27183
rect 79134 26213 93466 27263
rect 93546 26293 132854 27183
rect 132934 26213 147266 27263
rect 147346 26293 186654 27183
rect 186734 26213 202066 27263
rect 202146 26293 241454 27183
rect 241534 26213 255866 27263
rect 255946 26293 295254 27183
rect 295334 26213 310666 27263
rect 310746 26293 350054 27183
rect 350134 26213 365466 27263
rect 365546 26293 404854 27183
rect 404934 26213 420266 27263
rect 420346 26293 459654 27183
rect 459734 26213 475066 27263
rect 475146 26293 514454 27183
rect 514534 26213 529866 27263
rect 529946 26293 569254 27183
rect 569334 26213 583666 27263
rect 583746 26293 623054 27183
rect 623134 26213 637466 27263
rect 637546 26293 677054 27183
rect 677134 26213 717600 27263
rect 0 26073 47400 26213
rect 0 20920 39391 26073
rect 40000 25993 47400 26073
rect 71400 25993 78800 26213
rect 78993 26073 93607 26213
rect 39471 21000 79054 25993
rect 40000 20920 47400 21000
rect 0 20593 47400 20920
rect 71400 20593 78800 21000
rect 79134 20920 93466 26073
rect 93800 25993 101200 26213
rect 125200 25993 132600 26213
rect 132793 26073 147407 26213
rect 93546 21000 132854 25993
rect 0 5193 40000 20593
rect 0 4923 47400 5193
rect 0 0 39633 4923
rect 40000 4843 47400 4923
rect 71400 4843 78800 5193
rect 78993 4923 93607 20920
rect 93800 20593 101200 21000
rect 125200 20593 132600 21000
rect 132934 20920 147266 26073
rect 147600 25993 155000 26213
rect 179000 25993 186400 26213
rect 186606 26073 202207 26213
rect 147346 21000 186654 25993
rect 39713 0 79054 4843
rect 79134 0 93466 4923
rect 93800 4843 101200 5193
rect 125200 4843 132600 5193
rect 132793 4923 147407 20920
rect 147600 20593 155000 21000
rect 179000 20593 186400 21000
rect 186734 20920 202066 26073
rect 202400 25993 209800 26213
rect 233800 26073 263600 26213
rect 233800 25993 241200 26073
rect 202146 21000 241454 25993
rect 93546 0 132854 4843
rect 132934 0 147266 4923
rect 147600 4843 155000 5193
rect 179000 4843 186400 5193
rect 186606 4923 202207 20920
rect 202400 20593 209800 21000
rect 233800 20920 241200 21000
rect 241534 20920 255866 26073
rect 256200 25993 263600 26073
rect 287600 25993 295000 26213
rect 295206 26073 310807 26213
rect 255946 21000 295254 25993
rect 256200 20920 263600 21000
rect 233800 20593 263600 20920
rect 287600 20593 295000 21000
rect 295334 20920 310666 26073
rect 311000 25993 318400 26213
rect 342400 25993 349800 26213
rect 350006 26073 365607 26213
rect 310746 21000 350054 25993
rect 241200 5193 256200 20593
rect 147346 0 186654 4843
rect 186734 0 202066 4923
rect 202400 4843 209800 5193
rect 233800 4923 263600 5193
rect 233800 4850 241200 4923
rect 233800 4843 241243 4850
rect 202146 0 241454 4843
rect 241534 0 255866 4923
rect 256200 4843 263600 4923
rect 287600 4843 295000 5193
rect 295206 4923 310807 20920
rect 311000 20593 318400 21000
rect 342400 20593 349800 21000
rect 350134 20920 365466 26073
rect 365800 25993 373200 26213
rect 397200 25993 404600 26213
rect 404806 26073 420407 26213
rect 365546 21000 404854 25993
rect 255946 0 295254 4843
rect 295334 0 310666 4923
rect 311000 4843 318400 5193
rect 342400 4843 349800 5193
rect 350006 4923 365607 20920
rect 365800 20593 373200 21000
rect 397200 20593 404600 21000
rect 404934 20920 420266 26073
rect 420600 25993 428000 26213
rect 452000 25993 459400 26213
rect 459606 26073 475207 26213
rect 420346 21000 459654 25993
rect 310746 0 350054 4843
rect 350134 0 365466 4923
rect 365800 4843 373200 5193
rect 397200 4843 404600 5193
rect 404806 4923 420407 20920
rect 420600 20593 428000 21000
rect 452000 20593 459400 21000
rect 459734 20920 475066 26073
rect 475400 25993 482800 26213
rect 506800 25993 514200 26213
rect 514406 26073 530007 26213
rect 475146 21000 514454 25993
rect 365546 0 404854 4843
rect 404934 0 420266 4923
rect 420600 4843 428000 5193
rect 452000 4843 459400 5193
rect 459606 4923 475207 20920
rect 475400 20593 482800 21000
rect 506800 20593 514200 21000
rect 514534 20920 529866 26073
rect 530200 25993 537600 26213
rect 561600 25993 569000 26213
rect 569193 26073 583807 26213
rect 529946 21000 569254 25993
rect 420346 0 459654 4843
rect 459734 0 475066 4923
rect 475400 4843 482800 5193
rect 506800 4843 514200 5193
rect 514406 4923 530007 20920
rect 530200 20593 537600 21000
rect 561600 20593 569000 21000
rect 569334 20920 583666 26073
rect 584000 25993 591400 26213
rect 615400 25993 622800 26213
rect 622993 26073 637607 26213
rect 583746 21000 623054 25993
rect 475146 0 514454 4843
rect 514534 0 529866 4923
rect 530200 4843 537600 5193
rect 561600 4843 569000 5193
rect 569193 4923 583807 20920
rect 584000 20593 591400 21000
rect 615400 20593 622800 21000
rect 623134 20920 637466 26073
rect 637800 25993 645200 26213
rect 669200 25993 676800 26213
rect 677051 26073 717600 26213
rect 637546 21000 677171 25993
rect 529946 0 569254 4843
rect 569334 0 583666 4923
rect 584000 4843 591400 5193
rect 615400 4843 622800 5193
rect 622993 4923 637607 20920
rect 637800 20593 645200 21000
rect 669200 20593 676800 21000
rect 677251 20920 717600 26073
rect 583746 0 623054 4843
rect 623134 0 637466 4923
rect 637800 4843 645200 5193
rect 669200 4843 676800 5193
rect 677051 4923 717600 20920
rect 637546 0 677054 4843
rect 677134 0 717600 4923
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334620 1018402 347160 1030925
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 576820 1018402 589360 1030925
rect 628240 1018512 640760 1031002
rect 297746 1002787 333654 1003677
rect 348146 1002787 384054 1003677
rect 539946 1007147 575854 1008947
rect 539946 1004968 575854 1005617
rect 590346 1007147 626254 1008947
rect 590346 1004968 626254 1005617
rect 540200 1004967 575600 1004968
rect 590600 1004967 626000 1004968
rect 6598 956440 19088 968960
rect 37313 926746 38203 954454
rect 698512 952840 711002 965360
rect 6086 913863 19572 925191
rect 679397 922346 680287 951854
rect 37313 884546 38203 912254
rect 698028 909409 711514 920737
rect 679397 878146 680287 907854
rect 28653 842346 30453 870054
rect 31983 869800 32632 870054
rect 31983 842600 32633 869800
rect 31983 842346 32632 842600
rect 698512 863640 711002 876160
rect 6675 828820 19198 841360
rect 680607 833207 681257 862606
rect 28653 800146 30453 827854
rect 31983 827600 32632 827854
rect 31983 800400 32633 827600
rect 31983 800146 32632 800400
rect 698402 819640 710925 832180
rect 6598 786640 19088 799160
rect 680607 789007 681257 818593
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 36343 497807 36993 525393
rect 6675 484220 19198 496760
rect 30773 455546 31663 483254
rect 36343 455607 36993 483193
rect 685937 474546 686827 504054
rect 698028 461609 711514 472937
rect 6086 442663 19572 453991
rect 30773 413346 31663 441054
rect 685937 430346 686827 460054
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 6598 313440 19088 325960
rect 698512 326640 711002 339160
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 21003 124946 25993 125400
rect 35133 124946 36023 181854
rect 698512 146440 711002 158960
rect 6675 111420 19198 123960
rect 21003 109800 25993 110454
rect 35133 82746 36023 110454
rect 37313 82746 38203 110454
rect 698512 101240 711002 113760
rect 6086 69863 19572 81191
rect 37313 40546 38203 68254
rect 583807 36343 622993 36993
rect 637607 36343 677051 36993
rect 39733 32632 78800 32633
rect 93800 32632 132600 32633
rect 39733 31983 79054 32632
rect 35369 28653 79054 30453
rect 93546 31983 132854 32632
rect 93546 28653 132854 30453
rect 202146 30773 241454 31663
rect 255946 30773 295254 31663
rect 80040 6675 92580 19198
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243009 6086 254337 19572
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570240 6675 582780 19198
rect 624040 6675 636580 19198
<< obsm5 >>
rect 0 1032757 717600 1037600
rect 0 1016917 40800 1032757
rect 76200 1031322 92200 1032757
rect 76200 1018192 78120 1031322
rect 91280 1018192 92200 1031322
rect 76200 1016917 92200 1018192
rect 127600 1031322 143600 1032757
rect 127600 1018192 129520 1031322
rect 142680 1018192 143600 1031322
rect 127600 1016917 143600 1018192
rect 179000 1031322 195000 1032757
rect 179000 1018192 180920 1031322
rect 194080 1018192 195000 1031322
rect 179000 1016917 195000 1018192
rect 230400 1031322 246400 1032757
rect 230400 1018192 232320 1031322
rect 245480 1018192 246400 1031322
rect 230400 1016917 246400 1018192
rect 282000 1031322 298000 1032757
rect 282000 1018192 283920 1031322
rect 297080 1018192 298000 1031322
rect 282000 1016917 298000 1018192
rect 333400 1031245 348400 1032757
rect 333400 1018082 334300 1031245
rect 347480 1018082 348400 1031245
rect 333400 1016917 348400 1018082
rect 383800 1031322 399800 1032757
rect 383800 1018192 385720 1031322
rect 398880 1018192 399800 1031322
rect 383800 1016917 399800 1018192
rect 472800 1031322 488800 1032757
rect 472800 1018192 474720 1031322
rect 487880 1018192 488800 1031322
rect 472800 1016917 488800 1018192
rect 524200 1031322 540200 1032757
rect 524200 1018192 526120 1031322
rect 539280 1018192 540200 1031322
rect 524200 1016917 540200 1018192
rect 575600 1031245 590600 1032757
rect 575600 1018082 576500 1031245
rect 589680 1018082 590600 1031245
rect 575600 1016917 590600 1018082
rect 626000 1031322 642000 1032757
rect 626000 1018192 627920 1031322
rect 641080 1018192 642000 1031322
rect 626000 1016917 642000 1018192
rect 677600 1016917 717600 1032757
rect 0 1011287 40109 1016917
rect 40429 1011607 41000 1016597
rect 41320 1011607 44280 1016597
rect 44600 1011607 45000 1016597
rect 45320 1011607 48280 1016597
rect 48600 1011607 49000 1016597
rect 49320 1011607 52280 1016597
rect 52600 1011607 53000 1016597
rect 53320 1011607 56280 1016597
rect 56600 1011607 57000 1016597
rect 57320 1011607 60280 1016597
rect 60600 1011607 61000 1016597
rect 61320 1011607 64280 1016597
rect 64600 1011607 65000 1016597
rect 65320 1011607 68280 1016597
rect 68600 1011607 69000 1016597
rect 69320 1011607 72280 1016597
rect 72600 1011607 73000 1016597
rect 73320 1011607 74280 1016597
rect 74600 1011607 75000 1016597
rect 75600 1011607 76454 1016597
rect 0 1009267 40226 1011287
rect 40546 1010437 76454 1011287
rect 40546 1009267 76454 1010117
rect 0 1006827 35049 1009267
rect 35369 1007147 76454 1008947
rect 0 1002551 40226 1006827
rect 40546 1005937 76454 1006827
rect 40546 1004968 76454 1005617
rect 40800 1004967 76200 1004968
rect 40546 1003997 76454 1004647
rect 40546 1002787 76454 1003677
rect 0 998449 28333 1002551
rect 0 997600 20683 998449
rect 26313 998245 28333 998449
rect 26313 998216 27163 998245
rect 0 970200 4843 997600
rect 21003 997000 25993 998129
rect 21003 996000 25993 996400
rect 21003 994720 25993 995680
rect 21003 994000 25993 994400
rect 21003 990720 25993 993680
rect 21003 990000 25993 990400
rect 21003 986720 25993 989680
rect 21003 986000 25993 986400
rect 21003 982720 25993 985680
rect 21003 982000 25993 982400
rect 21003 978720 25993 981680
rect 21003 978000 25993 978400
rect 21003 974720 25993 977680
rect 21003 974000 25993 974400
rect 21003 970720 25993 973680
rect 0 969626 20683 970200
rect 21003 969946 25993 970400
rect 26313 969946 27163 997896
rect 27483 969946 28333 997925
rect 28653 969946 30453 1002231
rect 30773 1001257 40226 1002551
rect 40546 1001577 76454 1002467
rect 76774 1001257 91626 1016917
rect 91946 1011607 92400 1016597
rect 92720 1011607 95680 1016597
rect 96000 1011607 96400 1016597
rect 96720 1011607 99680 1016597
rect 100000 1011607 100400 1016597
rect 100720 1011607 103680 1016597
rect 104000 1011607 104400 1016597
rect 104720 1011607 107680 1016597
rect 108000 1011607 108400 1016597
rect 108720 1011607 111680 1016597
rect 112000 1011607 112400 1016597
rect 112720 1011607 115680 1016597
rect 116000 1011607 116400 1016597
rect 116720 1011607 119680 1016597
rect 120000 1011607 120400 1016597
rect 120720 1011607 123680 1016597
rect 124000 1011607 124400 1016597
rect 124720 1011607 125680 1016597
rect 126000 1011607 126400 1016597
rect 127000 1011607 127854 1016597
rect 91946 1010437 127854 1011287
rect 91946 1009267 127854 1010117
rect 91946 1007147 127854 1008947
rect 91946 1005937 127854 1006827
rect 91946 1004968 127854 1005617
rect 92200 1004967 127600 1004968
rect 91946 1003997 127854 1004647
rect 91946 1002787 127854 1003677
rect 91946 1001577 127854 1002467
rect 128174 1001257 143026 1016917
rect 143346 1011607 143800 1016597
rect 144120 1011607 147080 1016597
rect 147400 1011607 147800 1016597
rect 148120 1011607 151080 1016597
rect 151400 1011607 151800 1016597
rect 152120 1011607 155080 1016597
rect 155400 1011607 155800 1016597
rect 156120 1011607 159080 1016597
rect 159400 1011607 159800 1016597
rect 160120 1011607 163080 1016597
rect 163400 1011607 163800 1016597
rect 164120 1011607 167080 1016597
rect 167400 1011607 167800 1016597
rect 168120 1011607 171080 1016597
rect 171400 1011607 171800 1016597
rect 172120 1011607 175080 1016597
rect 175400 1011607 175800 1016597
rect 176120 1011607 177080 1016597
rect 177400 1011607 177800 1016597
rect 178400 1011607 179254 1016597
rect 143346 1010437 179254 1011287
rect 143346 1009267 179254 1010117
rect 143346 1007147 179254 1008947
rect 143346 1005937 179254 1006827
rect 143346 1004968 179254 1005617
rect 143600 1004967 179000 1004968
rect 143346 1003997 179254 1004647
rect 143346 1002787 179254 1003677
rect 143346 1001577 179254 1002467
rect 179574 1001257 194426 1016917
rect 194746 1011607 195200 1016597
rect 195520 1011607 198480 1016597
rect 198800 1011607 199200 1016597
rect 199520 1011607 202480 1016597
rect 202800 1011607 203200 1016597
rect 203520 1011607 206480 1016597
rect 206800 1011607 207200 1016597
rect 207520 1011607 210480 1016597
rect 210800 1011607 211200 1016597
rect 211520 1011607 214480 1016597
rect 214800 1011607 215200 1016597
rect 215520 1011607 218480 1016597
rect 218800 1011607 219200 1016597
rect 219520 1011607 222480 1016597
rect 222800 1011607 223200 1016597
rect 223520 1011607 226480 1016597
rect 226800 1011607 227200 1016597
rect 227520 1011607 228480 1016597
rect 228800 1011607 229200 1016597
rect 229800 1011607 230654 1016597
rect 194746 1010437 230654 1011287
rect 194746 1009267 230654 1010117
rect 194746 1007147 230654 1008947
rect 194746 1005937 230654 1006827
rect 194746 1004968 230654 1005617
rect 195000 1004967 230400 1004968
rect 194746 1003997 230654 1004647
rect 194746 1002787 230654 1003677
rect 194746 1001577 230654 1002467
rect 230974 1001257 245826 1016917
rect 246146 1011607 246600 1016597
rect 246920 1011607 249880 1016597
rect 250200 1011607 250600 1016597
rect 250920 1011607 253880 1016597
rect 254200 1011607 254600 1016597
rect 254920 1011607 257880 1016597
rect 258200 1011607 258600 1016597
rect 258920 1011607 261880 1016597
rect 262200 1011607 262600 1016597
rect 262920 1011607 265880 1016597
rect 266200 1011607 266600 1016597
rect 266920 1011607 269880 1016597
rect 270200 1011607 270600 1016597
rect 270920 1011607 273880 1016597
rect 274200 1011607 274600 1016597
rect 274920 1011607 277880 1016597
rect 278200 1011607 278600 1016597
rect 278920 1011607 279880 1016597
rect 280200 1011607 280600 1016597
rect 281200 1011607 282254 1016597
rect 246146 1010437 282254 1011287
rect 246146 1009267 282254 1010117
rect 246146 1007147 282254 1008947
rect 246146 1005937 282254 1006827
rect 246146 1004968 282254 1005617
rect 246400 1004967 282000 1004968
rect 246146 1003997 282254 1004647
rect 246146 1002787 282254 1003677
rect 246146 1001577 282254 1002467
rect 282574 1001257 297426 1016917
rect 297746 1011607 298200 1016597
rect 298520 1011607 301480 1016597
rect 301800 1011607 302200 1016597
rect 302520 1011607 305480 1016597
rect 305800 1011607 306200 1016597
rect 306520 1011607 309480 1016597
rect 309800 1011607 310200 1016597
rect 310520 1011607 313480 1016597
rect 313800 1011607 314200 1016597
rect 314520 1011607 317480 1016597
rect 317800 1011607 318200 1016597
rect 318520 1011607 321480 1016597
rect 321800 1011607 322200 1016597
rect 322520 1011607 325480 1016597
rect 325800 1011607 326200 1016597
rect 326520 1011607 329480 1016597
rect 329800 1011607 330200 1016597
rect 330520 1011607 331480 1016597
rect 331800 1011607 332200 1016597
rect 332800 1011607 333654 1016597
rect 297746 1010437 333654 1011287
rect 297746 1009267 333654 1010117
rect 297746 1007147 333654 1008947
rect 297746 1005937 333654 1006827
rect 297746 1004968 333654 1005617
rect 333974 1004968 347826 1016917
rect 348146 1011607 348600 1016597
rect 348920 1011607 351880 1016597
rect 352200 1011607 352600 1016597
rect 352920 1011607 355880 1016597
rect 356200 1011607 356600 1016597
rect 356920 1011607 359880 1016597
rect 360200 1011607 360600 1016597
rect 360920 1011607 363880 1016597
rect 364200 1011607 364600 1016597
rect 364920 1011607 367880 1016597
rect 368200 1011607 368600 1016597
rect 368920 1011607 371880 1016597
rect 372200 1011607 372600 1016597
rect 372920 1011607 375880 1016597
rect 376200 1011607 376600 1016597
rect 376920 1011607 379880 1016597
rect 380200 1011607 380600 1016597
rect 380920 1011607 381880 1016597
rect 382200 1011607 382600 1016597
rect 383200 1011607 384054 1016597
rect 348146 1010437 384054 1011287
rect 348146 1009267 384054 1010117
rect 348146 1007147 384054 1008947
rect 348146 1005937 384054 1006827
rect 348146 1004968 384054 1005617
rect 298000 1004967 383800 1004968
rect 297746 1003997 333654 1004647
rect 297746 1001577 333654 1002467
rect 333974 1001257 347826 1004967
rect 348146 1003997 384054 1004647
rect 348146 1001577 384054 1002467
rect 384374 1001257 399226 1016917
rect 399546 1011607 400000 1016597
rect 400320 1011607 403280 1016597
rect 403600 1011607 404000 1016597
rect 404320 1011607 407280 1016597
rect 407600 1011607 408000 1016597
rect 408320 1011607 411280 1016597
rect 411600 1011607 412000 1016597
rect 412320 1011607 415280 1016597
rect 415600 1011607 416000 1016597
rect 416320 1011607 419280 1016597
rect 419600 1011607 420000 1016597
rect 420320 1011607 423280 1016597
rect 423600 1011607 424000 1016597
rect 424320 1011607 427280 1016597
rect 427600 1011607 428000 1016597
rect 428320 1011607 431280 1016597
rect 431600 1011607 432000 1016597
rect 432320 1011607 433280 1016597
rect 433600 1011607 434000 1016597
rect 434600 1011607 437400 1016597
rect 437720 1011607 440680 1016597
rect 441000 1011607 441400 1016597
rect 441720 1011607 444680 1016597
rect 445000 1011607 445400 1016597
rect 445720 1011607 448680 1016597
rect 449000 1011607 449400 1016597
rect 449720 1011607 452680 1016597
rect 453000 1011607 453400 1016597
rect 453720 1011607 456680 1016597
rect 457000 1011607 457400 1016597
rect 457720 1011607 460680 1016597
rect 461000 1011607 461400 1016597
rect 461720 1011607 464680 1016597
rect 465000 1011607 465400 1016597
rect 465720 1011607 468680 1016597
rect 469000 1011607 469400 1016597
rect 469720 1011607 470680 1016597
rect 471000 1011607 471400 1016597
rect 472000 1011607 473054 1016597
rect 399546 1010437 473054 1011287
rect 399546 1009267 473054 1010117
rect 399546 1007147 435200 1008947
rect 436200 1007147 473054 1008947
rect 399546 1005937 436200 1006827
rect 437200 1005937 473054 1006827
rect 399546 1004968 435200 1005617
rect 399800 1004967 435200 1004968
rect 436200 1004968 473054 1005617
rect 436200 1004967 472800 1004968
rect 399546 1003997 473054 1004647
rect 399546 1002787 473054 1003677
rect 399546 1001577 473054 1002467
rect 473374 1001257 488226 1016917
rect 488546 1011607 489000 1016597
rect 489320 1011607 492280 1016597
rect 492600 1011607 493000 1016597
rect 493320 1011607 496280 1016597
rect 496600 1011607 497000 1016597
rect 497320 1011607 500280 1016597
rect 500600 1011607 501000 1016597
rect 501320 1011607 504280 1016597
rect 504600 1011607 505000 1016597
rect 505320 1011607 508280 1016597
rect 508600 1011607 509000 1016597
rect 509320 1011607 512280 1016597
rect 512600 1011607 513000 1016597
rect 513320 1011607 516280 1016597
rect 516600 1011607 517000 1016597
rect 517320 1011607 520280 1016597
rect 520600 1011607 521000 1016597
rect 521320 1011607 522280 1016597
rect 522600 1011607 523000 1016597
rect 523600 1011607 524454 1016597
rect 488546 1010437 524454 1011287
rect 488546 1009267 524454 1010117
rect 488546 1007147 524454 1008947
rect 488546 1005937 524454 1006827
rect 488546 1004968 524454 1005617
rect 488800 1004967 524200 1004968
rect 488546 1003997 524454 1004647
rect 488546 1002787 524454 1003677
rect 488546 1001577 524454 1002467
rect 524774 1001257 539626 1016917
rect 539946 1011607 540400 1016597
rect 540720 1011607 543680 1016597
rect 544000 1011607 544400 1016597
rect 544720 1011607 547680 1016597
rect 548000 1011607 548400 1016597
rect 548720 1011607 551680 1016597
rect 552000 1011607 552400 1016597
rect 552720 1011607 555680 1016597
rect 556000 1011607 556400 1016597
rect 556720 1011607 559680 1016597
rect 560000 1011607 560400 1016597
rect 560720 1011607 563680 1016597
rect 564000 1011607 564400 1016597
rect 564720 1011607 567680 1016597
rect 568000 1011607 568400 1016597
rect 568720 1011607 571680 1016597
rect 572000 1011607 572400 1016597
rect 572720 1011607 573680 1016597
rect 574000 1011607 574400 1016597
rect 575000 1011607 575854 1016597
rect 539946 1010437 575854 1011287
rect 539946 1009267 575854 1010117
rect 539946 1005937 575854 1006827
rect 576174 1004968 590026 1016917
rect 590346 1011607 590800 1016597
rect 591120 1011607 594080 1016597
rect 594400 1011607 594800 1016597
rect 595120 1011607 598080 1016597
rect 598400 1011607 598800 1016597
rect 599120 1011607 602080 1016597
rect 602400 1011607 602800 1016597
rect 603120 1011607 606080 1016597
rect 606400 1011607 606800 1016597
rect 607120 1011607 610080 1016597
rect 610400 1011607 610800 1016597
rect 611120 1011607 614080 1016597
rect 614400 1011607 614800 1016597
rect 615120 1011607 618080 1016597
rect 618400 1011607 618800 1016597
rect 619120 1011607 622080 1016597
rect 622400 1011607 622800 1016597
rect 623120 1011607 624080 1016597
rect 624400 1011607 624800 1016597
rect 625400 1011607 626254 1016597
rect 590346 1010437 626254 1011287
rect 590346 1009267 626254 1010117
rect 590346 1005937 626254 1006827
rect 575600 1004967 590600 1004968
rect 539946 1003997 575854 1004647
rect 539946 1002787 575854 1003677
rect 539946 1001577 575854 1002467
rect 576174 1001257 590026 1004967
rect 590346 1003997 626254 1004647
rect 590346 1002787 626254 1003677
rect 590346 1001577 626254 1002467
rect 626574 1001257 641426 1016917
rect 641746 1011607 642200 1016597
rect 642520 1011607 645480 1016597
rect 645800 1011607 646200 1016597
rect 646520 1011607 649480 1016597
rect 649800 1011607 650200 1016597
rect 650520 1011607 653480 1016597
rect 653800 1011607 654200 1016597
rect 654520 1011607 657480 1016597
rect 657800 1011607 658200 1016597
rect 658520 1011607 661480 1016597
rect 661800 1011607 662200 1016597
rect 662520 1011607 665480 1016597
rect 665800 1011607 666200 1016597
rect 666520 1011607 669480 1016597
rect 669800 1011607 670200 1016597
rect 670520 1011607 673480 1016597
rect 673800 1011607 674200 1016597
rect 674520 1011607 675480 1016597
rect 675800 1011607 676200 1016597
rect 676800 1011607 678129 1016597
rect 678449 1011287 717600 1016917
rect 641746 1010437 677896 1011287
rect 678216 1010437 717600 1011287
rect 641746 1009267 677925 1010117
rect 678245 1009267 717600 1010437
rect 641746 1007147 682231 1008947
rect 682551 1006827 717600 1009267
rect 641746 1005937 677895 1006827
rect 678215 1005617 717600 1006827
rect 641746 1004968 677867 1005617
rect 642000 1004967 677867 1004968
rect 678187 1004967 717600 1005617
rect 641746 1003997 677877 1004647
rect 678197 1003997 717600 1004967
rect 641746 1002787 677920 1003677
rect 678240 1002551 717600 1003997
rect 678240 1002467 686827 1002551
rect 641746 1001577 677905 1002467
rect 678225 1001257 686827 1002467
rect 30773 1000607 40229 1001257
rect 40549 1000607 76393 1001257
rect 76713 1000607 91674 1001257
rect 91994 1000607 127793 1001257
rect 128113 1000607 143074 1001257
rect 143394 1000607 179193 1001257
rect 179513 1000607 194474 1001257
rect 194794 1000607 230593 1001257
rect 230913 1000607 245874 1001257
rect 246194 1000607 282193 1001257
rect 282513 1000607 297474 1001257
rect 297794 1000607 333593 1001257
rect 333913 1000607 347887 1001257
rect 348207 1000607 383993 1001257
rect 384313 1000607 399274 1001257
rect 399594 1000607 435200 1001257
rect 436200 1000607 472993 1001257
rect 473313 1000607 488274 1001257
rect 488594 1000607 524393 1001257
rect 524713 1000607 539674 1001257
rect 539994 1000607 575793 1001257
rect 576113 1000607 590087 1001257
rect 590407 1000607 626193 1001257
rect 626513 1000607 641474 1001257
rect 641794 1000607 677894 1001257
rect 678214 1000607 686827 1001257
rect 30773 998677 40226 1000607
rect 40546 999397 76454 1000287
rect 30773 998240 36993 998677
rect 38523 998390 40226 998677
rect 30773 998215 33603 998240
rect 35133 998225 36993 998240
rect 31983 998197 33603 998215
rect 36343 998214 36993 998225
rect 31983 998187 32633 998197
rect 30773 969946 31663 997895
rect 31983 970200 32633 997867
rect 31983 969946 32632 970200
rect 32953 969946 33603 997877
rect 33923 969946 34813 997920
rect 35133 969946 36023 997905
rect 36343 969994 36993 997894
rect 37313 969946 38203 998357
rect 38523 998027 39573 998070
rect 39893 998027 40226 998390
rect 40546 998027 76454 999077
rect 76774 998027 91626 1000607
rect 91946 999397 127854 1000287
rect 91946 998027 127854 999077
rect 128174 998027 143026 1000607
rect 143346 999397 179254 1000287
rect 143346 998027 179254 999077
rect 179574 998027 194426 1000607
rect 194746 999397 230654 1000287
rect 194746 998027 230654 999077
rect 230974 998027 245826 1000607
rect 246146 999397 282254 1000287
rect 246146 998027 282254 999077
rect 282574 998027 297426 1000607
rect 297746 999397 333654 1000287
rect 297746 998027 333654 999077
rect 333974 998027 347826 1000607
rect 348146 999397 384054 1000287
rect 348146 998027 384054 999077
rect 384374 998027 399226 1000607
rect 399546 999397 436200 1000287
rect 437200 999397 473054 1000287
rect 399546 998027 473054 999077
rect 473374 998027 488226 1000607
rect 488546 999397 524454 1000287
rect 488546 998027 524454 999077
rect 524774 998027 539626 1000607
rect 539946 999397 575854 1000287
rect 539946 998027 575854 999077
rect 576174 998027 590026 1000607
rect 590346 999397 626254 1000287
rect 590346 998027 626254 999077
rect 626574 998027 641426 1000607
rect 641746 999397 678357 1000287
rect 678677 999077 686827 1000607
rect 641746 998027 678070 999077
rect 38523 997920 40226 998027
rect 38523 969946 39573 997920
tri 39573 997600 39893 997920 nw
rect 39893 997707 40226 997920
tri 677600 997707 677920 998027 ne
rect 677920 997707 678027 998027
rect 678390 997707 686827 999077
rect 39893 997600 40800 997707
rect 677600 997374 686827 997707
rect 677600 996800 677707 997374
rect 680607 997371 681257 997374
rect 36343 969626 36993 969674
rect 0 969280 39573 969626
rect 0 956120 6278 969280
rect 19408 956120 39573 969280
rect 678027 967346 679077 997054
rect 679397 967346 680287 997054
rect 680607 967407 681257 997051
rect 681577 967346 682467 997054
rect 682787 967346 683677 997054
rect 683997 967346 684647 997054
rect 684968 996800 685617 997054
rect 684967 967600 685617 996800
rect 684968 967346 685617 967600
rect 685937 967346 686827 997054
rect 687147 967346 688947 1002231
rect 689267 997491 717600 1002551
rect 689267 997374 691287 997491
rect 689267 967346 690117 997054
rect 690437 967346 691287 997054
rect 691607 996400 696597 997171
rect 696917 996800 717600 997491
rect 691607 995400 696597 995800
rect 691607 992120 696597 995080
rect 691607 991400 696597 991800
rect 691607 988120 696597 991080
rect 691607 987400 696597 987800
rect 691607 984120 696597 987080
rect 691607 983400 696597 983800
rect 691607 980120 696597 983080
rect 691607 979400 696597 979800
rect 691607 976120 696597 979080
rect 691607 975400 696597 975800
rect 691607 972120 696597 975080
rect 691607 971400 696597 971800
rect 691607 968120 696597 971080
rect 691607 967346 696597 967800
rect 712757 967600 717600 996800
rect 680607 967026 681257 967087
rect 696917 967026 717600 967600
rect 0 954774 39573 956120
rect 678027 965680 717600 967026
rect 0 954200 20683 954774
rect 36343 954713 36993 954774
rect 0 927000 4843 954200
rect 21003 953800 25993 954454
rect 21003 952800 25993 953200
rect 21003 951520 25993 952480
rect 21003 950800 25993 951200
rect 21003 947520 25993 950480
rect 21003 946800 25993 947200
rect 21003 943520 25993 946480
rect 21003 942800 25993 943200
rect 21003 939520 25993 942480
rect 21003 938800 25993 939200
rect 21003 935520 25993 938480
rect 21003 934800 25993 935200
rect 21003 931520 25993 934480
rect 21003 930800 25993 931200
rect 21003 927520 25993 930480
rect 0 926426 20683 927000
rect 21003 926746 25993 927200
rect 26313 926746 27163 954454
rect 27483 926746 28333 954454
rect 28653 926746 30453 954454
rect 30773 926746 31663 954454
rect 31983 954200 32632 954454
rect 31983 926746 32633 954200
rect 32953 926746 33603 954454
rect 33923 926746 34813 954454
rect 35133 926746 36023 954454
rect 36343 926807 36993 954393
rect 38523 926746 39573 954454
rect 678027 952520 698192 965680
rect 711322 952520 717600 965680
rect 678027 952174 717600 952520
rect 680607 952126 681257 952174
rect 32632 926426 32633 926746
rect 36343 926426 36993 926487
rect 0 925511 39573 926426
rect 0 913543 5766 925511
rect 19892 913543 39573 925511
rect 678027 922346 679077 951854
rect 680607 922407 681257 951806
rect 681577 922346 682467 951854
rect 682787 922346 683677 951854
rect 683997 922346 684647 951854
rect 684968 951600 685617 951854
rect 684967 922346 685617 951600
rect 685937 922346 686827 951854
rect 687147 922346 688947 951854
rect 689267 922346 690117 951854
rect 690437 922346 691287 951854
rect 691607 951400 696597 951854
rect 696917 951600 717600 952174
rect 691607 950400 696597 950800
rect 691607 947120 696597 950080
rect 691607 946400 696597 946800
rect 691607 943120 696597 946080
rect 691607 942400 696597 942800
rect 691607 939120 696597 942080
rect 691607 938400 696597 938800
rect 691607 935120 696597 938080
rect 691607 934400 696597 934800
rect 691607 931120 696597 934080
rect 691607 930400 696597 930800
rect 691607 927120 696597 930080
rect 691607 926400 696597 926800
rect 691607 923120 696597 926080
rect 691607 922346 696597 922800
rect 712757 922600 717600 951600
rect 680607 922026 681257 922087
rect 684967 922026 684968 922346
rect 696917 922026 717600 922600
rect 0 912574 39573 913543
rect 678027 921057 717600 922026
rect 0 912000 20683 912574
rect 32632 912254 32633 912574
rect 36343 912513 36993 912574
rect 0 884800 4843 912000
rect 21003 911600 25993 912254
rect 21003 910600 25993 911000
rect 21003 909320 25993 910280
rect 21003 908600 25993 909000
rect 21003 905320 25993 908280
rect 21003 904600 25993 905000
rect 21003 901320 25993 904280
rect 21003 900600 25993 901000
rect 21003 897320 25993 900280
rect 21003 896600 25993 897000
rect 21003 893320 25993 896280
rect 21003 892600 25993 893000
rect 21003 889320 25993 892280
rect 21003 888600 25993 889000
rect 21003 885320 25993 888280
rect 0 884226 20683 884800
rect 21003 884546 25993 885000
rect 26313 884546 27163 912254
rect 27483 884546 28333 912254
rect 28653 884546 30453 912254
rect 30773 884546 31663 912254
rect 31983 884546 32633 912254
rect 32953 884546 33603 912254
rect 33923 884546 34813 912254
rect 35133 884546 36023 912254
rect 36343 884607 36993 912193
rect 38523 884546 39573 912254
rect 678027 909089 697708 921057
rect 711834 909089 717600 921057
rect 678027 908174 717600 909089
rect 680607 908113 681257 908174
rect 684967 907854 684968 908174
rect 32632 884226 32633 884546
rect 36343 884226 36993 884287
rect 0 883880 39573 884226
rect 0 870700 6355 883880
rect 6675 871020 19198 883560
rect 19518 870700 39573 883880
rect 678027 878146 679077 907854
rect 680607 878207 681257 907793
rect 681577 878146 682467 907854
rect 682787 878146 683677 907854
rect 683997 878146 684647 907854
rect 684967 878400 685617 907854
rect 684968 878146 685617 878400
rect 685937 878146 686827 907854
rect 687147 878146 688947 907854
rect 689267 878146 690117 907854
rect 690437 878146 691287 907854
rect 691607 907200 696597 907854
rect 696917 907600 717600 908174
rect 691607 906200 696597 906600
rect 691607 902920 696597 905880
rect 691607 902200 696597 902600
rect 691607 898920 696597 901880
rect 691607 898200 696597 898600
rect 691607 894920 696597 897880
rect 691607 894200 696597 894600
rect 691607 890920 696597 893880
rect 691607 890200 696597 890600
rect 691607 886920 696597 889880
rect 691607 886200 696597 886600
rect 691607 882920 696597 885880
rect 691607 882200 696597 882600
rect 691607 878920 696597 881880
rect 691607 878146 696597 878600
rect 712757 878400 717600 907600
rect 680607 877826 681257 877887
rect 696917 877826 717600 878400
rect 0 870374 39573 870700
rect 678027 876480 717600 877826
rect 0 869800 20683 870374
rect 0 842600 4843 869800
rect 21003 869400 25993 870054
rect 21003 868400 25993 868800
rect 21003 867120 25993 868080
rect 21003 866400 25993 866800
rect 21003 863120 25993 866080
rect 21003 862400 25993 862800
rect 21003 859120 25993 862080
rect 21003 858400 25993 858800
rect 21003 855120 25993 858080
rect 21003 854400 25993 854800
rect 21003 851120 25993 854080
rect 21003 850400 25993 850800
rect 21003 847120 25993 850080
rect 21003 846400 25993 846800
rect 21003 843120 25993 846080
rect 0 842026 20683 842600
rect 21003 842346 25993 842800
rect 26313 842346 27163 870054
rect 27483 842346 28333 870054
rect 30773 842346 31663 870054
rect 32632 869800 32633 870374
rect 36343 870313 36993 870374
rect 32632 842026 32633 842600
rect 32953 842346 33603 870054
rect 33923 842346 34813 870054
rect 35133 842346 36023 870054
rect 36343 842407 36993 869993
rect 37313 842346 38203 870054
rect 38523 842346 39573 870054
rect 678027 863320 698192 876480
rect 711322 863320 717600 876480
rect 678027 862974 717600 863320
rect 680607 862926 681257 862974
rect 36343 842026 36993 842087
rect 0 841680 39573 842026
rect 0 828500 6355 841680
rect 19518 828500 39573 841680
rect 678027 833146 679077 862654
rect 679397 833146 680287 862654
rect 681577 833146 682467 862654
rect 682787 833146 683677 862654
rect 683997 833146 684647 862654
rect 684968 862400 685617 862654
rect 684967 833146 685617 862400
rect 685937 833146 686827 862654
rect 687147 833146 688947 862654
rect 689267 833146 690117 862654
rect 690437 833146 691287 862654
rect 691607 862200 696597 862654
rect 696917 862400 717600 862974
rect 691607 861200 696597 861600
rect 691607 857920 696597 860880
rect 691607 857200 696597 857600
rect 691607 853920 696597 856880
rect 691607 853200 696597 853600
rect 691607 849920 696597 852880
rect 691607 849200 696597 849600
rect 691607 845920 696597 848880
rect 691607 845200 696597 845600
rect 691607 841920 696597 844880
rect 691607 841200 696597 841600
rect 691607 837920 696597 840880
rect 691607 837200 696597 837600
rect 691607 833920 696597 836880
rect 691607 833146 696597 833600
rect 712757 833400 717600 862400
rect 680607 832826 681257 832887
rect 684967 832826 684968 833146
rect 696917 832826 717600 833400
rect 0 828174 39573 828500
rect 678027 832500 717600 832826
rect 0 827600 20683 828174
rect 0 800400 4843 827600
rect 21003 827200 25993 827854
rect 21003 826200 25993 826600
rect 21003 824920 25993 825880
rect 21003 824200 25993 824600
rect 21003 820920 25993 823880
rect 21003 820200 25993 820600
rect 21003 816920 25993 819880
rect 21003 816200 25993 816600
rect 21003 812920 25993 815880
rect 21003 812200 25993 812600
rect 21003 808920 25993 811880
rect 21003 808200 25993 808600
rect 21003 804920 25993 807880
rect 21003 804200 25993 804600
rect 21003 800920 25993 803880
rect 0 799826 20683 800400
rect 21003 800146 25993 800600
rect 26313 800146 27163 827854
rect 27483 800146 28333 827854
rect 30773 800146 31663 827854
rect 32632 827600 32633 828174
rect 36343 828113 36993 828174
rect 32953 800146 33603 827854
rect 33923 800146 34813 827854
rect 35133 800146 36023 827854
rect 36343 800194 36993 827793
rect 37313 800146 38203 827854
rect 38523 800146 39573 827854
rect 678027 819320 698082 832500
rect 711245 819320 717600 832500
rect 678027 818974 717600 819320
rect 680607 818913 681257 818974
rect 684967 818654 684968 818974
rect 36343 799826 36993 799874
rect 0 799480 39573 799826
rect 0 786320 6278 799480
rect 19408 786320 39573 799480
rect 678027 788946 679077 818654
rect 679397 788946 680287 818654
rect 681577 788946 682467 818654
rect 682787 788946 683677 818654
rect 683997 788946 684647 818654
rect 684967 789200 685617 818654
rect 684968 788946 685617 789200
rect 685937 788946 686827 818654
rect 687147 788946 688947 818654
rect 689267 788946 690117 818654
rect 690437 788946 691287 818654
rect 691607 818000 696597 818654
rect 696917 818400 717600 818974
rect 691607 817000 696597 817400
rect 691607 813720 696597 816680
rect 691607 813000 696597 813400
rect 691607 809720 696597 812680
rect 691607 809000 696597 809400
rect 691607 805720 696597 808680
rect 691607 805000 696597 805400
rect 691607 801720 696597 804680
rect 691607 801000 696597 801400
rect 691607 797720 696597 800680
rect 691607 797000 696597 797400
rect 691607 793720 696597 796680
rect 691607 793000 696597 793400
rect 691607 789720 696597 792680
rect 691607 788946 696597 789400
rect 712757 789200 717600 818400
rect 680607 788626 681257 788687
rect 696917 788626 717600 789200
rect 0 784974 39573 786320
rect 678027 787280 717600 788626
rect 0 784400 20683 784974
rect 36343 784913 36993 784974
rect 0 757200 4843 784400
rect 21003 784000 25993 784654
rect 21003 783000 25993 783400
rect 21003 781720 25993 782680
rect 21003 781000 25993 781400
rect 21003 777720 25993 780680
rect 21003 777000 25993 777400
rect 21003 773720 25993 776680
rect 21003 773000 25993 773400
rect 21003 769720 25993 772680
rect 21003 769000 25993 769400
rect 21003 765720 25993 768680
rect 21003 765000 25993 765400
rect 21003 761720 25993 764680
rect 21003 761000 25993 761400
rect 21003 757720 25993 760680
rect 0 756626 20683 757200
rect 21003 756946 25993 757400
rect 26313 756946 27163 784654
rect 27483 756946 28333 784654
rect 28653 756946 30453 784654
rect 30773 756946 31663 784654
rect 31983 784400 32632 784654
rect 31983 757200 32633 784400
rect 31983 756946 32632 757200
rect 32953 756946 33603 784654
rect 33923 756946 34813 784654
rect 35133 756946 36023 784654
rect 36343 756994 36993 784593
rect 37313 756946 38203 784654
rect 38523 756946 39573 784654
rect 678027 774120 698192 787280
rect 711322 774120 717600 787280
rect 678027 773774 717600 774120
rect 680607 773726 681257 773774
rect 36343 756626 36993 756674
rect 0 756280 39573 756626
rect 0 743120 6278 756280
rect 19408 743120 39573 756280
rect 678027 743946 679077 773454
rect 679397 743946 680287 773454
rect 680607 744007 681257 773406
rect 681577 743946 682467 773454
rect 682787 743946 683677 773454
rect 683997 743946 684647 773454
rect 684968 773200 685617 773454
rect 684967 744200 685617 773200
rect 684968 743946 685617 744200
rect 685937 743946 686827 773454
rect 687147 743946 688947 773454
rect 689267 743946 690117 773454
rect 690437 743946 691287 773454
rect 691607 773000 696597 773454
rect 696917 773200 717600 773774
rect 691607 772000 696597 772400
rect 691607 768720 696597 771680
rect 691607 768000 696597 768400
rect 691607 764720 696597 767680
rect 691607 764000 696597 764400
rect 691607 760720 696597 763680
rect 691607 760000 696597 760400
rect 691607 756720 696597 759680
rect 691607 756000 696597 756400
rect 691607 752720 696597 755680
rect 691607 752000 696597 752400
rect 691607 748720 696597 751680
rect 691607 748000 696597 748400
rect 691607 744720 696597 747680
rect 691607 743946 696597 744400
rect 712757 744200 717600 773200
rect 680607 743626 681257 743687
rect 696917 743626 717600 744200
rect 0 741774 39573 743120
rect 678027 742280 717600 743626
rect 0 741200 20683 741774
rect 36343 741713 36993 741774
rect 0 714000 4843 741200
rect 21003 740800 25993 741454
rect 21003 739800 25993 740200
rect 21003 738520 25993 739480
rect 21003 737800 25993 738200
rect 21003 734520 25993 737480
rect 21003 733800 25993 734200
rect 21003 730520 25993 733480
rect 21003 729800 25993 730200
rect 21003 726520 25993 729480
rect 21003 725800 25993 726200
rect 21003 722520 25993 725480
rect 21003 721800 25993 722200
rect 21003 718520 25993 721480
rect 21003 717800 25993 718200
rect 21003 714520 25993 717480
rect 0 713426 20683 714000
rect 21003 713746 25993 714200
rect 26313 713746 27163 741454
rect 27483 713746 28333 741454
rect 28653 713746 30453 741454
rect 30773 713746 31663 741454
rect 31983 741200 32632 741454
rect 31983 714000 32633 741200
rect 31983 713746 32632 714000
rect 32953 713746 33603 741454
rect 33923 713746 34813 741454
rect 35133 713746 36023 741454
rect 36343 713794 36993 741393
rect 37313 713746 38203 741454
rect 38523 713746 39573 741454
rect 678027 729120 698192 742280
rect 711322 729120 717600 742280
rect 678027 728774 717600 729120
rect 680607 728726 681257 728774
rect 36343 713426 36993 713474
rect 0 713080 39573 713426
rect 0 699920 6278 713080
rect 19408 699920 39573 713080
rect 0 698574 39573 699920
rect 678027 698946 679077 728454
rect 679397 698946 680287 728454
rect 680607 699007 681257 728406
rect 681577 698946 682467 728454
rect 682787 698946 683677 728454
rect 683997 698946 684647 728454
rect 684968 728200 685617 728454
rect 684967 699200 685617 728200
rect 684968 698946 685617 699200
rect 685937 698946 686827 728454
rect 687147 698946 688947 728454
rect 689267 698946 690117 728454
rect 690437 698946 691287 728454
rect 691607 728000 696597 728454
rect 696917 728200 717600 728774
rect 691607 727000 696597 727400
rect 691607 723720 696597 726680
rect 691607 723000 696597 723400
rect 691607 719720 696597 722680
rect 691607 719000 696597 719400
rect 691607 715720 696597 718680
rect 691607 715000 696597 715400
rect 691607 711720 696597 714680
rect 691607 711000 696597 711400
rect 691607 707720 696597 710680
rect 691607 707000 696597 707400
rect 691607 703720 696597 706680
rect 691607 703000 696597 703400
rect 691607 699720 696597 702680
rect 691607 698946 696597 699400
rect 712757 699200 717600 728200
rect 680607 698626 681257 698687
rect 696917 698626 717600 699200
rect 0 698000 20683 698574
rect 36343 698513 36993 698574
rect 0 670800 4843 698000
rect 21003 697600 25993 698254
rect 21003 696600 25993 697000
rect 21003 695320 25993 696280
rect 21003 694600 25993 695000
rect 21003 691320 25993 694280
rect 21003 690600 25993 691000
rect 21003 687320 25993 690280
rect 21003 686600 25993 687000
rect 21003 683320 25993 686280
rect 21003 682600 25993 683000
rect 21003 679320 25993 682280
rect 21003 678600 25993 679000
rect 21003 675320 25993 678280
rect 21003 674600 25993 675000
rect 21003 671320 25993 674280
rect 0 670226 20683 670800
rect 21003 670546 25993 671000
rect 26313 670546 27163 698254
rect 27483 670546 28333 698254
rect 28653 670546 30453 698254
rect 30773 670546 31663 698254
rect 31983 698000 32632 698254
rect 31983 670800 32633 698000
rect 31983 670546 32632 670800
rect 32953 670546 33603 698254
rect 33923 670546 34813 698254
rect 35133 670546 36023 698254
rect 36343 670594 36993 698193
rect 37313 670546 38203 698254
rect 38523 670546 39573 698254
rect 678027 697280 717600 698626
rect 678027 684120 698192 697280
rect 711322 684120 717600 697280
rect 678027 683774 717600 684120
rect 680607 683726 681257 683774
rect 36343 670226 36993 670274
rect 0 669880 39573 670226
rect 0 656720 6278 669880
rect 19408 656720 39573 669880
rect 0 655374 39573 656720
rect 0 654800 20683 655374
rect 36343 655313 36993 655374
rect 0 627600 4843 654800
rect 21003 654400 25993 655054
rect 21003 653400 25993 653800
rect 21003 652120 25993 653080
rect 21003 651400 25993 651800
rect 21003 648120 25993 651080
rect 21003 647400 25993 647800
rect 21003 644120 25993 647080
rect 21003 643400 25993 643800
rect 21003 640120 25993 643080
rect 21003 639400 25993 639800
rect 21003 636120 25993 639080
rect 21003 635400 25993 635800
rect 21003 632120 25993 635080
rect 21003 631400 25993 631800
rect 21003 628120 25993 631080
rect 0 627026 20683 627600
rect 21003 627346 25993 627800
rect 26313 627346 27163 655054
rect 27483 627346 28333 655054
rect 28653 627346 30453 655054
rect 30773 627346 31663 655054
rect 31983 654800 32632 655054
rect 31983 627600 32633 654800
rect 31983 627346 32632 627600
rect 32953 627346 33603 655054
rect 33923 627346 34813 655054
rect 35133 627346 36023 655054
rect 36343 627394 36993 654993
rect 37313 627346 38203 655054
rect 38523 627346 39573 655054
rect 678027 653746 679077 683454
rect 679397 653746 680287 683454
rect 680607 653807 681257 683406
rect 681577 653746 682467 683454
rect 682787 653746 683677 683454
rect 683997 653746 684647 683454
rect 684968 683200 685617 683454
rect 684967 654000 685617 683200
rect 684968 653746 685617 654000
rect 685937 653746 686827 683454
rect 687147 653746 688947 683454
rect 689267 653746 690117 683454
rect 690437 653746 691287 683454
rect 691607 682800 696597 683454
rect 696917 683200 717600 683774
rect 691607 681800 696597 682200
rect 691607 678520 696597 681480
rect 691607 677800 696597 678200
rect 691607 674520 696597 677480
rect 691607 673800 696597 674200
rect 691607 670520 696597 673480
rect 691607 669800 696597 670200
rect 691607 666520 696597 669480
rect 691607 665800 696597 666200
rect 691607 662520 696597 665480
rect 691607 661800 696597 662200
rect 691607 658520 696597 661480
rect 691607 657800 696597 658200
rect 691607 654520 696597 657480
rect 691607 653746 696597 654200
rect 712757 654000 717600 683200
rect 680607 653426 681257 653487
rect 696917 653426 717600 654000
rect 678027 652080 717600 653426
rect 678027 638920 698192 652080
rect 711322 638920 717600 652080
rect 678027 638574 717600 638920
rect 680607 638526 681257 638574
rect 36343 627026 36993 627074
rect 0 626680 39573 627026
rect 0 613520 6278 626680
rect 19408 613520 39573 626680
rect 0 612174 39573 613520
rect 0 611600 20683 612174
rect 36343 612113 36993 612174
rect 0 584400 4843 611600
rect 21003 611200 25993 611854
rect 21003 610200 25993 610600
rect 21003 608920 25993 609880
rect 21003 608200 25993 608600
rect 21003 604920 25993 607880
rect 21003 604200 25993 604600
rect 21003 600920 25993 603880
rect 21003 600200 25993 600600
rect 21003 596920 25993 599880
rect 21003 596200 25993 596600
rect 21003 592920 25993 595880
rect 21003 592200 25993 592600
rect 21003 588920 25993 591880
rect 21003 588200 25993 588600
rect 21003 584920 25993 587880
rect 0 583826 20683 584400
rect 21003 584146 25993 584600
rect 26313 584146 27163 611854
rect 27483 584146 28333 611854
rect 28653 584146 30453 611854
rect 30773 584146 31663 611854
rect 31983 611600 32632 611854
rect 31983 584400 32633 611600
rect 31983 584146 32632 584400
rect 32953 584146 33603 611854
rect 33923 584146 34813 611854
rect 35133 584146 36023 611854
rect 36343 584194 36993 611793
rect 37313 584146 38203 611854
rect 38523 584146 39573 611854
rect 678027 608746 679077 638254
rect 679397 608746 680287 638254
rect 680607 608807 681257 638206
rect 681577 608746 682467 638254
rect 682787 608746 683677 638254
rect 683997 608746 684647 638254
rect 684968 638000 685617 638254
rect 684967 609000 685617 638000
rect 684968 608746 685617 609000
rect 685937 608746 686827 638254
rect 687147 608746 688947 638254
rect 689267 608746 690117 638254
rect 690437 608746 691287 638254
rect 691607 637800 696597 638254
rect 696917 638000 717600 638574
rect 691607 636800 696597 637200
rect 691607 633520 696597 636480
rect 691607 632800 696597 633200
rect 691607 629520 696597 632480
rect 691607 628800 696597 629200
rect 691607 625520 696597 628480
rect 691607 624800 696597 625200
rect 691607 621520 696597 624480
rect 691607 620800 696597 621200
rect 691607 617520 696597 620480
rect 691607 616800 696597 617200
rect 691607 613520 696597 616480
rect 691607 612800 696597 613200
rect 691607 609520 696597 612480
rect 691607 608746 696597 609200
rect 712757 609000 717600 638000
rect 680607 608426 681257 608487
rect 696917 608426 717600 609000
rect 678027 607080 717600 608426
rect 678027 593920 698192 607080
rect 711322 593920 717600 607080
rect 678027 593574 717600 593920
rect 680607 593526 681257 593574
rect 36343 583826 36993 583874
rect 0 583480 39573 583826
rect 0 570320 6278 583480
rect 19408 570320 39573 583480
rect 0 568974 39573 570320
rect 0 568400 20683 568974
rect 36343 568913 36993 568974
rect 0 541200 4843 568400
rect 21003 568000 25993 568654
rect 21003 567000 25993 567400
rect 21003 565720 25993 566680
rect 21003 565000 25993 565400
rect 21003 561720 25993 564680
rect 21003 561000 25993 561400
rect 21003 557720 25993 560680
rect 21003 557000 25993 557400
rect 21003 553720 25993 556680
rect 21003 553000 25993 553400
rect 21003 549720 25993 552680
rect 21003 549000 25993 549400
rect 21003 545720 25993 548680
rect 21003 545000 25993 545400
rect 21003 541720 25993 544680
rect 0 540626 20683 541200
rect 21003 540946 25993 541400
rect 26313 540946 27163 568654
rect 27483 540946 28333 568654
rect 28653 540946 30453 568654
rect 30773 540946 31663 568654
rect 31983 568400 32632 568654
rect 31983 541200 32633 568400
rect 31983 540946 32632 541200
rect 32953 540946 33603 568654
rect 33923 540946 34813 568654
rect 35133 540946 36023 568654
rect 36343 540994 36993 568593
rect 37313 540946 38203 568654
rect 38523 540946 39573 568654
rect 678027 563546 679077 593254
rect 679397 563546 680287 593254
rect 680607 563607 681257 593206
rect 681577 563546 682467 593254
rect 682787 563546 683677 593254
rect 683997 563546 684647 593254
rect 684968 593000 685617 593254
rect 684967 563800 685617 593000
rect 684968 563546 685617 563800
rect 685937 563546 686827 593254
rect 687147 563546 688947 593254
rect 689267 563546 690117 593254
rect 690437 563546 691287 593254
rect 691607 592600 696597 593254
rect 696917 593000 717600 593574
rect 691607 591600 696597 592000
rect 691607 588320 696597 591280
rect 691607 587600 696597 588000
rect 691607 584320 696597 587280
rect 691607 583600 696597 584000
rect 691607 580320 696597 583280
rect 691607 579600 696597 580000
rect 691607 576320 696597 579280
rect 691607 575600 696597 576000
rect 691607 572320 696597 575280
rect 691607 571600 696597 572000
rect 691607 568320 696597 571280
rect 691607 567600 696597 568000
rect 691607 564320 696597 567280
rect 691607 563546 696597 564000
rect 712757 563800 717600 593000
rect 680607 563226 681257 563287
rect 696917 563226 717600 563800
rect 678027 561880 717600 563226
rect 678027 548720 698192 561880
rect 711322 548720 717600 561880
rect 678027 548374 717600 548720
rect 680607 548326 681257 548374
rect 36343 540626 36993 540674
rect 0 540280 39573 540626
rect 0 527120 6278 540280
rect 19408 527120 39573 540280
rect 0 525774 39573 527120
rect 0 525200 20683 525774
rect 36343 525713 36993 525774
rect 0 498000 4843 525200
rect 21003 524800 25993 525454
rect 21003 523800 25993 524200
rect 21003 522520 25993 523480
rect 21003 521800 25993 522200
rect 21003 518520 25993 521480
rect 21003 517800 25993 518200
rect 21003 514520 25993 517480
rect 21003 513800 25993 514200
rect 21003 510520 25993 513480
rect 21003 509800 25993 510200
rect 21003 506520 25993 509480
rect 21003 505800 25993 506200
rect 21003 502520 25993 505480
rect 21003 501800 25993 502200
rect 21003 498520 25993 501480
rect 0 497426 20683 498000
rect 21003 497746 25993 498200
rect 26313 497746 27163 525454
rect 27483 497746 28333 525454
rect 28653 497746 30453 525454
rect 30773 497746 31663 525454
rect 31983 525200 32632 525454
rect 31983 497746 32633 525200
rect 32953 497746 33603 525454
rect 33923 497746 34813 525454
rect 35133 497746 36023 525454
rect 37313 497746 38203 525454
rect 38523 497746 39573 525454
rect 678027 518546 679077 548054
rect 679397 518546 680287 548054
rect 680607 518607 681257 548006
rect 681577 518546 682467 548054
rect 682787 518546 683677 548054
rect 683997 518546 684647 548054
rect 684968 547800 685617 548054
rect 684967 518546 685617 547800
rect 685937 518546 686827 548054
rect 687147 518546 688947 548054
rect 689267 518546 690117 548054
rect 690437 518546 691287 548054
rect 691607 547600 696597 548054
rect 696917 547800 717600 548374
rect 691607 546600 696597 547000
rect 691607 543320 696597 546280
rect 691607 542600 696597 543000
rect 691607 539320 696597 542280
rect 691607 538600 696597 539000
rect 691607 535320 696597 538280
rect 691607 534600 696597 535000
rect 691607 531320 696597 534280
rect 691607 530600 696597 531000
rect 691607 527320 696597 530280
rect 691607 526600 696597 527000
rect 691607 523320 696597 526280
rect 691607 522600 696597 523000
rect 691607 519320 696597 522280
rect 691607 518546 696597 519000
rect 712757 518800 717600 547800
rect 680607 518226 681257 518287
rect 684967 518226 684968 518546
rect 696917 518226 717600 518800
rect 678027 517900 717600 518226
rect 678027 504720 698082 517900
rect 698402 505040 710925 517580
rect 711245 504720 717600 517900
rect 678027 504374 717600 504720
rect 680607 504313 681257 504374
rect 684967 504054 684968 504374
rect 32632 497426 32633 497746
rect 36343 497426 36993 497487
rect 0 497080 39573 497426
rect 0 483900 6355 497080
rect 19518 483900 39573 497080
rect 0 483574 39573 483900
rect 0 483000 20683 483574
rect 32632 483254 32633 483574
rect 36343 483513 36993 483574
rect 0 455800 4843 483000
rect 21003 482600 25993 483254
rect 21003 481600 25993 482000
rect 21003 480320 25993 481280
rect 21003 479600 25993 480000
rect 21003 476320 25993 479280
rect 21003 475600 25993 476000
rect 21003 472320 25993 475280
rect 21003 471600 25993 472000
rect 21003 468320 25993 471280
rect 21003 467600 25993 468000
rect 21003 464320 25993 467280
rect 21003 463600 25993 464000
rect 21003 460320 25993 463280
rect 21003 459600 25993 460000
rect 21003 456320 25993 459280
rect 0 455226 20683 455800
rect 21003 455546 25993 456000
rect 26313 455546 27163 483254
rect 27483 455546 28333 483254
rect 28653 455546 30453 483254
rect 31983 455546 32633 483254
rect 32953 455546 33603 483254
rect 33923 455546 34813 483254
rect 35133 455546 36023 483254
rect 37313 455546 38203 483254
rect 38523 455546 39573 483254
rect 678027 474546 679077 504054
rect 679397 474546 680287 504054
rect 680607 474607 681257 503993
rect 681577 474546 682467 504054
rect 682787 474546 683677 504054
rect 683997 474546 684647 504054
rect 684967 474546 685617 504054
rect 687147 474546 688947 504054
rect 689267 474546 690117 504054
rect 690437 474546 691287 504054
rect 691607 503600 696597 504054
rect 696917 503800 717600 504374
rect 691607 502600 696597 503000
rect 691607 499320 696597 502280
rect 691607 498600 696597 499000
rect 691607 495320 696597 498280
rect 691607 494600 696597 495000
rect 691607 491320 696597 494280
rect 691607 490600 696597 491000
rect 691607 487320 696597 490280
rect 691607 486600 696597 487000
rect 691607 483320 696597 486280
rect 691607 482600 696597 483000
rect 691607 479320 696597 482280
rect 691607 478600 696597 479000
rect 691607 475320 696597 478280
rect 691607 474546 696597 475000
rect 712757 474800 717600 503800
rect 680607 474226 681257 474287
rect 684967 474226 684968 474546
rect 696917 474226 717600 474800
rect 678027 473257 717600 474226
rect 678027 461289 697708 473257
rect 711834 461289 717600 473257
rect 678027 460374 717600 461289
rect 680607 460313 681257 460374
rect 684967 460054 684968 460374
rect 32632 455226 32633 455546
rect 36343 455226 36993 455287
rect 0 454311 39573 455226
rect 0 442343 5766 454311
rect 19892 442343 39573 454311
rect 0 441374 39573 442343
rect 0 440800 20683 441374
rect 32632 441054 32633 441374
rect 36343 441313 36993 441374
rect 0 413600 4843 440800
rect 21003 440400 25993 441054
rect 21003 439400 25993 439800
rect 21003 438120 25993 439080
rect 21003 437400 25993 437800
rect 21003 434120 25993 437080
rect 21003 433400 25993 433800
rect 21003 430120 25993 433080
rect 21003 429400 25993 429800
rect 21003 426120 25993 429080
rect 21003 425400 25993 425800
rect 21003 422120 25993 425080
rect 21003 421400 25993 421800
rect 21003 418120 25993 421080
rect 21003 417400 25993 417800
rect 21003 414120 25993 417080
rect 0 413026 20683 413600
rect 21003 413346 25993 413800
rect 26313 413346 27163 441054
rect 27483 413346 28333 441054
rect 28653 413346 30453 441054
rect 31983 413600 32633 441054
rect 31983 413346 32632 413600
rect 32953 413346 33603 441054
rect 33923 413346 34813 441054
rect 35133 413346 36023 441054
rect 36343 413394 36993 440993
rect 37313 413346 38203 441054
rect 38523 413346 39573 441054
rect 678027 430346 679077 460054
rect 679397 430346 680287 460054
rect 680607 430407 681257 459993
rect 681577 430346 682467 460054
rect 682787 430346 683677 460054
rect 683997 430346 684647 460054
rect 684967 430346 685617 460054
rect 687147 430346 688947 460054
rect 689267 430346 690117 460054
rect 690437 430346 691287 460054
rect 691607 459400 696597 460054
rect 696917 459800 717600 460374
rect 691607 458400 696597 458800
rect 691607 455120 696597 458080
rect 691607 454400 696597 454800
rect 691607 451120 696597 454080
rect 691607 450400 696597 450800
rect 691607 447120 696597 450080
rect 691607 446400 696597 446800
rect 691607 443120 696597 446080
rect 691607 442400 696597 442800
rect 691607 439120 696597 442080
rect 691607 438400 696597 438800
rect 691607 435120 696597 438080
rect 691607 434400 696597 434800
rect 691607 431120 696597 434080
rect 691607 430346 696597 430800
rect 712757 430600 717600 459800
rect 680607 430026 681257 430087
rect 684967 430026 684968 430346
rect 696917 430026 717600 430600
rect 678027 429700 717600 430026
rect 678027 416520 698082 429700
rect 698402 416840 710925 429380
rect 711245 416520 717600 429700
rect 678027 416174 717600 416520
rect 680607 416113 681257 416174
rect 684967 415854 684968 416174
rect 36343 413026 36993 413074
rect 0 412680 39573 413026
rect 0 399520 6278 412680
rect 19408 399520 39573 412680
rect 0 398174 39573 399520
rect 0 397600 20683 398174
rect 36343 398113 36993 398174
rect 0 370400 4843 397600
rect 21003 397200 25993 397854
rect 21003 396200 25993 396600
rect 21003 394920 25993 395880
rect 21003 394200 25993 394600
rect 21003 390920 25993 393880
rect 21003 390200 25993 390600
rect 21003 386920 25993 389880
rect 21003 386200 25993 386600
rect 21003 382920 25993 385880
rect 21003 382200 25993 382600
rect 21003 378920 25993 381880
rect 21003 378200 25993 378600
rect 21003 374920 25993 377880
rect 21003 374200 25993 374600
rect 21003 370920 25993 373880
rect 0 369826 20683 370400
rect 21003 370146 25993 370600
rect 26313 370146 27163 397854
rect 27483 370146 28333 397854
rect 28653 370146 30453 397854
rect 30773 370146 31663 397854
rect 31983 397600 32632 397854
rect 31983 370400 32633 397600
rect 31983 370146 32632 370400
rect 32953 370146 33603 397854
rect 33923 370146 34813 397854
rect 35133 370146 36023 397854
rect 36343 370194 36993 397793
rect 37313 370146 38203 397854
rect 38523 370146 39573 397854
rect 678027 386346 679077 415854
rect 679397 386346 680287 415854
rect 680607 386407 681257 415793
rect 681577 386346 682467 415854
rect 682787 386346 683677 415854
rect 683997 386346 684647 415854
rect 684967 386600 685617 415854
rect 684968 386346 685617 386600
rect 685937 386346 686827 415854
rect 687147 386346 688947 415854
rect 689267 386346 690117 415854
rect 690437 386346 691287 415854
rect 691607 415400 696597 415854
rect 696917 415600 717600 416174
rect 691607 414400 696597 414800
rect 691607 411120 696597 414080
rect 691607 410400 696597 410800
rect 691607 407120 696597 410080
rect 691607 406400 696597 406800
rect 691607 403120 696597 406080
rect 691607 402400 696597 402800
rect 691607 399120 696597 402080
rect 691607 398400 696597 398800
rect 691607 395120 696597 398080
rect 691607 394400 696597 394800
rect 691607 391120 696597 394080
rect 691607 390400 696597 390800
rect 691607 387120 696597 390080
rect 691607 386346 696597 386800
rect 712757 386600 717600 415600
rect 680607 386026 681257 386087
rect 696917 386026 717600 386600
rect 678027 384680 717600 386026
rect 678027 371520 698192 384680
rect 711322 371520 717600 384680
rect 678027 371174 717600 371520
rect 680607 371126 681257 371174
rect 36343 369826 36993 369874
rect 0 369480 39573 369826
rect 0 356320 6278 369480
rect 19408 356320 39573 369480
rect 0 354974 39573 356320
rect 0 354400 20683 354974
rect 36343 354913 36993 354974
rect 0 327200 4843 354400
rect 21003 354000 25993 354654
rect 21003 353000 25993 353400
rect 21003 351720 25993 352680
rect 21003 351000 25993 351400
rect 21003 347720 25993 350680
rect 21003 347000 25993 347400
rect 21003 343720 25993 346680
rect 21003 343000 25993 343400
rect 21003 339720 25993 342680
rect 21003 339000 25993 339400
rect 21003 335720 25993 338680
rect 21003 335000 25993 335400
rect 21003 331720 25993 334680
rect 21003 331000 25993 331400
rect 21003 327720 25993 330680
rect 0 326626 20683 327200
rect 21003 326946 25993 327400
rect 26313 326946 27163 354654
rect 27483 326946 28333 354654
rect 28653 326946 30453 354654
rect 30773 326946 31663 354654
rect 31983 354400 32632 354654
rect 31983 327200 32633 354400
rect 31983 326946 32632 327200
rect 32953 326946 33603 354654
rect 33923 326946 34813 354654
rect 35133 326946 36023 354654
rect 36343 326994 36993 354593
rect 37313 326946 38203 354654
rect 38523 326946 39573 354654
rect 678027 341146 679077 370854
rect 679397 341146 680287 370854
rect 680607 341207 681257 370806
rect 681577 341146 682467 370854
rect 682787 341146 683677 370854
rect 683997 341146 684647 370854
rect 684968 370600 685617 370854
rect 684967 341400 685617 370600
rect 684968 341146 685617 341400
rect 685937 341146 686827 370854
rect 687147 341146 688947 370854
rect 689267 341146 690117 370854
rect 690437 341146 691287 370854
rect 691607 370200 696597 370854
rect 696917 370600 717600 371174
rect 691607 369200 696597 369600
rect 691607 365920 696597 368880
rect 691607 365200 696597 365600
rect 691607 361920 696597 364880
rect 691607 361200 696597 361600
rect 691607 357920 696597 360880
rect 691607 357200 696597 357600
rect 691607 353920 696597 356880
rect 691607 353200 696597 353600
rect 691607 349920 696597 352880
rect 691607 349200 696597 349600
rect 691607 345920 696597 348880
rect 691607 345200 696597 345600
rect 691607 341920 696597 344880
rect 691607 341146 696597 341600
rect 712757 341400 717600 370600
rect 680607 340826 681257 340887
rect 696917 340826 717600 341400
rect 678027 339480 717600 340826
rect 36343 326626 36993 326674
rect 0 326280 39573 326626
rect 0 313120 6278 326280
rect 19408 313120 39573 326280
rect 678027 326320 698192 339480
rect 711322 326320 717600 339480
rect 678027 325974 717600 326320
rect 680607 325926 681257 325974
rect 0 311774 39573 313120
rect 0 311200 20683 311774
rect 36343 311713 36993 311774
rect 0 284000 4843 311200
rect 21003 310800 25993 311454
rect 21003 309800 25993 310200
rect 21003 308520 25993 309480
rect 21003 307800 25993 308200
rect 21003 304520 25993 307480
rect 21003 303800 25993 304200
rect 21003 300520 25993 303480
rect 21003 299800 25993 300200
rect 21003 296520 25993 299480
rect 21003 295800 25993 296200
rect 21003 292520 25993 295480
rect 21003 291800 25993 292200
rect 21003 288520 25993 291480
rect 21003 287800 25993 288200
rect 21003 284520 25993 287480
rect 0 283426 20683 284000
rect 21003 283746 25993 284200
rect 26313 283746 27163 311454
rect 27483 283746 28333 311454
rect 28653 283746 30453 311454
rect 30773 283746 31663 311454
rect 31983 311200 32632 311454
rect 31983 284000 32633 311200
rect 31983 283746 32632 284000
rect 32953 283746 33603 311454
rect 33923 283746 34813 311454
rect 35133 283746 36023 311454
rect 36343 283794 36993 311393
rect 37313 283746 38203 311454
rect 38523 283746 39573 311454
rect 678027 296146 679077 325654
rect 679397 296146 680287 325654
rect 680607 296207 681257 325606
rect 681577 296146 682467 325654
rect 682787 296146 683677 325654
rect 683997 296146 684647 325654
rect 684968 325400 685617 325654
rect 684967 296400 685617 325400
rect 684968 296146 685617 296400
rect 685937 296146 686827 325654
rect 687147 296146 688947 325654
rect 689267 296146 690117 325654
rect 690437 296146 691287 325654
rect 691607 325200 696597 325654
rect 696917 325400 717600 325974
rect 691607 324200 696597 324600
rect 691607 320920 696597 323880
rect 691607 320200 696597 320600
rect 691607 316920 696597 319880
rect 691607 316200 696597 316600
rect 691607 312920 696597 315880
rect 691607 312200 696597 312600
rect 691607 308920 696597 311880
rect 691607 308200 696597 308600
rect 691607 304920 696597 307880
rect 691607 304200 696597 304600
rect 691607 300920 696597 303880
rect 691607 300200 696597 300600
rect 691607 296920 696597 299880
rect 691607 296146 696597 296600
rect 712757 296400 717600 325400
rect 680607 295826 681257 295887
rect 696917 295826 717600 296400
rect 678027 294480 717600 295826
rect 36343 283426 36993 283474
rect 0 283080 39573 283426
rect 0 269920 6278 283080
rect 19408 269920 39573 283080
rect 678027 281320 698192 294480
rect 711322 281320 717600 294480
rect 678027 280974 717600 281320
rect 680607 280926 681257 280974
rect 0 268574 39573 269920
rect 0 268000 20683 268574
rect 36343 268513 36993 268574
rect 0 240800 4843 268000
rect 21003 267600 25993 268254
rect 21003 266600 25993 267000
rect 21003 265320 25993 266280
rect 21003 264600 25993 265000
rect 21003 261320 25993 264280
rect 21003 260600 25993 261000
rect 21003 257320 25993 260280
rect 21003 256600 25993 257000
rect 21003 253320 25993 256280
rect 21003 252600 25993 253000
rect 21003 249320 25993 252280
rect 21003 248600 25993 249000
rect 21003 245320 25993 248280
rect 21003 244600 25993 245000
rect 21003 241320 25993 244280
rect 0 240226 20683 240800
rect 21003 240546 25993 241000
rect 26313 240546 27163 268254
rect 27483 240546 28333 268254
rect 28653 240546 30453 268254
rect 30773 240546 31663 268254
rect 31983 268000 32632 268254
rect 31983 240800 32633 268000
rect 31983 240546 32632 240800
rect 32953 240546 33603 268254
rect 33923 240546 34813 268254
rect 35133 240546 36023 268254
rect 36343 240594 36993 268193
rect 37313 240546 38203 268254
rect 38523 240546 39573 268254
rect 678027 251146 679077 280654
rect 679397 251146 680287 280654
rect 680607 251207 681257 280606
rect 681577 251146 682467 280654
rect 682787 251146 683677 280654
rect 683997 251146 684647 280654
rect 684968 280400 685617 280654
rect 684967 251400 685617 280400
rect 684968 251146 685617 251400
rect 685937 251146 686827 280654
rect 687147 251146 688947 280654
rect 689267 251146 690117 280654
rect 690437 251146 691287 280654
rect 691607 280200 696597 280654
rect 696917 280400 717600 280974
rect 691607 279200 696597 279600
rect 691607 275920 696597 278880
rect 691607 275200 696597 275600
rect 691607 271920 696597 274880
rect 691607 271200 696597 271600
rect 691607 267920 696597 270880
rect 691607 267200 696597 267600
rect 691607 263920 696597 266880
rect 691607 263200 696597 263600
rect 691607 259920 696597 262880
rect 691607 259200 696597 259600
rect 691607 255920 696597 258880
rect 691607 255200 696597 255600
rect 691607 251920 696597 254880
rect 691607 251146 696597 251600
rect 712757 251400 717600 280400
rect 680607 250826 681257 250887
rect 696917 250826 717600 251400
rect 678027 249480 717600 250826
rect 36343 240226 36993 240274
rect 0 239880 39573 240226
rect 0 226720 6278 239880
rect 19408 226720 39573 239880
rect 678027 236320 698192 249480
rect 711322 236320 717600 249480
rect 678027 235974 717600 236320
rect 680607 235926 681257 235974
rect 0 225374 39573 226720
rect 0 224800 20683 225374
rect 36343 225313 36993 225374
rect 0 197600 4843 224800
rect 21003 224400 25993 225054
rect 21003 223400 25993 223800
rect 21003 222120 25993 223080
rect 21003 221400 25993 221800
rect 21003 218120 25993 221080
rect 21003 217400 25993 217800
rect 21003 214120 25993 217080
rect 21003 213400 25993 213800
rect 21003 210120 25993 213080
rect 21003 209400 25993 209800
rect 21003 206120 25993 209080
rect 21003 205400 25993 205800
rect 21003 202120 25993 205080
rect 21003 201400 25993 201800
rect 21003 198120 25993 201080
rect 0 197026 20683 197600
rect 21003 197346 25993 197800
rect 26313 197346 27163 225054
rect 27483 197346 28333 225054
rect 28653 197346 30453 225054
rect 30773 197346 31663 225054
rect 31983 224800 32632 225054
rect 31983 197600 32633 224800
rect 31983 197346 32632 197600
rect 32953 197346 33603 225054
rect 33923 197346 34813 225054
rect 35133 197346 36023 225054
rect 36343 197394 36993 224993
rect 37313 197346 38203 225054
rect 38523 197346 39573 225054
rect 678027 205946 679077 235654
rect 679397 205946 680287 235654
rect 680607 206007 681257 235606
rect 681577 205946 682467 235654
rect 682787 205946 683677 235654
rect 683997 205946 684647 235654
rect 684968 235400 685617 235654
rect 684967 206200 685617 235400
rect 684968 205946 685617 206200
rect 685937 205946 686827 235654
rect 687147 205946 688947 235654
rect 689267 205946 690117 235654
rect 690437 205946 691287 235654
rect 691607 235000 696597 235654
rect 696917 235400 717600 235974
rect 691607 234000 696597 234400
rect 691607 230720 696597 233680
rect 691607 230000 696597 230400
rect 691607 226720 696597 229680
rect 691607 226000 696597 226400
rect 691607 222720 696597 225680
rect 691607 222000 696597 222400
rect 691607 218720 696597 221680
rect 691607 218000 696597 218400
rect 691607 214720 696597 217680
rect 691607 214000 696597 214400
rect 691607 210720 696597 213680
rect 691607 210000 696597 210400
rect 691607 206720 696597 209680
rect 691607 205946 696597 206400
rect 712757 206200 717600 235400
rect 680607 205626 681257 205687
rect 696917 205626 717600 206200
rect 678027 204280 717600 205626
rect 36343 197026 36993 197074
rect 0 196680 39573 197026
rect 0 183520 6278 196680
rect 19408 183520 39573 196680
rect 678027 191120 698192 204280
rect 711322 191120 717600 204280
rect 678027 190774 717600 191120
rect 680607 190726 681257 190774
rect 0 182174 39573 183520
rect 0 181600 20683 182174
rect 36343 182113 36993 182174
rect 0 125200 4843 181600
rect 21003 181200 25993 181854
rect 21003 180200 25993 180600
rect 21003 178920 25993 179880
rect 21003 178200 25993 178600
rect 21003 174920 25993 177880
rect 21003 174200 25993 174600
rect 21003 170920 25993 173880
rect 21003 170200 25993 170600
rect 21003 166920 25993 169880
rect 21003 166200 25993 166600
rect 21003 162920 25993 165880
rect 21003 162200 25993 162600
rect 21003 158920 25993 161880
rect 21003 158200 25993 158600
rect 21003 154920 25993 157880
rect 21003 152000 25993 154600
rect 21003 151000 25993 151400
rect 21003 149720 25993 150680
rect 21003 149000 25993 149400
rect 21003 145720 25993 148680
rect 21003 145000 25993 145400
rect 21003 141720 25993 144680
rect 21003 141000 25993 141400
rect 21003 137720 25993 140680
rect 21003 137000 25993 137400
rect 21003 133720 25993 136680
rect 21003 133000 25993 133400
rect 21003 129720 25993 132680
rect 21003 129000 25993 129400
rect 21003 125720 25993 128680
rect 0 124626 20683 125200
rect 26313 124946 27163 181854
rect 27483 124946 28333 181854
rect 28653 153400 30453 181854
rect 30773 154400 31663 181854
rect 31983 181600 32632 181854
rect 31983 153400 32633 181600
rect 28653 124946 30453 152400
rect 30773 124946 31663 153400
rect 31983 124946 32633 152400
rect 32953 124946 33603 181854
rect 33923 124946 34813 181854
rect 36343 153400 36993 181793
rect 37313 154400 38203 181854
rect 36343 125007 36993 152400
rect 37313 124946 38203 153400
rect 38523 124946 39573 181854
rect 678027 160946 679077 190454
rect 679397 160946 680287 190454
rect 680607 161007 681257 190406
rect 681577 160946 682467 190454
rect 682787 160946 683677 190454
rect 683997 160946 684647 190454
rect 684968 190200 685617 190454
rect 684967 161200 685617 190200
rect 684968 160946 685617 161200
rect 685937 160946 686827 190454
rect 687147 160946 688947 190454
rect 689267 160946 690117 190454
rect 690437 160946 691287 190454
rect 691607 190000 696597 190454
rect 696917 190200 717600 190774
rect 691607 189000 696597 189400
rect 691607 185720 696597 188680
rect 691607 185000 696597 185400
rect 691607 181720 696597 184680
rect 691607 181000 696597 181400
rect 691607 177720 696597 180680
rect 691607 177000 696597 177400
rect 691607 173720 696597 176680
rect 691607 173000 696597 173400
rect 691607 169720 696597 172680
rect 691607 169000 696597 169400
rect 691607 165720 696597 168680
rect 691607 165000 696597 165400
rect 691607 161720 696597 164680
rect 691607 160946 696597 161400
rect 712757 161200 717600 190200
rect 680607 160626 681257 160687
rect 696917 160626 717600 161200
rect 678027 159280 717600 160626
rect 678027 146120 698192 159280
rect 711322 146120 717600 159280
rect 678027 145774 717600 146120
rect 680607 145726 681257 145774
rect 32632 124626 32633 124946
rect 36343 124626 36993 124687
rect 0 124280 39573 124626
rect 0 111100 6355 124280
rect 19518 111100 39573 124280
rect 678027 115746 679077 145454
rect 679397 115746 680287 145454
rect 680607 115807 681257 145406
rect 681577 115746 682467 145454
rect 682787 115746 683677 145454
rect 683997 115746 684647 145454
rect 684968 145200 685617 145454
rect 684967 116000 685617 145200
rect 684968 115746 685617 116000
rect 685937 115746 686827 145454
rect 687147 115746 688947 145454
rect 689267 115746 690117 145454
rect 690437 115746 691287 145454
rect 691607 144800 696597 145454
rect 696917 145200 717600 145774
rect 691607 143800 696597 144200
rect 691607 140520 696597 143480
rect 691607 139800 696597 140200
rect 691607 136520 696597 139480
rect 691607 135800 696597 136200
rect 691607 132520 696597 135480
rect 691607 131800 696597 132200
rect 691607 128520 696597 131480
rect 691607 127800 696597 128200
rect 691607 124520 696597 127480
rect 691607 123800 696597 124200
rect 691607 120520 696597 123480
rect 691607 119800 696597 120200
rect 691607 116520 696597 119480
rect 691607 115746 696597 116200
rect 712757 116000 717600 145200
rect 680607 115426 681257 115487
rect 696917 115426 717600 116000
rect 0 110774 39573 111100
rect 678027 114080 717600 115426
rect 0 110200 20683 110774
rect 32632 110454 32633 110774
rect 36343 110713 36993 110774
rect 0 83000 4843 110200
rect 21003 108800 25993 109200
rect 21003 107520 25993 108480
rect 21003 106800 25993 107200
rect 21003 103520 25993 106480
rect 21003 102800 25993 103200
rect 21003 99520 25993 102480
rect 21003 98800 25993 99200
rect 21003 95520 25993 98480
rect 21003 94800 25993 95200
rect 21003 91520 25993 94480
rect 21003 90800 25993 91200
rect 21003 87520 25993 90480
rect 21003 86800 25993 87200
rect 21003 83520 25993 86480
rect 0 82426 20683 83000
rect 21003 82746 25993 83200
rect 26313 82746 27163 110454
rect 27483 82746 28333 110454
rect 28653 82746 30453 110454
rect 30773 82746 31663 110454
rect 31983 83000 32633 110454
rect 31983 82746 32632 83000
rect 32953 82746 33603 110454
rect 33923 82746 34813 110454
rect 36343 82807 36993 110393
rect 38523 82746 39573 110454
rect 678027 100920 698192 114080
rect 711322 100920 717600 114080
rect 678027 100574 717600 100920
rect 680607 100526 681257 100574
rect 36343 82426 36993 82487
rect 0 81511 39573 82426
rect 0 69543 5766 81511
rect 19892 69543 39573 81511
rect 0 68574 39573 69543
rect 0 68000 20683 68574
rect 36343 68513 36993 68574
rect 0 40800 4843 68000
rect 21003 67600 25993 68254
rect 21003 66600 25993 67000
rect 21003 65320 25993 66280
rect 21003 64600 25993 65000
rect 21003 61320 25993 64280
rect 21003 60600 25993 61000
rect 21003 57320 25993 60280
rect 21003 56600 25993 57000
rect 21003 53320 25993 56280
rect 21003 52600 25993 53000
rect 21003 49320 25993 52280
rect 21003 48600 25993 49000
rect 21003 45320 25993 48280
rect 21003 44600 25993 45000
rect 21003 41320 25993 44280
rect 0 40109 20683 40800
rect 21003 40429 25993 41000
rect 26313 40546 27163 68254
rect 27483 40546 28333 68254
rect 26313 40109 28333 40226
rect 0 35049 28333 40109
rect 28653 35369 30453 68254
rect 30773 40546 31663 68254
rect 31983 68000 32632 68254
rect 31983 40800 32633 68000
rect 31983 40546 32632 40800
rect 32953 40546 33603 68254
rect 33923 40546 34813 68254
rect 35133 40546 36023 68254
rect 36343 40549 36993 68193
rect 38523 40546 39573 68254
rect 36343 40226 36993 40229
rect 39893 40226 40000 40800
rect 30773 39893 40000 40226
rect 676800 39893 677707 40000
rect 30773 38523 39210 39893
rect 39573 39573 39680 39893
tri 39680 39573 40000 39893 sw
rect 677374 39680 677707 39893
tri 677707 39680 678027 40000 se
rect 678027 39680 679077 100254
rect 679397 71000 680287 100254
rect 680607 70000 681257 100206
rect 677374 39573 679077 39680
rect 39530 38523 79054 39573
rect 30773 36993 38923 38523
rect 47400 38203 71400 38523
rect 39243 37313 79054 38203
rect 79374 36993 93226 39573
rect 93546 38523 132854 39573
rect 101200 38203 125200 38523
rect 93546 37313 132854 38203
rect 133174 36993 147026 39573
rect 147346 38523 186654 39573
rect 155000 38203 179000 38523
rect 147346 37313 186654 38203
rect 186974 36993 201826 39573
rect 202146 38523 241454 39573
rect 209800 38203 233800 38523
rect 202146 37313 241454 38203
rect 241774 36993 255626 39573
rect 255946 38523 295254 39573
rect 263600 38203 287600 38523
rect 255946 37313 295254 38203
rect 295574 36993 310426 39573
rect 310746 38523 350054 39573
rect 318400 38203 342400 38523
rect 310746 37313 350054 38203
rect 350374 36993 365226 39573
rect 365546 38523 404854 39573
rect 373200 38203 397200 38523
rect 365546 37313 404854 38203
rect 405174 36993 420026 39573
rect 420346 38523 459654 39573
rect 428000 38203 452000 38523
rect 420346 37313 459654 38203
rect 459974 36993 474826 39573
rect 475146 38523 514454 39573
rect 482800 38203 506800 38523
rect 475146 37313 514454 38203
rect 514774 36993 529626 39573
rect 529946 38523 569254 39573
rect 537600 38203 561600 38523
rect 529946 37313 569254 38203
rect 569574 36993 583426 39573
rect 583746 38523 623054 39573
rect 591400 38203 615400 38523
rect 583746 37313 623054 38203
rect 623374 36993 637226 39573
rect 637546 38523 677054 39573
rect 677374 39210 677707 39573
rect 678027 39530 679077 39573
rect 679397 39243 680287 70000
rect 680607 39706 681257 69000
rect 681577 39695 682467 100254
rect 682787 39680 683677 100254
rect 683997 39723 684647 100254
rect 684968 100000 685617 100254
rect 684967 70000 685617 100000
rect 685937 71000 686827 100254
rect 687147 70000 688947 100254
rect 684967 39733 685617 69000
rect 685937 39705 686827 70000
rect 684967 39403 685617 39413
rect 680607 39375 681257 39386
rect 683997 39385 685617 39403
rect 680607 39360 682467 39375
rect 683997 39360 686827 39385
rect 677374 38923 679077 39210
rect 680607 38923 686827 39360
rect 645200 38203 669200 38523
rect 637546 37313 677054 38203
rect 677374 36993 686827 38923
rect 30773 36343 39386 36993
rect 39706 36343 78993 36993
rect 79313 36343 93287 36993
rect 93607 36343 132793 36993
rect 133113 36343 147087 36993
rect 147407 36343 186606 36993
rect 186926 36343 201887 36993
rect 202207 36343 241393 36993
rect 241713 36343 255687 36993
rect 256007 36343 295206 36993
rect 295526 36343 310487 36993
rect 310807 36343 350006 36993
rect 350326 36343 365287 36993
rect 365607 36343 404806 36993
rect 405126 36343 420087 36993
rect 420407 36343 459606 36993
rect 459926 36343 474887 36993
rect 475207 36343 514406 36993
rect 514726 36343 529687 36993
rect 530007 36343 569193 36993
rect 569513 36343 583487 36993
rect 623313 36343 637287 36993
rect 677371 36343 686827 36993
rect 30773 35133 39375 36343
rect 39695 35133 79054 36023
rect 30773 35049 39360 35133
rect 0 33603 39360 35049
rect 39680 33923 79054 34813
rect 0 32633 39403 33603
rect 39723 32953 79054 33603
rect 79374 32633 93226 36343
rect 93546 35133 132854 36023
rect 93546 33923 132854 34813
rect 93546 32953 132854 33603
rect 0 31983 39413 32633
rect 78800 32632 93800 32633
rect 0 30773 39385 31983
rect 39705 30773 79054 31663
rect 0 28333 35049 30773
rect 0 27163 39355 28333
rect 39675 27483 79054 28333
rect 0 26313 39384 27163
rect 39704 26313 79054 27163
rect 0 20683 39151 26313
rect 39471 21003 40200 25993
rect 40520 21003 43480 25993
rect 43800 21003 44200 25993
rect 44520 21003 45480 25993
rect 45800 21003 46200 25993
rect 46800 21003 71600 25993
rect 71920 21003 74880 25993
rect 75200 21003 75600 25993
rect 75920 21003 76880 25993
rect 77200 21003 77600 25993
rect 78200 21003 79054 25993
rect 79374 20683 93226 32632
rect 93546 30773 132854 31663
rect 93546 27483 132854 28333
rect 93546 26313 132854 27163
rect 93546 21003 94000 25993
rect 94320 21003 97280 25993
rect 97600 21003 98000 25993
rect 98320 21003 99280 25993
rect 99600 21003 100000 25993
rect 100600 21003 125400 25993
rect 125720 21003 128680 25993
rect 129000 21003 129400 25993
rect 129720 21003 130680 25993
rect 131000 21003 131400 25993
rect 132000 21003 132854 25993
rect 133174 20683 147026 36343
rect 147346 35133 186654 36023
rect 147346 33923 186654 34813
rect 147346 32953 186654 33603
rect 147600 32632 186400 32633
rect 147346 31983 186654 32632
rect 147346 30773 186654 31663
rect 147346 28653 186654 30453
rect 147346 27483 186654 28333
rect 147346 26313 186654 27163
rect 147346 21003 147800 25993
rect 148120 21003 151080 25993
rect 151400 21003 151800 25993
rect 152120 21003 153080 25993
rect 153400 21003 153800 25993
rect 154400 21003 179200 25993
rect 179520 21003 182480 25993
rect 182800 21003 183200 25993
rect 183520 21003 184480 25993
rect 184800 21003 185200 25993
rect 185800 21003 186654 25993
rect 186974 20683 201826 36343
rect 202146 35133 241454 36023
rect 202146 33923 241454 34813
rect 202146 32953 241454 33603
rect 202400 32632 241200 32633
rect 202146 31983 241454 32632
rect 202146 28653 241454 30453
rect 202146 27483 241454 28333
rect 202146 26313 241454 27163
rect 202146 21003 202600 25993
rect 202920 21003 205880 25993
rect 206200 21003 206600 25993
rect 206920 21003 207880 25993
rect 208200 21003 208600 25993
rect 209200 21003 234000 25993
rect 234320 21003 237280 25993
rect 237600 21003 238000 25993
rect 238320 21003 239280 25993
rect 239600 21003 240000 25993
rect 240600 21003 241454 25993
rect 241774 20683 255626 36343
rect 255946 35133 295254 36023
rect 255946 33923 295254 34813
rect 255946 32953 295254 33603
rect 256200 32632 295000 32633
rect 255946 31983 295254 32632
rect 255946 28653 295254 30453
rect 255946 27483 295254 28333
rect 255946 26313 295254 27163
rect 255946 21003 256400 25993
rect 256720 21003 259680 25993
rect 260000 21003 260400 25993
rect 260720 21003 261680 25993
rect 262000 21003 262400 25993
rect 263000 21003 287800 25993
rect 288120 21003 291080 25993
rect 291400 21003 291800 25993
rect 292120 21003 293080 25993
rect 293400 21003 293800 25993
rect 294400 21003 295254 25993
rect 295574 20683 310426 36343
rect 310746 35133 350054 36023
rect 310746 33923 350054 34813
rect 310746 32953 350054 33603
rect 311000 32632 349800 32633
rect 310746 31983 350054 32632
rect 310746 30773 350054 31663
rect 310746 28653 350054 30453
rect 310746 27483 350054 28333
rect 310746 26313 350054 27163
rect 310746 21003 311200 25993
rect 311520 21003 314480 25993
rect 314800 21003 315200 25993
rect 315520 21003 316480 25993
rect 316800 21003 317200 25993
rect 317800 21003 342600 25993
rect 342920 21003 345880 25993
rect 346200 21003 346600 25993
rect 346920 21003 347880 25993
rect 348200 21003 348600 25993
rect 349200 21003 350054 25993
rect 350374 20683 365226 36343
rect 365546 35133 404854 36023
rect 365546 33923 404854 34813
rect 365546 32953 404854 33603
rect 365800 32632 404600 32633
rect 365546 31983 404854 32632
rect 365546 30773 404854 31663
rect 365546 28653 404854 30453
rect 365546 27483 404854 28333
rect 365546 26313 404854 27163
rect 365546 21003 366000 25993
rect 366320 21003 369280 25993
rect 369600 21003 370000 25993
rect 370320 21003 371280 25993
rect 371600 21003 372000 25993
rect 372600 21003 397400 25993
rect 397720 21003 400680 25993
rect 401000 21003 401400 25993
rect 401720 21003 402680 25993
rect 403000 21003 403400 25993
rect 404000 21003 404854 25993
rect 405174 20683 420026 36343
rect 420346 35133 459654 36023
rect 420346 33923 459654 34813
rect 420346 32953 459654 33603
rect 420600 32632 459400 32633
rect 420346 31983 459654 32632
rect 420346 30773 459654 31663
rect 420346 28653 459654 30453
rect 420346 27483 459654 28333
rect 420346 26313 459654 27163
rect 420346 21003 420800 25993
rect 421120 21003 424080 25993
rect 424400 21003 424800 25993
rect 425120 21003 426080 25993
rect 426400 21003 426800 25993
rect 427400 21003 452200 25993
rect 452520 21003 455480 25993
rect 455800 21003 456200 25993
rect 456520 21003 457480 25993
rect 457800 21003 458200 25993
rect 458800 21003 459654 25993
rect 459974 20683 474826 36343
rect 475146 35133 514454 36023
rect 475146 33923 514454 34813
rect 475146 32953 514454 33603
rect 475400 32632 514200 32633
rect 475146 31983 514454 32632
rect 475146 30773 514454 31663
rect 475146 28653 514454 30453
rect 475146 27483 514454 28333
rect 475146 26313 514454 27163
rect 475146 21003 475600 25993
rect 475920 21003 478880 25993
rect 479200 21003 479600 25993
rect 479920 21003 480880 25993
rect 481200 21003 481600 25993
rect 482200 21003 507000 25993
rect 507320 21003 510280 25993
rect 510600 21003 511000 25993
rect 511320 21003 512280 25993
rect 512600 21003 513000 25993
rect 513600 21003 514454 25993
rect 514774 20683 529626 36343
rect 529946 35133 569254 36023
rect 529946 33923 569254 34813
rect 529946 32953 569254 33603
rect 569574 32633 583426 36343
rect 583746 35133 623054 36023
rect 583746 33923 623054 34813
rect 583746 32953 623054 33603
rect 623374 32633 637226 36343
rect 637546 35133 677054 36023
rect 677374 35049 686827 36343
rect 687147 35369 688947 69000
rect 689267 39675 690117 100254
rect 690437 39704 691287 100254
rect 691607 99800 696597 100254
rect 696917 100000 717600 100574
rect 691607 98800 696597 99200
rect 691607 95520 696597 98480
rect 691607 94800 696597 95200
rect 691607 91520 696597 94480
rect 691607 90800 696597 91200
rect 691607 87520 696597 90480
rect 691607 86800 696597 87200
rect 691607 83520 696597 86480
rect 691607 82800 696597 83200
rect 691607 79520 696597 82480
rect 691607 78800 696597 79200
rect 691607 75520 696597 78480
rect 691607 74800 696597 75200
rect 691607 71520 696597 74480
rect 691607 68800 696597 71200
rect 691607 67800 696597 68200
rect 691607 64520 696597 67480
rect 691607 63800 696597 64200
rect 691607 60520 696597 63480
rect 691607 59800 696597 60200
rect 691607 56520 696597 59480
rect 691607 55800 696597 56200
rect 691607 52520 696597 55480
rect 691607 51800 696597 52200
rect 691607 48520 696597 51480
rect 691607 47800 696597 48200
rect 691607 44520 696597 47480
rect 691607 43800 696597 44200
rect 691607 40520 696597 43480
rect 691607 39471 696597 40200
rect 712757 40000 717600 100000
rect 690437 39355 691287 39384
rect 689267 39151 691287 39355
rect 696917 39151 717600 40000
rect 689267 35049 717600 39151
rect 637546 33923 677054 34813
rect 637546 32953 677054 33603
rect 530200 32632 676800 32633
rect 529946 31983 569254 32632
rect 529946 30773 569254 31663
rect 529946 28653 569254 30453
rect 529946 27483 569254 28333
rect 529946 26313 569254 27163
rect 529946 21003 530400 25993
rect 530720 21003 533680 25993
rect 534000 21003 534400 25993
rect 534720 21003 535680 25993
rect 536000 21003 536400 25993
rect 537000 21003 561800 25993
rect 562120 21003 565080 25993
rect 565400 21003 565800 25993
rect 566120 21003 567080 25993
rect 567400 21003 567800 25993
rect 568400 21003 569254 25993
rect 569574 20683 583426 32632
rect 583746 31983 623054 32632
rect 583746 30773 623054 31663
rect 583746 28653 623054 30453
rect 583746 27483 623054 28333
rect 583746 26313 623054 27163
rect 583746 21003 584200 25993
rect 584520 21003 587480 25993
rect 587800 21003 588200 25993
rect 588520 21003 589480 25993
rect 589800 21003 590200 25993
rect 590800 21003 615600 25993
rect 615920 21003 618880 25993
rect 619200 21003 619600 25993
rect 619920 21003 620880 25993
rect 621200 21003 621600 25993
rect 622200 21003 623054 25993
rect 623374 20683 637226 32632
rect 637546 31983 677054 32632
rect 637546 30773 677054 31663
rect 677374 30773 717600 35049
rect 637546 28653 682231 30453
rect 682551 28333 717600 30773
rect 637546 27483 677054 28333
rect 637546 26313 677054 27163
rect 677374 26313 717600 28333
rect 637546 21003 638000 25993
rect 638320 21003 641280 25993
rect 641600 21003 642000 25993
rect 642320 21003 643280 25993
rect 643600 21003 644000 25993
rect 644600 21003 669400 25993
rect 669720 21003 672680 25993
rect 673000 21003 673400 25993
rect 673720 21003 674680 25993
rect 675000 21003 675400 25993
rect 676000 21003 677171 25993
rect 677491 20683 717600 26313
rect 0 4843 40000 20683
rect 78800 19518 93800 20683
rect 78800 6355 79720 19518
rect 92900 6355 93800 19518
rect 78800 4843 93800 6355
rect 132600 18629 147600 20683
rect 132600 6823 136393 18629
rect 144470 6823 147600 18629
rect 132600 5163 147600 6823
rect 186400 19408 202400 20683
rect 186400 6278 187320 19408
rect 200480 6278 202400 19408
rect 0 0 132854 4843
rect 133174 0 147026 5163
rect 186400 4843 202400 6278
rect 241200 19892 256200 20683
rect 241200 5766 242689 19892
rect 254657 5766 256200 19892
rect 241200 4843 256200 5766
rect 295000 19408 311000 20683
rect 295000 6278 295920 19408
rect 309080 6278 311000 19408
rect 295000 4843 311000 6278
rect 349800 19408 365800 20683
rect 349800 6278 350720 19408
rect 363880 6278 365800 19408
rect 349800 4843 365800 6278
rect 404600 19408 420600 20683
rect 404600 6278 405520 19408
rect 418680 6278 420600 19408
rect 404600 4843 420600 6278
rect 459400 19408 475400 20683
rect 459400 6278 460320 19408
rect 473480 6278 475400 19408
rect 459400 4843 475400 6278
rect 514200 19408 530200 20683
rect 514200 6278 515120 19408
rect 528280 6278 530200 19408
rect 514200 4843 530200 6278
rect 569000 19518 584000 20683
rect 569000 6355 569920 19518
rect 583100 6355 584000 19518
rect 569000 4843 584000 6355
rect 622800 19518 637800 20683
rect 622800 6355 623720 19518
rect 636900 6355 637800 19518
rect 622800 4843 637800 6355
rect 676800 4843 717600 20683
rect 147346 0 717600 4843
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 1 nsew signal input
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 2 nsew signal output
rlabel metal2 s 194043 41713 194099 42193 6 por
port 3 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 4 nsew signal output
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 5 nsew signal input
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 6 nsew signal input
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 7 nsew signal input
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 8 nsew signal output
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 9 nsew signal input
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 10 nsew signal input
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 11 nsew signal input
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 12 nsew signal bidirectional
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 13 nsew signal output
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 14 nsew signal input
rlabel metal2 s 415371 41713 415427 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41754 415268 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415216 41806 415427 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412364 41754 412416 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41713 412299 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41806 412416 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409328 41754 409380 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41713 409263 41806 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41806 409380 41818 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415228 41818 415427 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41818 412404 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41818 409368 41834 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 415371 41834 415427 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 412243 41834 412299 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 409207 41834 409263 42193 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 415216 41760 415268 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 412364 41760 412416 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel via1 s 409328 41760 409380 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41760 415274 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41760 412422 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41760 409386 41772 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41772 415274 41800 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 415210 41800 415274 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 412358 41800 412422 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal1 s 409322 41800 409386 41812 6 flash_io0_ieb_core
port 15 nsew signal input
rlabel metal2 s 419695 41713 419751 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41713 411103 41820 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419695 41820 419764 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411047 41820 411116 42193 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419736 42193 419764 44202 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411088 42193 411116 44202 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 419724 44202 419776 44266 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal2 s 411076 44202 411128 44266 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via1 s 419724 44208 419776 44260 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel via1 s 411076 44208 411128 44260 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal1 s 419718 44208 419782 44220 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal1 s 411070 44208 411134 44220 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal1 s 411070 44220 419782 44248 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal1 s 419718 44248 419782 44260 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal1 s 411070 44248 411134 44260 6 flash_io0_oeb_core
port 16 nsew signal input
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 17 nsew signal bidirectional
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 18 nsew signal output
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 19 nsew signal input
rlabel metal2 s 470171 41713 470227 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41713 467099 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41713 464063 41806 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470060 41806 470227 41822 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41806 467236 41822 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41806 464200 41822 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41822 470227 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470171 41834 470227 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 470048 41834 470100 41886 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41822 467248 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467196 41834 467248 41886 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 467043 41834 467099 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41822 464212 41834 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464160 41834 464212 41886 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal2 s 464007 41834 464063 42193 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 470048 41828 470100 41880 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 467196 41828 467248 41880 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel via1 s 464160 41828 464212 41880 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41828 470106 41840 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41828 467254 41840 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41828 464218 41840 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41840 470106 41868 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 470042 41868 470106 41880 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 467190 41868 467254 41880 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal1 s 464154 41868 464218 41880 6 flash_io1_ieb_core
port 20 nsew signal input
rlabel metal3 s 474457 44235 474523 44238 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44235 465875 44238 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44238 474523 44298 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 474457 44298 474523 44301 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal3 s 465809 44298 465875 44301 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 474462 44240 474518 44296 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel via2 s 465814 44240 465870 44296 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474495 41713 474551 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465847 41713 465903 41806 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 41806 474551 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 41806 465903 42193 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474476 42193 474504 44231 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465828 42193 465856 44231 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 474462 44231 474518 44305 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal2 s 465814 44231 465870 44305 6 flash_io1_oeb_core
port 21 nsew signal input
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 22 nsew signal bidirectional
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 23 nsew signal output
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 24 nsew signal input
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 25 nsew signal input
rlabel metal3 s 524965 44235 525031 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44235 518867 44238 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44238 525031 44298 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 524965 44298 525031 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal3 s 518801 44298 518867 44301 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 524970 44240 525026 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel via2 s 518806 44240 518862 44296 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524971 41713 525027 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518807 41713 518863 42193 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524984 42193 525012 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518820 42193 518848 44231 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 524970 44231 525026 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 518806 44231 518862 44305 6 gpio_mode1_core
port 26 nsew signal input
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 27 nsew signal input
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 28 nsew signal input
rlabel metal4 s 37293 40546 38223 68254 6 vccd
port 29 nsew signal bidirectional
rlabel metal4 s 37293 82746 38223 110454 6 vccd
port 30 nsew signal bidirectional
rlabel metal5 s 37313 40546 38203 68254 6 vccd
port 31 nsew signal bidirectional
rlabel metal5 s 37313 82746 38203 110454 6 vccd
port 32 nsew signal bidirectional
rlabel metal3 s 38220 68100 39600 72900 6 vccd
port 33 nsew signal bidirectional
rlabel metal3 s 145816 36683 145934 36711 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145816 36711 146052 36741 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145962 36741 146052 36801 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145816 36741 145934 36801 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145816 36801 145962 36843 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145816 36843 145920 40000 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145820 40000 145898 40014 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 149605 40291 149671 40294 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145838 40014 145898 40294 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145790 40294 149671 40354 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 149605 40354 149671 40357 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 145790 40354 145850 40430 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 143533 40427 143599 40430 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 143533 40430 145850 40490 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 143533 40490 143599 40493 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 502057 44643 502123 44646 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 483013 44643 483079 44646 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 483013 44646 502123 44706 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 502057 44706 502123 44709 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 483013 44706 483079 44709 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 41413 78235 41479 78238 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 38220 78151 39600 78238 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 38220 78238 41479 78298 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 41413 78298 41479 78301 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 42701 80547 42767 80550 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 41413 80547 41479 80550 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 41413 80550 42767 80610 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 42701 80610 42767 80613 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 41413 80610 41479 80613 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 38220 78298 39600 82940 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 673821 154531 673887 154534 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 673637 154531 673703 154534 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 673637 154534 673887 154594 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 673821 154594 673887 154597 6 vccd
port 34 nsew signal bidirectional
rlabel metal3 s 673637 154594 673703 154597 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 149610 40296 149666 40352 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 143538 40432 143594 40488 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 502062 44648 502118 44704 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 483018 44648 483074 44704 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 41418 78240 41474 78296 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 42706 80552 42762 80608 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 41418 80552 41474 80608 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 673826 154536 673882 154592 6 vccd
port 34 nsew signal bidirectional
rlabel via2 s 673642 154536 673698 154592 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 149610 40287 149666 40361 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 516323 41713 516379 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 461523 41713 461579 41806 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 461504 41806 461579 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 406723 41713 406779 41820 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 516336 42193 516364 44474 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 502076 44390 502288 44418 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 502260 44418 502288 44474 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 516324 44474 516376 44538 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 502248 44474 502300 44538 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 516336 44538 516364 45494 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 502076 44418 502104 44639 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 469140 44526 469260 44542 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 461504 42193 461532 44542 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 406723 41820 406792 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 360571 41713 360627 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 354407 41713 354463 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 351923 41713 351979 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 305771 41713 305827 41806 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 299607 41713 299663 41806 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 297123 41713 297179 41806 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 305748 41806 305827 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 299584 41806 299663 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 297100 41806 297179 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 201495 41713 201551 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192847 41713 192903 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 188523 41713 188579 41942 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 149624 40361 149652 41754 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 143538 40423 143594 40497 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 187700 41754 187752 41818 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 149612 41754 149664 41818 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 187712 41818 187740 41890 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 188436 41890 188488 41942 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 188436 41942 188579 41954 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 187700 41890 187752 41954 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 188448 41954 188579 41970 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 188523 41970 188579 42193 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 444208 44390 444328 44418 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 444300 44418 444328 44474 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 444288 44474 444340 44538 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 469128 44542 469272 44554 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 469220 44554 469272 44606 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 469128 44554 469180 44606 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 461492 44542 461544 44606 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 483020 44610 483072 44639 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 502062 44639 502118 44713 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 483018 44639 483074 44713 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 444208 44418 444236 44678 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 406764 42193 406792 44474 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 360580 42193 360608 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 354416 42193 354444 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 351932 42193 351960 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 305748 42193 305776 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 299584 42193 299612 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 297100 42193 297128 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 201512 42193 201540 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192864 42193 192892 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 188540 42193 188568 44270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 399668 44270 399720 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 360568 44270 360620 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 354404 44270 354456 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 351920 44270 351972 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 305736 44270 305788 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 299572 44270 299624 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 297088 44270 297140 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 201500 44270 201552 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192852 44270 192904 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 188528 44270 188580 44334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 399680 44334 399708 44474 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 360580 44334 360608 44474 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 354416 44334 354444 44474 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 406752 44474 406804 44538 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 399668 44474 399720 44538 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 360568 44474 360620 44538 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 354404 44474 354456 44538 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 425060 44542 425112 44606 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 425072 44606 425100 44678 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 406764 44538 406792 44678 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 444196 44678 444248 44742 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 425060 44678 425112 44742 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 406752 44678 406804 44742 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 45494 673696 45558 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 516324 45494 516376 45558 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 102123 675887 102151 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 102151 675887 102179 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 102179 675432 102274 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673656 45558 673684 102274 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 143552 40497 143580 45562 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 143540 45562 143592 45626 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 45562 42760 45626 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 45626 42748 80543 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41418 78231 41474 78305 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41432 78305 41460 80543 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42706 80543 42762 80617 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41418 80543 41474 80617 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 80617 42748 91038 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 91038 42748 91066 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 102274 675444 102338 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675024 102274 675076 102338 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 102274 673696 102338 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675036 102338 675064 115806 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 91066 42564 110434 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 110434 42760 110498 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 110434 42576 110498 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675024 115806 675076 115870 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673828 115806 673880 115870 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673840 115870 673868 115942 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674012 115942 674064 116006 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673828 115942 673880 116006 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674024 116006 674052 140626 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 110498 42748 129662 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 129662 42748 129690 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675024 140626 675076 140690 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674012 140626 674064 140690 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675036 140690 675064 147086 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 147086 675444 147150 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675024 147086 675076 147150 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 147086 673696 147150 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 147150 675432 147323 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 147323 675887 147356 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 147356 675887 147379 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673656 147150 673684 154527 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 129690 42564 149058 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 149058 42760 149122 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 149058 42576 149122 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673826 154527 673882 154601 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673642 154527 673698 154601 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673840 154601 673868 173878 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674748 173878 674800 173942 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673828 173878 673880 173942 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674760 173942 674788 192102 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 149122 42748 185302 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 185302 42760 185366 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42432 185302 42484 185366 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 192102 675444 192166 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675208 192102 675260 192166 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674748 192102 674800 192166 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 192166 675432 192323 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 192323 675887 192372 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 192372 675887 192379 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675220 192166 675248 198698 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42444 185366 42472 194890 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42892 194890 42944 194954 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42432 194890 42484 194954 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 194890 41840 194954 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675208 198698 675260 198762 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674012 198698 674064 198762 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674024 198762 674052 212502 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42904 194954 42932 208354 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 194954 41828 195421 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 195421 42193 195477 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42892 208354 42944 208418 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42340 208354 42392 208418 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674288 212502 674340 212566 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674012 212502 674064 212566 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674300 212566 674328 231746 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674288 231746 674340 231810 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674104 231746 674156 231810 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674116 231810 674144 237322 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42352 208418 42380 232834 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42616 232834 42668 232898 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42340 232834 42392 232898 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 674104 237322 674156 237386 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673920 237322 673972 237386 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 237523 675887 237524 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 237524 675887 237579 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 237579 675432 237662 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673932 237386 673960 237662 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 237662 675444 237726 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673920 237662 673972 237726 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673932 237726 673960 244038 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42628 232898 42656 238070 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42892 238070 42944 238134 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42616 238070 42668 238134 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 238070 41840 238134 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673748 244038 673960 244066 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673748 244066 673776 282066 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42904 238134 42932 245550 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 238134 41828 238621 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 238621 42193 238677 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42892 245550 42944 245614 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42340 245550 42392 245614 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42352 245614 42380 275998 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42352 275998 42564 276026 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 282066 675444 282130 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673736 282066 673788 282130 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 282130 675432 282523 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 282523 675887 282540 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 282540 675887 282579 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 327523 675887 327556 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 327556 675887 327579 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 327579 675432 328034 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673748 282130 673776 328034 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 276026 42564 282270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 281821 42193 281877 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 281877 41828 282270 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 282270 42576 282334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 282270 41840 282334 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 282334 42564 283675 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42352 283675 42564 283703 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42352 283703 42380 314162 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 314162 42760 314226 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42340 314162 42392 314226 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 314226 42748 322798 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 322798 42760 322862 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42432 322866 42484 322930 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42444 322930 42472 325450 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 325021 42193 325077 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 325077 41828 325450 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 325450 42760 325514 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42432 325450 42484 325514 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 325450 41840 325514 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 328034 675444 328098 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673736 328034 673788 328098 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673748 328098 673776 372302 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 325514 42748 342230 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 342230 42840 342258 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42812 342258 42840 367696 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42812 367696 42932 367724 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42904 367724 42932 368630 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 368221 42193 368277 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 368277 41828 368630 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42892 368630 42944 368694 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 368630 41840 368694 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 372302 675444 372366 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673736 372302 673788 372366 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 372366 675432 372723 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 372723 675887 372751 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 372751 675887 372779 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42904 368694 42932 386310 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42892 386310 42944 386374 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42616 386310 42668 386374 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42628 386374 42656 391870 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 391870 42656 391898 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 391898 42564 411198 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 411198 42576 411262 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 411198 41840 411262 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 411262 42564 539446 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 411262 41828 411421 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 411421 42193 411477 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 539021 42193 539077 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 539077 41828 539446 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 539446 42576 539510 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 539446 41840 539510 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 539510 42564 540518 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42352 540518 42564 540546 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 549923 675887 549951 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 549951 675887 549979 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 549979 675432 550462 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 550462 675444 550526 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 550462 673696 550526 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673656 550526 673684 594866 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42352 540546 42380 574058 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42800 574058 42852 574122 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42340 574058 42392 574122 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42812 574122 42840 582626 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 582221 42193 582277 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 582277 41828 582626 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42800 582626 42852 582690 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 582626 41840 582690 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 594866 675444 594930 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673920 594866 673972 594930 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 594866 673696 594930 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 594930 675432 595123 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 595123 675887 595151 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 595151 675887 595179 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673932 594930 673960 639678 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42812 582690 42840 612614 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42800 612614 42852 612678 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42616 612614 42668 612678 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42628 612678 42656 612750 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42616 612750 42668 612814 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42800 612818 42852 612882 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42812 612882 42840 624922 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42800 624922 42852 624986 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 624922 41840 624986 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42812 624986 42840 631858 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 624986 41828 625421 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 625421 42193 625477 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42800 631858 42852 631922 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 631994 42576 632058 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 639678 675444 639742 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673920 639678 673972 639742 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673460 639678 673512 639742 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 639742 675432 640123 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 640123 675887 640151 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 640151 675887 640179 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673472 639742 673500 685170 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 632058 42564 669054 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 668621 42193 668677 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 668677 41828 669054 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 669054 42576 669118 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 669054 41840 669118 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 669118 42564 672166 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 672166 42656 672194 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42628 672194 42656 678422 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42628 678422 42748 678450 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 685170 675444 685234 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673460 685170 673512 685234 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 685234 675432 685323 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 685323 675887 685372 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 685372 675887 685379 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673472 685234 673500 730118 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 678450 42748 711282 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 711282 42760 711346 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42432 711282 42484 711346 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 711282 41840 711346 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 730118 675444 730182 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673460 730118 673512 730182 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 730182 675432 730323 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 730323 675887 730351 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 730351 675887 730379 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673472 730182 673500 774862 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42444 711346 42472 754462 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 711346 41828 711821 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 711821 42193 711877 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42432 754462 42484 754526 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 754462 41840 754526 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42444 754526 42472 767314 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 754526 41828 755021 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 755021 42193 755077 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 767314 42760 767378 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42432 767314 42484 767378 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 774862 675444 774926 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 774862 673696 774926 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673460 774862 673512 774926 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 774926 675432 775323 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 775323 675887 775351 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 775351 675887 775379 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673656 774926 673684 864418 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42720 767378 42748 797710 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42708 797710 42760 797774 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 797710 42576 797774 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 797710 41840 797774 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 864418 675444 864482 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 864418 673696 864482 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 864482 675432 864523 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 864523 675887 864551 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 864551 675887 864579 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673656 864482 673684 953294 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675392 953294 675444 953358 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 953294 673696 953358 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 953358 675432 953723 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675404 953723 675887 953751 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 675407 953751 675887 953779 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673656 953358 673684 990150 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 797774 42564 968458 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 797774 41828 798221 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 798221 42193 798277 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41713 968021 42193 968077 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41800 968077 41828 968458 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 968458 42576 968522 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 41788 968458 41840 968522 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42536 968522 42564 990014 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 42524 990014 42576 990078 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 89904 990082 89956 990134 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 89904 990134 90036 990146 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 673644 990150 673696 990214 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 639788 990150 639840 990214 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 89916 990146 90036 990162 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 639800 990214 639828 990762 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 194968 990422 195020 990486 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192852 990422 192904 990486 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 397460 990490 397512 990554 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 295800 990490 295852 990554 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 397472 990554 397500 990762 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 295812 990554 295840 990694 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 194980 990486 195008 990694 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192864 990486 192892 990694 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 90008 990162 90036 990694 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 295800 990694 295852 990758 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 244188 990694 244240 990758 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 194968 990694 195020 990758 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192852 990694 192904 990758 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 141424 990694 141476 990758 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 89996 990694 90048 990758 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 639788 990762 639840 990826 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 538036 990762 538088 990826 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 486608 990762 486660 990826 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 397644 990762 397696 990826 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 397460 990762 397512 990826 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 639800 990826 639828 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 538048 990826 538076 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 486620 990826 486648 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 639800 995407 639877 995466 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 639821 995466 639877 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 538021 995407 538077 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 486620 995407 486677 995452 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 397656 990826 397684 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 295812 990758 295840 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 244200 990758 244228 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 397621 995407 397684 995452 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 486621 995452 486677 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 397621 995452 397677 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 295812 995407 295877 995452 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 295821 995452 295877 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 244200 995407 244277 995466 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192864 990758 192892 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 141436 990758 141464 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 90008 990758 90036 995407 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192821 995407 192892 995466 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 244221 995466 244277 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 192821 995466 192877 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 141421 995407 141477 995887 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 90008 995407 90077 995452 6 vccd
port 34 nsew signal bidirectional
rlabel metal2 s 90021 995452 90077 995887 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 187700 41760 187752 41812 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 149612 41760 149664 41812 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 188436 41896 188488 41948 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 187700 41896 187752 41948 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 399668 44276 399720 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 360568 44276 360620 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 354404 44276 354456 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 351920 44276 351972 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 305736 44276 305788 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 299572 44276 299624 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 297088 44276 297140 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 201500 44276 201552 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 192852 44276 192904 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 188528 44276 188580 44328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 516324 44480 516376 44532 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 502248 44480 502300 44532 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 483020 44616 483072 44668 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 469220 44548 469272 44600 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 469128 44548 469180 44600 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 461492 44548 461544 44600 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 444288 44480 444340 44532 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 406752 44480 406804 44532 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 399668 44480 399720 44532 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 360568 44480 360620 44532 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 354404 44480 354456 44532 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 425060 44548 425112 44600 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 444196 44684 444248 44736 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 425060 44684 425112 44736 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 406752 44684 406804 44736 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 45500 673696 45552 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 516324 45500 516376 45552 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 143540 45568 143592 45620 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 45568 42760 45620 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 102280 675444 102332 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675024 102280 675076 102332 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 102280 673696 102332 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 110440 42760 110492 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 110440 42576 110492 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675024 115812 675076 115864 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673828 115812 673880 115864 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674012 115948 674064 116000 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673828 115948 673880 116000 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675024 140632 675076 140684 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674012 140632 674064 140684 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 147092 675444 147144 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675024 147092 675076 147144 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 147092 673696 147144 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 149064 42760 149116 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 149064 42576 149116 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674748 173884 674800 173936 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673828 173884 673880 173936 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 185308 42760 185360 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42432 185308 42484 185360 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 192108 675444 192160 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675208 192108 675260 192160 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674748 192108 674800 192160 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42892 194896 42944 194948 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42432 194896 42484 194948 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 194896 41840 194948 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675208 198704 675260 198756 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674012 198704 674064 198756 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42892 208360 42944 208412 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42340 208360 42392 208412 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674288 212508 674340 212560 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674012 212508 674064 212560 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674288 231752 674340 231804 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674104 231752 674156 231804 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42616 232840 42668 232892 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42340 232840 42392 232892 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 674104 237328 674156 237380 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673920 237328 673972 237380 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 237668 675444 237720 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673920 237668 673972 237720 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42892 238076 42944 238128 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42616 238076 42668 238128 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 238076 41840 238128 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42892 245556 42944 245608 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42340 245556 42392 245608 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 282072 675444 282124 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673736 282072 673788 282124 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 282276 42576 282328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 282276 41840 282328 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 314168 42760 314220 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42340 314168 42392 314220 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 322804 42760 322856 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42432 322872 42484 322924 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 325456 42760 325508 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42432 325456 42484 325508 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 325456 41840 325508 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 328040 675444 328092 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673736 328040 673788 328092 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42892 368636 42944 368688 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 368636 41840 368688 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 372308 675444 372360 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673736 372308 673788 372360 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42892 386316 42944 386368 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42616 386316 42668 386368 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 411204 42576 411256 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 411204 41840 411256 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 539452 42576 539504 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 539452 41840 539504 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 550468 675444 550520 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 550468 673696 550520 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42800 574064 42852 574116 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42340 574064 42392 574116 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42800 582632 42852 582684 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 582632 41840 582684 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 594872 675444 594924 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673920 594872 673972 594924 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 594872 673696 594924 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42800 612620 42852 612672 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42616 612620 42668 612672 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42616 612756 42668 612808 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42800 612824 42852 612876 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42800 624928 42852 624980 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 624928 41840 624980 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42800 631864 42852 631916 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 632000 42576 632052 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 639684 675444 639736 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673920 639684 673972 639736 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673460 639684 673512 639736 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 669060 42576 669112 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 669060 41840 669112 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 685176 675444 685228 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673460 685176 673512 685228 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 711288 42760 711340 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42432 711288 42484 711340 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 711288 41840 711340 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 730124 675444 730176 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673460 730124 673512 730176 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42432 754468 42484 754520 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 754468 41840 754520 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 767320 42760 767372 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42432 767320 42484 767372 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 774868 675444 774920 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 774868 673696 774920 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673460 774868 673512 774920 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42708 797716 42760 797768 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 797716 42576 797768 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 797716 41840 797768 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 864424 675444 864476 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 864424 673696 864476 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 675392 953300 675444 953352 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 953300 673696 953352 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 968464 42576 968516 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 41788 968464 41840 968516 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 42524 990020 42576 990072 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 89904 990088 89956 990140 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 673644 990156 673696 990208 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 639788 990156 639840 990208 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 194968 990428 195020 990480 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 192852 990428 192904 990480 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 397460 990496 397512 990548 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 295800 990496 295852 990548 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 295800 990700 295852 990752 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 244188 990700 244240 990752 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 194968 990700 195020 990752 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 192852 990700 192904 990752 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 141424 990700 141476 990752 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 89996 990700 90048 990752 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 639788 990768 639840 990820 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 538036 990768 538088 990820 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 486608 990768 486660 990820 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 397644 990768 397696 990820 6 vccd
port 34 nsew signal bidirectional
rlabel via1 s 397460 990768 397512 990820 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 187694 41760 187758 41772 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 149606 41760 149670 41772 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 149606 41772 187758 41800 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 187694 41800 187758 41812 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 149606 41800 149670 41812 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 188430 41896 188494 41908 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 187694 41896 187758 41908 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 187694 41908 188494 41936 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 188430 41936 188494 41948 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 187694 41936 187758 41948 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 399662 44276 399726 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 360562 44276 360626 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 360562 44288 399726 44316 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 399662 44316 399726 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 360562 44316 360626 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 354398 44276 354462 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 351914 44276 351978 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 305730 44276 305794 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 299566 44276 299630 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 297082 44276 297146 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 201494 44276 201558 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 192846 44276 192910 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 188522 44276 188586 44288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 188522 44288 354462 44316 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 354398 44316 354462 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 351914 44316 351978 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 305730 44316 305794 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 299566 44316 299630 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 297082 44316 297146 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 201494 44316 201558 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 192846 44316 192910 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 188522 44316 188586 44328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 516318 44480 516382 44492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 502352 44492 516382 44520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 516318 44520 516382 44532 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 502352 44520 502380 44560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 502242 44480 502306 44532 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 444282 44480 444346 44492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 444282 44492 449848 44520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 502260 44532 502288 44560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 469214 44548 469278 44560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 502260 44560 502380 44588 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 469214 44560 473308 44588 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 483014 44616 483078 44628 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 473280 44588 473308 44628 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 469214 44588 469278 44600 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 469122 44548 469186 44560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 461486 44548 461550 44560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 449820 44520 449848 44560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 444282 44520 444346 44532 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 406746 44480 406810 44492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 399662 44480 399726 44492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 399662 44492 406810 44520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 406746 44520 406810 44532 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 399662 44520 399726 44532 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 360562 44480 360626 44492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 354398 44480 354462 44492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 354398 44492 360626 44520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 360562 44520 360626 44532 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 354398 44520 354462 44532 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 449820 44560 469186 44588 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 425054 44548 425118 44560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 411272 44560 425118 44588 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 469122 44588 469186 44600 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 461486 44588 461550 44600 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 425054 44588 425118 44600 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 473280 44628 483078 44656 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 483014 44656 483078 44668 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 444190 44684 444254 44696 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 425054 44684 425118 44696 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 425054 44696 444254 44724 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 411272 44588 411300 44696 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 406746 44684 406810 44696 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 406746 44696 411300 44724 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 444190 44724 444254 44736 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 425054 44724 425118 44736 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 406746 44724 406810 44736 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 45500 673702 45512 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 516318 45500 516382 45512 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 516318 45512 673702 45540 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 45540 673702 45552 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 516318 45540 516382 45552 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 143534 45568 143598 45580 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 45568 42766 45580 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 45580 143598 45608 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 143534 45608 143598 45620 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 45608 42766 45620 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 102280 675450 102292 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 102280 675082 102292 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 102280 673702 102292 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 102292 675450 102320 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 102320 675450 102332 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 102320 675082 102332 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 102320 673702 102332 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 110440 42766 110452 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 110440 42582 110452 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 110452 42766 110480 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 110480 42766 110492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 110480 42582 110492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 115812 675082 115824 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 115812 673886 115824 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 115824 675082 115852 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 115852 675082 115864 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 115852 673886 115864 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 115948 674070 115960 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 115948 673886 115960 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 115960 674070 115988 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 115988 674070 116000 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 115988 673886 116000 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 140632 675082 140644 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 140632 674070 140644 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 140644 675082 140672 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 140672 675082 140684 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 140672 674070 140684 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 147092 675450 147104 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 147092 675082 147104 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 147092 673702 147104 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 147104 675450 147132 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 147132 675450 147144 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675018 147132 675082 147144 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 147132 673702 147144 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 149064 42766 149076 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 149064 42582 149076 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 149076 42766 149104 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 149104 42766 149116 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 149104 42582 149116 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674742 173884 674806 173896 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 173884 673886 173896 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 173896 674806 173924 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674742 173924 674806 173936 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673822 173924 673886 173936 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 185308 42766 185320 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 185308 42490 185320 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 185320 42766 185348 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 185348 42766 185360 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 185348 42490 185360 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 192108 675450 192120 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675202 192108 675266 192120 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674742 192108 674806 192120 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674742 192120 675450 192148 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 192148 675450 192160 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675202 192148 675266 192160 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674742 192148 674806 192160 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 194896 42950 194908 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 194896 42490 194908 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 194896 41846 194908 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 194908 42950 194936 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 194936 42950 194948 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 194936 42490 194948 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 194936 41846 194948 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675202 198704 675266 198716 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 198704 674070 198716 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 198716 675266 198744 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675202 198744 675266 198756 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 198744 674070 198756 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 208360 42950 208372 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 208360 42398 208372 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 208372 42950 208400 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 208400 42950 208412 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 208400 42398 208412 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674282 212508 674346 212520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 212508 674070 212520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 212520 674346 212548 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674282 212548 674346 212560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674006 212548 674070 212560 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674282 231752 674346 231764 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674098 231752 674162 231764 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674098 231764 674346 231792 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674282 231792 674346 231804 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674098 231792 674162 231804 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 232840 42674 232852 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 232840 42398 232852 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 232852 42674 232880 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 232880 42674 232892 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 232880 42398 232892 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674098 237328 674162 237340 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 237328 673978 237340 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 237340 674162 237368 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 674098 237368 674162 237380 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 237368 673978 237380 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 237668 675450 237680 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 237668 673978 237680 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 237680 675450 237708 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 237708 675450 237720 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 237708 673978 237720 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 238076 42950 238088 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 238076 42674 238088 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 238076 41846 238088 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 238088 42950 238116 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 238116 42950 238128 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 238116 42674 238128 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 238116 41846 238128 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 245556 42950 245568 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 245556 42398 245568 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 245568 42950 245596 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 245596 42950 245608 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 245596 42398 245608 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 282072 675450 282084 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 282072 673794 282084 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 282084 675450 282112 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 282112 675450 282124 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 282112 673794 282124 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 282276 42582 282288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 282276 41846 282288 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 282288 42582 282316 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 282316 42582 282328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 282316 41846 282328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 314168 42766 314180 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 314168 42398 314180 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 314180 42766 314208 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 314208 42766 314220 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 314208 42398 314220 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 322804 42766 322856 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42720 322856 42748 322884 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 322872 42490 322884 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 322884 42748 322912 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 322912 42490 322924 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 325456 42766 325468 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 325456 42490 325468 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 325456 41846 325468 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 325468 42766 325496 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 325496 42766 325508 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 325496 42490 325508 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 325496 41846 325508 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 328040 675450 328052 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 328040 673794 328052 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 328052 675450 328080 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 328080 675450 328092 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 328080 673794 328092 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 368636 42950 368648 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 368636 41846 368648 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 368648 42950 368676 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 368676 42950 368688 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 368676 41846 368688 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 372308 675450 372320 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 372308 673794 372320 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 372320 675450 372348 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 372348 675450 372360 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673730 372348 673794 372360 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 386316 42950 386328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 386316 42674 386328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 386328 42950 386356 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42886 386356 42950 386368 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 386356 42674 386368 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 411204 42582 411216 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 411204 41846 411216 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 411216 42582 411244 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 411244 42582 411256 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 411244 41846 411256 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 539452 42582 539464 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 539452 41846 539464 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 539464 42582 539492 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 539492 42582 539504 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 539492 41846 539504 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 550468 675450 550480 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 550468 673702 550480 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 550480 675450 550508 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 550508 675450 550520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 550508 673702 550520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 574064 42858 574076 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 574064 42398 574076 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 574076 42858 574104 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 574104 42858 574116 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42334 574104 42398 574116 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 582632 42858 582644 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 582632 41846 582644 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 582644 42858 582672 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 582672 42858 582684 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 582672 41846 582684 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 594872 675450 594884 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 594872 673978 594884 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 594872 673702 594884 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 594884 675450 594912 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 594912 675450 594924 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 594912 673978 594924 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 594912 673702 594924 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 612620 42858 612632 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 612620 42674 612632 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 612632 42858 612660 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 612660 42858 612672 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 612660 42674 612672 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 612756 42674 612768 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 612768 42840 612796 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42812 612796 42840 612824 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42610 612796 42674 612808 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 612824 42858 612876 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 624928 42858 624940 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 624928 41846 624940 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 624940 42858 624968 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 624968 42858 624980 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 624968 41846 624980 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 631864 42858 631876 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42536 631876 42858 631904 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42794 631904 42858 631916 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42536 631904 42564 632000 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 632000 42582 632052 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 639684 675450 639696 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 639684 673978 639696 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 639684 673518 639696 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 639696 675450 639724 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 639724 675450 639736 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673914 639724 673978 639736 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 639724 673518 639736 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 669060 42582 669072 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 669060 41846 669072 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 669072 42582 669100 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 669100 42582 669112 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 669100 41846 669112 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 685176 675450 685188 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 685176 673518 685188 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 685188 675450 685216 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 685216 675450 685228 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 685216 673518 685228 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 711288 42766 711300 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 711288 42490 711300 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 711288 41846 711300 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 711300 42766 711328 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 711328 42766 711340 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 711328 42490 711340 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 711328 41846 711340 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 730124 675450 730136 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 730124 673518 730136 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 730136 675450 730164 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 730164 675450 730176 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 730164 673518 730176 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 754468 42490 754480 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 754468 41846 754480 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 754480 42490 754508 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 754508 42490 754520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 754508 41846 754520 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 767320 42766 767332 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 767320 42490 767332 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 767332 42766 767360 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 767360 42766 767372 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42426 767360 42490 767372 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 774868 675450 774880 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 774868 673702 774880 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 774868 673518 774880 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 774880 675450 774908 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 774908 675450 774920 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 774908 673702 774920 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673454 774908 673518 774920 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 797716 42766 797728 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 797716 42582 797728 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 797716 41846 797728 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 797728 42766 797756 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42702 797756 42766 797768 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 797756 42582 797768 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 797756 41846 797768 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 864424 675450 864436 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 864424 673702 864436 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 864436 675450 864464 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 864464 675450 864476 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 864464 673702 864476 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 953300 675450 953312 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 953300 673702 953312 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 953312 675450 953340 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 675386 953340 675450 953352 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 953340 673702 953352 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 968464 42582 968476 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 968464 41846 968476 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 968476 42582 968504 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 968504 42582 968516 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 41782 968504 41846 968516 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 990020 42582 990032 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 990032 89944 990060 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 89916 990060 89944 990088 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 42518 990060 42582 990072 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 89898 990088 89962 990140 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 990156 673702 990168 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 639782 990156 639846 990168 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 639782 990168 673702 990196 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 673638 990196 673702 990208 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 639782 990196 639846 990208 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 194962 990428 195026 990440 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 192846 990428 192910 990440 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 192846 990440 195026 990468 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 194962 990468 195026 990480 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 192846 990468 192910 990480 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 397454 990496 397518 990508 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 295794 990496 295858 990508 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 295794 990508 397518 990536 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 397454 990536 397518 990548 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 295794 990536 295858 990548 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 295794 990700 295858 990712 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 244182 990700 244246 990712 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 194962 990700 195026 990712 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 194962 990712 295858 990740 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 295794 990740 295858 990752 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 244182 990740 244246 990752 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 194962 990740 195026 990752 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 192846 990700 192910 990712 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 141418 990700 141482 990712 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 89990 990700 90054 990712 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 89990 990712 192910 990740 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 192846 990740 192910 990752 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 141418 990740 141482 990752 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 89990 990740 90054 990752 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 639782 990768 639846 990780 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 538030 990768 538094 990780 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 486602 990768 486666 990780 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 397638 990768 397702 990780 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 397454 990768 397518 990780 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 397454 990780 639846 990808 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 639782 990808 639846 990820 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 538030 990808 538094 990820 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 486602 990808 486666 990820 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 397638 990808 397702 990820 6 vccd
port 34 nsew signal bidirectional
rlabel metal1 s 397454 990808 397518 990820 6 vccd
port 34 nsew signal bidirectional
rlabel metal5 s 6086 69863 19572 81191 6 vccd
port 35 nsew signal bidirectional
rlabel metal4 s 637607 36323 677051 37013 6 vdda
port 36 nsew signal bidirectional
rlabel metal4 s 583807 36323 622993 37013 6 vdda
port 37 nsew signal bidirectional
rlabel metal5 s 637607 36343 677051 36993 6 vdda
port 38 nsew signal bidirectional
rlabel metal5 s 583807 36343 622993 36993 6 vdda
port 39 nsew signal bidirectional
rlabel metal3 s 632921 37008 637701 40000 6 vdda
port 40 nsew signal bidirectional
rlabel metal3 s 622942 37008 627722 40000 6 vdda
port 41 nsew signal bidirectional
rlabel metal5 s 624040 6675 636580 19198 6 vdda
port 42 nsew signal bidirectional
rlabel metal4 s 21000 109800 25993 110454 6 vddio
port 43 nsew signal bidirectional
rlabel metal4 s 35113 82746 36043 110454 6 vddio
port 44 nsew signal bidirectional
rlabel metal4 s 21000 124946 25993 125400 6 vddio
port 45 nsew signal bidirectional
rlabel metal4 s 35113 124946 36043 181854 6 vddio
port 46 nsew signal bidirectional
rlabel metal5 s 35133 82746 36023 110454 6 vddio
port 47 nsew signal bidirectional
rlabel metal5 s 21003 109800 25993 110454 6 vddio
port 48 nsew signal bidirectional
rlabel metal5 s 35133 124946 36023 181854 6 vddio
port 49 nsew signal bidirectional
rlabel metal5 s 21003 124946 25993 125400 6 vddio
port 50 nsew signal bidirectional
rlabel metal3 s 405641 44507 405707 44510 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 386413 44507 386479 44510 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 386413 44510 405707 44570 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 405641 44570 405707 44573 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 386413 44570 386479 44573 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 44633 96595 44699 96598 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 42977 96595 43043 96598 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 42977 96598 44699 96658 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 44633 96658 44699 96661 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 42977 96658 43043 96661 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 42977 110331 43043 110334 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 36040 110299 40000 110334 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 36040 110334 43043 110394 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 42977 110394 43043 110397 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 36040 110394 40000 115079 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 42241 870027 42307 870030 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 36040 869899 40000 870030 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 36040 870030 42307 870090 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 42241 870090 42307 870093 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 36040 870090 40000 874679 6 vddio
port 51 nsew signal bidirectional
rlabel via2 s 405646 44512 405702 44568 6 vddio
port 51 nsew signal bidirectional
rlabel via2 s 386418 44512 386474 44568 6 vddio
port 51 nsew signal bidirectional
rlabel via2 s 44638 96600 44694 96656 6 vddio
port 51 nsew signal bidirectional
rlabel via2 s 42982 96600 43038 96656 6 vddio
port 51 nsew signal bidirectional
rlabel via2 s 42982 110336 43038 110392 6 vddio
port 51 nsew signal bidirectional
rlabel via2 s 42246 870032 42302 870088 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 523775 41713 523831 42193 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 468975 41713 469031 41806 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 468956 41806 469031 42193 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 414175 41713 414231 41820 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 523788 42193 523816 44202 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 468956 42193 468984 44202 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 414175 41820 414244 42193 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 359375 41713 359431 42193 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 304575 41713 304631 41806 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 304552 41806 304631 42193 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 195975 41713 196031 42193 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 523776 44202 523828 44266 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 468944 44202 468996 44266 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 419816 44202 419868 44266 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 419828 44266 419856 44406 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 414216 42193 414244 44406 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 359384 42193 359412 44338 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 360660 44338 360712 44402 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 359372 44338 359424 44402 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 419816 44406 419868 44470 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 414204 44406 414256 44470 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 360672 44402 360700 44474 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 411260 44474 411312 44538 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 386420 44474 386472 44503 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 411272 44538 411300 44746 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 405646 44503 405702 44577 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 386418 44503 386474 44577 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 360660 44474 360712 44538 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 405660 44577 405688 44746 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 359384 44402 359412 44678 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 304552 42193 304580 44406 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 195992 42193 196020 44406 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 304540 44406 304592 44470 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 195980 44406 196032 44470 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 359372 44678 359424 44742 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 411260 44746 411312 44810 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 405648 44746 405700 44810 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 195992 44470 196020 45494 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 195980 45494 196032 45558 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44916 45494 44968 45558 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44928 45558 44956 82606 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44836 82606 44956 82634 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44836 82634 44864 82758 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44824 82758 44876 82822 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44640 82826 44692 82890 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44652 82890 44680 96591 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44638 96591 44694 96665 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42982 96591 43038 96665 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42996 96665 43024 110327 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42982 110327 43038 110401 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42996 110401 43024 115874 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44732 115874 44784 115938 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42984 115874 43036 115938 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44744 115938 44772 121450 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 44732 121450 44784 121514 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42248 121450 42300 121514 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42260 121514 42288 870023 6 vddio
port 51 nsew signal bidirectional
rlabel metal2 s 42246 870023 42302 870097 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 523776 44208 523828 44260 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 468944 44208 468996 44260 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 419816 44208 419868 44260 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 360660 44344 360712 44396 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 359372 44344 359424 44396 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 419816 44412 419868 44464 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 414204 44412 414256 44464 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 411260 44480 411312 44532 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 386420 44480 386472 44532 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 360660 44480 360712 44532 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 359372 44684 359424 44736 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 304540 44412 304592 44464 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 195980 44412 196032 44464 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 411260 44752 411312 44804 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 405648 44752 405700 44804 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 195980 45500 196032 45552 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 44916 45500 44968 45552 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 44824 82764 44876 82816 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 44640 82832 44692 82884 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 44732 115880 44784 115932 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 42984 115880 43036 115932 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 44732 121456 44784 121508 6 vddio
port 51 nsew signal bidirectional
rlabel via1 s 42248 121456 42300 121508 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 523770 44208 523834 44220 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 468938 44208 469002 44220 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 419810 44208 419874 44220 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 419810 44220 523834 44248 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 523770 44248 523834 44260 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 468938 44248 469002 44260 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 419810 44248 419874 44260 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 360654 44344 360718 44356 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 359366 44344 359430 44356 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 359366 44356 360718 44384 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 360654 44384 360718 44396 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 359366 44384 359430 44396 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 419810 44412 419874 44424 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 414198 44412 414262 44424 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 304534 44412 304598 44424 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 195974 44412 196038 44424 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 414198 44424 419874 44452 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 419810 44452 419874 44464 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 414198 44452 414262 44464 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 195974 44424 342300 44452 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 414216 44464 414244 44492 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 411254 44480 411318 44492 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 411254 44492 414244 44520 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 411254 44520 411318 44532 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 386414 44480 386478 44492 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 360654 44480 360718 44492 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 360654 44492 386478 44520 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 386414 44520 386478 44532 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 360654 44520 360718 44532 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 359366 44684 359430 44696 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 342272 44452 342300 44696 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 304534 44452 304598 44464 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 195974 44452 196038 44464 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 342272 44696 359430 44724 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 359366 44724 359430 44736 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 411254 44752 411318 44764 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 405642 44752 405706 44764 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 405642 44764 411318 44792 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 411254 44792 411318 44804 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 405642 44792 405706 44804 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 195974 45500 196038 45512 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44910 45500 44974 45512 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44910 45512 196038 45540 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 195974 45540 196038 45552 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44910 45540 44974 45552 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44818 82764 44882 82776 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44652 82776 44882 82804 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44818 82804 44882 82816 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44652 82804 44680 82832 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44634 82832 44698 82884 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44726 115880 44790 115892 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 42978 115880 43042 115892 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 42978 115892 44790 115920 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44726 115920 44790 115932 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 42978 115920 43042 115932 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44726 121456 44790 121468 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 42242 121456 42306 121468 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 42242 121468 44790 121496 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 44726 121496 44790 121508 6 vddio
port 51 nsew signal bidirectional
rlabel metal1 s 42242 121496 42306 121508 6 vddio
port 51 nsew signal bidirectional
rlabel metal3 s 36040 120278 40000 125058 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6675 111420 19198 123960 6 vddio
port 53 nsew signal bidirectional
rlabel metal4 s 93546 31963 132854 32653 6 vssa
port 54 nsew signal bidirectional
rlabel metal4 s 93546 28653 192982 28719 6 vssa
port 55 nsew signal bidirectional
rlabel metal4 s 93546 29435 93800 29671 6 vssa
port 56 nsew signal bidirectional
rlabel metal4 s 93546 30387 192982 30453 6 vssa
port 57 nsew signal bidirectional
rlabel metal4 s 39733 31963 79054 32653 6 vssa
port 58 nsew signal bidirectional
rlabel metal4 s 36085 30387 79054 30453 6 vssa
port 59 nsew signal bidirectional
rlabel metal4 s 35365 28653 79054 28719 6 vssa
port 60 nsew signal bidirectional
rlabel metal4 s 78800 29435 79054 29671 6 vssa
port 61 nsew signal bidirectional
rlabel metal5 s 93546 31983 132854 32632 6 vssa
port 62 nsew signal bidirectional
rlabel metal5 s 93800 32632 132600 32633 6 vssa
port 62 nsew signal bidirectional
rlabel metal5 s 93546 28653 132854 30453 6 vssa
port 63 nsew signal bidirectional
rlabel metal5 s 39733 31983 79054 32632 6 vssa
port 64 nsew signal bidirectional
rlabel metal5 s 39733 32632 78800 32633 6 vssa
port 64 nsew signal bidirectional
rlabel metal5 s 35369 28653 79054 30453 6 vssa
port 65 nsew signal bidirectional
rlabel metal3 s 78942 32648 83722 40000 6 vssa
port 66 nsew signal bidirectional
rlabel metal3 s 88921 33497 93701 40000 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 93761 40155 93827 40158 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 91142 40000 91202 40158 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 91142 40158 93827 40218 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 93761 40218 93827 40221 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 362401 41787 362467 41790 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 349613 41787 349679 41790 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 349613 41790 362467 41850 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 362401 41850 362467 41853 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 349613 41850 349679 41853 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 386137 41923 386203 41926 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 367093 41923 367159 41926 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 367093 41926 386203 41986 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 386137 41986 386203 41989 6 vssa
port 67 nsew signal bidirectional
rlabel metal3 s 367093 41986 367159 41989 6 vssa
port 67 nsew signal bidirectional
rlabel via2 s 93766 40160 93822 40216 6 vssa
port 67 nsew signal bidirectional
rlabel via2 s 362406 41792 362462 41848 6 vssa
port 67 nsew signal bidirectional
rlabel via2 s 349618 41792 349674 41848 6 vssa
port 67 nsew signal bidirectional
rlabel via2 s 386142 41928 386198 41984 6 vssa
port 67 nsew signal bidirectional
rlabel via2 s 367098 41928 367154 41984 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 93766 40151 93822 40225 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 507768 41482 507820 41534 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 507768 41534 507900 41546 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 507780 41546 507900 41550 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 507780 41550 507912 41562 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 386156 41534 386368 41562 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 168288 41482 168340 41546 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 140688 41482 140740 41534 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 121276 41482 121328 41534 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 140688 41534 140912 41546 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 121276 41534 121592 41546 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 507860 41562 507912 41614 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 386340 41562 386368 41618 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 386328 41618 386380 41682 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 526811 41713 526867 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 526720 41754 526772 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 526720 41806 526867 41818 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 472011 41713 472067 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 471888 41754 471940 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 471888 41806 472067 41818 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 417211 41713 417267 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 417056 41754 417108 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 417056 41806 417267 41818 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 526732 41818 526867 41834 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 471900 41818 472067 41834 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 417068 41818 417267 41834 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 526811 41834 526867 42193 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 472011 41834 472067 42193 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 417211 41834 417267 42193 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 386156 41562 386184 41919 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 349620 41550 349672 41614 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 362411 41713 362467 41783 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 349632 41614 349660 41783 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 314660 41618 314712 41670 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 314568 41618 314620 41670 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 314568 41670 314712 41682 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 314580 41682 314700 41698 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 168300 41546 168328 41686 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 140700 41546 140912 41550 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 121288 41546 121592 41550 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 93780 40225 93808 41550 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 140700 41550 140924 41562 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 121288 41550 121604 41562 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 140872 41562 140924 41614 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 121552 41562 121604 41614 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 93768 41550 93820 41614 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 362406 41783 362467 41857 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 349618 41783 349674 41857 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 307611 41713 307667 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 199011 41713 199067 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 168288 41686 168340 41750 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 198832 41754 198884 41806 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 307496 41806 307667 41834 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 367100 41890 367152 41919 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 362500 41890 362552 41908 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 362411 41857 362467 41908 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 386142 41919 386198 41993 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 367098 41919 367154 41993 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 362411 41908 362552 41936 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 362500 41936 362552 41954 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 362411 41936 362467 42193 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 307611 41834 307667 42193 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 307496 41834 307524 41890 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 198832 41806 199067 41818 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 198844 41818 199067 41834 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 307484 41890 307536 41954 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 199011 41834 199067 42193 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 198936 41834 198964 41890 6 vssa
port 67 nsew signal bidirectional
rlabel metal2 s 198924 41890 198976 41954 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 507768 41488 507820 41540 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 507860 41556 507912 41608 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 349620 41556 349672 41608 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 526720 41760 526772 41812 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 471888 41760 471940 41812 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 386328 41624 386380 41676 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 314660 41624 314712 41676 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 314568 41624 314620 41676 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 417056 41760 417108 41812 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 367100 41896 367152 41948 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 362500 41896 362552 41948 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 307484 41896 307536 41948 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 198832 41760 198884 41812 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 168288 41488 168340 41540 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 140688 41488 140740 41540 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 140872 41556 140924 41608 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 121276 41488 121328 41540 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 121552 41556 121604 41608 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 93768 41556 93820 41608 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 168288 41692 168340 41744 6 vssa
port 67 nsew signal bidirectional
rlabel via1 s 198924 41896 198976 41948 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 391860 41432 417280 41460 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 507762 41488 507826 41500 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 521580 41500 526760 41528 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 526732 41528 526760 41760 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 521580 41528 521608 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 502352 41500 507826 41528 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 507762 41528 507826 41540 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 507854 41556 507918 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 507854 41568 521608 41596 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 502352 41528 502380 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 430500 41500 472112 41528 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 488460 41568 502380 41596 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 507854 41596 507918 41608 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 488460 41596 488488 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 472084 41528 472112 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 472084 41636 488488 41664 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 430500 41528 430528 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 417252 41460 417280 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 417252 41636 430528 41664 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 391860 41460 391888 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 168282 41488 168346 41500 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 333900 41500 334020 41528 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 349614 41556 349678 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 333992 41528 334020 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 333992 41568 349678 41596 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 333900 41528 333928 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 168282 41500 198780 41528 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 328380 41568 333928 41596 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 349614 41596 349678 41608 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 386322 41624 386386 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 386322 41636 391888 41664 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 328380 41596 328408 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 314654 41624 314718 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 314654 41636 328408 41664 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 526714 41760 526778 41812 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 472084 41664 472112 41772 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 471882 41760 471946 41772 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 471882 41772 472112 41800 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 417252 41664 417280 41772 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 386322 41664 386386 41676 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 314654 41664 314718 41676 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 314562 41624 314626 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 309152 41636 314626 41664 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 314562 41664 314626 41676 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 309152 41664 309180 41704 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 307404 41704 309180 41732 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 417050 41760 417114 41772 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 417050 41772 417280 41800 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 471882 41800 471946 41812 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 417050 41800 417114 41812 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 367094 41896 367158 41908 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 362494 41896 362558 41908 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 362494 41908 367158 41936 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 367094 41936 367158 41948 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 362494 41936 362558 41948 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 307478 41896 307542 41908 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 307404 41732 307432 41908 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 198826 41760 198890 41772 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 198752 41528 198780 41772 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 168282 41528 168346 41540 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 140682 41488 140746 41500 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 121270 41488 121334 41500 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 135272 41500 140746 41528 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 140682 41528 140746 41540 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 140866 41556 140930 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 140866 41568 154528 41596 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 135272 41528 135300 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 102152 41500 121334 41528 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 121270 41528 121334 41540 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 121546 41556 121610 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 121546 41568 135300 41596 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 102152 41528 102180 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 93762 41556 93826 41568 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 93762 41568 102180 41596 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 154500 41596 154528 41636 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 140866 41596 140930 41608 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 121546 41596 121610 41608 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 93762 41596 93826 41608 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 154500 41636 160048 41664 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 168282 41692 168346 41704 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 160020 41664 160048 41704 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 160020 41704 168346 41732 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 168282 41732 168346 41744 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 198752 41772 198890 41800 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 198826 41800 198890 41812 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 198918 41896 198982 41908 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 198918 41908 307542 41936 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 307478 41936 307542 41948 6 vssa
port 67 nsew signal bidirectional
rlabel metal1 s 198918 41936 198982 41948 6 vssa
port 67 nsew signal bidirectional
rlabel metal5 s 80040 6675 92580 19198 6 vssa
port 68 nsew signal bidirectional
rlabel metal4 s 255946 30753 295254 31683 6 vssd
port 69 nsew signal bidirectional
rlabel metal4 s 202146 30753 241454 31683 6 vssd
port 70 nsew signal bidirectional
rlabel metal5 s 255946 30773 295254 31663 6 vssd
port 71 nsew signal bidirectional
rlabel metal5 s 202146 30773 241454 31663 6 vssd
port 72 nsew signal bidirectional
rlabel metal3 s 251300 31680 256100 39600 6 vssd
port 73 nsew signal bidirectional
rlabel metal3 s 241260 31680 246049 39600 6 vssd
port 74 nsew signal bidirectional
rlabel metal3 s 241286 39600 241346 39883 6 vssd
port 74 nsew signal bidirectional
rlabel metal3 s 241286 39883 241395 39946 6 vssd
port 74 nsew signal bidirectional
rlabel metal3 s 241329 39946 241395 39949 6 vssd
port 74 nsew signal bidirectional
rlabel via2 s 241334 39888 241390 39944 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 241334 39879 241390 39953 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 528651 41713 528707 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 528007 41713 528063 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 525615 41713 525671 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 524327 41713 524383 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 521291 41713 521347 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 520003 41713 520059 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 527928 41806 528707 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 525536 41806 525671 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 524248 41806 524383 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 521212 41806 521347 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 520003 41806 520136 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 527916 41822 528707 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 528651 41834 528707 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 528007 41834 528063 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 527916 41834 527968 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 525524 41822 525671 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 525615 41834 525671 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 525524 41834 525576 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 524236 41822 524383 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 524327 41834 524383 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 524236 41834 524288 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 521200 41822 521347 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 521291 41834 521347 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 521200 41834 521252 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 520003 41822 520148 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 520096 41834 520148 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 520003 41834 520059 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 516967 41713 517023 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473851 41713 473907 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473207 41713 473263 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 470815 41713 470871 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473096 41806 473907 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 470815 41806 471008 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 469680 41754 469732 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 469527 41713 469583 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 469527 41806 469732 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473084 41822 473907 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473832 41834 473907 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473207 41834 473263 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473084 41834 473136 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 470815 41822 471020 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 469527 41818 469720 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 470968 41834 471020 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 470815 41834 470871 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 469527 41834 469583 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 466491 41713 466547 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 466368 41754 466420 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 466368 41806 466547 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 465356 41754 465408 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 465203 41713 465259 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 462167 41713 462223 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 419051 41713 419107 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 418407 41713 418463 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 416015 41713 416071 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 414727 41713 414783 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 411691 41713 411747 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 410403 41713 410459 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 465184 41806 465408 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 466380 41818 466547 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 465184 41818 465396 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 466491 41834 466547 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 465184 41834 465259 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 462148 41806 462223 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 418407 41806 419107 41820 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 520016 42193 520044 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 516980 42193 517008 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473832 42193 473860 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 465184 42193 465212 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 462148 42193 462176 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 418407 41820 419120 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 416015 41806 416176 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 414727 41806 414888 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 411691 41806 411852 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 410403 41806 410564 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 407367 41713 407423 41820 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 419051 41834 419120 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 418528 41834 418580 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 418540 41886 418568 41917 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 418407 41834 418463 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 416015 41822 416188 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 416136 41834 416188 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 416015 41834 416071 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 414727 41822 414900 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 414848 41834 414900 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 414727 41834 414783 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 411691 41822 411864 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 411812 41834 411864 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 411691 41834 411747 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 410403 41822 410576 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 410524 41834 410576 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 410403 41834 410472 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 407367 41820 407436 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 364251 41713 364307 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 363607 41713 363663 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 361215 41713 361271 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 359927 41713 359983 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 363524 41806 364307 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 361132 41806 361271 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 359927 41806 360056 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 363512 41822 364307 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 364251 41834 364307 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 363607 41834 363663 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 363512 41834 363564 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 361120 41822 361271 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 361215 41834 361271 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 361120 41834 361172 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 359927 41822 360068 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 360016 41834 360068 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 359927 41834 359983 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 356891 41713 356947 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 356247 41713 356303 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355603 41713 355659 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355603 41806 356947 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 356891 41834 356947 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 356247 41834 356303 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355603 41834 355659 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 352567 41713 352623 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 309451 41713 309507 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 308807 41713 308863 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 308807 41806 309507 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 309428 41834 309507 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 308807 41834 308863 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 306415 41713 306471 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 306288 41754 306340 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 306288 41806 306471 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 305127 41713 305183 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 305000 41754 305052 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 305000 41806 305183 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 302240 41754 302292 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 302091 41713 302147 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 301447 41713 301503 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 300803 41713 300859 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 297767 41713 297823 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 300688 41806 302292 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 306300 41818 306471 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 305012 41818 305183 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 300688 41818 302280 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 297652 41806 297823 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 300676 41822 302280 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 306392 41834 306471 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 305127 41834 305183 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 302091 41834 302147 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 301447 41834 301503 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 300803 41834 300859 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 300676 41834 300728 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 297640 41822 297823 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 297767 41834 297823 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 297640 41834 297692 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 255228 41822 255280 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 255240 41886 255268 42026 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 255228 42026 255280 42090 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 251088 42026 251140 42090 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 419092 42193 419120 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 410444 42193 410472 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 407408 42193 407436 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 364260 42193 364288 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 359936 42193 359964 44202 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355612 42193 355640 44202 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 359924 44202 359976 44266 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355600 44202 355652 44254 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355428 44254 355652 44266 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355428 44266 355640 44282 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355428 44282 355456 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 352576 42193 352604 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 309428 42193 309456 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 306392 42193 306420 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 251100 42090 251128 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 241348 39953 241376 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200851 41713 200907 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200207 41713 200263 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 198367 41713 198423 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 197815 41713 197871 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 197171 41713 197227 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 196527 41713 196583 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 196440 41754 196492 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200132 41806 200907 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 196440 41806 198504 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 193588 41754 193640 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 193491 41713 193547 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 193491 41806 193640 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 192300 41754 192352 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 192203 41713 192259 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 192203 41806 192352 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 191104 41754 191156 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 191007 41713 191063 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 191007 41806 191156 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 189264 41754 189316 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 189167 41713 189223 41806 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 189167 41806 189316 41818 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 196452 41818 198504 41822 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200120 41822 200907 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200851 41834 200907 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200207 41834 200263 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200120 41834 200172 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 196452 41822 198516 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 193491 41818 193628 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 192203 41818 192340 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 191007 41818 191144 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 189167 41818 189304 41834 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 198464 41834 198516 41886 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 198367 41834 198423 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 197815 41834 197871 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 197171 41834 197227 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 196527 41834 196583 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 193491 41834 193547 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 192203 41834 192259 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 191007 41834 191063 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 189167 41834 189223 42193 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200868 42193 200896 44338 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 520004 44338 520056 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 516968 44338 517020 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 473820 44338 473872 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 465172 44338 465224 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 462136 44338 462188 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 419080 44338 419132 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 410432 44338 410484 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 407396 44338 407448 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 364248 44338 364300 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 355416 44338 355468 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 352564 44338 352616 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 309416 44338 309468 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 306380 44338 306432 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 251088 44338 251140 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 241336 44338 241388 44402 6 vssd
port 74 nsew signal bidirectional
rlabel metal2 s 200856 44338 200908 44402 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 527916 41828 527968 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 525524 41828 525576 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 524236 41828 524288 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 521200 41828 521252 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 520096 41828 520148 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 473084 41828 473136 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 470968 41828 471020 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 469680 41760 469732 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 466368 41760 466420 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 465356 41760 465408 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 306288 41760 306340 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 305000 41760 305052 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 302240 41760 302292 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 196440 41760 196492 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 193588 41760 193640 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 192300 41760 192352 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 191104 41760 191156 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 189264 41760 189316 41812 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 418528 41828 418580 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 416136 41828 416188 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 414848 41828 414900 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 411812 41828 411864 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 410524 41828 410576 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 363512 41828 363564 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 361120 41828 361172 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 360016 41828 360068 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 300676 41828 300728 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 297640 41828 297692 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 255228 41828 255280 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 200120 41828 200172 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 198464 41828 198516 41880 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 255228 42032 255280 42084 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 251088 42032 251140 42084 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 359924 44208 359976 44260 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 355600 44208 355652 44260 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 520004 44344 520056 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 516968 44344 517020 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 473820 44344 473872 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 465172 44344 465224 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 462136 44344 462188 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 419080 44344 419132 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 410432 44344 410484 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 407396 44344 407448 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 364248 44344 364300 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 355416 44344 355468 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 352564 44344 352616 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 309416 44344 309468 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 306380 44344 306432 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 251088 44344 251140 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 241336 44344 241388 44396 6 vssd
port 74 nsew signal bidirectional
rlabel via1 s 200856 44344 200908 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 469674 41760 469738 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 466362 41760 466426 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 465350 41760 465414 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 465350 41772 470180 41800 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 527910 41828 527974 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 525518 41828 525582 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 524230 41828 524294 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 521194 41828 521258 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 520090 41828 520154 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 520090 41840 527974 41868 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 527910 41868 527974 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 525518 41868 525582 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 524230 41868 524294 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 521194 41868 521258 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 520090 41868 520154 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 473078 41828 473142 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 470962 41828 471026 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 470152 41800 470180 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 469674 41800 469738 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 466362 41800 466426 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 465350 41800 465414 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 306282 41760 306346 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 304994 41760 305058 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 302234 41760 302298 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 302234 41772 306346 41800 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 306282 41800 306346 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 304994 41800 305058 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 302234 41800 302298 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 196434 41760 196498 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 193582 41760 193646 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 192294 41760 192358 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 191098 41760 191162 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 189258 41760 189322 41772 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 189258 41772 196498 41800 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 196434 41800 196498 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 193582 41800 193646 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 192294 41800 192358 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 191098 41800 191162 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 189258 41800 189322 41812 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 470152 41840 473142 41868 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 418522 41828 418586 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 416130 41828 416194 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 414842 41828 414906 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 411806 41828 411870 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 410518 41828 410582 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 410518 41840 418586 41868 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 473078 41868 473142 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 470962 41868 471026 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 418522 41868 418586 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 416130 41868 416194 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 414842 41868 414906 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 411806 41868 411870 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 410518 41868 410582 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 363506 41828 363570 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 361114 41828 361178 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 360010 41828 360074 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 360010 41840 363570 41868 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 363506 41868 363570 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 361114 41868 361178 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 360010 41868 360074 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 300670 41828 300734 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 297634 41828 297698 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 255222 41828 255286 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 255222 41840 300734 41868 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 300670 41868 300734 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 297634 41868 297698 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 255222 41868 255286 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 200114 41828 200178 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 198458 41828 198522 41840 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 198458 41840 200178 41868 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 200114 41868 200178 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 198458 41868 198522 41880 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 255222 42032 255286 42044 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 251082 42032 251146 42044 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 251082 42044 255286 42072 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 255222 42072 255286 42084 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 251082 42072 251146 42084 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 359918 44208 359982 44220 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 355594 44208 355658 44220 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 355594 44220 359982 44248 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 359918 44248 359982 44260 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 355594 44248 355658 44260 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 519998 44344 520062 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 516962 44344 517026 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 473814 44344 473878 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 473814 44356 520062 44384 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 519998 44384 520062 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 516962 44384 517026 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 473814 44384 473878 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 465166 44344 465230 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 462130 44344 462194 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 419074 44344 419138 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 419074 44356 465230 44384 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 465166 44384 465230 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 462130 44384 462194 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 419074 44384 419138 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 410426 44344 410490 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 407390 44344 407454 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 364242 44344 364306 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 364242 44356 410490 44384 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 410426 44384 410490 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 407390 44384 407454 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 364242 44384 364306 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 355410 44344 355474 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 352558 44344 352622 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 309410 44344 309474 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 306374 44344 306438 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 306374 44356 355474 44384 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 355410 44384 355474 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 352558 44384 352622 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 309410 44384 309474 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 306374 44384 306438 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 251082 44344 251146 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 241330 44344 241394 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 200850 44344 200914 44356 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 200850 44356 251146 44384 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 251082 44384 251146 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 241330 44384 241394 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal1 s 200850 44384 200914 44396 6 vssd
port 74 nsew signal bidirectional
rlabel metal5 s 243009 6086 254337 19572 6 vssd
port 75 nsew signal bidirectional
rlabel metal4 s 297746 1002767 333654 1003697 6 vssio
port 76 nsew signal bidirectional
rlabel metal5 s 570240 6675 582780 19198 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 579121 34830 583901 40000 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 569142 34830 573922 40000 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143332 38317 143388 38373 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143388 38373 143585 38420 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143062 38373 143355 38420 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143062 38420 143585 38666 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143355 38666 143585 40000 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 569174 40000 569234 40155 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 569125 40155 569234 40218 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143398 40000 143458 40158 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143073 40155 143139 40158 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143073 40158 143458 40218 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 569125 40218 569191 40221 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 143073 40218 143139 40221 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 674005 521595 674071 521598 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 673729 521595 673795 521598 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 673729 521598 674071 521658 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 674005 521658 674071 521661 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 673729 521658 673795 521661 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 131021 990387 131087 990390 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 121269 990387 121335 990390 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 121269 990390 131087 990450 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 131021 990450 131087 990453 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 121269 990450 121335 990453 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 342159 997409 342229 997418 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 342159 997418 343650 997478 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 343590 997478 343650 997600 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 342159 997478 342229 997479 6 vssio
port 76 nsew signal bidirectional
rlabel metal3 s 343478 997600 348258 1002770 6 vssio
port 76 nsew signal bidirectional
rlabel via2 s 569130 40160 569186 40216 6 vssio
port 76 nsew signal bidirectional
rlabel via2 s 143078 40160 143134 40216 6 vssio
port 76 nsew signal bidirectional
rlabel via2 s 674010 521600 674066 521656 6 vssio
port 76 nsew signal bidirectional
rlabel via2 s 673734 521600 673790 521656 6 vssio
port 76 nsew signal bidirectional
rlabel via2 s 131026 990392 131082 990448 6 vssio
port 76 nsew signal bidirectional
rlabel via2 s 121274 990392 121330 990448 6 vssio
port 76 nsew signal bidirectional
rlabel via2 s 342164 997414 342224 997474 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141475 35901 141527 36730 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141475 36730 141601 36804 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141601 36804 141646 36821 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141527 36804 141594 36821 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141527 36821 141646 36871 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141594 36871 141646 37693 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141594 37693 141720 37767 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141720 37767 141736 37783 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141646 37767 141684 37783 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141646 37783 141736 37805 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141684 37805 141736 38906 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141684 38906 141784 38928 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141736 38928 141784 38954 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141684 38928 141710 38954 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141784 38954 141850 38969 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141710 38954 141776 38969 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141710 38969 141850 39011 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141784 39011 141850 39020 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141710 39011 141776 39020 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141850 39020 141869 39039 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141776 39020 141847 39039 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141776 39039 144497 39049 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144423 39049 144497 39063 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143068 39049 143128 39063 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141776 39049 141847 39063 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141776 39063 144497 39091 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144401 39091 144497 39113 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144423 39113 144571 39187 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143011 39091 143188 39148 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143068 39148 143188 39151 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144571 39187 144625 39205 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144497 39187 144551 39205 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 145414 39214 145461 39219 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 145414 39219 145530 39247 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144497 39205 144625 39233 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144571 39233 144625 39241 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144497 39233 144551 39241 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 145464 39247 145530 39271 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 145414 39247 145461 39261 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144625 39241 144645 39261 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144551 39241 144623 39261 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144551 39261 145436 39271 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144551 39271 145530 39285 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144551 39285 145464 39313 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144573 39803 144689 40000 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143068 39151 143128 40000 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140996 39872 141048 40000 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144656 40000 144684 40054 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143092 40000 143120 40054 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141008 40000 141036 40054 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144644 40054 144696 40118 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143080 40054 143132 40118 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140996 40054 141048 40118 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 569130 40151 569186 40225 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 569144 40225 569172 41958 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144656 40118 144684 40734 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143092 40118 143120 40151 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 143078 40151 143134 40225 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 141008 40118 141036 40174 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140976 40174 141036 40202 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 146300 40734 146352 40798 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 144644 40734 144696 40798 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 146312 40798 146340 41958 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 576768 41958 576820 42022 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 569132 41958 569184 42022 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 146300 41958 146352 42022 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 576780 42022 576808 42706 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673460 42706 673512 42770 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 576768 42706 576820 42770 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673472 42770 673500 112066 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140976 40202 141004 45698 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140964 45698 141016 45762 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42340 45698 42392 45762 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 112066 675444 112130 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673460 112066 673512 112130 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 112130 675432 112611 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 112611 675887 112639 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 112639 675887 112667 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673472 112130 673500 157286 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 157286 675444 157350 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673460 157286 673512 157350 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 157350 675432 157811 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 157811 675887 157828 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 157828 675887 157867 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 202811 675887 202844 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 202844 675887 202867 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 202867 675432 203322 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673472 157350 673500 203238 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42352 45762 42380 185438 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 184933 42193 184989 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 184989 41828 185438 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 185438 42760 185502 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42340 185438 42392 185502 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 185438 41840 185502 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673472 203238 673684 203266 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673656 203266 673684 203322 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 203322 675444 203386 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673644 203322 673696 203386 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673656 203386 673684 247454 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 185502 42748 228618 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 228133 42193 228189 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 228189 41828 228618 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 228618 42760 228682 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 228618 41840 228682 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 247454 675444 247518 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673920 247454 673972 247518 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673644 247454 673696 247518 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 247518 675432 248011 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 248011 675887 248039 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 248039 675887 248067 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 293011 675887 293012 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 293012 675887 293067 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 293067 675432 293558 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673932 247518 673960 293558 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 228682 42748 271866 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 271333 42193 271389 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 271389 41828 271866 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 271866 42760 271930 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 271866 41840 271930 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 293558 675444 293622 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673920 293558 673972 293622 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673644 293558 673696 293622 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673656 293622 673684 337486 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 271930 42748 314026 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 314026 42760 314090 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42524 314026 42576 314090 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 314026 41840 314090 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 337486 675444 337550 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673644 337486 673696 337550 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 337550 675432 338011 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 338011 675887 338028 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 338028 675887 338067 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675312 383142 675340 383182 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673656 337550 673684 383182 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42536 314090 42564 358226 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 314090 41828 314533 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 314533 42193 314589 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 357733 42193 357789 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 357789 41828 358226 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42524 358226 42576 358290 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 358226 41840 358290 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42536 358290 42564 367814 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42800 367814 42852 367878 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42524 367814 42576 367878 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42812 367878 42840 372574 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42984 372574 43036 372638 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42800 372574 42852 372638 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 383211 675887 383225 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675300 383182 675352 383225 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675300 383225 675887 383246 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673644 383182 673696 383246 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675312 383246 675887 383253 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 383253 675887 383267 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675312 383253 675340 401542 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42996 372638 43024 401254 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 400933 42193 400989 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42904 401254 43024 401282 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42904 401282 42932 401338 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 400989 41828 401338 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42892 401338 42944 401402 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 401338 41840 401402 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675300 401542 675352 401606 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673828 401542 673880 401606 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673840 401606 673868 420718 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42904 401402 42932 405690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42892 405690 42944 405754 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 405690 42668 405754 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673828 420718 673880 420782 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673644 420718 673696 420782 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673656 420782 673684 420974 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673656 420974 673776 421002 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673748 421002 673776 444314 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42628 405754 42656 422282 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 422282 42760 422346 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 422282 42668 422346 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 422346 42748 441526 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42800 441526 42852 441590 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 441526 42760 441590 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42812 441590 42840 444314 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674012 444314 674064 444378 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673736 444314 673788 444378 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42800 444314 42852 444378 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 444314 42668 444378 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674024 444378 674052 463626 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674012 463626 674064 463690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673736 463626 673788 463690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673748 463690 673776 469134 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673736 469134 673788 469198 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673828 469270 673880 469334 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673840 469334 673868 488430 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673840 488430 673960 488458 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673932 488458 673960 502318 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673920 502318 673972 502382 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673736 502318 673788 502382 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673748 502382 673776 521591 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674010 521591 674066 521665 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673734 521591 673790 521665 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674024 521665 674052 559914 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42628 444378 42656 528022 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 528022 42668 528086 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 528022 41840 528086 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42628 528086 42656 554746 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 528086 41828 528533 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 528533 42193 528589 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42800 554746 42852 554810 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 554746 42668 554810 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 559914 675444 559978 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674380 559914 674432 559978 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674012 559914 674064 559978 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 559978 675432 560411 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 560411 675887 560439 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 560439 675887 560467 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674392 559978 674420 575418 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42812 554810 42840 571202 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42800 571202 42852 571254 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 571254 42852 571266 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 571202 41840 571266 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 571266 42840 571282 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 674380 575418 674432 575482 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673736 575418 673788 575482 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673748 575482 673776 594730 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675024 594730 675076 594794 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673736 594730 673788 594794 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 605611 675887 605639 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 605639 675887 605667 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 605667 675432 606154 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675036 594794 675064 606154 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 606154 675444 606218 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675024 606154 675076 606218 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 606154 673604 606218 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 650611 675887 650639 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 650639 675887 650667 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 650667 675432 651102 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673564 606218 673592 651102 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 571282 42748 612734 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 571266 41828 571733 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 571733 42193 571789 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 612734 43024 612762 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42996 612762 43024 615470 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 614933 42193 614989 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 614989 41828 615470 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42984 615470 43036 615534 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 615470 41840 615534 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42996 615534 43024 631994 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42984 631994 43036 632058 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 631994 42760 632058 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 651102 675444 651166 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 651102 673604 651166 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673564 651166 673592 695302 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42720 632058 42748 658650 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 658133 42193 658189 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 658189 41828 658650 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42708 658650 42760 658714 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42432 658650 42484 658714 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 658650 41840 658714 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42444 658714 42472 676126 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42984 676126 43036 676190 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42432 676126 42484 676190 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42996 676190 43024 678506 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42984 678506 43036 678570 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 678506 42668 678570 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 695302 675444 695366 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 695302 673604 695366 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 695366 675432 695811 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 695811 675887 695844 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 695844 675887 695867 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673564 695366 673592 740658 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42628 678570 42656 700946 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 700946 42668 701010 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 700946 41840 701010 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42628 701010 42656 739570 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 701010 41828 701333 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 701333 42193 701389 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 739570 42668 739634 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42340 739570 42392 739634 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 740658 675444 740722 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 740658 673604 740722 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 740722 675432 740811 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 740811 675887 740860 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 740860 675887 740867 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 785811 675887 785839 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 785839 675887 785867 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 785867 675432 786354 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673564 740722 673592 786354 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42352 739634 42380 744126 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 744126 42668 744190 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42340 744126 42392 744190 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 744126 41840 744190 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 786354 675444 786418 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 786354 673604 786418 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673564 786418 673592 874482 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42628 744190 42656 787238 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 744190 41828 744533 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 744533 42193 744589 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42616 787238 42668 787302 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 787238 41840 787302 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 787302 41828 787733 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 787733 42193 787789 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 874482 675444 874546 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 874482 673604 874546 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 874546 675432 875011 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 875011 675887 875039 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 875039 675887 875067 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675407 964211 675887 964239 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 964239 675887 964267 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675404 964267 675432 964718 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673564 874546 673592 964718 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41713 957533 42193 957589 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41800 957589 41828 958054 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42340 958054 42392 958118 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 41788 958054 41840 958118 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 675392 964718 675444 964782 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 964718 673604 964782 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673564 964782 673592 990082 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42352 958118 42380 990082 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 673552 990082 673604 990146 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 631232 990082 631284 990146 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 79508 990082 79560 990146 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 42340 990082 42392 990146 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 631244 990146 631272 990694 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 173900 990218 173952 990282 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140780 990218 140832 990270 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140700 990270 140832 990282 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 131028 990218 131080 990282 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 173912 990282 173940 990354 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140700 990282 140820 990286 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 160008 990286 160060 990350 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140688 990286 140820 990298 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 140688 990298 140740 990350 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 182456 990354 182508 990418 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 173900 990354 173952 990418 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 160020 990350 160048 990406 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 131040 990282 131068 990383 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 400128 990422 400180 990486 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 387156 990422 387208 990486 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 386420 990422 386472 990486 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 477408 990490 477460 990554 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 476120 990490 476172 990554 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 458180 990490 458232 990554 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 438768 990490 438820 990554 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 419540 990490 419592 990554 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 477420 990554 477448 990694 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 631232 990694 631284 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 629300 990694 629352 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 527548 990694 527600 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 477408 990694 477460 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 629312 990758 629340 995407 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 527560 990758 527588 995407 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 476132 990554 476160 995407 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 458192 990554 458220 990694 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 438780 990554 438808 990694 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 419552 990554 419580 990694 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 400140 990486 400168 990694 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 458180 990694 458232 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 438768 990694 438820 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 419540 990694 419592 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 400128 990694 400180 990758 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 629312 995407 629389 995466 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 629333 995466 629389 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 527533 995407 527589 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 476132 995407 476189 995452 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 387168 990486 387196 995407 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 386432 990486 386460 990626 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 386420 990626 386472 990690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 345020 990626 345072 990644 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 345020 990644 345152 990672 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 345124 990672 345152 990762 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 345020 990672 345072 990690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 342168 990626 342220 990690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 285312 990626 285364 990690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 233700 990626 233752 990690 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 372620 990762 372672 990814 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 372528 990762 372580 990814 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 372528 990814 372672 990826 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 345112 990762 345164 990826 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 372540 990826 372660 990842 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 387133 995407 387196 995452 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 476133 995452 476189 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 387133 995452 387189 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 342180 990690 342208 997405 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 285324 990690 285352 995407 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 233712 990690 233740 995407 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 285324 995407 285389 995452 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 285333 995452 285389 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 233712 995407 233789 995466 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 182468 990418 182496 995438 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 160020 990406 160232 990422 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 160020 990422 160244 990434 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 160192 990434 160244 990486 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 131026 990383 131082 990457 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 121274 990383 121330 990457 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 182333 995407 182389 995438 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 182333 995438 182496 995466 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 131040 990457 131068 995438 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 121288 990457 121316 990558 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 121276 990558 121328 990622 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 79520 990146 79548 995407 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 130933 995407 130989 995438 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 130933 995438 131068 995466 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 233733 995466 233789 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 182333 995466 182389 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 130933 995466 130989 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 79520 995407 79589 995452 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 79533 995452 79589 995887 6 vssio
port 76 nsew signal bidirectional
rlabel metal2 s 342164 997405 342224 997483 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 144644 40060 144696 40112 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 143080 40060 143132 40112 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 140996 40060 141048 40112 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 146300 40740 146352 40792 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 144644 40740 144696 40792 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 576768 41964 576820 42016 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 569132 41964 569184 42016 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 146300 41964 146352 42016 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673460 42712 673512 42764 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 576768 42712 576820 42764 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 140964 45704 141016 45756 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42340 45704 42392 45756 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 112072 675444 112124 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673460 112072 673512 112124 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 157292 675444 157344 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673460 157292 673512 157344 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 185444 42760 185496 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42340 185444 42392 185496 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 185444 41840 185496 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 203328 675444 203380 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673644 203328 673696 203380 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 228624 42760 228676 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 228624 41840 228676 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 247460 675444 247512 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673920 247460 673972 247512 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673644 247460 673696 247512 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 271872 42760 271924 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 271872 41840 271924 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 293564 675444 293616 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673920 293564 673972 293616 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673644 293564 673696 293616 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 314032 42760 314084 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42524 314032 42576 314084 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 314032 41840 314084 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 337492 675444 337544 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673644 337492 673696 337544 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42524 358232 42576 358284 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 358232 41840 358284 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42800 367820 42852 367872 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42524 367820 42576 367872 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42984 372580 43036 372632 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42800 372580 42852 372632 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675300 383188 675352 383240 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673644 383188 673696 383240 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42892 401344 42944 401396 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 401344 41840 401396 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675300 401548 675352 401600 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673828 401548 673880 401600 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42892 405696 42944 405748 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 405696 42668 405748 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673828 420724 673880 420776 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673644 420724 673696 420776 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 422288 42760 422340 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 422288 42668 422340 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42800 441532 42852 441584 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 441532 42760 441584 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 674012 444320 674064 444372 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673736 444320 673788 444372 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42800 444320 42852 444372 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 444320 42668 444372 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 674012 463632 674064 463684 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673736 463632 673788 463684 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673736 469140 673788 469192 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673828 469276 673880 469328 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673920 502324 673972 502376 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673736 502324 673788 502376 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 528028 42668 528080 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 528028 41840 528080 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42800 554752 42852 554804 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 554752 42668 554804 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 559920 675444 559972 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 674380 559920 674432 559972 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 674012 559920 674064 559972 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42800 571208 42852 571260 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 571208 41840 571260 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 674380 575424 674432 575476 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673736 575424 673788 575476 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675024 594736 675076 594788 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673736 594736 673788 594788 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 606160 675444 606212 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675024 606160 675076 606212 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 606160 673604 606212 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42984 615476 43036 615528 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 615476 41840 615528 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42984 632000 43036 632052 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 632000 42760 632052 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 651108 675444 651160 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 651108 673604 651160 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42708 658656 42760 658708 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42432 658656 42484 658708 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 658656 41840 658708 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42984 676132 43036 676184 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42432 676132 42484 676184 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42984 678512 43036 678564 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 678512 42668 678564 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 695308 675444 695360 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 695308 673604 695360 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 700952 42668 701004 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 700952 41840 701004 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 739576 42668 739628 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42340 739576 42392 739628 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 740664 675444 740716 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 740664 673604 740716 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 744132 42668 744184 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42340 744132 42392 744184 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 744132 41840 744184 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 786360 675444 786412 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 786360 673604 786412 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42616 787244 42668 787296 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 787244 41840 787296 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 874488 675444 874540 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 874488 673604 874540 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42340 958060 42392 958112 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 41788 958060 41840 958112 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 675392 964724 675444 964776 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 964724 673604 964776 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 673552 990088 673604 990140 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 631232 990088 631284 990140 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 173900 990224 173952 990276 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 160008 990292 160060 990344 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 140780 990224 140832 990276 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 140688 990292 140740 990344 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 131028 990224 131080 990276 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 79508 990088 79560 990140 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 42340 990088 42392 990140 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 400128 990428 400180 990480 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 387156 990428 387208 990480 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 386420 990428 386472 990480 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 477408 990496 477460 990548 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 476120 990496 476172 990548 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 458180 990496 458232 990548 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 438768 990496 438820 990548 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 419540 990496 419592 990548 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 386420 990632 386472 990684 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 631232 990700 631284 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 629300 990700 629352 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 527548 990700 527600 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 477408 990700 477460 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 458180 990700 458232 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 438768 990700 438820 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 419540 990700 419592 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 400128 990700 400180 990752 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 345020 990632 345072 990684 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 342168 990632 342220 990684 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 285312 990632 285364 990684 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 233700 990632 233752 990684 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 182456 990360 182508 990412 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 173900 990360 173952 990412 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 160192 990428 160244 990480 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 121276 990564 121328 990616 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 372620 990768 372672 990820 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 372528 990768 372580 990820 6 vssio
port 76 nsew signal bidirectional
rlabel via1 s 345112 990768 345164 990820 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 142573 38005 142619 40000 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 144638 40060 144702 40072 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 143074 40060 143138 40072 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 142586 40000 142614 40072 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140990 40060 141054 40072 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140990 40072 144702 40100 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 144638 40100 144702 40112 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 143074 40100 143138 40112 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140990 40100 141054 40112 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 146294 40740 146358 40752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 144638 40740 144702 40752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 144638 40752 146358 40780 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 146294 40780 146358 40792 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 144638 40780 144702 40792 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 576762 41964 576826 41976 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 569126 41964 569190 41976 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 146294 41964 146358 41976 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 146294 41976 576826 42004 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 576762 42004 576826 42016 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 569126 42004 569190 42016 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 146294 42004 146358 42016 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 42712 673518 42724 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 576762 42712 576826 42724 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 576762 42724 673518 42752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 42752 673518 42764 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 576762 42752 576826 42764 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140958 45704 141022 45716 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 45704 42398 45716 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 45716 141022 45744 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140958 45744 141022 45756 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 45744 42398 45756 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 112072 675450 112084 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 112072 673518 112084 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 112084 675450 112112 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 112112 675450 112124 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 112112 673518 112124 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 157292 675450 157304 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 157292 673518 157304 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 157304 675450 157332 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 157332 675450 157344 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673454 157332 673518 157344 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 185444 42766 185456 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 185444 42398 185456 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 185444 41846 185456 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 185456 42766 185484 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 185484 42766 185496 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 185484 42398 185496 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 185484 41846 185496 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 203328 675450 203340 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 203328 673702 203340 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 203340 675450 203368 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 203368 675450 203380 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 203368 673702 203380 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 228624 42766 228636 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 228624 41846 228636 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 228636 42766 228664 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 228664 42766 228676 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 228664 41846 228676 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 247460 675450 247472 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673914 247460 673978 247472 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 247460 673702 247472 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 247472 675450 247500 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 247500 675450 247512 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673914 247500 673978 247512 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 247500 673702 247512 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 271872 42766 271884 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 271872 41846 271884 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 271884 42766 271912 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 271912 42766 271924 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 271912 41846 271924 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 293564 675450 293576 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673914 293564 673978 293576 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 293564 673702 293576 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 293576 675450 293604 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 293604 675450 293616 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673914 293604 673978 293616 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 293604 673702 293616 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 314032 42766 314044 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42518 314032 42582 314044 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 314032 41846 314044 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 314044 42766 314072 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 314072 42766 314084 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42518 314072 42582 314084 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 314072 41846 314084 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 337492 675450 337504 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 337492 673702 337504 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 337504 675450 337532 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 337532 675450 337544 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 337532 673702 337544 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42518 358232 42582 358244 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 358232 41846 358244 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 358244 42582 358272 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42518 358272 42582 358284 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 358272 41846 358284 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 367820 42858 367832 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42518 367820 42582 367832 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42518 367832 42858 367860 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 367860 42858 367872 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42518 367860 42582 367872 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 372580 43042 372592 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 372580 42858 372592 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 372592 43042 372620 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 372620 43042 372632 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 372620 42858 372632 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675294 383188 675358 383200 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 383188 673702 383200 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 383200 675358 383228 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675294 383228 675358 383240 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 383228 673702 383240 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42886 401344 42950 401356 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 401344 41846 401356 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 401356 42950 401384 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42886 401384 42950 401396 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 401384 41846 401396 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675294 401548 675358 401560 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673822 401548 673886 401560 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673822 401560 675358 401588 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675294 401588 675358 401600 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673822 401588 673886 401600 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42886 405696 42950 405708 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 405696 42674 405708 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 405708 42950 405736 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42886 405736 42950 405748 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 405736 42674 405748 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673822 420724 673886 420736 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 420724 673702 420736 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 420736 673886 420764 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673822 420764 673886 420776 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673638 420764 673702 420776 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 422288 42766 422300 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 422288 42674 422300 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 422300 42766 422328 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 422328 42766 422340 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 422328 42674 422340 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 441532 42858 441544 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 441532 42766 441544 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 441544 42858 441572 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 441572 42858 441584 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 441572 42766 441584 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674006 444320 674070 444332 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 444320 673794 444332 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 444332 674070 444360 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674006 444360 674070 444372 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 444360 673794 444372 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 444320 42858 444332 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 444320 42674 444332 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 444332 42858 444360 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 444360 42858 444372 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 444360 42674 444372 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674006 463632 674070 463644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 463632 673794 463644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 463644 674070 463672 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674006 463672 674070 463684 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 463672 673794 463684 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 469140 673794 469192 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673822 469276 673886 469288 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673748 469192 673776 469288 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673748 469288 673886 469316 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673822 469316 673886 469328 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673914 502324 673978 502336 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 502324 673794 502336 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 502336 673978 502364 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673914 502364 673978 502376 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 502364 673794 502376 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 528028 42674 528040 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 528028 41846 528040 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 528040 42674 528068 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 528068 42674 528080 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 528068 41846 528080 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 554752 42858 554764 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 554752 42674 554764 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 554764 42858 554792 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 554792 42858 554804 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 554792 42674 554804 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 559920 675450 559932 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674374 559920 674438 559932 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674006 559920 674070 559932 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674006 559932 675450 559960 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 559960 675450 559972 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674374 559960 674438 559972 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674006 559960 674070 559972 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 571208 42858 571220 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 571208 41846 571220 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 571220 42858 571248 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42794 571248 42858 571260 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 571248 41846 571260 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674374 575424 674438 575436 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 575424 673794 575436 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 575436 674438 575464 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 674374 575464 674438 575476 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 575464 673794 575476 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675018 594736 675082 594748 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 594736 673794 594748 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 594748 675082 594776 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675018 594776 675082 594788 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673730 594776 673794 594788 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 606160 675450 606172 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675018 606160 675082 606172 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 606160 673610 606172 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 606172 675450 606200 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 606200 675450 606212 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675018 606200 675082 606212 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 606200 673610 606212 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 615476 43042 615488 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 615476 41846 615488 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 615488 43042 615516 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 615516 43042 615528 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 615516 41846 615528 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 632000 43042 632012 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 632000 42766 632012 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 632012 43042 632040 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 632040 43042 632052 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 632040 42766 632052 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 651108 675450 651120 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 651108 673610 651120 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 651120 675450 651148 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 651148 675450 651160 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 651148 673610 651160 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 658656 42766 658668 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42426 658656 42490 658668 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 658656 41846 658668 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 658668 42766 658696 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42702 658696 42766 658708 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42426 658696 42490 658708 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 658696 41846 658708 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 676132 43042 676144 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42426 676132 42490 676144 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42426 676144 43042 676172 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 676172 43042 676184 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42426 676172 42490 676184 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 678512 43042 678524 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 678512 42674 678524 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 678524 43042 678552 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42978 678552 43042 678564 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 678552 42674 678564 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 695308 675450 695320 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 695308 673610 695320 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 695320 675450 695348 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 695348 675450 695360 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 695348 673610 695360 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 700952 42674 700964 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 700952 41846 700964 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 700964 42674 700992 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 700992 42674 701004 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 700992 41846 701004 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 739576 42674 739588 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 739576 42398 739588 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 739588 42674 739616 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 739616 42674 739628 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 739616 42398 739628 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 740664 675450 740676 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 740664 673610 740676 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 740676 675450 740704 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 740704 675450 740716 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 740704 673610 740716 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 744132 42674 744144 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 744132 42398 744144 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 744132 41846 744144 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 744144 42674 744172 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 744172 42674 744184 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 744172 42398 744184 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 744172 41846 744184 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 786360 675450 786372 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 786360 673610 786372 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 786372 675450 786400 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 786400 675450 786412 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 786400 673610 786412 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 787244 42674 787256 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 787244 41846 787256 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 787256 42674 787284 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42610 787284 42674 787296 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 787284 41846 787296 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 874488 675450 874500 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 874488 673610 874500 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 874500 675450 874528 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 874528 675450 874540 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 874528 673610 874540 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 958060 42398 958072 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 958060 41846 958072 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 958072 42398 958100 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 958100 42398 958112 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 41782 958100 41846 958112 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 964724 675450 964736 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 964724 673610 964736 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 964736 675450 964764 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 675386 964764 675450 964776 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 964764 673610 964776 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 990088 673610 990100 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 631226 990088 631290 990100 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 79502 990088 79566 990100 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 990088 42398 990100 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 631226 990100 673610 990128 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 673546 990128 673610 990140 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 631226 990128 631290 990140 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 990100 84424 990128 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 173894 990224 173958 990236 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140774 990224 140838 990236 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 131022 990224 131086 990236 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 84396 990128 84424 990236 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 79502 990128 79566 990140 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 42334 990128 42398 990140 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 173894 990236 182496 990264 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 182468 990264 182496 990360 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 173894 990264 173958 990276 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140774 990236 154528 990264 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 160002 990292 160066 990304 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 154500 990264 154528 990304 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140774 990264 140838 990276 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 131022 990236 135300 990264 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 154500 990304 160066 990332 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140682 990292 140746 990304 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 135272 990264 135300 990304 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 131022 990264 131086 990276 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 84396 990236 96568 990264 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 135272 990304 140746 990332 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 160002 990332 160066 990344 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 140682 990332 140746 990344 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 182450 990360 182514 990372 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 182450 990372 195100 990400 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 400122 990428 400186 990440 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 387150 990428 387214 990440 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 386414 990428 386478 990440 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 386414 990440 400186 990468 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 400122 990468 400186 990480 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 387150 990468 387214 990480 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 386414 990468 386478 990480 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 477402 990496 477466 990508 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 476114 990496 476178 990508 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 458174 990496 458238 990508 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 458174 990508 477466 990536 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 477402 990536 477466 990548 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 476114 990536 476178 990548 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 458174 990536 458238 990548 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 438762 990496 438826 990508 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 419534 990496 419598 990508 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 419534 990508 438826 990536 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 438762 990536 438826 990548 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 419534 990536 419598 990548 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 386414 990632 386478 990644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 345014 990632 345078 990644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 342162 990632 342226 990644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 285306 990632 285370 990644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 233694 990632 233758 990644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 195072 990400 195100 990644 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 182450 990400 182514 990412 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 173894 990360 173958 990412 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 173912 990412 173940 990440 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 160186 990428 160250 990440 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 160186 990440 173940 990468 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 160186 990468 160250 990480 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 96540 990264 96568 990508 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 96540 990508 102088 990536 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 121270 990564 121334 990576 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 102060 990536 102088 990576 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 102060 990576 121334 990604 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 121270 990604 121334 990616 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 383580 990644 386478 990672 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 386414 990672 386478 990684 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 631226 990700 631290 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 629294 990700 629358 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 527542 990700 527606 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 477402 990700 477466 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 477402 990712 631290 990740 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 631226 990740 631290 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 629294 990740 629358 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 527542 990740 527606 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 477402 990740 477466 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 458174 990700 458238 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 438762 990700 438826 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 438762 990712 458238 990740 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 458174 990740 458238 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 438762 990740 438826 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 419534 990700 419598 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 400122 990700 400186 990712 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 400122 990712 419598 990740 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 419534 990740 419598 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 400122 990740 400186 990752 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 383580 990672 383608 990780 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 195072 990644 345078 990672 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 345014 990672 345078 990684 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 342162 990672 342226 990684 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 285306 990672 285370 990684 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 233694 990672 233758 990684 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 372614 990768 372678 990780 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 372614 990780 383608 990808 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 372614 990808 372678 990820 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 372522 990768 372586 990780 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 345106 990768 345170 990780 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 345106 990780 372586 990808 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 372522 990808 372586 990820 6 vssio
port 76 nsew signal bidirectional
rlabel metal1 s 345106 990808 345170 990820 6 vssio
port 76 nsew signal bidirectional
rlabel metal4 s 333400 1032757 333654 1037600 6 vssio
port 77 nsew signal bidirectional
rlabel metal4 s 348146 1032757 348400 1037600 6 vssio
port 78 nsew signal bidirectional
rlabel metal4 s 348146 1002767 384054 1003697 6 vssio
port 79 nsew signal bidirectional
rlabel metal5 s 297746 1002787 333654 1003677 6 vssio
port 80 nsew signal bidirectional
rlabel metal5 s 348146 1002787 384054 1003677 6 vssio
port 81 nsew signal bidirectional
rlabel metal3 s 333499 997600 338279 1002770 6 vssio
port 82 nsew signal bidirectional
rlabel metal5 s 334620 1018402 347160 1030925 6 vssio
port 83 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 84 nsew signal bidirectional
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 85 nsew signal input
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 86 nsew signal input
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 87 nsew signal input
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 88 nsew signal input
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 89 nsew signal input
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 90 nsew signal input
rlabel metal2 s 675407 108931 675887 108987 6 mprj_io_enh[0]
port 91 nsew signal input
rlabel metal2 s 675407 109575 675887 109631 6 mprj_io_hldh_n[0]
port 92 nsew signal input
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 93 nsew signal input
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 94 nsew signal input
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 95 nsew signal input
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 96 nsew signal input
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 97 nsew signal input
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 98 nsew signal input
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 99 nsew signal input
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 100 nsew signal output
rlabel metal2 s 675407 686611 675887 686667 6 mprj_analog_io[3]
port 101 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 102 nsew signal bidirectional
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 103 nsew signal input
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 104 nsew signal input
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 105 nsew signal input
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 106 nsew signal input
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 107 nsew signal input
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 108 nsew signal input
rlabel metal2 s 675407 692131 675887 692187 6 mprj_io_enh[10]
port 109 nsew signal input
rlabel metal2 s 675407 692775 675887 692831 6 mprj_io_hldh_n[10]
port 110 nsew signal input
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 111 nsew signal input
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 112 nsew signal input
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 113 nsew signal input
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 114 nsew signal input
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 115 nsew signal input
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 116 nsew signal input
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 117 nsew signal input
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 118 nsew signal output
rlabel metal2 s 675407 731611 675887 731667 6 mprj_analog_io[4]
port 119 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 120 nsew signal bidirectional
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 121 nsew signal input
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 122 nsew signal input
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 123 nsew signal input
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 124 nsew signal input
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 125 nsew signal input
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 126 nsew signal input
rlabel metal2 s 675407 737131 675887 737187 6 mprj_io_enh[11]
port 127 nsew signal input
rlabel metal2 s 675407 737775 675887 737831 6 mprj_io_hldh_n[11]
port 128 nsew signal input
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 129 nsew signal input
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 130 nsew signal input
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 131 nsew signal input
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 132 nsew signal input
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 133 nsew signal input
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 134 nsew signal input
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 135 nsew signal input
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 136 nsew signal output
rlabel metal2 s 675407 776611 675887 776667 6 mprj_analog_io[5]
port 137 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 138 nsew signal bidirectional
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 139 nsew signal input
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 140 nsew signal input
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 141 nsew signal input
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 142 nsew signal input
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 143 nsew signal input
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 144 nsew signal input
rlabel metal2 s 675407 782131 675887 782187 6 mprj_io_enh[12]
port 145 nsew signal input
rlabel metal2 s 675407 782775 675887 782831 6 mprj_io_hldh_n[12]
port 146 nsew signal input
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 147 nsew signal input
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 148 nsew signal input
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 149 nsew signal input
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 150 nsew signal input
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 151 nsew signal input
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 152 nsew signal input
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 153 nsew signal input
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 154 nsew signal output
rlabel metal2 s 675407 865811 675887 865867 6 mprj_analog_io[6]
port 155 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 156 nsew signal bidirectional
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 157 nsew signal input
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 158 nsew signal input
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 159 nsew signal input
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 160 nsew signal input
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 161 nsew signal input
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 162 nsew signal input
rlabel metal2 s 675407 871331 675887 871387 6 mprj_io_enh[13]
port 163 nsew signal input
rlabel metal2 s 675407 871975 675887 872031 6 mprj_io_hldh_n[13]
port 164 nsew signal input
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 165 nsew signal input
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 166 nsew signal input
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 167 nsew signal input
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 168 nsew signal input
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 169 nsew signal input
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 170 nsew signal input
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 171 nsew signal input
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 172 nsew signal output
rlabel metal2 s 675407 955011 675887 955067 6 mprj_analog_io[7]
port 173 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 174 nsew signal bidirectional
rlabel metal2 s 675407 957403 675887 957459 6 mprj_io_analog_en[14]
port 175 nsew signal input
rlabel metal2 s 675407 958691 675887 958747 6 mprj_io_analog_pol[14]
port 176 nsew signal input
rlabel metal2 s 675407 961727 675887 961783 6 mprj_io_analog_sel[14]
port 177 nsew signal input
rlabel metal2 s 675407 958047 675887 958103 6 mprj_io_dm[42]
port 178 nsew signal input
rlabel metal2 s 675407 956207 675887 956263 6 mprj_io_dm[43]
port 179 nsew signal input
rlabel metal2 s 675407 962371 675887 962427 6 mprj_io_dm[44]
port 180 nsew signal input
rlabel metal2 s 675407 960531 675887 960587 6 mprj_io_enh[14]
port 181 nsew signal input
rlabel metal2 s 675407 961175 675887 961231 6 mprj_io_hldh_n[14]
port 182 nsew signal input
rlabel metal2 s 675407 963015 675887 963071 6 mprj_io_holdover[14]
port 183 nsew signal input
rlabel metal2 s 675407 966051 675887 966107 6 mprj_io_ib_mode_sel[14]
port 184 nsew signal input
rlabel metal2 s 675407 959243 675887 959299 6 mprj_io_inp_dis[14]
port 185 nsew signal input
rlabel metal2 s 675407 966695 675887 966751 6 mprj_io_oeb[14]
port 186 nsew signal input
rlabel metal2 s 675407 963567 675887 963623 6 mprj_io_out[14]
port 187 nsew signal input
rlabel metal2 s 675407 954367 675887 954423 6 mprj_io_slow_sel[14]
port 188 nsew signal input
rlabel metal2 s 675407 965407 675887 965463 6 mprj_io_vtrip_sel[14]
port 189 nsew signal input
rlabel metal2 s 675407 952527 675887 952583 6 mprj_io_in[14]
port 190 nsew signal output
rlabel metal2 s 638533 995407 638589 995887 6 mprj_analog_io[8]
port 191 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 192 nsew signal bidirectional
rlabel metal2 s 636141 995407 636197 995887 6 mprj_io_analog_en[15]
port 193 nsew signal input
rlabel metal2 s 634853 995407 634909 995887 6 mprj_io_analog_pol[15]
port 194 nsew signal input
rlabel metal2 s 631817 995407 631873 995887 6 mprj_io_analog_sel[15]
port 195 nsew signal input
rlabel metal2 s 635497 995407 635553 995887 6 mprj_io_dm[45]
port 196 nsew signal input
rlabel metal2 s 637337 995407 637393 995887 6 mprj_io_dm[46]
port 197 nsew signal input
rlabel metal2 s 631173 995407 631229 995887 6 mprj_io_dm[47]
port 198 nsew signal input
rlabel metal2 s 633013 995407 633069 995887 6 mprj_io_enh[15]
port 199 nsew signal input
rlabel metal2 s 632369 995407 632425 995887 6 mprj_io_hldh_n[15]
port 200 nsew signal input
rlabel metal2 s 630529 995407 630585 995887 6 mprj_io_holdover[15]
port 201 nsew signal input
rlabel metal2 s 627493 995407 627549 995887 6 mprj_io_ib_mode_sel[15]
port 202 nsew signal input
rlabel metal2 s 634301 995407 634357 995887 6 mprj_io_inp_dis[15]
port 203 nsew signal input
rlabel metal2 s 626849 995407 626905 995887 6 mprj_io_oeb[15]
port 204 nsew signal input
rlabel metal2 s 629977 995407 630033 995887 6 mprj_io_out[15]
port 205 nsew signal input
rlabel metal2 s 639177 995407 639233 995887 6 mprj_io_slow_sel[15]
port 206 nsew signal input
rlabel metal2 s 628137 995407 628193 995887 6 mprj_io_vtrip_sel[15]
port 207 nsew signal input
rlabel metal2 s 641017 995407 641073 995887 6 mprj_io_in[15]
port 208 nsew signal output
rlabel metal2 s 536733 995407 536789 995887 6 mprj_analog_io[9]
port 209 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 210 nsew signal bidirectional
rlabel metal2 s 534341 995407 534397 995887 6 mprj_io_analog_en[16]
port 211 nsew signal input
rlabel metal2 s 533053 995407 533109 995887 6 mprj_io_analog_pol[16]
port 212 nsew signal input
rlabel metal2 s 530017 995407 530073 995887 6 mprj_io_analog_sel[16]
port 213 nsew signal input
rlabel metal2 s 533697 995407 533753 995887 6 mprj_io_dm[48]
port 214 nsew signal input
rlabel metal2 s 535537 995407 535593 995887 6 mprj_io_dm[49]
port 215 nsew signal input
rlabel metal2 s 529373 995407 529429 995887 6 mprj_io_dm[50]
port 216 nsew signal input
rlabel metal2 s 531213 995407 531269 995887 6 mprj_io_enh[16]
port 217 nsew signal input
rlabel metal2 s 530569 995407 530625 995887 6 mprj_io_hldh_n[16]
port 218 nsew signal input
rlabel metal2 s 528729 995407 528785 995887 6 mprj_io_holdover[16]
port 219 nsew signal input
rlabel metal2 s 525693 995407 525749 995887 6 mprj_io_ib_mode_sel[16]
port 220 nsew signal input
rlabel metal2 s 532501 995407 532557 995887 6 mprj_io_inp_dis[16]
port 221 nsew signal input
rlabel metal2 s 525049 995407 525105 995887 6 mprj_io_oeb[16]
port 222 nsew signal input
rlabel metal2 s 528177 995407 528233 995887 6 mprj_io_out[16]
port 223 nsew signal input
rlabel metal2 s 537377 995407 537433 995887 6 mprj_io_slow_sel[16]
port 224 nsew signal input
rlabel metal2 s 526337 995407 526393 995887 6 mprj_io_vtrip_sel[16]
port 225 nsew signal input
rlabel metal2 s 539217 995407 539273 995887 6 mprj_io_in[16]
port 226 nsew signal output
rlabel metal2 s 485333 995407 485389 995887 6 mprj_analog_io[10]
port 227 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 228 nsew signal bidirectional
rlabel metal2 s 482941 995407 482997 995887 6 mprj_io_analog_en[17]
port 229 nsew signal input
rlabel metal2 s 481653 995407 481709 995887 6 mprj_io_analog_pol[17]
port 230 nsew signal input
rlabel metal2 s 478617 995407 478673 995887 6 mprj_io_analog_sel[17]
port 231 nsew signal input
rlabel metal2 s 482297 995407 482353 995887 6 mprj_io_dm[51]
port 232 nsew signal input
rlabel metal2 s 484137 995407 484193 995887 6 mprj_io_dm[52]
port 233 nsew signal input
rlabel metal2 s 477973 995407 478029 995887 6 mprj_io_dm[53]
port 234 nsew signal input
rlabel metal2 s 479813 995407 479869 995887 6 mprj_io_enh[17]
port 235 nsew signal input
rlabel metal2 s 479169 995407 479225 995887 6 mprj_io_hldh_n[17]
port 236 nsew signal input
rlabel metal2 s 477329 995407 477385 995887 6 mprj_io_holdover[17]
port 237 nsew signal input
rlabel metal2 s 474293 995407 474349 995887 6 mprj_io_ib_mode_sel[17]
port 238 nsew signal input
rlabel metal2 s 481101 995407 481157 995887 6 mprj_io_inp_dis[17]
port 239 nsew signal input
rlabel metal2 s 473649 995407 473705 995887 6 mprj_io_oeb[17]
port 240 nsew signal input
rlabel metal2 s 476777 995407 476833 995887 6 mprj_io_out[17]
port 241 nsew signal input
rlabel metal2 s 485977 995407 486033 995887 6 mprj_io_slow_sel[17]
port 242 nsew signal input
rlabel metal2 s 474937 995407 474993 995887 6 mprj_io_vtrip_sel[17]
port 243 nsew signal input
rlabel metal2 s 487817 995407 487873 995887 6 mprj_io_in[17]
port 244 nsew signal output
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 245 nsew signal bidirectional
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 246 nsew signal input
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 247 nsew signal input
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 248 nsew signal input
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 249 nsew signal input
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 250 nsew signal input
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 251 nsew signal input
rlabel metal2 s 675407 154131 675887 154187 6 mprj_io_enh[1]
port 252 nsew signal input
rlabel metal2 s 675407 154775 675887 154831 6 mprj_io_hldh_n[1]
port 253 nsew signal input
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 254 nsew signal input
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 255 nsew signal input
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 256 nsew signal input
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 257 nsew signal input
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 258 nsew signal input
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 259 nsew signal input
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 260 nsew signal input
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 261 nsew signal output
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 262 nsew signal bidirectional
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 263 nsew signal input
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 264 nsew signal input
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 265 nsew signal input
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 266 nsew signal input
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 267 nsew signal input
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 268 nsew signal input
rlabel metal2 s 675407 199131 675887 199187 6 mprj_io_enh[2]
port 269 nsew signal input
rlabel metal2 s 675407 199775 675887 199831 6 mprj_io_hldh_n[2]
port 270 nsew signal input
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 271 nsew signal input
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 272 nsew signal input
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 273 nsew signal input
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 274 nsew signal input
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 275 nsew signal input
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 276 nsew signal input
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 277 nsew signal input
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 278 nsew signal output
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 279 nsew signal bidirectional
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 280 nsew signal input
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 281 nsew signal input
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 282 nsew signal input
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 283 nsew signal input
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 284 nsew signal input
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 285 nsew signal input
rlabel metal2 s 675407 244331 675887 244387 6 mprj_io_enh[3]
port 286 nsew signal input
rlabel metal2 s 675407 244975 675887 245031 6 mprj_io_hldh_n[3]
port 287 nsew signal input
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 288 nsew signal input
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 289 nsew signal input
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 290 nsew signal input
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 291 nsew signal input
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 292 nsew signal input
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 293 nsew signal input
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 294 nsew signal input
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 295 nsew signal output
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 296 nsew signal bidirectional
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 297 nsew signal input
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 298 nsew signal input
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 299 nsew signal input
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 300 nsew signal input
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 301 nsew signal input
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 302 nsew signal input
rlabel metal2 s 675407 289331 675887 289387 6 mprj_io_enh[4]
port 303 nsew signal input
rlabel metal2 s 675407 289975 675887 290031 6 mprj_io_hldh_n[4]
port 304 nsew signal input
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 305 nsew signal input
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 306 nsew signal input
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 307 nsew signal input
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 308 nsew signal input
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 309 nsew signal input
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 310 nsew signal input
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 311 nsew signal input
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 312 nsew signal output
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 313 nsew signal bidirectional
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 314 nsew signal input
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 315 nsew signal input
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 316 nsew signal input
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 317 nsew signal input
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 318 nsew signal input
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 319 nsew signal input
rlabel metal2 s 675407 334331 675887 334387 6 mprj_io_enh[5]
port 320 nsew signal input
rlabel metal2 s 675407 334975 675887 335031 6 mprj_io_hldh_n[5]
port 321 nsew signal input
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 322 nsew signal input
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 323 nsew signal input
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 324 nsew signal input
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 325 nsew signal input
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 326 nsew signal input
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 327 nsew signal input
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 328 nsew signal input
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 329 nsew signal output
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 330 nsew signal bidirectional
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 331 nsew signal input
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 332 nsew signal input
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 333 nsew signal input
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 334 nsew signal input
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 335 nsew signal input
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 336 nsew signal input
rlabel metal2 s 675407 379531 675887 379587 6 mprj_io_enh[6]
port 337 nsew signal input
rlabel metal2 s 675407 380175 675887 380231 6 mprj_io_hldh_n[6]
port 338 nsew signal input
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 339 nsew signal input
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 340 nsew signal input
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 341 nsew signal input
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 342 nsew signal input
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 343 nsew signal input
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 344 nsew signal input
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 345 nsew signal input
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 346 nsew signal output
rlabel metal2 s 675407 551211 675887 551267 6 mprj_analog_io[0]
port 347 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 348 nsew signal bidirectional
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 349 nsew signal input
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 350 nsew signal input
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 351 nsew signal input
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 352 nsew signal input
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 353 nsew signal input
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 354 nsew signal input
rlabel metal2 s 675407 556731 675887 556787 6 mprj_io_enh[7]
port 355 nsew signal input
rlabel metal2 s 675407 557375 675887 557431 6 mprj_io_hldh_n[7]
port 356 nsew signal input
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 357 nsew signal input
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 358 nsew signal input
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 359 nsew signal input
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 360 nsew signal input
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 361 nsew signal input
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 362 nsew signal input
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 363 nsew signal input
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 364 nsew signal output
rlabel metal2 s 675407 596411 675887 596467 6 mprj_analog_io[1]
port 365 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 366 nsew signal bidirectional
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 367 nsew signal input
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 368 nsew signal input
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 369 nsew signal input
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 370 nsew signal input
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 371 nsew signal input
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 372 nsew signal input
rlabel metal2 s 675407 601931 675887 601987 6 mprj_io_enh[8]
port 373 nsew signal input
rlabel metal2 s 675407 602575 675887 602631 6 mprj_io_hldh_n[8]
port 374 nsew signal input
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 375 nsew signal input
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 376 nsew signal input
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 377 nsew signal input
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 378 nsew signal input
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 379 nsew signal input
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 380 nsew signal input
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 381 nsew signal input
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 382 nsew signal output
rlabel metal2 s 675407 641411 675887 641467 6 mprj_analog_io[2]
port 383 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 384 nsew signal bidirectional
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 385 nsew signal input
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 386 nsew signal input
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 387 nsew signal input
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 388 nsew signal input
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 389 nsew signal input
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 390 nsew signal input
rlabel metal2 s 675407 646931 675887 646987 6 mprj_io_enh[9]
port 391 nsew signal input
rlabel metal2 s 675407 647575 675887 647631 6 mprj_io_hldh_n[9]
port 392 nsew signal input
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 393 nsew signal input
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 394 nsew signal input
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 395 nsew signal input
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 396 nsew signal input
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 397 nsew signal input
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 398 nsew signal input
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 399 nsew signal input
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 400 nsew signal output
rlabel metal2 s 396333 995407 396389 995887 6 mprj_analog_io[11]
port 401 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 402 nsew signal bidirectional
rlabel metal2 s 393941 995407 393997 995887 6 mprj_io_analog_en[18]
port 403 nsew signal input
rlabel metal2 s 392653 995407 392709 995887 6 mprj_io_analog_pol[18]
port 404 nsew signal input
rlabel metal2 s 389617 995407 389673 995887 6 mprj_io_analog_sel[18]
port 405 nsew signal input
rlabel metal2 s 393297 995407 393353 995887 6 mprj_io_dm[54]
port 406 nsew signal input
rlabel metal2 s 395137 995407 395193 995887 6 mprj_io_dm[55]
port 407 nsew signal input
rlabel metal2 s 388973 995407 389029 995887 6 mprj_io_dm[56]
port 408 nsew signal input
rlabel metal2 s 390813 995407 390869 995887 6 mprj_io_enh[18]
port 409 nsew signal input
rlabel metal2 s 390169 995407 390225 995887 6 mprj_io_hldh_n[18]
port 410 nsew signal input
rlabel metal2 s 388329 995407 388385 995887 6 mprj_io_holdover[18]
port 411 nsew signal input
rlabel metal2 s 385293 995407 385349 995887 6 mprj_io_ib_mode_sel[18]
port 412 nsew signal input
rlabel metal2 s 392101 995407 392157 995887 6 mprj_io_inp_dis[18]
port 413 nsew signal input
rlabel metal2 s 384649 995407 384705 995887 6 mprj_io_oeb[18]
port 414 nsew signal input
rlabel metal2 s 387777 995407 387833 995887 6 mprj_io_out[18]
port 415 nsew signal input
rlabel metal2 s 396977 995407 397033 995887 6 mprj_io_slow_sel[18]
port 416 nsew signal input
rlabel metal2 s 385937 995407 385993 995887 6 mprj_io_vtrip_sel[18]
port 417 nsew signal input
rlabel metal2 s 398817 995407 398873 995887 6 mprj_io_in[18]
port 418 nsew signal output
rlabel metal2 s 41713 667333 42193 667389 6 mprj_analog_io[21]
port 419 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 420 nsew signal bidirectional
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[28]
port 421 nsew signal input
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[28]
port 422 nsew signal input
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[28]
port 423 nsew signal input
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[84]
port 424 nsew signal input
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[85]
port 425 nsew signal input
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[86]
port 426 nsew signal input
rlabel metal2 s 41713 661813 42193 661869 6 mprj_io_enh[28]
port 427 nsew signal input
rlabel metal2 s 41713 661169 42193 661225 6 mprj_io_hldh_n[28]
port 428 nsew signal input
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[28]
port 429 nsew signal input
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[28]
port 430 nsew signal input
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[28]
port 431 nsew signal input
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[28]
port 432 nsew signal input
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[28]
port 433 nsew signal input
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[28]
port 434 nsew signal input
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[28]
port 435 nsew signal input
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[28]
port 436 nsew signal output
rlabel metal2 s 41713 624133 42193 624189 6 mprj_analog_io[22]
port 437 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 438 nsew signal bidirectional
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[29]
port 439 nsew signal input
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[29]
port 440 nsew signal input
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[29]
port 441 nsew signal input
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[87]
port 442 nsew signal input
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[88]
port 443 nsew signal input
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[89]
port 444 nsew signal input
rlabel metal2 s 41713 618613 42193 618669 6 mprj_io_enh[29]
port 445 nsew signal input
rlabel metal2 s 41713 617969 42193 618025 6 mprj_io_hldh_n[29]
port 446 nsew signal input
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[29]
port 447 nsew signal input
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[29]
port 448 nsew signal input
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[29]
port 449 nsew signal input
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[29]
port 450 nsew signal input
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[29]
port 451 nsew signal input
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[29]
port 452 nsew signal input
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[29]
port 453 nsew signal input
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[29]
port 454 nsew signal output
rlabel metal2 s 41713 580933 42193 580989 6 mprj_analog_io[23]
port 455 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 456 nsew signal bidirectional
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[30]
port 457 nsew signal input
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[30]
port 458 nsew signal input
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[30]
port 459 nsew signal input
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[90]
port 460 nsew signal input
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[91]
port 461 nsew signal input
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[92]
port 462 nsew signal input
rlabel metal2 s 41713 575413 42193 575469 6 mprj_io_enh[30]
port 463 nsew signal input
rlabel metal2 s 41713 574769 42193 574825 6 mprj_io_hldh_n[30]
port 464 nsew signal input
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[30]
port 465 nsew signal input
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[30]
port 466 nsew signal input
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[30]
port 467 nsew signal input
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[30]
port 468 nsew signal input
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[30]
port 469 nsew signal input
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[30]
port 470 nsew signal input
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[30]
port 471 nsew signal input
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[30]
port 472 nsew signal output
rlabel metal2 s 41713 537733 42193 537789 6 mprj_analog_io[24]
port 473 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 474 nsew signal bidirectional
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[31]
port 475 nsew signal input
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[31]
port 476 nsew signal input
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[31]
port 477 nsew signal input
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[93]
port 478 nsew signal input
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[94]
port 479 nsew signal input
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[95]
port 480 nsew signal input
rlabel metal2 s 41713 532213 42193 532269 6 mprj_io_enh[31]
port 481 nsew signal input
rlabel metal2 s 41713 531569 42193 531625 6 mprj_io_hldh_n[31]
port 482 nsew signal input
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[31]
port 483 nsew signal input
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[31]
port 484 nsew signal input
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[31]
port 485 nsew signal input
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[31]
port 486 nsew signal input
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[31]
port 487 nsew signal input
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[31]
port 488 nsew signal input
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[31]
port 489 nsew signal input
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[31]
port 490 nsew signal output
rlabel metal2 s 41713 410133 42193 410189 6 mprj_analog_io[25]
port 491 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 492 nsew signal bidirectional
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[32]
port 493 nsew signal input
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[32]
port 494 nsew signal input
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[32]
port 495 nsew signal input
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[96]
port 496 nsew signal input
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[97]
port 497 nsew signal input
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[98]
port 498 nsew signal input
rlabel metal2 s 41713 404613 42193 404669 6 mprj_io_enh[32]
port 499 nsew signal input
rlabel metal2 s 41713 403969 42193 404025 6 mprj_io_hldh_n[32]
port 500 nsew signal input
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[32]
port 501 nsew signal input
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[32]
port 502 nsew signal input
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[32]
port 503 nsew signal input
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[32]
port 504 nsew signal input
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[32]
port 505 nsew signal input
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[32]
port 506 nsew signal input
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[32]
port 507 nsew signal input
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[32]
port 508 nsew signal output
rlabel metal2 s 41713 366933 42193 366989 6 mprj_analog_io[26]
port 509 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 510 nsew signal bidirectional
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[33]
port 511 nsew signal input
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[33]
port 512 nsew signal input
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[33]
port 513 nsew signal input
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[100]
port 514 nsew signal input
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[101]
port 515 nsew signal input
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[99]
port 516 nsew signal input
rlabel metal2 s 41713 361413 42193 361469 6 mprj_io_enh[33]
port 517 nsew signal input
rlabel metal2 s 41713 360769 42193 360825 6 mprj_io_hldh_n[33]
port 518 nsew signal input
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[33]
port 519 nsew signal input
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[33]
port 520 nsew signal input
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[33]
port 521 nsew signal input
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[33]
port 522 nsew signal input
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[33]
port 523 nsew signal input
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[33]
port 524 nsew signal input
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[33]
port 525 nsew signal input
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[33]
port 526 nsew signal output
rlabel metal2 s 41713 323733 42193 323789 6 mprj_analog_io[27]
port 527 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 528 nsew signal bidirectional
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[34]
port 529 nsew signal input
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[34]
port 530 nsew signal input
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[34]
port 531 nsew signal input
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[102]
port 532 nsew signal input
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[103]
port 533 nsew signal input
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[104]
port 534 nsew signal input
rlabel metal2 s 41713 318213 42193 318269 6 mprj_io_enh[34]
port 535 nsew signal input
rlabel metal2 s 41713 317569 42193 317625 6 mprj_io_hldh_n[34]
port 536 nsew signal input
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[34]
port 537 nsew signal input
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[34]
port 538 nsew signal input
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[34]
port 539 nsew signal input
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[34]
port 540 nsew signal input
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[34]
port 541 nsew signal input
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[34]
port 542 nsew signal input
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[34]
port 543 nsew signal input
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[34]
port 544 nsew signal output
rlabel metal2 s 41713 280533 42193 280589 6 mprj_analog_io[28]
port 545 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 546 nsew signal bidirectional
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[35]
port 547 nsew signal input
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[35]
port 548 nsew signal input
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[35]
port 549 nsew signal input
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[105]
port 550 nsew signal input
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[106]
port 551 nsew signal input
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[107]
port 552 nsew signal input
rlabel metal2 s 41713 275013 42193 275069 6 mprj_io_enh[35]
port 553 nsew signal input
rlabel metal2 s 41713 274369 42193 274425 6 mprj_io_hldh_n[35]
port 554 nsew signal input
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[35]
port 555 nsew signal input
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[35]
port 556 nsew signal input
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[35]
port 557 nsew signal input
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[35]
port 558 nsew signal input
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[35]
port 559 nsew signal input
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[35]
port 560 nsew signal input
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[35]
port 561 nsew signal input
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[35]
port 562 nsew signal output
rlabel metal2 s 41713 237333 42193 237389 6 mprj_analog_io[29]
port 563 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 564 nsew signal bidirectional
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[36]
port 565 nsew signal input
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[36]
port 566 nsew signal input
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[36]
port 567 nsew signal input
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[108]
port 568 nsew signal input
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[109]
port 569 nsew signal input
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[110]
port 570 nsew signal input
rlabel metal2 s 41713 231813 42193 231869 6 mprj_io_enh[36]
port 571 nsew signal input
rlabel metal2 s 41713 231169 42193 231225 6 mprj_io_hldh_n[36]
port 572 nsew signal input
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[36]
port 573 nsew signal input
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[36]
port 574 nsew signal input
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[36]
port 575 nsew signal input
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[36]
port 576 nsew signal input
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[36]
port 577 nsew signal input
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[36]
port 578 nsew signal input
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[36]
port 579 nsew signal input
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[36]
port 580 nsew signal output
rlabel metal2 s 41713 194133 42193 194189 6 mprj_analog_io[30]
port 581 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 582 nsew signal bidirectional
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[37]
port 583 nsew signal input
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[37]
port 584 nsew signal input
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[37]
port 585 nsew signal input
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[111]
port 586 nsew signal input
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[112]
port 587 nsew signal input
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[113]
port 588 nsew signal input
rlabel metal2 s 41713 188613 42193 188669 6 mprj_io_enh[37]
port 589 nsew signal input
rlabel metal2 s 41713 187969 42193 188025 6 mprj_io_hldh_n[37]
port 590 nsew signal input
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[37]
port 591 nsew signal input
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[37]
port 592 nsew signal input
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[37]
port 593 nsew signal input
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[37]
port 594 nsew signal input
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[37]
port 595 nsew signal input
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[37]
port 596 nsew signal input
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[37]
port 597 nsew signal input
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[37]
port 598 nsew signal output
rlabel metal2 s 294533 995407 294589 995887 6 mprj_analog_io[12]
port 599 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 600 nsew signal bidirectional
rlabel metal2 s 292141 995407 292197 995887 6 mprj_io_analog_en[19]
port 601 nsew signal input
rlabel metal2 s 290853 995407 290909 995887 6 mprj_io_analog_pol[19]
port 602 nsew signal input
rlabel metal2 s 287817 995407 287873 995887 6 mprj_io_analog_sel[19]
port 603 nsew signal input
rlabel metal2 s 291497 995407 291553 995887 6 mprj_io_dm[57]
port 604 nsew signal input
rlabel metal2 s 293337 995407 293393 995887 6 mprj_io_dm[58]
port 605 nsew signal input
rlabel metal2 s 287173 995407 287229 995887 6 mprj_io_dm[59]
port 606 nsew signal input
rlabel metal2 s 289013 995407 289069 995887 6 mprj_io_enh[19]
port 607 nsew signal input
rlabel metal2 s 288369 995407 288425 995887 6 mprj_io_hldh_n[19]
port 608 nsew signal input
rlabel metal2 s 286529 995407 286585 995887 6 mprj_io_holdover[19]
port 609 nsew signal input
rlabel metal2 s 283493 995407 283549 995887 6 mprj_io_ib_mode_sel[19]
port 610 nsew signal input
rlabel metal2 s 290301 995407 290357 995887 6 mprj_io_inp_dis[19]
port 611 nsew signal input
rlabel metal2 s 282849 995407 282905 995887 6 mprj_io_oeb[19]
port 612 nsew signal input
rlabel metal2 s 285977 995407 286033 995887 6 mprj_io_out[19]
port 613 nsew signal input
rlabel metal2 s 295177 995407 295233 995887 6 mprj_io_slow_sel[19]
port 614 nsew signal input
rlabel metal2 s 284137 995407 284193 995887 6 mprj_io_vtrip_sel[19]
port 615 nsew signal input
rlabel metal2 s 297017 995407 297073 995887 6 mprj_io_in[19]
port 616 nsew signal output
rlabel metal2 s 242933 995407 242989 995887 6 mprj_analog_io[13]
port 617 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 618 nsew signal bidirectional
rlabel metal2 s 240541 995407 240597 995887 6 mprj_io_analog_en[20]
port 619 nsew signal input
rlabel metal2 s 239253 995407 239309 995887 6 mprj_io_analog_pol[20]
port 620 nsew signal input
rlabel metal2 s 236217 995407 236273 995887 6 mprj_io_analog_sel[20]
port 621 nsew signal input
rlabel metal2 s 239897 995407 239953 995887 6 mprj_io_dm[60]
port 622 nsew signal input
rlabel metal2 s 241737 995407 241793 995887 6 mprj_io_dm[61]
port 623 nsew signal input
rlabel metal2 s 235573 995407 235629 995887 6 mprj_io_dm[62]
port 624 nsew signal input
rlabel metal2 s 237413 995407 237469 995887 6 mprj_io_enh[20]
port 625 nsew signal input
rlabel metal2 s 236769 995407 236825 995887 6 mprj_io_hldh_n[20]
port 626 nsew signal input
rlabel metal2 s 234929 995407 234985 995887 6 mprj_io_holdover[20]
port 627 nsew signal input
rlabel metal2 s 231893 995407 231949 995887 6 mprj_io_ib_mode_sel[20]
port 628 nsew signal input
rlabel metal2 s 238701 995407 238757 995887 6 mprj_io_inp_dis[20]
port 629 nsew signal input
rlabel metal2 s 231249 995407 231305 995887 6 mprj_io_oeb[20]
port 630 nsew signal input
rlabel metal2 s 234377 995407 234433 995887 6 mprj_io_out[20]
port 631 nsew signal input
rlabel metal2 s 243577 995407 243633 995887 6 mprj_io_slow_sel[20]
port 632 nsew signal input
rlabel metal2 s 232537 995407 232593 995887 6 mprj_io_vtrip_sel[20]
port 633 nsew signal input
rlabel metal2 s 245417 995407 245473 995887 6 mprj_io_in[20]
port 634 nsew signal output
rlabel metal2 s 191533 995407 191589 995887 6 mprj_analog_io[14]
port 635 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 636 nsew signal bidirectional
rlabel metal2 s 189141 995407 189197 995887 6 mprj_io_analog_en[21]
port 637 nsew signal input
rlabel metal2 s 187853 995407 187909 995887 6 mprj_io_analog_pol[21]
port 638 nsew signal input
rlabel metal2 s 184817 995407 184873 995887 6 mprj_io_analog_sel[21]
port 639 nsew signal input
rlabel metal2 s 188497 995407 188553 995887 6 mprj_io_dm[63]
port 640 nsew signal input
rlabel metal2 s 190337 995407 190393 995887 6 mprj_io_dm[64]
port 641 nsew signal input
rlabel metal2 s 184173 995407 184229 995887 6 mprj_io_dm[65]
port 642 nsew signal input
rlabel metal2 s 186013 995407 186069 995887 6 mprj_io_enh[21]
port 643 nsew signal input
rlabel metal2 s 185369 995407 185425 995887 6 mprj_io_hldh_n[21]
port 644 nsew signal input
rlabel metal2 s 183529 995407 183585 995887 6 mprj_io_holdover[21]
port 645 nsew signal input
rlabel metal2 s 180493 995407 180549 995887 6 mprj_io_ib_mode_sel[21]
port 646 nsew signal input
rlabel metal2 s 187301 995407 187357 995887 6 mprj_io_inp_dis[21]
port 647 nsew signal input
rlabel metal2 s 179849 995407 179905 995887 6 mprj_io_oeb[21]
port 648 nsew signal input
rlabel metal2 s 182977 995407 183033 995887 6 mprj_io_out[21]
port 649 nsew signal input
rlabel metal2 s 192177 995407 192233 995887 6 mprj_io_slow_sel[21]
port 650 nsew signal input
rlabel metal2 s 181137 995407 181193 995887 6 mprj_io_vtrip_sel[21]
port 651 nsew signal input
rlabel metal2 s 194017 995407 194073 995887 6 mprj_io_in[21]
port 652 nsew signal output
rlabel metal2 s 140133 995407 140189 995887 6 mprj_analog_io[15]
port 653 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 654 nsew signal bidirectional
rlabel metal2 s 137741 995407 137797 995887 6 mprj_io_analog_en[22]
port 655 nsew signal input
rlabel metal2 s 136453 995407 136509 995887 6 mprj_io_analog_pol[22]
port 656 nsew signal input
rlabel metal2 s 133417 995407 133473 995887 6 mprj_io_analog_sel[22]
port 657 nsew signal input
rlabel metal2 s 137097 995407 137153 995887 6 mprj_io_dm[66]
port 658 nsew signal input
rlabel metal2 s 138937 995407 138993 995887 6 mprj_io_dm[67]
port 659 nsew signal input
rlabel metal2 s 132773 995407 132829 995887 6 mprj_io_dm[68]
port 660 nsew signal input
rlabel metal2 s 134613 995407 134669 995887 6 mprj_io_enh[22]
port 661 nsew signal input
rlabel metal2 s 133969 995407 134025 995887 6 mprj_io_hldh_n[22]
port 662 nsew signal input
rlabel metal2 s 132129 995407 132185 995887 6 mprj_io_holdover[22]
port 663 nsew signal input
rlabel metal2 s 129093 995407 129149 995887 6 mprj_io_ib_mode_sel[22]
port 664 nsew signal input
rlabel metal2 s 135901 995407 135957 995887 6 mprj_io_inp_dis[22]
port 665 nsew signal input
rlabel metal2 s 128449 995407 128505 995887 6 mprj_io_oeb[22]
port 666 nsew signal input
rlabel metal2 s 131577 995407 131633 995887 6 mprj_io_out[22]
port 667 nsew signal input
rlabel metal2 s 140777 995407 140833 995887 6 mprj_io_slow_sel[22]
port 668 nsew signal input
rlabel metal2 s 129737 995407 129793 995887 6 mprj_io_vtrip_sel[22]
port 669 nsew signal input
rlabel metal2 s 142617 995407 142673 995887 6 mprj_io_in[22]
port 670 nsew signal output
rlabel metal2 s 88733 995407 88789 995887 6 mprj_analog_io[16]
port 671 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 672 nsew signal bidirectional
rlabel metal2 s 86341 995407 86397 995887 6 mprj_io_analog_en[23]
port 673 nsew signal input
rlabel metal2 s 85053 995407 85109 995887 6 mprj_io_analog_pol[23]
port 674 nsew signal input
rlabel metal2 s 82017 995407 82073 995887 6 mprj_io_analog_sel[23]
port 675 nsew signal input
rlabel metal2 s 85697 995407 85753 995887 6 mprj_io_dm[69]
port 676 nsew signal input
rlabel metal2 s 87537 995407 87593 995887 6 mprj_io_dm[70]
port 677 nsew signal input
rlabel metal2 s 81373 995407 81429 995887 6 mprj_io_dm[71]
port 678 nsew signal input
rlabel metal2 s 83213 995407 83269 995887 6 mprj_io_enh[23]
port 679 nsew signal input
rlabel metal2 s 82569 995407 82625 995887 6 mprj_io_hldh_n[23]
port 680 nsew signal input
rlabel metal2 s 80729 995407 80785 995887 6 mprj_io_holdover[23]
port 681 nsew signal input
rlabel metal2 s 77693 995407 77749 995887 6 mprj_io_ib_mode_sel[23]
port 682 nsew signal input
rlabel metal2 s 84501 995407 84557 995887 6 mprj_io_inp_dis[23]
port 683 nsew signal input
rlabel metal2 s 77049 995407 77105 995887 6 mprj_io_oeb[23]
port 684 nsew signal input
rlabel metal2 s 80177 995407 80233 995887 6 mprj_io_out[23]
port 685 nsew signal input
rlabel metal2 s 89377 995407 89433 995887 6 mprj_io_slow_sel[23]
port 686 nsew signal input
rlabel metal2 s 78337 995407 78393 995887 6 mprj_io_vtrip_sel[23]
port 687 nsew signal input
rlabel metal2 s 91217 995407 91273 995887 6 mprj_io_in[23]
port 688 nsew signal output
rlabel metal2 s 41713 966733 42193 966789 6 mprj_analog_io[17]
port 689 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 690 nsew signal bidirectional
rlabel metal2 s 41713 964341 42193 964397 6 mprj_io_analog_en[24]
port 691 nsew signal input
rlabel metal2 s 41713 963053 42193 963109 6 mprj_io_analog_pol[24]
port 692 nsew signal input
rlabel metal2 s 41713 960017 42193 960073 6 mprj_io_analog_sel[24]
port 693 nsew signal input
rlabel metal2 s 41713 963697 42193 963753 6 mprj_io_dm[72]
port 694 nsew signal input
rlabel metal2 s 41713 965537 42193 965593 6 mprj_io_dm[73]
port 695 nsew signal input
rlabel metal2 s 41713 959373 42193 959429 6 mprj_io_dm[74]
port 696 nsew signal input
rlabel metal2 s 41713 961213 42193 961269 6 mprj_io_enh[24]
port 697 nsew signal input
rlabel metal2 s 41713 960569 42193 960625 6 mprj_io_hldh_n[24]
port 698 nsew signal input
rlabel metal2 s 41713 958729 42193 958785 6 mprj_io_holdover[24]
port 699 nsew signal input
rlabel metal2 s 41713 955693 42193 955749 6 mprj_io_ib_mode_sel[24]
port 700 nsew signal input
rlabel metal2 s 41713 962501 42193 962557 6 mprj_io_inp_dis[24]
port 701 nsew signal input
rlabel metal2 s 41713 955049 42193 955105 6 mprj_io_oeb[24]
port 702 nsew signal input
rlabel metal2 s 41713 958177 42193 958233 6 mprj_io_out[24]
port 703 nsew signal input
rlabel metal2 s 41713 967377 42193 967433 6 mprj_io_slow_sel[24]
port 704 nsew signal input
rlabel metal2 s 41713 956337 42193 956393 6 mprj_io_vtrip_sel[24]
port 705 nsew signal input
rlabel metal2 s 41713 969217 42193 969273 6 mprj_io_in[24]
port 706 nsew signal output
rlabel metal2 s 41713 796933 42193 796989 6 mprj_analog_io[18]
port 707 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 708 nsew signal bidirectional
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[25]
port 709 nsew signal input
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[25]
port 710 nsew signal input
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[25]
port 711 nsew signal input
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[75]
port 712 nsew signal input
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[76]
port 713 nsew signal input
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[77]
port 714 nsew signal input
rlabel metal2 s 41713 791413 42193 791469 6 mprj_io_enh[25]
port 715 nsew signal input
rlabel metal2 s 41713 790769 42193 790825 6 mprj_io_hldh_n[25]
port 716 nsew signal input
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[25]
port 717 nsew signal input
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[25]
port 718 nsew signal input
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[25]
port 719 nsew signal input
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[25]
port 720 nsew signal input
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[25]
port 721 nsew signal input
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[25]
port 722 nsew signal input
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[25]
port 723 nsew signal input
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[25]
port 724 nsew signal output
rlabel metal2 s 41713 753733 42193 753789 6 mprj_analog_io[19]
port 725 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 726 nsew signal bidirectional
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[26]
port 727 nsew signal input
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[26]
port 728 nsew signal input
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[26]
port 729 nsew signal input
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[78]
port 730 nsew signal input
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[79]
port 731 nsew signal input
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[80]
port 732 nsew signal input
rlabel metal2 s 41713 748213 42193 748269 6 mprj_io_enh[26]
port 733 nsew signal input
rlabel metal2 s 41713 747569 42193 747625 6 mprj_io_hldh_n[26]
port 734 nsew signal input
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[26]
port 735 nsew signal input
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[26]
port 736 nsew signal input
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[26]
port 737 nsew signal input
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[26]
port 738 nsew signal input
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[26]
port 739 nsew signal input
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[26]
port 740 nsew signal input
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[26]
port 741 nsew signal input
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[26]
port 742 nsew signal output
rlabel metal2 s 41713 710533 42193 710589 6 mprj_analog_io[20]
port 743 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 744 nsew signal bidirectional
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[27]
port 745 nsew signal input
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[27]
port 746 nsew signal input
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[27]
port 747 nsew signal input
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[81]
port 748 nsew signal input
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[82]
port 749 nsew signal input
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[83]
port 750 nsew signal input
rlabel metal2 s 41713 705013 42193 705069 6 mprj_io_enh[27]
port 751 nsew signal input
rlabel metal2 s 41713 704369 42193 704425 6 mprj_io_hldh_n[27]
port 752 nsew signal input
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[27]
port 753 nsew signal input
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[27]
port 754 nsew signal input
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[27]
port 755 nsew signal input
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[27]
port 756 nsew signal input
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[27]
port 757 nsew signal input
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[27]
port 758 nsew signal input
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[27]
port 759 nsew signal input
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[27]
port 760 nsew signal output
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 761 nsew signal input
rlabel metal2 s 145103 40000 145131 40174 6 porb_h
port 761 nsew signal input
rlabel metal2 s 145103 40174 145144 40202 6 porb_h
port 761 nsew signal input
rlabel metal2 s 527455 41713 527511 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 523131 41713 523187 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 472655 41713 472711 41806 6 porb_h
port 761 nsew signal input
rlabel metal2 s 468331 41713 468387 41806 6 porb_h
port 761 nsew signal input
rlabel metal2 s 472636 41806 472711 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 468312 41806 468387 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 417855 41713 417911 41820 6 porb_h
port 761 nsew signal input
rlabel metal2 s 413531 41713 413587 41820 6 porb_h
port 761 nsew signal input
rlabel metal2 s 527468 42193 527496 44134 6 porb_h
port 761 nsew signal input
rlabel metal2 s 523144 42193 523172 44134 6 porb_h
port 761 nsew signal input
rlabel metal2 s 527456 44134 527508 44198 6 porb_h
port 761 nsew signal input
rlabel metal2 s 523132 44134 523184 44198 6 porb_h
port 761 nsew signal input
rlabel metal2 s 527468 44198 527496 45562 6 porb_h
port 761 nsew signal input
rlabel metal2 s 523144 44198 523172 44270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 472636 42193 472664 44270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 468312 42193 468340 44270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 417855 41820 417924 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 413531 41820 413600 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 363055 41713 363111 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 358731 41713 358787 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 308255 41713 308311 41806 6 porb_h
port 761 nsew signal input
rlabel metal2 s 303931 41713 303987 41806 6 porb_h
port 761 nsew signal input
rlabel metal2 s 308232 41806 308311 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 303908 41806 303987 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 199655 41713 199711 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 195331 41713 195387 42193 6 porb_h
port 761 nsew signal input
rlabel metal2 s 417896 42193 417924 44270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 413572 42193 413600 44270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 363064 42193 363092 44202 6 porb_h
port 761 nsew signal input
rlabel metal2 s 358740 42193 358768 44134 6 porb_h
port 761 nsew signal input
rlabel metal2 s 358728 44134 358780 44198 6 porb_h
port 761 nsew signal input
rlabel metal2 s 363052 44202 363104 44266 6 porb_h
port 761 nsew signal input
rlabel metal2 s 358740 44198 358768 44270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 308232 42193 308260 44202 6 porb_h
port 761 nsew signal input
rlabel metal2 s 303908 42193 303936 44202 6 porb_h
port 761 nsew signal input
rlabel metal2 s 199672 42193 199700 44202 6 porb_h
port 761 nsew signal input
rlabel metal2 s 308220 44202 308272 44266 6 porb_h
port 761 nsew signal input
rlabel metal2 s 303896 44202 303948 44266 6 porb_h
port 761 nsew signal input
rlabel metal2 s 199660 44202 199712 44266 6 porb_h
port 761 nsew signal input
rlabel metal2 s 523132 44270 523184 44334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 472624 44270 472676 44334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 468300 44270 468352 44334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 417884 44270 417936 44334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 413560 44270 413612 44334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 358728 44270 358780 44334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 199672 44266 199700 44338 6 porb_h
port 761 nsew signal input
rlabel metal2 s 195348 42193 195376 44338 6 porb_h
port 761 nsew signal input
rlabel metal2 s 145116 40202 145144 44338 6 porb_h
port 761 nsew signal input
rlabel metal2 s 199660 44338 199712 44402 6 porb_h
port 761 nsew signal input
rlabel metal2 s 195336 44338 195388 44402 6 porb_h
port 761 nsew signal input
rlabel metal2 s 145104 44338 145156 44402 6 porb_h
port 761 nsew signal input
rlabel metal2 s 143632 44338 143684 44402 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 45562 673604 45626 6 porb_h
port 761 nsew signal input
rlabel metal2 s 527456 45562 527508 45626 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 45626 673592 112746 6 porb_h
port 761 nsew signal input
rlabel metal2 s 143644 44402 143672 45630 6 porb_h
port 761 nsew signal input
rlabel metal2 s 143632 45630 143684 45694 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 45630 42484 45694 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 112746 675444 112810 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 112746 673604 112810 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 112810 675432 113255 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 113255 675887 113283 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 113283 675887 113311 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 112810 673592 158306 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 158306 675444 158370 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 158306 673604 158370 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 158370 675432 158455 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 158455 675887 158508 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 158508 675887 158511 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 158370 673592 203102 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42444 45694 42472 184826 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 184289 42193 184345 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 184345 41828 184826 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42616 184826 42668 184890 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 184826 42484 184890 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 184826 41840 184890 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 203102 673776 203130 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 203455 675887 203483 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 203483 675887 203511 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 203511 675432 203866 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673748 203130 673776 203866 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 203866 675444 203930 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673736 203866 673788 203930 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673748 203930 673776 212502 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 212502 673880 212566 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673736 212502 673788 212566 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673840 212566 673868 217942 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 217942 673880 218006 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 218078 673880 218142 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673840 218142 673868 243782 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42628 184890 42656 228006 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 227489 42193 227545 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 227545 41828 228006 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 228006 42852 228070 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42616 228006 42668 228070 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 228006 41840 228070 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675300 243782 675352 243846 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 243782 673880 243846 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 248655 675887 248662 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675312 243846 675340 248662 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42812 228070 42840 245482 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 245482 42852 245546 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 245482 42576 245546 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675312 248662 675887 248678 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675300 248678 675887 248690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 248690 675887 248711 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675300 248690 675352 248742 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673460 248678 673512 248742 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675312 248742 675340 248773 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673472 248742 673500 264930 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 264930 673696 264994 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673460 264930 673512 264994 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 264994 673684 293422 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42536 245546 42564 271186 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 270689 42193 270745 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 270745 41828 271186 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 271186 42852 271250 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 271186 42576 271250 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 271186 41840 271250 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675300 293422 675352 293486 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 293422 673696 293486 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 293655 675887 293678 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675312 293486 675340 293678 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675312 293678 675887 293706 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 293706 675887 293711 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675312 293706 675340 303554 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675300 303554 675352 303618 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 303554 673604 303618 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 303618 673592 338098 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42812 271250 42840 313398 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42812 313398 42932 313414 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 313414 42932 313426 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42904 313426 42932 322730 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 313426 42852 313478 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 313482 41840 313546 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 313546 41828 313889 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 313889 42193 313945 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42892 322730 42944 322794 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42616 322798 42668 322862 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 338098 675444 338162 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 338098 673604 338162 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 338162 675432 338655 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 338655 675887 338708 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 338708 675887 338711 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 338162 673592 380870 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42628 322862 42656 357614 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 357089 42193 357145 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 357145 41828 357614 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42616 357614 42668 357678 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 357614 42484 357678 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 357614 41840 357678 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673736 380870 673788 380934 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 380870 673604 380934 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 383855 675887 383860 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 383860 675887 383911 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 383911 675432 384270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673748 380934 673776 384270 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 384270 675444 384334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673736 384270 673788 384334 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673748 384334 673776 420838 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42444 357678 42472 400794 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 400289 42193 400345 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 400345 41828 400794 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 400794 42484 400858 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 400794 41840 400858 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673748 420838 673868 420866 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673840 420866 673868 449550 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 449550 673880 449614 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 449550 673604 449614 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 449614 673592 498170 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 498170 673880 498234 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 498170 673604 498234 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673840 498234 673868 546314 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42444 400858 42472 527478 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42708 527478 42760 527542 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 527478 42484 527542 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 527478 41840 527542 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 546314 673880 546378 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 546382 673604 546446 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 546446 673592 560526 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 560526 675444 560590 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 560526 673880 560590 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 560526 673604 560590 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 560590 675432 561055 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 561055 675887 561068 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 561068 675887 561111 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673840 560590 673868 585142 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42720 527542 42748 570658 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 527542 41828 527889 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 527889 42193 527945 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42708 570658 42760 570722 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 570658 42576 570722 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 570658 41840 570722 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 585142 673880 585206 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673552 585142 673604 585206 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 585206 673592 595054 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673564 595054 673684 595082 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 606255 675887 606283 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 606283 675887 606311 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 606311 675432 606698 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 595082 673684 606698 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 606698 675444 606762 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 606698 673696 606762 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 651255 675887 651283 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 651283 675887 651311 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 651311 675432 651714 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 606762 673684 651714 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42536 570722 42564 614790 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 570722 41828 571089 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 571089 42193 571145 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 614289 42193 614345 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 614345 41828 614790 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 614790 42576 614854 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 614790 41840 614854 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42536 614854 42564 631910 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42444 631910 42564 631938 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42444 631938 42472 651374 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 651374 42852 651438 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 651374 42484 651438 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 651714 675444 651778 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 651714 673696 651778 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 651778 673684 695846 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42812 651438 42840 658038 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 657489 42193 657545 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 657545 41828 658038 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 658038 42852 658102 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 658038 41840 658102 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42812 658102 42840 681566 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 681566 42852 681630 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 681634 42484 681698 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42444 681698 42472 695506 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42892 695506 42944 695570 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42432 695506 42484 695570 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 695846 673696 695910 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 695914 675444 695978 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 695978 675432 696455 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 696455 675887 696483 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 696483 675887 696511 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 695910 673684 701014 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42904 695570 42932 700810 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 700689 42193 700745 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 700745 41828 700810 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42892 700810 42944 700874 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 700810 41840 700874 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673828 701014 673880 701078 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 701014 673696 701078 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673840 701078 673868 720310 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 720310 673868 720338 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42904 700874 42932 720326 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 720338 673684 739638 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42892 720326 42944 720390 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 720326 42576 720390 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42536 720390 42564 734130 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42984 734130 43036 734194 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 734130 42576 734194 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 739638 673696 739702 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 739774 673696 739838 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 741455 675887 741483 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 741483 675887 741511 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 741511 675432 741882 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 741882 675444 741946 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673656 739838 673684 741950 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673920 741950 673972 742014 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673644 741950 673696 742014 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673932 742014 673960 753510 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42996 734194 43024 743990 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 743889 42193 743945 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 743945 41828 743990 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42984 743990 43036 744054 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 743990 42576 744054 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 743990 41840 744054 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42536 744054 42564 753442 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 753442 42852 753506 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 753442 42576 753506 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673920 753510 673972 753574 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673736 753510 673788 753574 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673748 753574 673776 772754 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42812 753506 42840 758950 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42800 758950 42852 759014 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 758950 42576 759014 6 porb_h
port 761 nsew signal input
rlabel metal2 s 674012 772754 674064 772818 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673736 772754 673788 772818 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 786455 675887 786483 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 786483 675887 786511 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 786511 675432 786558 6 porb_h
port 761 nsew signal input
rlabel metal2 s 674024 772818 674052 786558 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 786558 675444 786622 6 porb_h
port 761 nsew signal input
rlabel metal2 s 674012 786558 674064 786622 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673460 786558 673512 786622 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673472 786622 673500 875162 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42536 759014 42564 786626 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42524 786626 42576 786690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41788 786626 41840 786690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41800 786690 41828 787089 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 787089 42193 787145 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 875162 675444 875226 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673460 875162 673512 875226 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 875226 675432 875655 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 875655 675887 875683 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 875683 675887 875711 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675407 964855 675887 964883 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 964883 675887 964911 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675404 964911 675432 965262 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673472 875226 673500 965262 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 956889 42193 956903 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 956903 42288 956931 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42260 956931 42288 957510 6 porb_h
port 761 nsew signal input
rlabel metal2 s 41713 956931 42193 956945 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42248 957510 42300 957574 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42248 957714 42300 957778 6 porb_h
port 761 nsew signal input
rlabel metal2 s 675392 965262 675444 965326 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673460 965262 673512 965326 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673472 965326 673500 990014 6 porb_h
port 761 nsew signal input
rlabel metal2 s 673460 990014 673512 990078 6 porb_h
port 761 nsew signal input
rlabel metal2 s 628656 990082 628708 990146 6 porb_h
port 761 nsew signal input
rlabel metal2 s 626540 990082 626592 990146 6 porb_h
port 761 nsew signal input
rlabel metal2 s 628668 990146 628696 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 626552 990146 626580 990626 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42260 957778 42288 990150 6 porb_h
port 761 nsew signal input
rlabel metal2 s 78864 990150 78916 990214 6 porb_h
port 761 nsew signal input
rlabel metal2 s 42248 990150 42300 990214 6 porb_h
port 761 nsew signal input
rlabel metal2 s 286968 990558 287020 990622 6 porb_h
port 761 nsew signal input
rlabel metal2 s 626540 990626 626592 990690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 526904 990626 526956 990690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 475476 990626 475528 990690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 386512 990626 386564 990690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 526916 990690 526944 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 475488 990690 475516 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 628668 995407 628745 995466 6 porb_h
port 761 nsew signal input
rlabel metal2 s 628689 995466 628745 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 526889 995407 526945 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 475488 995407 475545 995452 6 porb_h
port 761 nsew signal input
rlabel metal2 s 386524 990690 386552 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 286980 990622 287008 990762 6 porb_h
port 761 nsew signal input
rlabel metal2 s 181720 990626 181772 990690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 130292 990626 130344 990690 6 porb_h
port 761 nsew signal input
rlabel metal2 s 286968 990762 287020 990826 6 porb_h
port 761 nsew signal input
rlabel metal2 s 284668 990762 284720 990826 6 porb_h
port 761 nsew signal input
rlabel metal2 s 233056 990762 233108 990826 6 porb_h
port 761 nsew signal input
rlabel metal2 s 284680 990826 284708 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 233068 990826 233096 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 386489 995407 386552 995452 6 porb_h
port 761 nsew signal input
rlabel metal2 s 475489 995452 475545 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 386489 995452 386545 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 284680 995407 284745 995452 6 porb_h
port 761 nsew signal input
rlabel metal2 s 284689 995452 284745 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 233068 995407 233145 995466 6 porb_h
port 761 nsew signal input
rlabel metal2 s 181732 990690 181760 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 130304 990690 130332 990762 6 porb_h
port 761 nsew signal input
rlabel metal2 s 78876 990214 78904 990762 6 porb_h
port 761 nsew signal input
rlabel metal2 s 130292 990762 130344 990826 6 porb_h
port 761 nsew signal input
rlabel metal2 s 78864 990762 78916 990826 6 porb_h
port 761 nsew signal input
rlabel metal2 s 130304 990826 130332 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 78876 990826 78904 995407 6 porb_h
port 761 nsew signal input
rlabel metal2 s 181689 995407 181760 995466 6 porb_h
port 761 nsew signal input
rlabel metal2 s 233089 995466 233145 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 181689 995466 181745 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 130289 995407 130345 995887 6 porb_h
port 761 nsew signal input
rlabel metal2 s 78876 995407 78945 995452 6 porb_h
port 761 nsew signal input
rlabel metal2 s 78889 995452 78945 995887 6 porb_h
port 761 nsew signal input
rlabel via1 s 527456 44140 527508 44192 6 porb_h
port 761 nsew signal input
rlabel via1 s 523132 44140 523184 44192 6 porb_h
port 761 nsew signal input
rlabel via1 s 358728 44140 358780 44192 6 porb_h
port 761 nsew signal input
rlabel via1 s 523132 44276 523184 44328 6 porb_h
port 761 nsew signal input
rlabel via1 s 472624 44276 472676 44328 6 porb_h
port 761 nsew signal input
rlabel via1 s 468300 44276 468352 44328 6 porb_h
port 761 nsew signal input
rlabel via1 s 417884 44276 417936 44328 6 porb_h
port 761 nsew signal input
rlabel via1 s 413560 44276 413612 44328 6 porb_h
port 761 nsew signal input
rlabel via1 s 363052 44208 363104 44260 6 porb_h
port 761 nsew signal input
rlabel via1 s 358728 44276 358780 44328 6 porb_h
port 761 nsew signal input
rlabel via1 s 308220 44208 308272 44260 6 porb_h
port 761 nsew signal input
rlabel via1 s 303896 44208 303948 44260 6 porb_h
port 761 nsew signal input
rlabel via1 s 199660 44208 199712 44260 6 porb_h
port 761 nsew signal input
rlabel via1 s 199660 44344 199712 44396 6 porb_h
port 761 nsew signal input
rlabel via1 s 195336 44344 195388 44396 6 porb_h
port 761 nsew signal input
rlabel via1 s 145104 44344 145156 44396 6 porb_h
port 761 nsew signal input
rlabel via1 s 143632 44344 143684 44396 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 45568 673604 45620 6 porb_h
port 761 nsew signal input
rlabel via1 s 527456 45568 527508 45620 6 porb_h
port 761 nsew signal input
rlabel via1 s 143632 45636 143684 45688 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 45636 42484 45688 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 112752 675444 112804 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 112752 673604 112804 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 158312 675444 158364 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 158312 673604 158364 6 porb_h
port 761 nsew signal input
rlabel via1 s 42616 184832 42668 184884 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 184832 42484 184884 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 184832 41840 184884 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 203872 675444 203924 6 porb_h
port 761 nsew signal input
rlabel via1 s 673736 203872 673788 203924 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 212508 673880 212560 6 porb_h
port 761 nsew signal input
rlabel via1 s 673736 212508 673788 212560 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 217948 673880 218000 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 218084 673880 218136 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 228012 42852 228064 6 porb_h
port 761 nsew signal input
rlabel via1 s 42616 228012 42668 228064 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 228012 41840 228064 6 porb_h
port 761 nsew signal input
rlabel via1 s 675300 243788 675352 243840 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 243788 673880 243840 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 245488 42852 245540 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 245488 42576 245540 6 porb_h
port 761 nsew signal input
rlabel via1 s 675300 248684 675352 248736 6 porb_h
port 761 nsew signal input
rlabel via1 s 673460 248684 673512 248736 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 264936 673696 264988 6 porb_h
port 761 nsew signal input
rlabel via1 s 673460 264936 673512 264988 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 271192 42852 271244 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 271192 42576 271244 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 271192 41840 271244 6 porb_h
port 761 nsew signal input
rlabel via1 s 675300 293428 675352 293480 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 293428 673696 293480 6 porb_h
port 761 nsew signal input
rlabel via1 s 675300 303560 675352 303612 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 303560 673604 303612 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 313420 42852 313472 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 313488 41840 313540 6 porb_h
port 761 nsew signal input
rlabel via1 s 42892 322736 42944 322788 6 porb_h
port 761 nsew signal input
rlabel via1 s 42616 322804 42668 322856 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 338104 675444 338156 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 338104 673604 338156 6 porb_h
port 761 nsew signal input
rlabel via1 s 42616 357620 42668 357672 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 357620 42484 357672 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 357620 41840 357672 6 porb_h
port 761 nsew signal input
rlabel via1 s 673736 380876 673788 380928 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 380876 673604 380928 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 384276 675444 384328 6 porb_h
port 761 nsew signal input
rlabel via1 s 673736 384276 673788 384328 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 400800 42484 400852 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 400800 41840 400852 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 449556 673880 449608 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 449556 673604 449608 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 498176 673880 498228 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 498176 673604 498228 6 porb_h
port 761 nsew signal input
rlabel via1 s 42708 527484 42760 527536 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 527484 42484 527536 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 527484 41840 527536 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 546320 673880 546372 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 546388 673604 546440 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 560532 675444 560584 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 560532 673880 560584 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 560532 673604 560584 6 porb_h
port 761 nsew signal input
rlabel via1 s 42708 570664 42760 570716 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 570664 42576 570716 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 570664 41840 570716 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 585148 673880 585200 6 porb_h
port 761 nsew signal input
rlabel via1 s 673552 585148 673604 585200 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 606704 675444 606756 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 606704 673696 606756 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 614796 42576 614848 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 614796 41840 614848 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 651380 42852 651432 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 651380 42484 651432 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 651720 675444 651772 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 651720 673696 651772 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 658044 42852 658096 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 658044 41840 658096 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 681572 42852 681624 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 681640 42484 681692 6 porb_h
port 761 nsew signal input
rlabel via1 s 42892 695512 42944 695564 6 porb_h
port 761 nsew signal input
rlabel via1 s 42432 695512 42484 695564 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 695852 673696 695904 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 695920 675444 695972 6 porb_h
port 761 nsew signal input
rlabel via1 s 42892 700816 42944 700868 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 700816 41840 700868 6 porb_h
port 761 nsew signal input
rlabel via1 s 673828 701020 673880 701072 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 701020 673696 701072 6 porb_h
port 761 nsew signal input
rlabel via1 s 42892 720332 42944 720384 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 720332 42576 720384 6 porb_h
port 761 nsew signal input
rlabel via1 s 42984 734136 43036 734188 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 734136 42576 734188 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 739644 673696 739696 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 739780 673696 739832 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 741888 675444 741940 6 porb_h
port 761 nsew signal input
rlabel via1 s 673920 741956 673972 742008 6 porb_h
port 761 nsew signal input
rlabel via1 s 673644 741956 673696 742008 6 porb_h
port 761 nsew signal input
rlabel via1 s 42984 743996 43036 744048 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 743996 42576 744048 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 743996 41840 744048 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 753448 42852 753500 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 753448 42576 753500 6 porb_h
port 761 nsew signal input
rlabel via1 s 673920 753516 673972 753568 6 porb_h
port 761 nsew signal input
rlabel via1 s 673736 753516 673788 753568 6 porb_h
port 761 nsew signal input
rlabel via1 s 42800 758956 42852 759008 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 758956 42576 759008 6 porb_h
port 761 nsew signal input
rlabel via1 s 674012 772760 674064 772812 6 porb_h
port 761 nsew signal input
rlabel via1 s 673736 772760 673788 772812 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 786564 675444 786616 6 porb_h
port 761 nsew signal input
rlabel via1 s 674012 786564 674064 786616 6 porb_h
port 761 nsew signal input
rlabel via1 s 673460 786564 673512 786616 6 porb_h
port 761 nsew signal input
rlabel via1 s 42524 786632 42576 786684 6 porb_h
port 761 nsew signal input
rlabel via1 s 41788 786632 41840 786684 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 875168 675444 875220 6 porb_h
port 761 nsew signal input
rlabel via1 s 673460 875168 673512 875220 6 porb_h
port 761 nsew signal input
rlabel via1 s 42248 957516 42300 957568 6 porb_h
port 761 nsew signal input
rlabel via1 s 42248 957720 42300 957772 6 porb_h
port 761 nsew signal input
rlabel via1 s 675392 965268 675444 965320 6 porb_h
port 761 nsew signal input
rlabel via1 s 673460 965268 673512 965320 6 porb_h
port 761 nsew signal input
rlabel via1 s 673460 990020 673512 990072 6 porb_h
port 761 nsew signal input
rlabel via1 s 628656 990088 628708 990140 6 porb_h
port 761 nsew signal input
rlabel via1 s 626540 990088 626592 990140 6 porb_h
port 761 nsew signal input
rlabel via1 s 78864 990156 78916 990208 6 porb_h
port 761 nsew signal input
rlabel via1 s 42248 990156 42300 990208 6 porb_h
port 761 nsew signal input
rlabel via1 s 286968 990564 287020 990616 6 porb_h
port 761 nsew signal input
rlabel via1 s 626540 990632 626592 990684 6 porb_h
port 761 nsew signal input
rlabel via1 s 526904 990632 526956 990684 6 porb_h
port 761 nsew signal input
rlabel via1 s 475476 990632 475528 990684 6 porb_h
port 761 nsew signal input
rlabel via1 s 386512 990632 386564 990684 6 porb_h
port 761 nsew signal input
rlabel via1 s 286968 990768 287020 990820 6 porb_h
port 761 nsew signal input
rlabel via1 s 284668 990768 284720 990820 6 porb_h
port 761 nsew signal input
rlabel via1 s 233056 990768 233108 990820 6 porb_h
port 761 nsew signal input
rlabel via1 s 181720 990632 181772 990684 6 porb_h
port 761 nsew signal input
rlabel via1 s 130292 990632 130344 990684 6 porb_h
port 761 nsew signal input
rlabel via1 s 130292 990768 130344 990820 6 porb_h
port 761 nsew signal input
rlabel via1 s 78864 990768 78916 990820 6 porb_h
port 761 nsew signal input
rlabel metal1 s 527450 44140 527514 44152 6 porb_h
port 761 nsew signal input
rlabel metal1 s 523126 44140 523190 44152 6 porb_h
port 761 nsew signal input
rlabel metal1 s 358722 44140 358786 44152 6 porb_h
port 761 nsew signal input
rlabel metal1 s 523126 44152 527514 44180 6 porb_h
port 761 nsew signal input
rlabel metal1 s 527450 44180 527514 44192 6 porb_h
port 761 nsew signal input
rlabel metal1 s 523126 44180 523190 44192 6 porb_h
port 761 nsew signal input
rlabel metal1 s 358722 44152 363092 44180 6 porb_h
port 761 nsew signal input
rlabel metal1 s 363064 44180 363092 44208 6 porb_h
port 761 nsew signal input
rlabel metal1 s 358722 44180 358786 44192 6 porb_h
port 761 nsew signal input
rlabel metal1 s 363046 44208 363110 44220 6 porb_h
port 761 nsew signal input
rlabel metal1 s 308214 44208 308278 44220 6 porb_h
port 761 nsew signal input
rlabel metal1 s 303890 44208 303954 44220 6 porb_h
port 761 nsew signal input
rlabel metal1 s 199654 44208 199718 44220 6 porb_h
port 761 nsew signal input
rlabel metal1 s 363046 44220 399800 44248 6 porb_h
port 761 nsew signal input
rlabel metal1 s 523126 44276 523190 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 472618 44276 472682 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 468294 44276 468358 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 417878 44276 417942 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 413554 44276 413618 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 399772 44248 399800 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 363046 44248 363110 44260 6 porb_h
port 761 nsew signal input
rlabel metal1 s 199654 44220 355548 44248 6 porb_h
port 761 nsew signal input
rlabel metal1 s 399772 44288 523190 44316 6 porb_h
port 761 nsew signal input
rlabel metal1 s 358722 44276 358786 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 355520 44248 355548 44288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 308214 44248 308278 44260 6 porb_h
port 761 nsew signal input
rlabel metal1 s 303890 44248 303954 44260 6 porb_h
port 761 nsew signal input
rlabel metal1 s 199654 44248 199718 44260 6 porb_h
port 761 nsew signal input
rlabel metal1 s 355520 44288 358786 44316 6 porb_h
port 761 nsew signal input
rlabel metal1 s 523126 44316 523190 44328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 472618 44316 472682 44328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 468294 44316 468358 44328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 417878 44316 417942 44328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 413554 44316 413618 44328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 358722 44316 358786 44328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 199654 44344 199718 44356 6 porb_h
port 761 nsew signal input
rlabel metal1 s 195330 44344 195394 44356 6 porb_h
port 761 nsew signal input
rlabel metal1 s 145098 44344 145162 44356 6 porb_h
port 761 nsew signal input
rlabel metal1 s 143626 44344 143690 44356 6 porb_h
port 761 nsew signal input
rlabel metal1 s 143626 44356 199718 44384 6 porb_h
port 761 nsew signal input
rlabel metal1 s 199654 44384 199718 44396 6 porb_h
port 761 nsew signal input
rlabel metal1 s 195330 44384 195394 44396 6 porb_h
port 761 nsew signal input
rlabel metal1 s 145098 44384 145162 44396 6 porb_h
port 761 nsew signal input
rlabel metal1 s 143626 44384 143690 44396 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 45568 673610 45580 6 porb_h
port 761 nsew signal input
rlabel metal1 s 527450 45568 527514 45580 6 porb_h
port 761 nsew signal input
rlabel metal1 s 527450 45580 673610 45608 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 45608 673610 45620 6 porb_h
port 761 nsew signal input
rlabel metal1 s 527450 45608 527514 45620 6 porb_h
port 761 nsew signal input
rlabel metal1 s 143626 45636 143690 45648 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 45636 42490 45648 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 45648 143690 45676 6 porb_h
port 761 nsew signal input
rlabel metal1 s 143626 45676 143690 45688 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 45676 42490 45688 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 112752 675450 112764 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 112752 673610 112764 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 112764 675450 112792 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 112792 675450 112804 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 112792 673610 112804 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 158312 675450 158324 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 158312 673610 158324 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 158324 675450 158352 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 158352 675450 158364 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 158352 673610 158364 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42610 184832 42674 184844 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 184832 42490 184844 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 184832 41846 184844 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 184844 42674 184872 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42610 184872 42674 184884 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 184872 42490 184884 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 184872 41846 184884 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 203872 675450 203884 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 203872 673794 203884 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 203884 675450 203912 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 203912 675450 203924 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 203912 673794 203924 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 212508 673886 212520 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 212508 673794 212520 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 212520 673886 212548 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 212548 673886 212560 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 212548 673794 212560 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 217948 673886 218000 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673840 218000 673868 218084 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 218084 673886 218136 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 228012 42858 228024 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42610 228012 42674 228024 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 228012 41846 228024 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 228024 42858 228052 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 228052 42858 228064 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42610 228052 42674 228064 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 228052 41846 228064 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 243788 675358 243800 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 243788 673886 243800 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 243800 675358 243828 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 243828 675358 243840 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 243828 673886 243840 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 245488 42858 245500 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 245488 42582 245500 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 245500 42858 245528 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 245528 42858 245540 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 245528 42582 245540 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 248684 675358 248696 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 248684 673518 248696 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 248696 675358 248724 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 248724 675358 248736 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 248724 673518 248736 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 264936 673702 264948 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 264936 673518 264948 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 264948 673702 264976 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 264976 673702 264988 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 264976 673518 264988 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 271192 42858 271204 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 271192 42582 271204 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 271192 41846 271204 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 271204 42858 271232 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 271232 42858 271244 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 271232 42582 271244 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 271232 41846 271244 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 293428 675358 293440 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 293428 673702 293440 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 293440 675358 293468 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 293468 675358 293480 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 293468 673702 293480 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 303560 675358 303572 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 303560 673610 303572 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 303572 675358 303600 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675294 303600 675358 303612 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 303600 673610 303612 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 313420 42858 313432 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41800 313432 42858 313460 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 313460 42858 313472 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41800 313460 41828 313488 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 313488 41846 313540 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 322736 42950 322748 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42628 322748 42950 322776 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 322776 42950 322788 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42628 322776 42656 322804 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42610 322804 42674 322856 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 338104 675450 338116 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 338104 673610 338116 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 338116 675450 338144 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 338144 675450 338156 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 338144 673610 338156 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42610 357620 42674 357632 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 357620 42490 357632 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 357620 41846 357632 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 357632 42674 357660 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42610 357660 42674 357672 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 357660 42490 357672 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 357660 41846 357672 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 380876 673794 380888 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 380876 673610 380888 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 380888 673794 380916 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 380916 673794 380928 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 380916 673610 380928 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 384276 675450 384288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 384276 673794 384288 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 384288 675450 384316 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 384316 675450 384328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 384316 673794 384328 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 400800 42490 400812 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 400800 41846 400812 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 400812 42490 400840 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 400840 42490 400852 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 400840 41846 400852 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 449556 673886 449568 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 449556 673610 449568 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 449568 673886 449596 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 449596 673886 449608 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 449596 673610 449608 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 498176 673886 498188 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 498176 673610 498188 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 498188 673886 498216 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 498216 673886 498228 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 498216 673610 498228 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42702 527484 42766 527496 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 527484 42490 527496 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 527484 41846 527496 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 527496 42766 527524 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42702 527524 42766 527536 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 527524 42490 527536 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 527524 41846 527536 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 546320 673886 546332 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673564 546332 673886 546360 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 546360 673886 546372 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673564 546360 673592 546388 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 546388 673610 546440 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 560532 675450 560544 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 560532 673886 560544 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 560532 673610 560544 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 560544 675450 560572 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 560572 675450 560584 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 560572 673886 560584 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 560572 673610 560584 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42702 570664 42766 570676 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 570664 42582 570676 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 570664 41846 570676 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 570676 42766 570704 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42702 570704 42766 570716 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 570704 42582 570716 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 570704 41846 570716 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 585148 673886 585160 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 585148 673610 585160 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 585160 673886 585188 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 585188 673886 585200 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673546 585188 673610 585200 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 606704 675450 606716 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 606704 673702 606716 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 606716 675450 606744 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 606744 675450 606756 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 606744 673702 606756 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 614796 42582 614808 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 614796 41846 614808 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 614808 42582 614836 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 614836 42582 614848 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 614836 41846 614848 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 651380 42858 651392 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 651380 42490 651392 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 651392 42858 651420 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 651420 42858 651432 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 651420 42490 651432 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 651720 675450 651732 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 651720 673702 651732 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 651732 675450 651760 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 651760 675450 651772 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 651760 673702 651772 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 658044 42858 658056 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 658044 41846 658056 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 658056 42858 658084 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 658084 42858 658096 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 658084 41846 658096 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 681572 42858 681584 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42444 681584 42858 681612 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 681612 42858 681624 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42444 681612 42472 681640 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 681640 42490 681692 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 695512 42950 695524 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 695512 42490 695524 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 695524 42950 695552 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 695552 42950 695564 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42426 695552 42490 695564 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 695852 673702 695864 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 695864 675432 695892 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675404 695892 675432 695920 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 695892 673702 695904 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 695920 675450 695972 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 700816 42950 700828 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 700816 41846 700828 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 700828 42950 700856 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 700856 42950 700868 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 700856 41846 700868 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 701020 673886 701032 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 701020 673702 701032 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 701032 673886 701060 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673822 701060 673886 701072 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 701060 673702 701072 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 720332 42950 720344 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 720332 42582 720344 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 720344 42950 720372 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42886 720372 42950 720384 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 720372 42582 720384 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42978 734136 43042 734148 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 734136 42582 734148 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 734148 43042 734176 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42978 734176 43042 734188 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 734176 42582 734188 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 739644 673702 739696 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673656 739696 673684 739780 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 739780 673702 739832 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 741888 675450 741940 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675404 741940 675432 741968 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673914 741956 673978 741968 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 741956 673702 741968 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 741968 675432 741996 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673914 741996 673978 742008 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673638 741996 673702 742008 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42978 743996 43042 744008 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 743996 42582 744008 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 743996 41846 744008 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 744008 43042 744036 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42978 744036 43042 744048 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 744036 42582 744048 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 744036 41846 744048 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 753448 42858 753460 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 753448 42582 753460 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 753460 42858 753488 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 753488 42858 753500 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 753488 42582 753500 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673914 753516 673978 753528 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 753516 673794 753528 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 753528 673978 753556 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673914 753556 673978 753568 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 753556 673794 753568 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 758956 42858 758968 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 758956 42582 758968 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 758968 42858 758996 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42794 758996 42858 759008 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 758996 42582 759008 6 porb_h
port 761 nsew signal input
rlabel metal1 s 674006 772760 674070 772772 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 772760 673794 772772 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 772772 674070 772800 6 porb_h
port 761 nsew signal input
rlabel metal1 s 674006 772800 674070 772812 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673730 772800 673794 772812 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 786564 675450 786576 6 porb_h
port 761 nsew signal input
rlabel metal1 s 674006 786564 674070 786576 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 786564 673518 786576 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 786576 675450 786604 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 786604 675450 786616 6 porb_h
port 761 nsew signal input
rlabel metal1 s 674006 786604 674070 786616 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 786604 673518 786616 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 786632 42582 786644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 786632 41846 786644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 786644 42582 786672 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42518 786672 42582 786684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 41782 786672 41846 786684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 875168 675450 875180 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 875168 673518 875180 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 875180 675450 875208 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 875208 675450 875220 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 875208 673518 875220 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42242 957516 42306 957568 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42260 957568 42288 957720 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42242 957720 42306 957772 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 965268 675450 965280 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 965268 673518 965280 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 965280 675450 965308 6 porb_h
port 761 nsew signal input
rlabel metal1 s 675386 965308 675450 965320 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 965308 673518 965320 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 990020 673518 990032 6 porb_h
port 761 nsew signal input
rlabel metal1 s 626552 990032 673518 990060 6 porb_h
port 761 nsew signal input
rlabel metal1 s 673454 990060 673518 990072 6 porb_h
port 761 nsew signal input
rlabel metal1 s 628668 990060 628696 990088 6 porb_h
port 761 nsew signal input
rlabel metal1 s 626552 990060 626580 990088 6 porb_h
port 761 nsew signal input
rlabel metal1 s 628650 990088 628714 990140 6 porb_h
port 761 nsew signal input
rlabel metal1 s 626534 990088 626598 990140 6 porb_h
port 761 nsew signal input
rlabel metal1 s 78858 990156 78922 990168 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42242 990156 42306 990168 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42242 990168 78922 990196 6 porb_h
port 761 nsew signal input
rlabel metal1 s 78858 990196 78922 990208 6 porb_h
port 761 nsew signal input
rlabel metal1 s 42242 990196 42306 990208 6 porb_h
port 761 nsew signal input
rlabel metal1 s 286962 990564 287026 990576 6 porb_h
port 761 nsew signal input
rlabel metal1 s 286962 990576 386552 990604 6 porb_h
port 761 nsew signal input
rlabel metal1 s 386524 990604 386552 990632 6 porb_h
port 761 nsew signal input
rlabel metal1 s 286962 990604 287026 990616 6 porb_h
port 761 nsew signal input
rlabel metal1 s 626534 990632 626598 990644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 526898 990632 526962 990644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 475470 990632 475534 990644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 386506 990632 386570 990644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 181714 990632 181778 990644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 130286 990632 130350 990644 6 porb_h
port 761 nsew signal input
rlabel metal1 s 386506 990644 626598 990672 6 porb_h
port 761 nsew signal input
rlabel metal1 s 626534 990672 626598 990684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 526898 990672 526962 990684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 475470 990672 475534 990684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 386506 990672 386570 990684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 130286 990644 194732 990672 6 porb_h
port 761 nsew signal input
rlabel metal1 s 286962 990768 287026 990780 6 porb_h
port 761 nsew signal input
rlabel metal1 s 284662 990768 284726 990780 6 porb_h
port 761 nsew signal input
rlabel metal1 s 233050 990768 233114 990780 6 porb_h
port 761 nsew signal input
rlabel metal1 s 194704 990672 194732 990780 6 porb_h
port 761 nsew signal input
rlabel metal1 s 181714 990672 181778 990684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 130286 990672 130350 990684 6 porb_h
port 761 nsew signal input
rlabel metal1 s 194704 990780 287026 990808 6 porb_h
port 761 nsew signal input
rlabel metal1 s 130286 990768 130350 990780 6 porb_h
port 761 nsew signal input
rlabel metal1 s 78858 990768 78922 990780 6 porb_h
port 761 nsew signal input
rlabel metal1 s 78858 990780 130350 990808 6 porb_h
port 761 nsew signal input
rlabel metal1 s 286962 990808 287026 990820 6 porb_h
port 761 nsew signal input
rlabel metal1 s 284662 990808 284726 990820 6 porb_h
port 761 nsew signal input
rlabel metal1 s 233050 990808 233114 990820 6 porb_h
port 761 nsew signal input
rlabel metal1 s 130286 990808 130350 990820 6 porb_h
port 761 nsew signal input
rlabel metal1 s 78858 990808 78922 990820 6 porb_h
port 761 nsew signal input
rlabel metal1 s 145091 39934 145143 40000 6 porb_h
port 762 nsew signal input
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 763 nsew signal input
rlabel metal3 s 141820 37046 141966 37818 6 resetb_core_h
port 764 nsew signal output
rlabel metal3 s 141667 37818 141966 37911 6 resetb_core_h
port 764 nsew signal output
rlabel metal3 s 141873 37911 141966 37971 6 resetb_core_h
port 764 nsew signal output
rlabel metal3 s 141667 37911 141820 37971 6 resetb_core_h
port 764 nsew signal output
rlabel metal3 s 141667 37971 141873 38031 6 resetb_core_h
port 764 nsew signal output
rlabel metal3 s 141667 38031 141813 40000 6 resetb_core_h
port 764 nsew signal output
rlabel metal2 s 141667 39934 141813 40000 6 resetb_core_h
port 765 nsew signal output
rlabel metal4 s 679377 922346 680307 951854 6 vccd1
port 766 nsew signal bidirectional
rlabel metal4 s 679377 878146 680307 907854 6 vccd1
port 767 nsew signal bidirectional
rlabel metal5 s 679397 922346 680287 951854 6 vccd1
port 768 nsew signal bidirectional
rlabel metal5 s 679397 878146 680287 907854 6 vccd1
port 769 nsew signal bidirectional
rlabel metal3 s 678000 917700 679380 922500 6 vccd1
port 770 nsew signal bidirectional
rlabel metal3 s 678000 907660 679380 912449 6 vccd1
port 771 nsew signal bidirectional
rlabel metal5 s 698028 909409 711514 920737 6 vccd1
port 772 nsew signal bidirectional
rlabel metal4 s 680587 833207 681277 862606 6 vdda1
port 773 nsew signal bidirectional
rlabel metal4 s 680587 789007 681277 818593 6 vdda1
port 774 nsew signal bidirectional
rlabel metal5 s 680607 833207 681257 862606 6 vdda1
port 775 nsew signal bidirectional
rlabel metal5 s 680607 789007 681257 818593 6 vdda1
port 776 nsew signal bidirectional
rlabel metal3 s 677600 828521 680592 833301 6 vdda1
port 777 nsew signal bidirectional
rlabel metal3 s 677685 513707 677751 513710 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677685 513710 677794 513773 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677734 513773 677794 513921 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677600 513921 680592 518701 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677501 818347 677567 818350 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677501 818350 677794 818410 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677734 818410 677794 818542 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677501 818410 677567 818413 6 vdda1
port 778 nsew signal bidirectional
rlabel metal3 s 677600 818542 680592 823322 6 vdda1
port 778 nsew signal bidirectional
rlabel via2 s 677690 513712 677746 513768 6 vdda1
port 778 nsew signal bidirectional
rlabel via2 s 677506 818352 677562 818408 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 677690 513703 677746 513777 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 677692 513777 677744 513806 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675300 513742 675352 513806 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675312 513806 675340 548270 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 548270 675340 548298 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 548298 675248 556158 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 556158 675340 556186 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675312 556186 675340 593166 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675300 593166 675352 593230 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675300 593370 675352 593434 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675312 593434 675340 645730 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675300 645730 675352 645794 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675208 646002 675260 646066 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 646066 675248 646870 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 646870 675340 646898 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675312 646898 675340 683318 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 683318 675340 683346 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 683346 675248 691614 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 691614 675340 691642 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675312 691642 675340 728334 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 728334 675340 728362 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 728362 675248 736630 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675220 736630 675340 736658 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675312 736658 675340 781390 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675300 781390 675352 781454 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675300 781594 675352 781658 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675312 781658 675340 818314 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 677508 818314 677560 818343 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 677506 818343 677562 818417 6 vdda1
port 778 nsew signal bidirectional
rlabel metal2 s 675300 818314 675352 818378 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 677692 513748 677744 513800 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675300 513748 675352 513800 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675300 593172 675352 593224 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675300 593376 675352 593428 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675300 645736 675352 645788 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675208 646008 675260 646060 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675300 781396 675352 781448 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675300 781600 675352 781652 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 677508 818320 677560 818372 6 vdda1
port 778 nsew signal bidirectional
rlabel via1 s 675300 818320 675352 818372 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 677686 513748 677750 513760 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 513748 675358 513760 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 513760 677750 513788 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 677686 513788 677750 513800 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 513788 675358 513800 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 593172 675358 593224 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675312 593224 675340 593376 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 593376 675358 593428 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 645736 675358 645748 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675220 645748 675358 645776 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 645776 675358 645788 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675220 645776 675248 646008 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675202 646008 675266 646060 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 781396 675358 781448 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675312 781448 675340 781600 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 781600 675358 781652 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 677502 818320 677566 818332 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 818320 675358 818332 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 818332 677566 818360 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 677502 818360 677566 818372 6 vdda1
port 778 nsew signal bidirectional
rlabel metal1 s 675294 818360 675358 818372 6 vdda1
port 778 nsew signal bidirectional
rlabel metal5 s 698402 819640 710925 832180 6 vdda1
port 779 nsew signal bidirectional
rlabel metal4 s 539946 1004947 575854 1005637 6 vssa1
port 780 nsew signal bidirectional
rlabel metal4 s 533618 1008881 575854 1008947 6 vssa1
port 781 nsew signal bidirectional
rlabel metal4 s 575600 1007929 575854 1008165 6 vssa1
port 782 nsew signal bidirectional
rlabel metal4 s 533618 1007147 575854 1007213 6 vssa1
port 783 nsew signal bidirectional
rlabel metal4 s 590346 1004947 626254 1005637 6 vssa1
port 784 nsew signal bidirectional
rlabel metal4 s 590346 1007147 626522 1007213 6 vssa1
port 785 nsew signal bidirectional
rlabel metal4 s 590346 1008881 626522 1008947 6 vssa1
port 786 nsew signal bidirectional
rlabel metal4 s 590346 1007929 590600 1008165 6 vssa1
port 787 nsew signal bidirectional
rlabel metal5 s 540200 1004967 575600 1004968 6 vssa1
port 788 nsew signal bidirectional
rlabel metal5 s 539946 1004968 575854 1005617 6 vssa1
port 788 nsew signal bidirectional
rlabel metal5 s 539946 1007147 575854 1008947 6 vssa1
port 789 nsew signal bidirectional
rlabel metal5 s 590600 1004967 626000 1004968 6 vssa1
port 790 nsew signal bidirectional
rlabel metal5 s 590346 1004968 626254 1005617 6 vssa1
port 790 nsew signal bidirectional
rlabel metal5 s 590346 1007147 626254 1008947 6 vssa1
port 791 nsew signal bidirectional
rlabel metal3 s 677600 425721 684103 427792 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 677315 427787 677385 427792 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 677315 427792 684103 427852 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 677600 427852 684103 430501 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 677315 427852 677385 427857 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 585039 997383 585109 997386 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 585039 997386 585794 997446 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 585734 997446 585794 997600 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 585039 997446 585109 997453 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 585678 997600 590458 1004952 6 vssa1
port 792 nsew signal bidirectional
rlabel via2 s 677320 427792 677380 427852 6 vssa1
port 792 nsew signal bidirectional
rlabel via2 s 585044 997388 585104 997448 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 677311 427792 677389 427808 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 677124 427790 677176 427808 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 677124 427808 677389 427836 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 677311 427836 677389 427852 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 677124 427836 677176 427854 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 674748 427790 674800 427854 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 674760 427854 674788 992190 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 674748 992190 674800 992254 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 585048 992190 585100 992254 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 585060 992254 585088 997379 6 vssa1
port 792 nsew signal bidirectional
rlabel metal2 s 585044 997379 585104 997457 6 vssa1
port 792 nsew signal bidirectional
rlabel via1 s 677124 427796 677176 427848 6 vssa1
port 792 nsew signal bidirectional
rlabel via1 s 674748 427796 674800 427848 6 vssa1
port 792 nsew signal bidirectional
rlabel via1 s 674748 992196 674800 992248 6 vssa1
port 792 nsew signal bidirectional
rlabel via1 s 585048 992196 585100 992248 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 677118 427796 677182 427808 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 674742 427796 674806 427808 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 674742 427808 677182 427836 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 677118 427836 677182 427848 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 674742 427836 674806 427848 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 674742 992196 674806 992208 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 585042 992196 585106 992208 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 585042 992208 674806 992236 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 674742 992236 674806 992248 6 vssa1
port 792 nsew signal bidirectional
rlabel metal1 s 585042 992236 585106 992248 6 vssa1
port 792 nsew signal bidirectional
rlabel metal3 s 575699 997600 580479 1004103 6 vssa1
port 793 nsew signal bidirectional
rlabel metal5 s 576820 1018402 589360 1030925 6 vssa1
port 794 nsew signal bidirectional
rlabel metal4 s 685917 474546 686847 504054 6 vssd1
port 795 nsew signal bidirectional
rlabel metal4 s 685917 430346 686847 460054 6 vssd1
port 796 nsew signal bidirectional
rlabel metal5 s 685937 474546 686827 504054 6 vssd1
port 797 nsew signal bidirectional
rlabel metal5 s 685937 430346 686827 460054 6 vssd1
port 798 nsew signal bidirectional
rlabel metal3 s 678000 469900 685920 474700 6 vssd1
port 799 nsew signal bidirectional
rlabel metal3 s 678000 459860 685920 464649 6 vssd1
port 800 nsew signal bidirectional
rlabel metal5 s 698028 461609 711514 472937 6 vssd1
port 801 nsew signal bidirectional
rlabel metal4 s 37293 884546 38223 912254 6 vccd2
port 802 nsew signal bidirectional
rlabel metal4 s 37293 926746 38223 954454 6 vccd2
port 803 nsew signal bidirectional
rlabel metal5 s 37313 884546 38203 912254 6 vccd2
port 804 nsew signal bidirectional
rlabel metal5 s 37313 926746 38203 954454 6 vccd2
port 805 nsew signal bidirectional
rlabel metal3 s 38220 912100 39600 916900 6 vccd2
port 806 nsew signal bidirectional
rlabel metal3 s 38220 922151 39600 926940 6 vccd2
port 807 nsew signal bidirectional
rlabel metal5 s 6086 913863 19572 925191 6 vccd2
port 808 nsew signal bidirectional
rlabel metal4 s 36323 455607 37013 483193 6 vdda2
port 809 nsew signal bidirectional
rlabel metal4 s 36323 497807 37013 525393 6 vdda2
port 810 nsew signal bidirectional
rlabel metal5 s 36343 455607 36993 483193 6 vdda2
port 811 nsew signal bidirectional
rlabel metal5 s 36343 497807 36993 525393 6 vdda2
port 812 nsew signal bidirectional
rlabel metal3 s 37008 483099 40000 487879 6 vdda2
port 813 nsew signal bidirectional
rlabel metal3 s 37008 493078 40000 497858 6 vdda2
port 814 nsew signal bidirectional
rlabel metal5 s 6675 484220 19198 496760 6 vdda2
port 815 nsew signal bidirectional
rlabel metal4 s 31963 800146 32653 827854 6 vssa2
port 816 nsew signal bidirectional
rlabel metal4 s 28653 793818 28719 827854 6 vssa2
port 817 nsew signal bidirectional
rlabel metal4 s 29435 827600 29671 827854 6 vssa2
port 818 nsew signal bidirectional
rlabel metal4 s 30387 793818 30453 827854 6 vssa2
port 819 nsew signal bidirectional
rlabel metal4 s 31963 842346 32653 870054 6 vssa2
port 820 nsew signal bidirectional
rlabel metal4 s 30387 842346 30453 954722 6 vssa2
port 821 nsew signal bidirectional
rlabel metal4 s 28653 842346 28719 954722 6 vssa2
port 822 nsew signal bidirectional
rlabel metal4 s 29435 842346 29671 842600 6 vssa2
port 823 nsew signal bidirectional
rlabel metal5 s 31983 800146 32632 800400 6 vssa2
port 824 nsew signal bidirectional
rlabel metal5 s 31983 800400 32633 827600 6 vssa2
port 824 nsew signal bidirectional
rlabel metal5 s 31983 827600 32632 827854 6 vssa2
port 824 nsew signal bidirectional
rlabel metal5 s 28653 800146 30453 827854 6 vssa2
port 825 nsew signal bidirectional
rlabel metal5 s 31983 842346 32632 842600 6 vssa2
port 826 nsew signal bidirectional
rlabel metal5 s 31983 842600 32633 869800 6 vssa2
port 826 nsew signal bidirectional
rlabel metal5 s 31983 869800 32632 870054 6 vssa2
port 826 nsew signal bidirectional
rlabel metal5 s 28653 842346 30453 870054 6 vssa2
port 827 nsew signal bidirectional
rlabel metal3 s 32648 837678 40000 842458 6 vssa2
port 828 nsew signal bidirectional
rlabel metal3 s 33497 827699 40000 832479 6 vssa2
port 829 nsew signal bidirectional
rlabel metal5 s 6675 828820 19198 841360 6 vssa2
port 830 nsew signal bidirectional
rlabel metal4 s 30753 413346 31683 441054 6 vssd2
port 831 nsew signal bidirectional
rlabel metal4 s 30753 455546 31683 483254 6 vssd2
port 832 nsew signal bidirectional
rlabel metal5 s 30773 413346 31663 441054 6 vssd2
port 833 nsew signal bidirectional
rlabel metal5 s 30773 455546 31663 483254 6 vssd2
port 834 nsew signal bidirectional
rlabel metal3 s 31680 440900 39600 445700 6 vssd2
port 835 nsew signal bidirectional
rlabel metal3 s 31680 450951 39600 455740 6 vssd2
port 836 nsew signal bidirectional
rlabel metal5 s 6086 442663 19572 453991 6 vssd2
port 837 nsew signal bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 717600 1037600
string LEFview TRUE
string GDS_FILE ../gds/chip_io.gds
string GDS_END 36571046
string GDS_START 36076602
<< end >>
