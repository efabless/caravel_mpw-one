magic
tech sky130A
magscale 1 2
timestamp 1623348512
<< checkpaint >>
rect -1260 -1260 1930 2648
<< nwell >>
rect 0 0 670 1388
<< pmos >>
rect 171 189 201 1199
rect 257 189 307 1199
rect 363 189 413 1199
rect 469 189 499 1199
<< pdiff >>
rect 111 1187 171 1199
rect 111 1153 126 1187
rect 160 1153 171 1187
rect 111 1119 171 1153
rect 111 1085 126 1119
rect 160 1085 171 1119
rect 111 1051 171 1085
rect 111 1017 126 1051
rect 160 1017 171 1051
rect 111 983 171 1017
rect 111 949 126 983
rect 160 949 171 983
rect 111 915 171 949
rect 111 881 126 915
rect 160 881 171 915
rect 111 847 171 881
rect 111 813 126 847
rect 160 813 171 847
rect 111 779 171 813
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 1187 257 1199
rect 201 1153 212 1187
rect 246 1153 257 1187
rect 201 1119 257 1153
rect 201 1085 212 1119
rect 246 1085 257 1119
rect 201 1051 257 1085
rect 201 1017 212 1051
rect 246 1017 257 1051
rect 201 983 257 1017
rect 201 949 212 983
rect 246 949 257 983
rect 201 915 257 949
rect 201 881 212 915
rect 246 881 257 915
rect 201 847 257 881
rect 201 813 212 847
rect 246 813 257 847
rect 201 779 257 813
rect 201 745 212 779
rect 246 745 257 779
rect 201 711 257 745
rect 201 677 212 711
rect 246 677 257 711
rect 201 643 257 677
rect 201 609 212 643
rect 246 609 257 643
rect 201 575 257 609
rect 201 541 212 575
rect 246 541 257 575
rect 201 507 257 541
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 307 1187 363 1199
rect 307 1153 318 1187
rect 352 1153 363 1187
rect 307 1119 363 1153
rect 307 1085 318 1119
rect 352 1085 363 1119
rect 307 1051 363 1085
rect 307 1017 318 1051
rect 352 1017 363 1051
rect 307 983 363 1017
rect 307 949 318 983
rect 352 949 363 983
rect 307 915 363 949
rect 307 881 318 915
rect 352 881 363 915
rect 307 847 363 881
rect 307 813 318 847
rect 352 813 363 847
rect 307 779 363 813
rect 307 745 318 779
rect 352 745 363 779
rect 307 711 363 745
rect 307 677 318 711
rect 352 677 363 711
rect 307 643 363 677
rect 307 609 318 643
rect 352 609 363 643
rect 307 575 363 609
rect 307 541 318 575
rect 352 541 363 575
rect 307 507 363 541
rect 307 473 318 507
rect 352 473 363 507
rect 307 439 363 473
rect 307 405 318 439
rect 352 405 363 439
rect 307 371 363 405
rect 307 337 318 371
rect 352 337 363 371
rect 307 303 363 337
rect 307 269 318 303
rect 352 269 363 303
rect 307 235 363 269
rect 307 201 318 235
rect 352 201 363 235
rect 307 189 363 201
rect 413 1187 469 1199
rect 413 1153 424 1187
rect 458 1153 469 1187
rect 413 1119 469 1153
rect 413 1085 424 1119
rect 458 1085 469 1119
rect 413 1051 469 1085
rect 413 1017 424 1051
rect 458 1017 469 1051
rect 413 983 469 1017
rect 413 949 424 983
rect 458 949 469 983
rect 413 915 469 949
rect 413 881 424 915
rect 458 881 469 915
rect 413 847 469 881
rect 413 813 424 847
rect 458 813 469 847
rect 413 779 469 813
rect 413 745 424 779
rect 458 745 469 779
rect 413 711 469 745
rect 413 677 424 711
rect 458 677 469 711
rect 413 643 469 677
rect 413 609 424 643
rect 458 609 469 643
rect 413 575 469 609
rect 413 541 424 575
rect 458 541 469 575
rect 413 507 469 541
rect 413 473 424 507
rect 458 473 469 507
rect 413 439 469 473
rect 413 405 424 439
rect 458 405 469 439
rect 413 371 469 405
rect 413 337 424 371
rect 458 337 469 371
rect 413 303 469 337
rect 413 269 424 303
rect 458 269 469 303
rect 413 235 469 269
rect 413 201 424 235
rect 458 201 469 235
rect 413 189 469 201
rect 499 1187 559 1199
rect 499 1153 510 1187
rect 544 1153 559 1187
rect 499 1119 559 1153
rect 499 1085 510 1119
rect 544 1085 559 1119
rect 499 1051 559 1085
rect 499 1017 510 1051
rect 544 1017 559 1051
rect 499 983 559 1017
rect 499 949 510 983
rect 544 949 559 983
rect 499 915 559 949
rect 499 881 510 915
rect 544 881 559 915
rect 499 847 559 881
rect 499 813 510 847
rect 544 813 559 847
rect 499 779 559 813
rect 499 745 510 779
rect 544 745 559 779
rect 499 711 559 745
rect 499 677 510 711
rect 544 677 559 711
rect 499 643 559 677
rect 499 609 510 643
rect 544 609 559 643
rect 499 575 559 609
rect 499 541 510 575
rect 544 541 559 575
rect 499 507 559 541
rect 499 473 510 507
rect 544 473 559 507
rect 499 439 559 473
rect 499 405 510 439
rect 544 405 559 439
rect 499 371 559 405
rect 499 337 510 371
rect 544 337 559 371
rect 499 303 559 337
rect 499 269 510 303
rect 544 269 559 303
rect 499 235 559 269
rect 499 201 510 235
rect 544 201 559 235
rect 499 189 559 201
<< pdiffc >>
rect 126 1153 160 1187
rect 126 1085 160 1119
rect 126 1017 160 1051
rect 126 949 160 983
rect 126 881 160 915
rect 126 813 160 847
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 1153 246 1187
rect 212 1085 246 1119
rect 212 1017 246 1051
rect 212 949 246 983
rect 212 881 246 915
rect 212 813 246 847
rect 212 745 246 779
rect 212 677 246 711
rect 212 609 246 643
rect 212 541 246 575
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 318 1153 352 1187
rect 318 1085 352 1119
rect 318 1017 352 1051
rect 318 949 352 983
rect 318 881 352 915
rect 318 813 352 847
rect 318 745 352 779
rect 318 677 352 711
rect 318 609 352 643
rect 318 541 352 575
rect 318 473 352 507
rect 318 405 352 439
rect 318 337 352 371
rect 318 269 352 303
rect 318 201 352 235
rect 424 1153 458 1187
rect 424 1085 458 1119
rect 424 1017 458 1051
rect 424 949 458 983
rect 424 881 458 915
rect 424 813 458 847
rect 424 745 458 779
rect 424 677 458 711
rect 424 609 458 643
rect 424 541 458 575
rect 424 473 458 507
rect 424 405 458 439
rect 424 337 458 371
rect 424 269 458 303
rect 424 201 458 235
rect 510 1153 544 1187
rect 510 1085 544 1119
rect 510 1017 544 1051
rect 510 949 544 983
rect 510 881 544 915
rect 510 813 544 847
rect 510 745 544 779
rect 510 677 544 711
rect 510 609 544 643
rect 510 541 544 575
rect 510 473 544 507
rect 510 405 544 439
rect 510 337 544 371
rect 510 269 544 303
rect 510 201 544 235
<< nsubdiff >>
rect 41 1187 111 1199
rect 41 1153 58 1187
rect 92 1153 111 1187
rect 41 1119 111 1153
rect 41 1085 58 1119
rect 92 1085 111 1119
rect 41 1051 111 1085
rect 41 1017 58 1051
rect 92 1017 111 1051
rect 41 983 111 1017
rect 41 949 58 983
rect 92 949 111 983
rect 41 915 111 949
rect 41 881 58 915
rect 92 881 111 915
rect 41 847 111 881
rect 41 813 58 847
rect 92 813 111 847
rect 41 779 111 813
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 559 1187 629 1199
rect 559 1153 578 1187
rect 612 1153 629 1187
rect 559 1119 629 1153
rect 559 1085 578 1119
rect 612 1085 629 1119
rect 559 1051 629 1085
rect 559 1017 578 1051
rect 612 1017 629 1051
rect 559 983 629 1017
rect 559 949 578 983
rect 612 949 629 983
rect 559 915 629 949
rect 559 881 578 915
rect 612 881 629 915
rect 559 847 629 881
rect 559 813 578 847
rect 612 813 629 847
rect 559 779 629 813
rect 559 745 578 779
rect 612 745 629 779
rect 559 711 629 745
rect 559 677 578 711
rect 612 677 629 711
rect 559 643 629 677
rect 559 609 578 643
rect 612 609 629 643
rect 559 575 629 609
rect 559 541 578 575
rect 612 541 629 575
rect 559 507 629 541
rect 559 473 578 507
rect 612 473 629 507
rect 559 439 629 473
rect 559 405 578 439
rect 612 405 629 439
rect 559 371 629 405
rect 559 337 578 371
rect 612 337 629 371
rect 559 303 629 337
rect 559 269 578 303
rect 612 269 629 303
rect 559 235 629 269
rect 559 201 578 235
rect 612 201 629 235
rect 559 189 629 201
<< nsubdiffcont >>
rect 58 1153 92 1187
rect 58 1085 92 1119
rect 58 1017 92 1051
rect 58 949 92 983
rect 58 881 92 915
rect 58 813 92 847
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 578 1153 612 1187
rect 578 1085 612 1119
rect 578 1017 612 1051
rect 578 949 612 983
rect 578 881 612 915
rect 578 813 612 847
rect 578 745 612 779
rect 578 677 612 711
rect 578 609 612 643
rect 578 541 612 575
rect 578 473 612 507
rect 578 405 612 439
rect 578 337 612 371
rect 578 269 612 303
rect 578 201 612 235
<< poly >>
rect 243 1367 427 1388
rect 243 1333 278 1367
rect 312 1333 358 1367
rect 392 1333 427 1367
rect 243 1299 427 1333
rect 120 1281 201 1297
rect 120 1247 136 1281
rect 170 1247 201 1281
rect 243 1265 278 1299
rect 312 1265 358 1299
rect 392 1265 427 1299
rect 243 1249 427 1265
rect 469 1281 550 1297
rect 120 1231 201 1247
rect 171 1199 201 1231
rect 257 1199 307 1249
rect 363 1199 413 1249
rect 469 1247 500 1281
rect 534 1247 550 1281
rect 469 1231 550 1247
rect 469 1199 499 1231
rect 171 157 201 189
rect 120 141 201 157
rect 120 107 136 141
rect 170 107 201 141
rect 257 139 307 189
rect 363 139 413 189
rect 469 157 499 189
rect 469 141 550 157
rect 120 91 201 107
rect 243 123 427 139
rect 243 89 278 123
rect 312 89 358 123
rect 392 89 427 123
rect 469 107 500 141
rect 534 107 550 141
rect 469 91 550 107
rect 243 55 427 89
rect 243 21 278 55
rect 312 21 358 55
rect 392 21 427 55
rect 243 0 427 21
<< polycont >>
rect 278 1333 312 1367
rect 358 1333 392 1367
rect 136 1247 170 1281
rect 278 1265 312 1299
rect 358 1265 392 1299
rect 500 1247 534 1281
rect 136 107 170 141
rect 278 89 312 123
rect 358 89 392 123
rect 500 107 534 141
rect 278 21 312 55
rect 358 21 392 55
<< locali >>
rect 248 1369 422 1388
rect 248 1335 276 1369
rect 310 1367 360 1369
rect 248 1333 278 1335
rect 312 1333 358 1367
rect 394 1335 422 1369
rect 392 1333 422 1335
rect 248 1299 422 1333
rect 248 1297 278 1299
rect 120 1281 186 1297
rect 120 1247 136 1281
rect 170 1247 186 1281
rect 248 1263 276 1297
rect 312 1265 358 1299
rect 392 1297 422 1299
rect 310 1263 360 1265
rect 394 1263 422 1297
rect 248 1249 422 1263
rect 484 1281 550 1297
rect 120 1231 186 1247
rect 484 1247 500 1281
rect 534 1247 550 1281
rect 484 1231 550 1247
rect 120 1203 160 1231
rect 510 1203 550 1231
rect 41 1187 160 1203
rect 41 1153 58 1187
rect 92 1179 126 1187
rect 94 1153 126 1179
rect 41 1145 60 1153
rect 94 1145 160 1153
rect 41 1119 160 1145
rect 41 1085 58 1119
rect 92 1107 126 1119
rect 94 1085 126 1107
rect 41 1073 60 1085
rect 94 1073 160 1085
rect 41 1051 160 1073
rect 41 1017 58 1051
rect 92 1035 126 1051
rect 94 1017 126 1035
rect 41 1001 60 1017
rect 94 1001 160 1017
rect 41 983 160 1001
rect 41 949 58 983
rect 92 963 126 983
rect 94 949 126 963
rect 41 929 60 949
rect 94 929 160 949
rect 41 915 160 929
rect 41 881 58 915
rect 92 891 126 915
rect 94 881 126 891
rect 41 857 60 881
rect 94 857 160 881
rect 41 847 160 857
rect 41 813 58 847
rect 92 819 126 847
rect 94 813 126 819
rect 41 785 60 813
rect 94 785 160 813
rect 41 779 160 785
rect 41 745 58 779
rect 92 747 126 779
rect 94 745 126 747
rect 41 713 60 745
rect 94 713 160 745
rect 41 711 160 713
rect 41 677 58 711
rect 92 677 126 711
rect 41 675 160 677
rect 41 643 60 675
rect 94 643 160 675
rect 41 609 58 643
rect 94 641 126 643
rect 92 609 126 641
rect 41 603 160 609
rect 41 575 60 603
rect 94 575 160 603
rect 41 541 58 575
rect 94 569 126 575
rect 92 541 126 569
rect 41 531 160 541
rect 41 507 60 531
rect 94 507 160 531
rect 41 473 58 507
rect 94 497 126 507
rect 92 473 126 497
rect 41 459 160 473
rect 41 439 60 459
rect 94 439 160 459
rect 41 405 58 439
rect 94 425 126 439
rect 92 405 126 425
rect 41 387 160 405
rect 41 371 60 387
rect 94 371 160 387
rect 41 337 58 371
rect 94 353 126 371
rect 92 337 126 353
rect 41 315 160 337
rect 41 303 60 315
rect 94 303 160 315
rect 41 269 58 303
rect 94 281 126 303
rect 92 269 126 281
rect 41 243 160 269
rect 41 235 60 243
rect 94 235 160 243
rect 41 201 58 235
rect 94 209 126 235
rect 92 201 126 209
rect 41 185 160 201
rect 212 1187 246 1203
rect 212 1119 246 1145
rect 212 1051 246 1073
rect 212 983 246 1001
rect 212 915 246 929
rect 212 847 246 857
rect 212 779 246 785
rect 212 711 246 713
rect 212 675 246 677
rect 212 603 246 609
rect 212 531 246 541
rect 212 459 246 473
rect 212 387 246 405
rect 212 315 246 337
rect 212 243 246 269
rect 212 185 246 201
rect 318 1187 352 1203
rect 318 1119 352 1145
rect 318 1051 352 1073
rect 318 983 352 1001
rect 318 915 352 929
rect 318 847 352 857
rect 318 779 352 785
rect 318 711 352 713
rect 318 675 352 677
rect 318 603 352 609
rect 318 531 352 541
rect 318 459 352 473
rect 318 387 352 405
rect 318 315 352 337
rect 318 243 352 269
rect 318 185 352 201
rect 424 1187 458 1203
rect 424 1119 458 1145
rect 424 1051 458 1073
rect 424 983 458 1001
rect 424 915 458 929
rect 424 847 458 857
rect 424 779 458 785
rect 424 711 458 713
rect 424 675 458 677
rect 424 603 458 609
rect 424 531 458 541
rect 424 459 458 473
rect 424 387 458 405
rect 424 315 458 337
rect 424 243 458 269
rect 424 185 458 201
rect 510 1187 629 1203
rect 544 1179 578 1187
rect 544 1153 576 1179
rect 612 1153 629 1187
rect 510 1145 576 1153
rect 610 1145 629 1153
rect 510 1119 629 1145
rect 544 1107 578 1119
rect 544 1085 576 1107
rect 612 1085 629 1119
rect 510 1073 576 1085
rect 610 1073 629 1085
rect 510 1051 629 1073
rect 544 1035 578 1051
rect 544 1017 576 1035
rect 612 1017 629 1051
rect 510 1001 576 1017
rect 610 1001 629 1017
rect 510 983 629 1001
rect 544 963 578 983
rect 544 949 576 963
rect 612 949 629 983
rect 510 929 576 949
rect 610 929 629 949
rect 510 915 629 929
rect 544 891 578 915
rect 544 881 576 891
rect 612 881 629 915
rect 510 857 576 881
rect 610 857 629 881
rect 510 847 629 857
rect 544 819 578 847
rect 544 813 576 819
rect 612 813 629 847
rect 510 785 576 813
rect 610 785 629 813
rect 510 779 629 785
rect 544 747 578 779
rect 544 745 576 747
rect 612 745 629 779
rect 510 713 576 745
rect 610 713 629 745
rect 510 711 629 713
rect 544 677 578 711
rect 612 677 629 711
rect 510 675 629 677
rect 510 643 576 675
rect 610 643 629 675
rect 544 641 576 643
rect 544 609 578 641
rect 612 609 629 643
rect 510 603 629 609
rect 510 575 576 603
rect 610 575 629 603
rect 544 569 576 575
rect 544 541 578 569
rect 612 541 629 575
rect 510 531 629 541
rect 510 507 576 531
rect 610 507 629 531
rect 544 497 576 507
rect 544 473 578 497
rect 612 473 629 507
rect 510 459 629 473
rect 510 439 576 459
rect 610 439 629 459
rect 544 425 576 439
rect 544 405 578 425
rect 612 405 629 439
rect 510 387 629 405
rect 510 371 576 387
rect 610 371 629 387
rect 544 353 576 371
rect 544 337 578 353
rect 612 337 629 371
rect 510 315 629 337
rect 510 303 576 315
rect 610 303 629 315
rect 544 281 576 303
rect 544 269 578 281
rect 612 269 629 303
rect 510 243 629 269
rect 510 235 576 243
rect 610 235 629 243
rect 544 209 576 235
rect 544 201 578 209
rect 612 201 629 235
rect 510 185 629 201
rect 120 157 160 185
rect 510 157 550 185
rect 120 141 186 157
rect 120 107 136 141
rect 170 107 186 141
rect 484 141 550 157
rect 120 91 186 107
rect 248 125 422 139
rect 248 91 276 125
rect 310 123 360 125
rect 248 89 278 91
rect 312 89 358 123
rect 394 91 422 125
rect 484 107 500 141
rect 534 107 550 141
rect 484 91 550 107
rect 392 89 422 91
rect 248 55 422 89
rect 248 53 278 55
rect 248 19 276 53
rect 312 21 358 55
rect 392 53 422 55
rect 310 19 360 21
rect 394 19 422 53
rect 248 0 422 19
<< viali >>
rect 276 1367 310 1369
rect 360 1367 394 1369
rect 276 1335 278 1367
rect 278 1335 310 1367
rect 360 1335 392 1367
rect 392 1335 394 1367
rect 276 1265 278 1297
rect 278 1265 310 1297
rect 360 1265 392 1297
rect 392 1265 394 1297
rect 276 1263 310 1265
rect 360 1263 394 1265
rect 60 1153 92 1179
rect 92 1153 94 1179
rect 60 1145 94 1153
rect 60 1085 92 1107
rect 92 1085 94 1107
rect 60 1073 94 1085
rect 60 1017 92 1035
rect 92 1017 94 1035
rect 60 1001 94 1017
rect 60 949 92 963
rect 92 949 94 963
rect 60 929 94 949
rect 60 881 92 891
rect 92 881 94 891
rect 60 857 94 881
rect 60 813 92 819
rect 92 813 94 819
rect 60 785 94 813
rect 60 745 92 747
rect 92 745 94 747
rect 60 713 94 745
rect 60 643 94 675
rect 60 641 92 643
rect 92 641 94 643
rect 60 575 94 603
rect 60 569 92 575
rect 92 569 94 575
rect 60 507 94 531
rect 60 497 92 507
rect 92 497 94 507
rect 60 439 94 459
rect 60 425 92 439
rect 92 425 94 439
rect 60 371 94 387
rect 60 353 92 371
rect 92 353 94 371
rect 60 303 94 315
rect 60 281 92 303
rect 92 281 94 303
rect 60 235 94 243
rect 60 209 92 235
rect 92 209 94 235
rect 212 1153 246 1179
rect 212 1145 246 1153
rect 212 1085 246 1107
rect 212 1073 246 1085
rect 212 1017 246 1035
rect 212 1001 246 1017
rect 212 949 246 963
rect 212 929 246 949
rect 212 881 246 891
rect 212 857 246 881
rect 212 813 246 819
rect 212 785 246 813
rect 212 745 246 747
rect 212 713 246 745
rect 212 643 246 675
rect 212 641 246 643
rect 212 575 246 603
rect 212 569 246 575
rect 212 507 246 531
rect 212 497 246 507
rect 212 439 246 459
rect 212 425 246 439
rect 212 371 246 387
rect 212 353 246 371
rect 212 303 246 315
rect 212 281 246 303
rect 212 235 246 243
rect 212 209 246 235
rect 318 1153 352 1179
rect 318 1145 352 1153
rect 318 1085 352 1107
rect 318 1073 352 1085
rect 318 1017 352 1035
rect 318 1001 352 1017
rect 318 949 352 963
rect 318 929 352 949
rect 318 881 352 891
rect 318 857 352 881
rect 318 813 352 819
rect 318 785 352 813
rect 318 745 352 747
rect 318 713 352 745
rect 318 643 352 675
rect 318 641 352 643
rect 318 575 352 603
rect 318 569 352 575
rect 318 507 352 531
rect 318 497 352 507
rect 318 439 352 459
rect 318 425 352 439
rect 318 371 352 387
rect 318 353 352 371
rect 318 303 352 315
rect 318 281 352 303
rect 318 235 352 243
rect 318 209 352 235
rect 424 1153 458 1179
rect 424 1145 458 1153
rect 424 1085 458 1107
rect 424 1073 458 1085
rect 424 1017 458 1035
rect 424 1001 458 1017
rect 424 949 458 963
rect 424 929 458 949
rect 424 881 458 891
rect 424 857 458 881
rect 424 813 458 819
rect 424 785 458 813
rect 424 745 458 747
rect 424 713 458 745
rect 424 643 458 675
rect 424 641 458 643
rect 424 575 458 603
rect 424 569 458 575
rect 424 507 458 531
rect 424 497 458 507
rect 424 439 458 459
rect 424 425 458 439
rect 424 371 458 387
rect 424 353 458 371
rect 424 303 458 315
rect 424 281 458 303
rect 424 235 458 243
rect 424 209 458 235
rect 576 1153 578 1179
rect 578 1153 610 1179
rect 576 1145 610 1153
rect 576 1085 578 1107
rect 578 1085 610 1107
rect 576 1073 610 1085
rect 576 1017 578 1035
rect 578 1017 610 1035
rect 576 1001 610 1017
rect 576 949 578 963
rect 578 949 610 963
rect 576 929 610 949
rect 576 881 578 891
rect 578 881 610 891
rect 576 857 610 881
rect 576 813 578 819
rect 578 813 610 819
rect 576 785 610 813
rect 576 745 578 747
rect 578 745 610 747
rect 576 713 610 745
rect 576 643 610 675
rect 576 641 578 643
rect 578 641 610 643
rect 576 575 610 603
rect 576 569 578 575
rect 578 569 610 575
rect 576 507 610 531
rect 576 497 578 507
rect 578 497 610 507
rect 576 439 610 459
rect 576 425 578 439
rect 578 425 610 439
rect 576 371 610 387
rect 576 353 578 371
rect 578 353 610 371
rect 576 303 610 315
rect 576 281 578 303
rect 578 281 610 303
rect 576 235 610 243
rect 576 209 578 235
rect 578 209 610 235
rect 276 123 310 125
rect 360 123 394 125
rect 276 91 278 123
rect 278 91 310 123
rect 360 91 392 123
rect 392 91 394 123
rect 276 21 278 53
rect 278 21 310 53
rect 360 21 392 53
rect 392 21 394 53
rect 276 19 310 21
rect 360 19 394 21
<< metal1 >>
rect 250 1369 420 1388
rect 250 1335 276 1369
rect 310 1335 360 1369
rect 394 1335 420 1369
rect 250 1297 420 1335
rect 250 1263 276 1297
rect 310 1263 360 1297
rect 394 1263 420 1297
rect 250 1251 420 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 203 1179 255 1191
rect 203 1145 212 1179
rect 246 1145 255 1179
rect 203 1107 255 1145
rect 203 1073 212 1107
rect 246 1073 255 1107
rect 203 1035 255 1073
rect 203 1001 212 1035
rect 246 1001 255 1035
rect 203 963 255 1001
rect 203 929 212 963
rect 246 929 255 963
rect 203 891 255 929
rect 203 857 212 891
rect 246 857 255 891
rect 203 819 255 857
rect 203 785 212 819
rect 246 785 255 819
rect 203 747 255 785
rect 203 713 212 747
rect 246 713 255 747
rect 203 675 255 713
rect 203 641 212 675
rect 246 641 255 675
rect 203 639 255 641
rect 203 575 212 587
rect 246 575 255 587
rect 203 511 212 523
rect 246 511 255 523
rect 203 447 212 459
rect 246 447 255 459
rect 203 387 255 395
rect 203 383 212 387
rect 246 383 255 387
rect 203 319 255 331
rect 203 255 255 267
rect 203 197 255 203
rect 309 1185 361 1191
rect 309 1121 361 1133
rect 309 1057 361 1069
rect 309 1001 318 1005
rect 352 1001 361 1005
rect 309 993 361 1001
rect 309 929 318 941
rect 352 929 361 941
rect 309 865 318 877
rect 352 865 361 877
rect 309 801 318 813
rect 352 801 361 813
rect 309 747 361 749
rect 309 713 318 747
rect 352 713 361 747
rect 309 675 361 713
rect 309 641 318 675
rect 352 641 361 675
rect 309 603 361 641
rect 309 569 318 603
rect 352 569 361 603
rect 309 531 361 569
rect 309 497 318 531
rect 352 497 361 531
rect 309 459 361 497
rect 309 425 318 459
rect 352 425 361 459
rect 309 387 361 425
rect 309 353 318 387
rect 352 353 361 387
rect 309 315 361 353
rect 309 281 318 315
rect 352 281 361 315
rect 309 243 361 281
rect 309 209 318 243
rect 352 209 361 243
rect 309 197 361 209
rect 415 1179 467 1191
rect 415 1145 424 1179
rect 458 1145 467 1179
rect 415 1107 467 1145
rect 415 1073 424 1107
rect 458 1073 467 1107
rect 415 1035 467 1073
rect 415 1001 424 1035
rect 458 1001 467 1035
rect 415 963 467 1001
rect 415 929 424 963
rect 458 929 467 963
rect 415 891 467 929
rect 415 857 424 891
rect 458 857 467 891
rect 415 819 467 857
rect 415 785 424 819
rect 458 785 467 819
rect 415 747 467 785
rect 415 713 424 747
rect 458 713 467 747
rect 415 675 467 713
rect 415 641 424 675
rect 458 641 467 675
rect 415 639 467 641
rect 415 575 424 587
rect 458 575 467 587
rect 415 511 424 523
rect 458 511 467 523
rect 415 447 424 459
rect 458 447 467 459
rect 415 387 467 395
rect 415 383 424 387
rect 458 383 467 387
rect 415 319 467 331
rect 415 255 467 267
rect 415 197 467 203
rect 570 1179 629 1191
rect 570 1145 576 1179
rect 610 1145 629 1179
rect 570 1107 629 1145
rect 570 1073 576 1107
rect 610 1073 629 1107
rect 570 1035 629 1073
rect 570 1001 576 1035
rect 610 1001 629 1035
rect 570 963 629 1001
rect 570 929 576 963
rect 610 929 629 963
rect 570 891 629 929
rect 570 857 576 891
rect 610 857 629 891
rect 570 819 629 857
rect 570 785 576 819
rect 610 785 629 819
rect 570 747 629 785
rect 570 713 576 747
rect 610 713 629 747
rect 570 675 629 713
rect 570 641 576 675
rect 610 641 629 675
rect 570 603 629 641
rect 570 569 576 603
rect 610 569 629 603
rect 570 531 629 569
rect 570 497 576 531
rect 610 497 629 531
rect 570 459 629 497
rect 570 425 576 459
rect 610 425 629 459
rect 570 387 629 425
rect 570 353 576 387
rect 610 353 629 387
rect 570 315 629 353
rect 570 281 576 315
rect 610 281 629 315
rect 570 243 629 281
rect 570 209 576 243
rect 610 209 629 243
rect 570 197 629 209
rect 250 125 420 137
rect 250 91 276 125
rect 310 91 360 125
rect 394 91 420 125
rect 250 53 420 91
rect 250 19 276 53
rect 310 19 360 53
rect 394 19 420 53
rect 250 0 420 19
<< via1 >>
rect 203 603 255 639
rect 203 587 212 603
rect 212 587 246 603
rect 246 587 255 603
rect 203 569 212 575
rect 212 569 246 575
rect 246 569 255 575
rect 203 531 255 569
rect 203 523 212 531
rect 212 523 246 531
rect 246 523 255 531
rect 203 497 212 511
rect 212 497 246 511
rect 246 497 255 511
rect 203 459 255 497
rect 203 425 212 447
rect 212 425 246 447
rect 246 425 255 447
rect 203 395 255 425
rect 203 353 212 383
rect 212 353 246 383
rect 246 353 255 383
rect 203 331 255 353
rect 203 315 255 319
rect 203 281 212 315
rect 212 281 246 315
rect 246 281 255 315
rect 203 267 255 281
rect 203 243 255 255
rect 203 209 212 243
rect 212 209 246 243
rect 246 209 255 243
rect 203 203 255 209
rect 309 1179 361 1185
rect 309 1145 318 1179
rect 318 1145 352 1179
rect 352 1145 361 1179
rect 309 1133 361 1145
rect 309 1107 361 1121
rect 309 1073 318 1107
rect 318 1073 352 1107
rect 352 1073 361 1107
rect 309 1069 361 1073
rect 309 1035 361 1057
rect 309 1005 318 1035
rect 318 1005 352 1035
rect 352 1005 361 1035
rect 309 963 361 993
rect 309 941 318 963
rect 318 941 352 963
rect 352 941 361 963
rect 309 891 361 929
rect 309 877 318 891
rect 318 877 352 891
rect 352 877 361 891
rect 309 857 318 865
rect 318 857 352 865
rect 352 857 361 865
rect 309 819 361 857
rect 309 813 318 819
rect 318 813 352 819
rect 352 813 361 819
rect 309 785 318 801
rect 318 785 352 801
rect 352 785 361 801
rect 309 749 361 785
rect 415 603 467 639
rect 415 587 424 603
rect 424 587 458 603
rect 458 587 467 603
rect 415 569 424 575
rect 424 569 458 575
rect 458 569 467 575
rect 415 531 467 569
rect 415 523 424 531
rect 424 523 458 531
rect 458 523 467 531
rect 415 497 424 511
rect 424 497 458 511
rect 458 497 467 511
rect 415 459 467 497
rect 415 425 424 447
rect 424 425 458 447
rect 458 425 467 447
rect 415 395 467 425
rect 415 353 424 383
rect 424 353 458 383
rect 458 353 467 383
rect 415 331 467 353
rect 415 315 467 319
rect 415 281 424 315
rect 424 281 458 315
rect 458 281 467 315
rect 415 267 467 281
rect 415 243 467 255
rect 415 209 424 243
rect 424 209 458 243
rect 458 209 467 243
rect 415 203 467 209
<< metal2 >>
rect 14 1185 656 1191
rect 14 1133 309 1185
rect 361 1133 656 1185
rect 14 1121 656 1133
rect 14 1069 309 1121
rect 361 1069 656 1121
rect 14 1057 656 1069
rect 14 1005 309 1057
rect 361 1005 656 1057
rect 14 993 656 1005
rect 14 941 309 993
rect 361 941 656 993
rect 14 929 656 941
rect 14 877 309 929
rect 361 877 656 929
rect 14 865 656 877
rect 14 813 309 865
rect 361 813 656 865
rect 14 801 656 813
rect 14 749 309 801
rect 361 749 656 801
rect 14 719 656 749
rect 14 639 656 669
rect 14 587 203 639
rect 255 587 415 639
rect 467 587 656 639
rect 14 575 656 587
rect 14 523 203 575
rect 255 523 415 575
rect 467 523 656 575
rect 14 511 656 523
rect 14 459 203 511
rect 255 459 415 511
rect 467 459 656 511
rect 14 447 656 459
rect 14 395 203 447
rect 255 395 415 447
rect 467 395 656 447
rect 14 383 656 395
rect 14 331 203 383
rect 255 331 415 383
rect 467 331 656 383
rect 14 319 656 331
rect 14 267 203 319
rect 255 267 415 319
rect 467 267 656 319
rect 14 255 656 267
rect 14 203 203 255
rect 255 203 415 255
rect 467 203 656 255
rect 14 197 656 203
<< labels >>
flabel comment s 182 664 182 664 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 482 668 482 668 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 1288 414 1339 0 FreeSans 200 0 0 0 GATE
port 3 nsew
flabel metal1 s 255 44 414 95 0 FreeSans 200 0 0 0 GATE
port 3 nsew
flabel metal1 s 570 683 629 713 0 FreeSans 200 90 0 0 BULK
port 1 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 BULK
port 1 nsew
flabel metal2 s 14 384 35 512 7 FreeSans 300 180 0 0 SOURCE
port 4 nsew
flabel metal2 s 14 908 35 1036 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9687804
string GDS_START 9667720
<< end >>
