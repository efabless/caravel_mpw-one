magic
tech micross
magscale 1 2
timestamp 1611856895
<< checkpaint >>
rect -27000 -27000 27000 27000
<< rdl >>
tri -4689 26590 0 27000 se
rect 0 26590 27000 27000
tri -9235 25372 -4689 26590 se
rect -4689 25372 27000 26590
tri -13500 23383 -9235 25372 se
rect -9235 23383 27000 25372
tri -15475 22000 -13500 23383 se
rect -13500 22000 27000 23383
tri -15951 21666 -15475 22000 se
rect -15475 21666 -3820 22000
tri -3820 21666 0 22000 nw
tri 0 21666 3820 22000 ne
rect 3820 21666 27000 22000
tri -17355 20683 -15951 21666 se
rect -15951 20683 -7487 21666
tri -7487 20683 -3820 21666 nw
tri 3820 20683 7487 21666 ne
rect 7487 20683 27000 21666
tri -17365 20673 -17355 20683 se
rect -17355 20673 -7524 20683
tri -7524 20673 -7487 20683 nw
tri 7487 20673 7524 20683 ne
rect 7524 20673 27000 20683
tri -18985 19053 -17365 20673 se
rect -17365 19053 -11000 20673
tri -11000 19053 -7524 20673 nw
tri 7524 19053 11000 20673 ne
rect 11000 19053 27000 20673
tri -20683 17355 -18985 19053 se
rect -18985 17355 -13424 19053
tri -13424 17355 -11000 19053 nw
tri 11000 17355 13424 19053 ne
rect 13424 17355 27000 19053
tri -21035 16853 -20683 17355 se
rect -20683 16853 -14141 17355
tri -14141 16853 -13424 17355 nw
tri 13424 16853 14141 17355 ne
rect 14141 16853 27000 17355
tri -22934 14141 -21035 16852 se
rect -21035 14141 -16853 16853
tri -16853 14141 -14141 16853 nw
tri 14141 14141 16853 16853 ne
rect 16853 14141 27000 16853
tri -23383 13500 -22934 14141 se
rect -22934 13500 -17302 14141
tri -17302 13500 -16853 14141 nw
tri 16853 13500 17302 14141 ne
rect 17302 13500 27000 14141
tri -24549 11000 -23383 13500 se
rect -23383 11000 -19053 13500
tri -19053 11000 -17302 13500 nw
tri 17302 11000 19053 13500 ne
rect 19053 11000 27000 13500
tri -25372 9235 -24549 11000 se
rect -24549 9235 -19876 11000
tri -19876 9235 -19053 11000 nw
tri 19053 9235 19876 11000 ne
rect 19876 9235 27000 11000
tri -25830 7526 -25372 9235 se
rect -25372 7526 -20673 9235
rect -25830 7524 -20673 7526
tri -20673 7524 -19876 9235 nw
tri 19876 7524 20673 9235 ne
rect 20673 7524 27000 9235
tri -26590 4689 -25830 7524 se
rect -25830 4689 -21433 7524
tri -21433 4689 -20673 7524 nw
tri 20673 4689 21433 7524 ne
rect 21433 4689 27000 7524
tri -26666 3820 -26590 4689 se
rect -26590 3820 -21666 4689
tri -21666 3820 -21433 4689 nw
tri 21433 3820 21666 4689 ne
rect 21666 3820 27000 4689
tri -27000 0 -26666 3820 se
tri -27000 -3820 -26666 0 ne
rect -26666 -3820 -22000 3820
tri -22000 0 -21666 3820 nw
tri -22000 -3820 -21666 0 sw
tri 21666 0 22000 3820 ne
rect 22000 0 27000 3820
tri 21666 -3820 22000 0 se
rect 22000 -3820 26666 0
tri 26666 -3820 27000 0 nw
tri -26666 -4688 -26590 -3820 ne
rect -26590 -4688 -21666 -3820
tri -21666 -4688 -21433 -3820 sw
tri -26590 -7522 -25831 -4688 ne
rect -25831 -7524 -21433 -4688
tri 21433 -4688 21666 -3820 se
rect 21666 -4688 26590 -3820
rect 21433 -4689 26590 -4688
tri 26590 -4689 26666 -3820 nw
tri -21433 -7524 -20673 -4689 sw
tri 20673 -7524 21433 -4689 se
rect 21433 -7524 25830 -4689
tri 25830 -7524 26590 -4689 nw
tri -25831 -9235 -25372 -7524 ne
rect -25372 -9235 -20673 -7524
tri -20673 -9235 -19876 -7524 sw
tri 19876 -9235 20673 -7524 se
rect 20673 -7526 25830 -7524
rect 20673 -9235 25372 -7526
tri 25372 -9235 25830 -7526 nw
tri -25372 -11000 -24549 -9235 ne
rect -24549 -11000 -19876 -9235
tri -19876 -11000 -19053 -9235 sw
tri 19053 -11000 19876 -9235 se
rect 19876 -11000 24549 -9235
tri 24549 -11000 25372 -9235 nw
tri -24549 -13500 -23383 -11000 ne
rect -23383 -13500 -19053 -11000
tri -19053 -13500 -17302 -11000 sw
tri 17302 -13500 19053 -11000 se
rect 19053 -13500 23383 -11000
tri 23383 -13500 24549 -11000 nw
tri -23383 -14140 -22935 -13500 ne
rect -22935 -14141 -17302 -13500
tri -17302 -14141 -16853 -13500 sw
tri 16853 -14141 17302 -13500 se
rect 17302 -14141 22934 -13500
tri 22934 -14141 23383 -13500 nw
tri -22935 -16853 -21035 -14141 ne
rect -21035 -16853 -16853 -14141
tri -16853 -16853 -14141 -14141 sw
tri 14141 -16853 16853 -14141 se
rect 16853 -16853 21035 -14141
tri 21035 -16852 22934 -14141 nw
tri -21035 -17355 -20683 -16853 ne
rect -20683 -17355 -14141 -16853
tri -14141 -17355 -13424 -16853 sw
tri 13424 -17355 14141 -16853 se
rect 14141 -17355 20683 -16853
tri 20683 -17355 21035 -16853 nw
tri -20683 -19053 -18985 -17355 ne
rect -18985 -19053 -13424 -17355
tri -13424 -19053 -11000 -17355 sw
tri 11000 -19053 13424 -17355 se
rect 13424 -19053 18985 -17355
tri 18985 -19053 20683 -17355 nw
tri -18985 -20673 -17365 -19053 ne
rect -17365 -20673 -11000 -19053
tri -11000 -20673 -7524 -19053 sw
tri 7524 -20673 11000 -19053 se
rect 11000 -20673 17365 -19053
tri 17365 -20673 18985 -19053 nw
tri -17365 -20683 -17355 -20673 ne
rect -17355 -20683 -7524 -20673
tri -7524 -20683 -7487 -20673 sw
tri 7487 -20683 7524 -20673 se
rect 7524 -20683 17355 -20673
tri 17355 -20683 17365 -20673 nw
tri -17355 -21666 -15952 -20683 ne
rect -15952 -21666 -7487 -20683
tri -7487 -21666 -3820 -20683 sw
tri 3820 -21666 7487 -20683 se
rect 7487 -21666 15951 -20683
tri 15951 -21666 17355 -20683 nw
tri -15952 -22000 -15475 -21666 ne
rect -15475 -22000 -3820 -21666
tri -3820 -22000 0 -21666 sw
tri 0 -22000 3820 -21666 se
rect 3820 -22000 15475 -21666
tri 15475 -22000 15951 -21666 nw
tri -15475 -23383 -13500 -22000 ne
rect -13500 -23383 13500 -22000
tri 13500 -23383 15475 -22000 nw
tri -13500 -25372 -9235 -23383 ne
rect -9235 -25372 9235 -23383
tri 9235 -25372 13500 -23383 nw
tri -9235 -26590 -4689 -25372 ne
rect -4689 -26590 4688 -25372
tri 4688 -26590 9235 -25372 nw
tri -4689 -27000 0 -26590 ne
tri 0 -27000 4688 -26590 nw
<< pi2 >>
tri -3820 21666 0 22000 se
tri 0 21666 3820 22000 sw
tri -7487 20683 -3820 21666 se
rect -3820 20683 3820 21666
tri 3820 20683 7487 21666 sw
tri -7524 20673 -7487 20683 se
rect -7487 20673 7487 20683
tri 7487 20673 7524 20683 sw
tri -11000 19053 -7524 20673 se
rect -7524 19053 7524 20673
tri 7524 19053 11000 20673 sw
tri -13424 17355 -11000 19053 se
rect -11000 17355 11000 19053
tri 11000 17355 13424 19053 sw
tri -14141 16853 -13424 17355 se
rect -13424 16853 13424 17355
tri 13424 16853 14141 17355 sw
tri -16853 14141 -14141 16853 se
rect -14141 14141 14141 16853
tri 14141 14141 16853 16853 sw
tri -17302 13500 -16853 14141 se
rect -16853 13500 16853 14141
tri 16853 13500 17302 14141 sw
tri -19053 11000 -17302 13500 se
rect -17302 11000 17302 13500
tri 17302 11000 19053 13500 sw
tri -19876 9235 -19053 11000 se
rect -19053 9235 19053 11000
tri 19053 9235 19876 11000 sw
tri -20673 7524 -19876 9235 se
rect -19876 7524 19876 9235
tri 19876 7524 20673 9235 sw
tri -21433 4689 -20673 7524 se
rect -20673 4689 20673 7524
tri 20673 4689 21433 7524 sw
tri -21666 3820 -21433 4689 se
rect -21433 3820 21433 4689
tri 21433 3820 21666 4689 sw
tri -22000 0 -21666 3820 se
tri -22000 -3820 -21666 0 ne
rect -21666 -3820 21666 3820
tri 21666 0 22000 3820 sw
tri 21666 -3820 22000 0 nw
tri -21666 -4688 -21433 -3820 ne
rect -21433 -4689 21433 -3820
tri 21433 -4688 21666 -3820 nw
tri -21433 -7524 -20673 -4689 ne
rect -20673 -7524 20673 -4689
tri 20673 -7524 21433 -4689 nw
tri -20673 -9235 -19876 -7524 ne
rect -19876 -9235 19876 -7524
tri 19876 -9235 20673 -7524 nw
tri -19876 -11000 -19053 -9235 ne
rect -19053 -11000 19053 -9235
tri 19053 -11000 19876 -9235 nw
tri -19053 -13500 -17302 -11000 ne
rect -17302 -13500 17302 -11000
tri 17302 -13500 19053 -11000 nw
tri -17302 -14141 -16853 -13500 ne
rect -16853 -14141 16853 -13500
tri 16853 -14141 17302 -13500 nw
tri -16853 -16853 -14141 -14141 ne
rect -14141 -16853 14141 -14141
tri 14141 -16853 16853 -14141 nw
tri -14141 -17355 -13424 -16853 ne
rect -13424 -17355 13424 -16853
tri 13424 -17355 14141 -16853 nw
tri -13424 -19053 -11000 -17355 ne
rect -11000 -19053 11000 -17355
tri 11000 -19053 13424 -17355 nw
tri -11000 -20673 -7524 -19053 ne
rect -7524 -20673 7524 -19053
tri 7524 -20673 11000 -19053 nw
tri -7524 -20683 -7487 -20673 ne
rect -7487 -20683 7487 -20673
tri 7487 -20683 7524 -20673 nw
tri -7487 -21666 -3820 -20683 ne
rect -3820 -21666 3820 -20683
tri 3820 -21666 7487 -20683 nw
tri -3820 -22000 0 -21666 ne
tri 0 -22000 3820 -21666 nw
<< ubm >>
tri -4341 24620 0 25000 se
tri 0 24620 4341 25000 sw
tri -8551 23492 -4341 24620 se
rect -4341 23492 4341 24620
tri 4341 23492 8551 24620 sw
tri -12500 21651 -8551 23492 se
rect -8551 22000 8551 23492
rect -8551 21666 -3820 22000
tri -3820 21666 0 22000 nw
tri 0 21666 3820 22000 ne
rect 3820 21666 8551 22000
rect -8551 21651 -3876 21666
tri -3876 21651 -3820 21666 nw
tri 3820 21651 3875 21666 ne
rect 3875 21651 8551 21666
tri 8551 21651 12500 23492 sw
tri -16070 19151 -12500 21651 se
rect -12500 20673 -7524 21651
tri -7524 20673 -3876 21651 nw
tri 3875 20673 7524 21651 ne
rect 7524 20673 12500 21651
rect -12500 19151 -10790 20673
tri -10790 19151 -7524 20673 nw
tri 7524 19151 10789 20673 ne
rect 10789 19151 12500 20673
tri 12500 19151 16070 21651 sw
tri -18368 16853 -16070 19151 se
rect -16070 19053 -11000 19151
tri -11000 19053 -10790 19151 nw
tri 10789 19053 11000 19151 ne
rect 11000 19053 16070 19151
rect -16070 16853 -14141 19053
tri -14141 16853 -11000 19053 nw
tri 11000 16853 14141 19053 ne
rect 14141 16853 16070 19053
tri 16070 16853 18368 19151 sw
tri -19151 16070 -18368 16853 se
rect -18368 16070 -14924 16853
tri -14924 16070 -14141 16853 nw
tri 14141 16070 14924 16853 ne
rect 14924 16070 18368 16853
tri 18368 16070 19151 16853 sw
tri -21651 12500 -19151 16070 se
rect -19151 14141 -16853 16070
tri -16853 14141 -14924 16070 nw
tri 14924 14141 16853 16070 ne
rect 16853 14141 19151 16070
rect -19151 12500 -18002 14141
tri -18002 12501 -16853 14141 nw
tri 16853 12500 18002 14141 ne
rect 18002 12500 19151 14141
tri 19151 12500 21651 16070 sw
tri -23492 8551 -21651 12500 se
rect -21651 11000 -19053 12500
tri -19053 11000 -18002 12500 nw
tri 18002 11000 19053 12500 ne
rect 19053 11000 21651 12500
rect -21651 8551 -20194 11000
tri -20194 8552 -19053 11000 nw
tri 19053 8551 20194 11000 ne
rect 20194 8551 21651 11000
tri 21651 8551 23492 12500 sw
tri -24620 4341 -23492 8551 se
rect -23492 7524 -20673 8551
tri -20673 7524 -20194 8551 nw
tri 20194 7524 20673 8551 ne
rect 20673 7524 23492 8551
rect -23492 4341 -21526 7524
tri -21526 4342 -20673 7524 nw
tri 20673 4342 21526 7524 ne
tri -25000 0 -24620 4341 se
rect -24620 3820 -21666 4341
tri -21666 3820 -21526 4341 nw
rect 21526 4341 23492 7524
tri 23492 4341 24620 8551 sw
tri 21526 3820 21666 4341 ne
rect 21666 3820 24620 4341
tri -25000 -4341 -24620 0 ne
rect -24620 -3820 -22000 3820
tri -22000 0 -21666 3820 nw
tri -22000 -3820 -21666 0 sw
tri 21666 0 22000 3820 ne
tri 21666 -3820 22000 0 se
rect 22000 -3820 24620 3820
tri 24620 0 25000 4341 sw
rect -24620 -4339 -21666 -3820
tri -21666 -4339 -21527 -3820 sw
rect -24620 -4341 -21527 -4339
tri 21526 -4341 21666 -3820 se
rect 21666 -4341 24620 -3820
tri 24620 -4341 25000 0 nw
tri -24620 -8551 -23492 -4341 ne
rect -23492 -7524 -21527 -4341
tri -21527 -7524 -20673 -4341 sw
tri 20673 -7524 21526 -4342 se
rect 21526 -7524 23492 -4341
rect -23492 -8550 -20673 -7524
tri -20673 -8550 -20195 -7524 sw
rect -23492 -8551 -20195 -8550
tri 20194 -8551 20673 -7524 se
rect 20673 -8551 23492 -7524
tri 23492 -8551 24620 -4341 nw
tri -23492 -12500 -21651 -8551 ne
rect -21651 -11000 -20195 -8551
tri -20195 -11000 -19053 -8551 sw
tri 19053 -11000 20194 -8552 se
rect 20194 -11000 21651 -8551
rect -21651 -12500 -19053 -11000
tri -19053 -12500 -18003 -11000 sw
tri 18002 -12500 19053 -11000 se
rect 19053 -12500 21651 -11000
tri 21651 -12500 23492 -8551 nw
tri -21651 -16070 -19151 -12500 ne
rect -19151 -14141 -18003 -12500
tri -18003 -14141 -16853 -12500 sw
tri 16853 -14141 18002 -12501 se
rect 18002 -14141 19151 -12500
rect -19151 -16070 -16853 -14141
tri -16853 -16070 -14924 -14141 sw
tri 14924 -16070 16853 -14141 se
rect 16853 -16070 19151 -14141
tri 19151 -16070 21651 -12500 nw
tri -19151 -16853 -18368 -16070 ne
rect -18368 -16853 -14924 -16070
tri -14924 -16853 -14141 -16070 sw
tri 14141 -16853 14924 -16070 se
rect 14924 -16853 18368 -16070
tri 18368 -16853 19151 -16070 nw
tri -18368 -19151 -16070 -16853 ne
rect -16070 -19053 -14141 -16853
tri -14141 -19053 -11000 -16853 sw
tri 11000 -19053 14141 -16853 se
rect 14141 -19053 16070 -16853
rect -16070 -19151 -11000 -19053
tri -11000 -19151 -10790 -19053 sw
tri 10790 -19151 11000 -19053 se
rect 11000 -19151 16070 -19053
tri 16070 -19151 18368 -16853 nw
tri -16070 -21651 -12500 -19151 ne
rect -12500 -20673 -10790 -19151
tri -10790 -20673 -7524 -19151 sw
tri 7524 -20673 10790 -19151 se
rect 10790 -20673 12500 -19151
rect -12500 -21651 -7524 -20673
tri -7524 -21651 -3876 -20673 sw
tri 3876 -21651 7524 -20673 se
rect 7524 -21651 12500 -20673
tri 12500 -21651 16070 -19151 nw
tri -12500 -23492 -8551 -21651 ne
rect -8551 -21666 -3876 -21651
tri -3876 -21666 -3820 -21651 sw
tri 3820 -21666 3876 -21651 se
rect 3876 -21666 8551 -21651
rect -8551 -22000 -3820 -21666
tri -3820 -22000 0 -21666 sw
tri 0 -22000 3820 -21666 se
rect 3820 -22000 8551 -21666
rect -8551 -23492 8551 -22000
tri 8551 -23492 12500 -21651 nw
tri -8551 -24620 -4341 -23492 ne
rect -4341 -24620 4341 -23492
tri 4341 -24620 8551 -23492 nw
tri -4341 -25000 0 -24620 ne
tri 0 -25000 4341 -24620 nw
<< properties >>
string FIXED_BBOX -27000 -27000 27000 27000
<< end >>
