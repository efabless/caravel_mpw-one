magic
tech sky130A
magscale 12 1
timestamp 1598786148
<< metal5 >>
rect 0 75 30 105
rect 60 85 75 105
rect 55 80 75 85
rect 50 75 75 80
rect 45 70 70 75
rect 45 65 65 70
rect 40 60 60 65
rect 25 55 60 60
rect 20 50 55 55
rect 15 45 50 50
rect 15 40 35 45
rect 10 35 30 40
rect 5 30 30 35
rect 0 25 25 30
rect 0 20 20 25
rect 0 0 15 20
rect 45 0 75 30
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
