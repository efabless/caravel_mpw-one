magic
tech sky130A
magscale 12 1
timestamp 1598777283
<< metal5 >>
rect 10 70 45 75
rect 5 65 45 70
rect 0 60 45 65
rect 0 45 20 60
rect 0 40 35 45
rect 5 35 40 40
rect 10 30 45 35
rect 25 15 45 30
rect 0 10 45 15
rect 0 5 40 10
rect 0 0 35 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
