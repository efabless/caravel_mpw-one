magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1288 -1260 1700 1527
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_1
timestamp 1623348570
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_0
timestamp 1623348570
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_1
timestamp 1623348570
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1623348570
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 440 267 440 267 0 FreeSans 300 0 0 0 D
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48701544
string GDS_START 48699594
<< end >>
