magic
tech sky130A
magscale 1 2
timestamp 1606789654
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< pdiff >>
rect 77289 1034726 77323 1034752
rect 78523 1034726 78557 1034752
rect 128689 1034726 128723 1034752
rect 129923 1034726 129957 1034752
rect 180089 1034726 180123 1034752
rect 181323 1034726 181357 1034752
rect 231489 1034726 231523 1034752
rect 232723 1034726 232757 1034752
rect 283089 1034726 283123 1034752
rect 284323 1034726 284357 1034752
rect 384889 1034726 384923 1034752
rect 386123 1034726 386157 1034752
rect 473889 1034726 473923 1034752
rect 475123 1034726 475157 1034752
rect 525289 1034726 525323 1034752
rect 526523 1034726 526557 1034752
rect 627089 1034726 627123 1034752
rect 628323 1034726 628357 1034752
rect 82571 1032409 89682 1032431
rect 91517 1031619 91531 1032463
rect 133971 1032409 141082 1032431
rect 142917 1031619 142931 1032463
rect 185371 1032409 192482 1032431
rect 194317 1031619 194331 1032463
rect 236771 1032409 243882 1032431
rect 245717 1031619 245731 1032463
rect 288371 1032409 295482 1032431
rect 297317 1031619 297331 1032463
rect 390171 1032409 397282 1032431
rect 399117 1031619 399131 1032463
rect 479171 1032409 486282 1032431
rect 488117 1031619 488131 1032463
rect 530571 1032409 537682 1032431
rect 539517 1031619 539531 1032463
rect 632371 1032409 639482 1032431
rect 641317 1031619 641331 1032463
rect 91507 1031605 91531 1031619
rect 142907 1031605 142931 1031619
rect 194307 1031605 194331 1031619
rect 245707 1031605 245731 1031619
rect 297307 1031605 297331 1031619
rect 399107 1031605 399131 1031619
rect 488107 1031605 488131 1031619
rect 539507 1031605 539531 1031619
rect 641307 1031605 641331 1031619
rect 77501 1031579 89682 1031595
rect 89725 1031579 91531 1031605
rect 128901 1031579 141082 1031595
rect 141125 1031579 142931 1031605
rect 180301 1031579 192482 1031595
rect 192525 1031579 194331 1031605
rect 231701 1031579 243882 1031595
rect 243925 1031579 245731 1031605
rect 283301 1031579 295482 1031595
rect 295525 1031579 297331 1031605
rect 385101 1031579 397282 1031595
rect 397325 1031579 399131 1031605
rect 474101 1031579 486282 1031595
rect 486325 1031579 488131 1031605
rect 525501 1031579 537682 1031595
rect 537725 1031579 539531 1031605
rect 627301 1031579 639482 1031595
rect 639525 1031579 641331 1031605
rect 78136 1029211 78298 1030211
rect 90422 1029211 90463 1030211
rect 90984 1029211 91194 1030211
rect 129536 1029211 129698 1030211
rect 141822 1029211 141863 1030211
rect 142384 1029211 142594 1030211
rect 180936 1029211 181098 1030211
rect 193222 1029211 193263 1030211
rect 193784 1029211 193994 1030211
rect 232336 1029211 232498 1030211
rect 244622 1029211 244663 1030211
rect 245184 1029211 245394 1030211
rect 283936 1029211 284098 1030211
rect 296222 1029211 296263 1030211
rect 296784 1029211 296994 1030211
rect 385736 1029211 385898 1030211
rect 398022 1029211 398063 1030211
rect 398584 1029211 398794 1030211
rect 474736 1029211 474898 1030211
rect 487022 1029211 487063 1030211
rect 487584 1029211 487794 1030211
rect 526136 1029211 526298 1030211
rect 538422 1029211 538463 1030211
rect 538984 1029211 539194 1030211
rect 627936 1029211 628098 1030211
rect 640222 1029211 640263 1030211
rect 640784 1029211 640994 1030211
rect 78159 1027610 78299 1028610
rect 90422 1027610 90463 1028610
rect 90984 1027610 91194 1028610
rect 129559 1027610 129699 1028610
rect 141822 1027610 141863 1028610
rect 142384 1027610 142594 1028610
rect 180959 1027610 181099 1028610
rect 193222 1027610 193263 1028610
rect 193784 1027610 193994 1028610
rect 232359 1027610 232499 1028610
rect 244622 1027610 244663 1028610
rect 245184 1027610 245394 1028610
rect 283959 1027610 284099 1028610
rect 296222 1027610 296263 1028610
rect 296784 1027610 296994 1028610
rect 385759 1027610 385899 1028610
rect 398022 1027610 398063 1028610
rect 398584 1027610 398794 1028610
rect 474759 1027610 474899 1028610
rect 487022 1027610 487063 1028610
rect 487584 1027610 487794 1028610
rect 526159 1027610 526299 1028610
rect 538422 1027610 538463 1028610
rect 538984 1027610 539194 1028610
rect 627959 1027610 628099 1028610
rect 640222 1027610 640263 1028610
rect 640784 1027610 640994 1028610
rect 77035 1018110 77183 1022856
rect 77700 1020922 77726 1021922
rect 77771 1020922 77873 1021922
rect 90939 1020922 91094 1021922
rect 91264 1020922 91419 1021922
rect 77700 1019322 77726 1020322
rect 77771 1019322 77873 1020322
rect 90939 1019322 91094 1020322
rect 91264 1019322 91419 1020322
rect 128435 1018110 128583 1022856
rect 129100 1020922 129126 1021922
rect 129171 1020922 129273 1021922
rect 142339 1020922 142494 1021922
rect 142664 1020922 142819 1021922
rect 129100 1019322 129126 1020322
rect 129171 1019322 129273 1020322
rect 142339 1019322 142494 1020322
rect 142664 1019322 142819 1020322
rect 179835 1018110 179983 1022856
rect 180500 1020922 180526 1021922
rect 180571 1020922 180673 1021922
rect 193739 1020922 193894 1021922
rect 194064 1020922 194219 1021922
rect 180500 1019322 180526 1020322
rect 180571 1019322 180673 1020322
rect 193739 1019322 193894 1020322
rect 194064 1019322 194219 1020322
rect 231235 1018110 231383 1022856
rect 231900 1020922 231926 1021922
rect 231971 1020922 232073 1021922
rect 245139 1020922 245294 1021922
rect 245464 1020922 245619 1021922
rect 231900 1019322 231926 1020322
rect 231971 1019322 232073 1020322
rect 245139 1019322 245294 1020322
rect 245464 1019322 245619 1020322
rect 282835 1018110 282983 1022856
rect 283500 1020922 283526 1021922
rect 283571 1020922 283673 1021922
rect 296739 1020922 296894 1021922
rect 297064 1020922 297219 1021922
rect 283500 1019322 283526 1020322
rect 283571 1019322 283673 1020322
rect 296739 1019322 296894 1020322
rect 297064 1019322 297219 1020322
rect 384635 1018110 384783 1022856
rect 385300 1020922 385326 1021922
rect 385371 1020922 385473 1021922
rect 398539 1020922 398694 1021922
rect 398864 1020922 399019 1021922
rect 385300 1019322 385326 1020322
rect 385371 1019322 385473 1020322
rect 398539 1019322 398694 1020322
rect 398864 1019322 399019 1020322
rect 473635 1018110 473783 1022856
rect 474300 1020922 474326 1021922
rect 474371 1020922 474473 1021922
rect 487539 1020922 487694 1021922
rect 487864 1020922 488019 1021922
rect 474300 1019322 474326 1020322
rect 474371 1019322 474473 1020322
rect 487539 1019322 487694 1020322
rect 487864 1019322 488019 1020322
rect 525035 1018110 525183 1022856
rect 525700 1020922 525726 1021922
rect 525771 1020922 525873 1021922
rect 538939 1020922 539094 1021922
rect 539264 1020922 539419 1021922
rect 525700 1019322 525726 1020322
rect 525771 1019322 525873 1020322
rect 538939 1019322 539094 1020322
rect 539264 1019322 539419 1020322
rect 626835 1018110 626983 1022856
rect 627500 1020922 627526 1021922
rect 627571 1020922 627673 1021922
rect 640739 1020922 640894 1021922
rect 641064 1020922 641219 1021922
rect 627500 1019322 627526 1020322
rect 627571 1019322 627673 1020322
rect 640739 1019322 640894 1020322
rect 641064 1019322 641219 1020322
rect 77209 1018053 84133 1018084
rect 128609 1018053 135533 1018084
rect 180009 1018053 186933 1018084
rect 231409 1018053 238333 1018084
rect 283009 1018053 289933 1018084
rect 384809 1018053 391733 1018084
rect 473809 1018053 480733 1018084
rect 525209 1018053 532133 1018084
rect 627009 1018053 633933 1018084
rect 84137 1016817 85342 1016821
rect 135537 1016817 136742 1016821
rect 186937 1016817 188142 1016821
rect 238337 1016817 239542 1016821
rect 289937 1016817 291142 1016821
rect 391737 1016817 392942 1016821
rect 480737 1016817 481942 1016821
rect 532137 1016817 533342 1016821
rect 633937 1016817 635142 1016821
rect 77918 1016779 77974 1016791
rect 129318 1016779 129374 1016791
rect 180718 1016779 180774 1016791
rect 232118 1016779 232174 1016791
rect 283718 1016779 283774 1016791
rect 385518 1016779 385574 1016791
rect 474518 1016779 474574 1016791
rect 525918 1016779 525974 1016791
rect 627718 1016779 627774 1016791
rect 84763 1007758 85211 1007764
rect 87809 1007758 88283 1007764
rect 136163 1007758 136611 1007764
rect 139209 1007758 139683 1007764
rect 187563 1007758 188011 1007764
rect 190609 1007758 191083 1007764
rect 238963 1007758 239411 1007764
rect 242009 1007758 242483 1007764
rect 290563 1007758 291011 1007764
rect 293609 1007758 294083 1007764
rect 392363 1007758 392811 1007764
rect 395409 1007758 395883 1007764
rect 481363 1007758 481811 1007764
rect 484409 1007758 484883 1007764
rect 532763 1007758 533211 1007764
rect 535809 1007758 536283 1007764
rect 634563 1007758 635011 1007764
rect 637609 1007758 638083 1007764
rect 82935 1007645 88488 1007648
rect 134335 1007645 139888 1007648
rect 185735 1007645 191288 1007648
rect 237135 1007645 242688 1007648
rect 288735 1007645 294288 1007648
rect 390535 1007645 396088 1007648
rect 479535 1007645 485088 1007648
rect 530935 1007645 536488 1007648
rect 632735 1007645 638288 1007648
rect 83728 1007573 89477 1007585
rect 135128 1007573 140877 1007585
rect 186528 1007573 192277 1007585
rect 237928 1007573 243677 1007585
rect 289528 1007573 295277 1007585
rect 391328 1007573 397077 1007585
rect 480328 1007573 486077 1007585
rect 531728 1007573 537477 1007585
rect 633528 1007573 639277 1007585
rect 83728 1006882 83754 1007573
rect 135128 1006882 135154 1007573
rect 186528 1006882 186554 1007573
rect 237928 1006882 237954 1007573
rect 289528 1006882 289554 1007573
rect 391328 1006882 391354 1007573
rect 480328 1006882 480354 1007573
rect 531728 1006882 531754 1007573
rect 633528 1006882 633554 1007573
rect 83744 1006879 83754 1006882
rect 135144 1006879 135154 1006882
rect 186544 1006879 186554 1006882
rect 237944 1006879 237954 1006882
rect 289544 1006879 289554 1006882
rect 391344 1006879 391354 1006882
rect 480344 1006879 480354 1006882
rect 531744 1006879 531754 1006882
rect 633544 1006879 633554 1006882
rect 79916 1005803 79932 1006119
rect 81120 1005803 81138 1006119
rect 131316 1005803 131332 1006119
rect 132520 1005803 132538 1006119
rect 182716 1005803 182732 1006119
rect 183920 1005803 183938 1006119
rect 234116 1005803 234132 1006119
rect 235320 1005803 235338 1006119
rect 285716 1005803 285732 1006119
rect 286920 1005803 286938 1006119
rect 387516 1005803 387532 1006119
rect 388720 1005803 388738 1006119
rect 476516 1005803 476532 1006119
rect 477720 1005803 477738 1006119
rect 527916 1005803 527932 1006119
rect 529120 1005803 529138 1006119
rect 629716 1005803 629732 1006119
rect 630920 1005803 630938 1006119
rect 79916 1005777 79920 1005803
rect 131316 1005777 131320 1005803
rect 182716 1005777 182720 1005803
rect 234116 1005777 234120 1005803
rect 285716 1005777 285720 1005803
rect 387516 1005777 387520 1005803
rect 476516 1005777 476520 1005803
rect 527916 1005777 527920 1005803
rect 629716 1005777 629720 1005803
rect 79882 1005539 79920 1005777
rect 81140 1005539 81172 1005777
rect 131282 1005539 131320 1005777
rect 132540 1005539 132572 1005777
rect 182682 1005539 182720 1005777
rect 183940 1005539 183972 1005777
rect 234082 1005539 234120 1005777
rect 235340 1005539 235372 1005777
rect 285682 1005539 285720 1005777
rect 286940 1005539 286972 1005777
rect 387482 1005539 387520 1005777
rect 388740 1005539 388772 1005777
rect 476482 1005539 476520 1005777
rect 477740 1005539 477772 1005777
rect 527882 1005539 527920 1005777
rect 529140 1005539 529172 1005777
rect 629682 1005539 629720 1005777
rect 630940 1005539 630972 1005777
rect 80705 1001502 81195 1001529
rect 132105 1001502 132595 1001529
rect 183505 1001502 183995 1001529
rect 234905 1001502 235395 1001529
rect 286505 1001502 286995 1001529
rect 388305 1001502 388795 1001529
rect 477305 1001502 477795 1001529
rect 528705 1001502 529195 1001529
rect 630505 1001502 630995 1001529
rect 85213 998646 85239 998654
rect 88423 998646 88448 998654
rect 136613 998646 136639 998654
rect 139823 998646 139848 998654
rect 188013 998646 188039 998654
rect 191223 998646 191248 998654
rect 239413 998646 239439 998654
rect 242623 998646 242648 998654
rect 291013 998646 291039 998654
rect 294223 998646 294248 998654
rect 392813 998646 392839 998654
rect 396023 998646 396048 998654
rect 481813 998646 481839 998654
rect 485023 998646 485048 998654
rect 533213 998646 533239 998654
rect 536423 998646 536448 998654
rect 635013 998646 635039 998654
rect 638223 998646 638248 998654
rect 5137 969517 6021 969531
rect 5981 969507 6021 969517
rect 5995 967725 6021 969507
rect 15678 969264 16678 969419
rect 17278 969264 18278 969419
rect 7389 968984 8389 969194
rect 8990 968984 9990 969194
rect 15678 968939 16678 969094
rect 17278 968939 18278 969094
rect 7389 968422 8389 968463
rect 8990 968422 9990 968463
rect 5169 960571 5191 967682
rect 2848 956523 2874 956557
rect 6005 955501 6021 967682
rect 29836 965809 29842 966283
rect 20779 962137 20783 963342
rect 29836 962763 29842 963211
rect 7389 956136 8389 956298
rect 8990 956159 9990 956299
rect 15678 955771 16678 955873
rect 17278 955771 18278 955873
rect 15678 955700 16678 955726
rect 17278 955700 18278 955726
rect 2848 955289 2874 955323
rect 19516 955209 19547 962133
rect 29952 960935 29955 966488
rect 30015 961754 30027 967477
rect 698110 966617 702856 966765
rect 38946 966423 38954 966448
rect 696779 965826 696791 965882
rect 685539 963884 685777 963918
rect 685539 963880 686119 963884
rect 685803 963868 686119 963880
rect 38946 963213 38954 963239
rect 681502 962605 681529 963095
rect 685803 962662 686119 962680
rect 685539 962628 685777 962660
rect 30015 961744 30721 961754
rect 30015 961728 30718 961744
rect 686882 960056 687585 960072
rect 686879 960046 687585 960056
rect 31823 959140 32061 959172
rect 31481 959120 31797 959138
rect 36071 958705 36098 959195
rect 678646 958561 678654 958587
rect 31481 957920 31797 957932
rect 31481 957916 32061 957920
rect 31823 957882 32061 957916
rect 20809 955918 20821 955974
rect 678646 955352 678654 955377
rect 14744 955035 19490 955183
rect 687573 954323 687585 960046
rect 687645 955312 687648 960865
rect 698053 959667 698084 966591
rect 714726 966477 714752 966511
rect 699322 966074 700322 966100
rect 700922 966074 701922 966100
rect 699322 965927 700322 966029
rect 700922 965927 701922 966029
rect 707610 965501 708610 965641
rect 709211 965502 710211 965664
rect 687758 958589 687764 959037
rect 696817 958458 696821 959663
rect 687758 955517 687764 955991
rect 711579 954118 711595 966299
rect 714726 965243 714752 965277
rect 712409 954118 712431 961229
rect 707610 953337 708610 953378
rect 709211 953337 710211 953378
rect 699322 952706 700322 952861
rect 700922 952706 701922 952861
rect 707610 952606 708610 952816
rect 709211 952606 710211 952816
rect 699322 952381 700322 952536
rect 700922 952381 701922 952536
rect 711579 952293 711605 954075
rect 711579 952283 711619 952293
rect 711579 952269 712463 952283
rect 35930 919315 39318 919329
rect 678282 919187 681670 919245
rect 35930 915355 39318 915413
rect 678282 915271 681670 915285
rect 698110 877417 702856 877565
rect 696779 876626 696791 876682
rect 685539 874684 685777 874718
rect 685539 874680 686119 874684
rect 685803 874668 686119 874680
rect 681502 873405 681529 873895
rect 685803 873462 686119 873480
rect 685539 873428 685777 873460
rect 686882 870856 687585 870872
rect 686879 870846 687585 870856
rect 678646 869361 678654 869387
rect 678646 866152 678654 866177
rect 687573 865123 687585 870846
rect 687645 866112 687648 871665
rect 698053 870467 698084 877391
rect 714726 877277 714752 877311
rect 699322 876874 700322 876900
rect 700922 876874 701922 876900
rect 699322 876727 700322 876829
rect 700922 876727 701922 876829
rect 707610 876301 708610 876441
rect 709211 876302 710211 876464
rect 687758 869389 687764 869837
rect 696817 869258 696821 870463
rect 687758 866317 687764 866791
rect 711579 864918 711595 877099
rect 714726 876043 714752 876077
rect 712409 864918 712431 872029
rect 707610 864137 708610 864178
rect 709211 864137 710211 864178
rect 699322 863506 700322 863661
rect 700922 863506 701922 863661
rect 707610 863406 708610 863616
rect 709211 863406 710211 863616
rect 699322 863181 700322 863336
rect 700922 863181 701922 863336
rect 711579 863093 711605 864875
rect 711579 863083 711619 863093
rect 711579 863069 712463 863083
rect 5137 799717 6021 799731
rect 5981 799707 6021 799717
rect 5995 797925 6021 799707
rect 15678 799464 16678 799619
rect 17278 799464 18278 799619
rect 7389 799184 8389 799394
rect 8990 799184 9990 799394
rect 15678 799139 16678 799294
rect 17278 799139 18278 799294
rect 7389 798622 8389 798663
rect 8990 798622 9990 798663
rect 5169 790771 5191 797882
rect 2848 786723 2874 786757
rect 6005 785701 6021 797882
rect 29836 796009 29842 796483
rect 20779 792337 20783 793542
rect 29836 792963 29842 793411
rect 7389 786336 8389 786498
rect 8990 786359 9990 786499
rect 15678 785971 16678 786073
rect 17278 785971 18278 786073
rect 15678 785900 16678 785926
rect 17278 785900 18278 785926
rect 2848 785489 2874 785523
rect 19516 785409 19547 792333
rect 29952 791135 29955 796688
rect 30015 791954 30027 797677
rect 38946 796623 38954 796648
rect 38946 793413 38954 793439
rect 30015 791944 30721 791954
rect 30015 791928 30718 791944
rect 31823 789340 32061 789372
rect 31481 789320 31797 789338
rect 36071 788905 36098 789395
rect 698110 788217 702856 788365
rect 31481 788120 31797 788132
rect 31481 788116 32061 788120
rect 31823 788082 32061 788116
rect 696779 787426 696791 787482
rect 20809 786118 20821 786174
rect 685539 785484 685777 785518
rect 685539 785480 686119 785484
rect 685803 785468 686119 785480
rect 14744 785235 19490 785383
rect 681502 784205 681529 784695
rect 685803 784262 686119 784280
rect 685539 784228 685777 784260
rect 686882 781656 687585 781672
rect 686879 781646 687585 781656
rect 678646 780161 678654 780187
rect 678646 776952 678654 776977
rect 687573 775923 687585 781646
rect 687645 776912 687648 782465
rect 698053 781267 698084 788191
rect 714726 788077 714752 788111
rect 699322 787674 700322 787700
rect 700922 787674 701922 787700
rect 699322 787527 700322 787629
rect 700922 787527 701922 787629
rect 707610 787101 708610 787241
rect 709211 787102 710211 787264
rect 687758 780189 687764 780637
rect 696817 780058 696821 781263
rect 687758 777117 687764 777591
rect 711579 775718 711595 787899
rect 714726 786843 714752 786877
rect 712409 775718 712431 782829
rect 707610 774937 708610 774978
rect 709211 774937 710211 774978
rect 699322 774306 700322 774461
rect 700922 774306 701922 774461
rect 707610 774206 708610 774416
rect 709211 774206 710211 774416
rect 699322 773981 700322 774136
rect 700922 773981 701922 774136
rect 711579 773893 711605 775675
rect 711579 773883 711619 773893
rect 711579 773869 712463 773883
rect 5137 756517 6021 756531
rect 5981 756507 6021 756517
rect 5995 754725 6021 756507
rect 15678 756264 16678 756419
rect 17278 756264 18278 756419
rect 7389 755984 8389 756194
rect 8990 755984 9990 756194
rect 15678 755939 16678 756094
rect 17278 755939 18278 756094
rect 7389 755422 8389 755463
rect 8990 755422 9990 755463
rect 5169 747571 5191 754682
rect 2848 743523 2874 743557
rect 6005 742501 6021 754682
rect 29836 752809 29842 753283
rect 20779 749137 20783 750342
rect 29836 749763 29842 750211
rect 7389 743136 8389 743298
rect 8990 743159 9990 743299
rect 15678 742771 16678 742873
rect 17278 742771 18278 742873
rect 15678 742700 16678 742726
rect 17278 742700 18278 742726
rect 2848 742289 2874 742323
rect 19516 742209 19547 749133
rect 29952 747935 29955 753488
rect 30015 748754 30027 754477
rect 38946 753423 38954 753448
rect 38946 750213 38954 750239
rect 30015 748744 30721 748754
rect 30015 748728 30718 748744
rect 31823 746140 32061 746172
rect 31481 746120 31797 746138
rect 36071 745705 36098 746195
rect 31481 744920 31797 744932
rect 31481 744916 32061 744920
rect 31823 744882 32061 744916
rect 698110 743217 702856 743365
rect 20809 742918 20821 742974
rect 696779 742426 696791 742482
rect 14744 742035 19490 742183
rect 685539 740484 685777 740518
rect 685539 740480 686119 740484
rect 685803 740468 686119 740480
rect 681502 739205 681529 739695
rect 685803 739262 686119 739280
rect 685539 739228 685777 739260
rect 686882 736656 687585 736672
rect 686879 736646 687585 736656
rect 678646 735161 678654 735187
rect 678646 731952 678654 731977
rect 687573 730923 687585 736646
rect 687645 731912 687648 737465
rect 698053 736267 698084 743191
rect 714726 743077 714752 743111
rect 699322 742674 700322 742700
rect 700922 742674 701922 742700
rect 699322 742527 700322 742629
rect 700922 742527 701922 742629
rect 707610 742101 708610 742241
rect 709211 742102 710211 742264
rect 687758 735189 687764 735637
rect 696817 735058 696821 736263
rect 687758 732117 687764 732591
rect 711579 730718 711595 742899
rect 714726 741843 714752 741877
rect 712409 730718 712431 737829
rect 707610 729937 708610 729978
rect 709211 729937 710211 729978
rect 699322 729306 700322 729461
rect 700922 729306 701922 729461
rect 707610 729206 708610 729416
rect 709211 729206 710211 729416
rect 699322 728981 700322 729136
rect 700922 728981 701922 729136
rect 711579 728893 711605 730675
rect 711579 728883 711619 728893
rect 711579 728869 712463 728883
rect 5137 713317 6021 713331
rect 5981 713307 6021 713317
rect 5995 711525 6021 713307
rect 15678 713064 16678 713219
rect 17278 713064 18278 713219
rect 7389 712784 8389 712994
rect 8990 712784 9990 712994
rect 15678 712739 16678 712894
rect 17278 712739 18278 712894
rect 7389 712222 8389 712263
rect 8990 712222 9990 712263
rect 5169 704371 5191 711482
rect 2848 700323 2874 700357
rect 6005 699301 6021 711482
rect 29836 709609 29842 710083
rect 20779 705937 20783 707142
rect 29836 706563 29842 707011
rect 7389 699936 8389 700098
rect 8990 699959 9990 700099
rect 15678 699571 16678 699673
rect 17278 699571 18278 699673
rect 15678 699500 16678 699526
rect 17278 699500 18278 699526
rect 2848 699089 2874 699123
rect 19516 699009 19547 705933
rect 29952 704735 29955 710288
rect 30015 705554 30027 711277
rect 38946 710223 38954 710248
rect 38946 707013 38954 707039
rect 30015 705544 30721 705554
rect 30015 705528 30718 705544
rect 31823 702940 32061 702972
rect 31481 702920 31797 702938
rect 36071 702505 36098 702995
rect 31481 701720 31797 701732
rect 31481 701716 32061 701720
rect 31823 701682 32061 701716
rect 20809 699718 20821 699774
rect 14744 698835 19490 698983
rect 698110 698217 702856 698365
rect 696779 697426 696791 697482
rect 685539 695484 685777 695518
rect 685539 695480 686119 695484
rect 685803 695468 686119 695480
rect 681502 694205 681529 694695
rect 685803 694262 686119 694280
rect 685539 694228 685777 694260
rect 686882 691656 687585 691672
rect 686879 691646 687585 691656
rect 678646 690161 678654 690187
rect 678646 686952 678654 686977
rect 687573 685923 687585 691646
rect 687645 686912 687648 692465
rect 698053 691267 698084 698191
rect 714726 698077 714752 698111
rect 699322 697674 700322 697700
rect 700922 697674 701922 697700
rect 699322 697527 700322 697629
rect 700922 697527 701922 697629
rect 707610 697101 708610 697241
rect 709211 697102 710211 697264
rect 687758 690189 687764 690637
rect 696817 690058 696821 691263
rect 687758 687117 687764 687591
rect 711579 685718 711595 697899
rect 714726 696843 714752 696877
rect 712409 685718 712431 692829
rect 707610 684937 708610 684978
rect 709211 684937 710211 684978
rect 699322 684306 700322 684461
rect 700922 684306 701922 684461
rect 707610 684206 708610 684416
rect 709211 684206 710211 684416
rect 699322 683981 700322 684136
rect 700922 683981 701922 684136
rect 711579 683893 711605 685675
rect 711579 683883 711619 683893
rect 711579 683869 712463 683883
rect 5137 670117 6021 670131
rect 5981 670107 6021 670117
rect 5995 668325 6021 670107
rect 15678 669864 16678 670019
rect 17278 669864 18278 670019
rect 7389 669584 8389 669794
rect 8990 669584 9990 669794
rect 15678 669539 16678 669694
rect 17278 669539 18278 669694
rect 7389 669022 8389 669063
rect 8990 669022 9990 669063
rect 5169 661171 5191 668282
rect 2848 657123 2874 657157
rect 6005 656101 6021 668282
rect 29836 666409 29842 666883
rect 20779 662737 20783 663942
rect 29836 663363 29842 663811
rect 7389 656736 8389 656898
rect 8990 656759 9990 656899
rect 15678 656371 16678 656473
rect 17278 656371 18278 656473
rect 15678 656300 16678 656326
rect 17278 656300 18278 656326
rect 2848 655889 2874 655923
rect 19516 655809 19547 662733
rect 29952 661535 29955 667088
rect 30015 662354 30027 668077
rect 38946 667023 38954 667048
rect 38946 663813 38954 663839
rect 30015 662344 30721 662354
rect 30015 662328 30718 662344
rect 31823 659740 32061 659772
rect 31481 659720 31797 659738
rect 36071 659305 36098 659795
rect 31481 658520 31797 658532
rect 31481 658516 32061 658520
rect 31823 658482 32061 658516
rect 20809 656518 20821 656574
rect 14744 655635 19490 655783
rect 698110 653017 702856 653165
rect 696779 652226 696791 652282
rect 685539 650284 685777 650318
rect 685539 650280 686119 650284
rect 685803 650268 686119 650280
rect 681502 649005 681529 649495
rect 685803 649062 686119 649080
rect 685539 649028 685777 649060
rect 686882 646456 687585 646472
rect 686879 646446 687585 646456
rect 678646 644961 678654 644987
rect 678646 641752 678654 641777
rect 687573 640723 687585 646446
rect 687645 641712 687648 647265
rect 698053 646067 698084 652991
rect 714726 652877 714752 652911
rect 699322 652474 700322 652500
rect 700922 652474 701922 652500
rect 699322 652327 700322 652429
rect 700922 652327 701922 652429
rect 707610 651901 708610 652041
rect 709211 651902 710211 652064
rect 687758 644989 687764 645437
rect 696817 644858 696821 646063
rect 687758 641917 687764 642391
rect 711579 640518 711595 652699
rect 714726 651643 714752 651677
rect 712409 640518 712431 647629
rect 707610 639737 708610 639778
rect 709211 639737 710211 639778
rect 699322 639106 700322 639261
rect 700922 639106 701922 639261
rect 707610 639006 708610 639216
rect 709211 639006 710211 639216
rect 699322 638781 700322 638936
rect 700922 638781 701922 638936
rect 711579 638693 711605 640475
rect 711579 638683 711619 638693
rect 711579 638669 712463 638683
rect 5137 626917 6021 626931
rect 5981 626907 6021 626917
rect 5995 625125 6021 626907
rect 15678 626664 16678 626819
rect 17278 626664 18278 626819
rect 7389 626384 8389 626594
rect 8990 626384 9990 626594
rect 15678 626339 16678 626494
rect 17278 626339 18278 626494
rect 7389 625822 8389 625863
rect 8990 625822 9990 625863
rect 5169 617971 5191 625082
rect 2848 613923 2874 613957
rect 6005 612901 6021 625082
rect 29836 623209 29842 623683
rect 20779 619537 20783 620742
rect 29836 620163 29842 620611
rect 7389 613536 8389 613698
rect 8990 613559 9990 613699
rect 15678 613171 16678 613273
rect 17278 613171 18278 613273
rect 15678 613100 16678 613126
rect 17278 613100 18278 613126
rect 2848 612689 2874 612723
rect 19516 612609 19547 619533
rect 29952 618335 29955 623888
rect 30015 619154 30027 624877
rect 38946 623823 38954 623848
rect 38946 620613 38954 620639
rect 30015 619144 30721 619154
rect 30015 619128 30718 619144
rect 31823 616540 32061 616572
rect 31481 616520 31797 616538
rect 36071 616105 36098 616595
rect 31481 615320 31797 615332
rect 31481 615316 32061 615320
rect 31823 615282 32061 615316
rect 20809 613318 20821 613374
rect 14744 612435 19490 612583
rect 698110 608017 702856 608165
rect 696779 607226 696791 607282
rect 685539 605284 685777 605318
rect 685539 605280 686119 605284
rect 685803 605268 686119 605280
rect 681502 604005 681529 604495
rect 685803 604062 686119 604080
rect 685539 604028 685777 604060
rect 686882 601456 687585 601472
rect 686879 601446 687585 601456
rect 678646 599961 678654 599987
rect 678646 596752 678654 596777
rect 687573 595723 687585 601446
rect 687645 596712 687648 602265
rect 698053 601067 698084 607991
rect 714726 607877 714752 607911
rect 699322 607474 700322 607500
rect 700922 607474 701922 607500
rect 699322 607327 700322 607429
rect 700922 607327 701922 607429
rect 707610 606901 708610 607041
rect 709211 606902 710211 607064
rect 687758 599989 687764 600437
rect 696817 599858 696821 601063
rect 687758 596917 687764 597391
rect 711579 595518 711595 607699
rect 714726 606643 714752 606677
rect 712409 595518 712431 602629
rect 707610 594737 708610 594778
rect 709211 594737 710211 594778
rect 699322 594106 700322 594261
rect 700922 594106 701922 594261
rect 707610 594006 708610 594216
rect 709211 594006 710211 594216
rect 699322 593781 700322 593936
rect 700922 593781 701922 593936
rect 711579 593693 711605 595475
rect 711579 593683 711619 593693
rect 711579 593669 712463 593683
rect 5137 583717 6021 583731
rect 5981 583707 6021 583717
rect 5995 581925 6021 583707
rect 15678 583464 16678 583619
rect 17278 583464 18278 583619
rect 7389 583184 8389 583394
rect 8990 583184 9990 583394
rect 15678 583139 16678 583294
rect 17278 583139 18278 583294
rect 7389 582622 8389 582663
rect 8990 582622 9990 582663
rect 5169 574771 5191 581882
rect 2848 570723 2874 570757
rect 6005 569701 6021 581882
rect 29836 580009 29842 580483
rect 20779 576337 20783 577542
rect 29836 576963 29842 577411
rect 7389 570336 8389 570498
rect 8990 570359 9990 570499
rect 15678 569971 16678 570073
rect 17278 569971 18278 570073
rect 15678 569900 16678 569926
rect 17278 569900 18278 569926
rect 2848 569489 2874 569523
rect 19516 569409 19547 576333
rect 29952 575135 29955 580688
rect 30015 575954 30027 581677
rect 38946 580623 38954 580648
rect 38946 577413 38954 577439
rect 30015 575944 30721 575954
rect 30015 575928 30718 575944
rect 31823 573340 32061 573372
rect 31481 573320 31797 573338
rect 36071 572905 36098 573395
rect 31481 572120 31797 572132
rect 31481 572116 32061 572120
rect 31823 572082 32061 572116
rect 20809 570118 20821 570174
rect 14744 569235 19490 569383
rect 698110 562817 702856 562965
rect 696779 562026 696791 562082
rect 685539 560084 685777 560118
rect 685539 560080 686119 560084
rect 685803 560068 686119 560080
rect 681502 558805 681529 559295
rect 685803 558862 686119 558880
rect 685539 558828 685777 558860
rect 686882 556256 687585 556272
rect 686879 556246 687585 556256
rect 678646 554761 678654 554787
rect 678646 551552 678654 551577
rect 687573 550523 687585 556246
rect 687645 551512 687648 557065
rect 698053 555867 698084 562791
rect 714726 562677 714752 562711
rect 699322 562274 700322 562300
rect 700922 562274 701922 562300
rect 699322 562127 700322 562229
rect 700922 562127 701922 562229
rect 707610 561701 708610 561841
rect 709211 561702 710211 561864
rect 687758 554789 687764 555237
rect 696817 554658 696821 555863
rect 687758 551717 687764 552191
rect 711579 550318 711595 562499
rect 714726 561443 714752 561477
rect 712409 550318 712431 557429
rect 707610 549537 708610 549578
rect 709211 549537 710211 549578
rect 699322 548906 700322 549061
rect 700922 548906 701922 549061
rect 707610 548806 708610 549016
rect 709211 548806 710211 549016
rect 699322 548581 700322 548736
rect 700922 548581 701922 548736
rect 711579 548493 711605 550275
rect 711579 548483 711619 548493
rect 711579 548469 712463 548483
rect 5137 540517 6021 540531
rect 5981 540507 6021 540517
rect 5995 538725 6021 540507
rect 15678 540264 16678 540419
rect 17278 540264 18278 540419
rect 7389 539984 8389 540194
rect 8990 539984 9990 540194
rect 15678 539939 16678 540094
rect 17278 539939 18278 540094
rect 7389 539422 8389 539463
rect 8990 539422 9990 539463
rect 5169 531571 5191 538682
rect 2848 527523 2874 527557
rect 6005 526501 6021 538682
rect 29836 536809 29842 537283
rect 20779 533137 20783 534342
rect 29836 533763 29842 534211
rect 7389 527136 8389 527298
rect 8990 527159 9990 527299
rect 15678 526771 16678 526873
rect 17278 526771 18278 526873
rect 15678 526700 16678 526726
rect 17278 526700 18278 526726
rect 2848 526289 2874 526323
rect 19516 526209 19547 533133
rect 29952 531935 29955 537488
rect 30015 532754 30027 538477
rect 38946 537423 38954 537448
rect 38946 534213 38954 534239
rect 30015 532744 30721 532754
rect 30015 532728 30718 532744
rect 31823 530140 32061 530172
rect 31481 530120 31797 530138
rect 36071 529705 36098 530195
rect 31481 528920 31797 528932
rect 31481 528916 32061 528920
rect 31823 528882 32061 528916
rect 20809 526918 20821 526974
rect 14744 526035 19490 526183
rect 678282 471387 681670 471445
rect 678282 467471 681670 467485
rect 35930 448115 39318 448129
rect 35930 444155 39318 444213
rect 5137 412917 6021 412931
rect 5981 412907 6021 412917
rect 5995 411125 6021 412907
rect 15678 412664 16678 412819
rect 17278 412664 18278 412819
rect 7389 412384 8389 412594
rect 8990 412384 9990 412594
rect 15678 412339 16678 412494
rect 17278 412339 18278 412494
rect 7389 411822 8389 411863
rect 8990 411822 9990 411863
rect 5169 403971 5191 411082
rect 2848 399923 2874 399957
rect 6005 398901 6021 411082
rect 29836 409209 29842 409683
rect 20779 405537 20783 406742
rect 29836 406163 29842 406611
rect 7389 399536 8389 399698
rect 8990 399559 9990 399699
rect 15678 399171 16678 399273
rect 17278 399171 18278 399273
rect 15678 399100 16678 399126
rect 17278 399100 18278 399126
rect 2848 398689 2874 398723
rect 19516 398609 19547 405533
rect 29952 404335 29955 409888
rect 30015 405154 30027 410877
rect 38946 409823 38954 409848
rect 38946 406613 38954 406639
rect 30015 405144 30721 405154
rect 30015 405128 30718 405144
rect 31823 402540 32061 402572
rect 31481 402520 31797 402538
rect 36071 402105 36098 402595
rect 31481 401320 31797 401332
rect 31481 401316 32061 401320
rect 31823 401282 32061 401316
rect 20809 399318 20821 399374
rect 14744 398435 19490 398583
rect 698110 385617 702856 385765
rect 696779 384826 696791 384882
rect 685539 382884 685777 382918
rect 685539 382880 686119 382884
rect 685803 382868 686119 382880
rect 681502 381605 681529 382095
rect 685803 381662 686119 381680
rect 685539 381628 685777 381660
rect 686882 379056 687585 379072
rect 686879 379046 687585 379056
rect 678646 377561 678654 377587
rect 678646 374352 678654 374377
rect 687573 373323 687585 379046
rect 687645 374312 687648 379865
rect 698053 378667 698084 385591
rect 714726 385477 714752 385511
rect 699322 385074 700322 385100
rect 700922 385074 701922 385100
rect 699322 384927 700322 385029
rect 700922 384927 701922 385029
rect 707610 384501 708610 384641
rect 709211 384502 710211 384664
rect 687758 377589 687764 378037
rect 696817 377458 696821 378663
rect 687758 374517 687764 374991
rect 711579 373118 711595 385299
rect 714726 384243 714752 384277
rect 712409 373118 712431 380229
rect 707610 372337 708610 372378
rect 709211 372337 710211 372378
rect 699322 371706 700322 371861
rect 700922 371706 701922 371861
rect 707610 371606 708610 371816
rect 709211 371606 710211 371816
rect 699322 371381 700322 371536
rect 700922 371381 701922 371536
rect 711579 371293 711605 373075
rect 711579 371283 711619 371293
rect 711579 371269 712463 371283
rect 5137 369717 6021 369731
rect 5981 369707 6021 369717
rect 5995 367925 6021 369707
rect 15678 369464 16678 369619
rect 17278 369464 18278 369619
rect 7389 369184 8389 369394
rect 8990 369184 9990 369394
rect 15678 369139 16678 369294
rect 17278 369139 18278 369294
rect 7389 368622 8389 368663
rect 8990 368622 9990 368663
rect 5169 360771 5191 367882
rect 2848 356723 2874 356757
rect 6005 355701 6021 367882
rect 29836 366009 29842 366483
rect 20779 362337 20783 363542
rect 29836 362963 29842 363411
rect 7389 356336 8389 356498
rect 8990 356359 9990 356499
rect 15678 355971 16678 356073
rect 17278 355971 18278 356073
rect 15678 355900 16678 355926
rect 17278 355900 18278 355926
rect 2848 355489 2874 355523
rect 19516 355409 19547 362333
rect 29952 361135 29955 366688
rect 30015 361954 30027 367677
rect 38946 366623 38954 366648
rect 38946 363413 38954 363439
rect 30015 361944 30721 361954
rect 30015 361928 30718 361944
rect 31823 359340 32061 359372
rect 31481 359320 31797 359338
rect 36071 358905 36098 359395
rect 31481 358120 31797 358132
rect 31481 358116 32061 358120
rect 31823 358082 32061 358116
rect 20809 356118 20821 356174
rect 14744 355235 19490 355383
rect 698110 340417 702856 340565
rect 696779 339626 696791 339682
rect 685539 337684 685777 337718
rect 685539 337680 686119 337684
rect 685803 337668 686119 337680
rect 681502 336405 681529 336895
rect 685803 336462 686119 336480
rect 685539 336428 685777 336460
rect 686882 333856 687585 333872
rect 686879 333846 687585 333856
rect 678646 332361 678654 332387
rect 678646 329152 678654 329177
rect 687573 328123 687585 333846
rect 687645 329112 687648 334665
rect 698053 333467 698084 340391
rect 714726 340277 714752 340311
rect 699322 339874 700322 339900
rect 700922 339874 701922 339900
rect 699322 339727 700322 339829
rect 700922 339727 701922 339829
rect 707610 339301 708610 339441
rect 709211 339302 710211 339464
rect 687758 332389 687764 332837
rect 696817 332258 696821 333463
rect 687758 329317 687764 329791
rect 711579 327918 711595 340099
rect 714726 339043 714752 339077
rect 712409 327918 712431 335029
rect 707610 327137 708610 327178
rect 709211 327137 710211 327178
rect 5137 326517 6021 326531
rect 5981 326507 6021 326517
rect 5995 324725 6021 326507
rect 699322 326506 700322 326661
rect 700922 326506 701922 326661
rect 15678 326264 16678 326419
rect 17278 326264 18278 326419
rect 707610 326406 708610 326616
rect 709211 326406 710211 326616
rect 7389 325984 8389 326194
rect 8990 325984 9990 326194
rect 699322 326181 700322 326336
rect 700922 326181 701922 326336
rect 15678 325939 16678 326094
rect 17278 325939 18278 326094
rect 711579 326093 711605 327875
rect 711579 326083 711619 326093
rect 711579 326069 712463 326083
rect 7389 325422 8389 325463
rect 8990 325422 9990 325463
rect 5169 317571 5191 324682
rect 2848 313523 2874 313557
rect 6005 312501 6021 324682
rect 29836 322809 29842 323283
rect 20779 319137 20783 320342
rect 29836 319763 29842 320211
rect 7389 313136 8389 313298
rect 8990 313159 9990 313299
rect 15678 312771 16678 312873
rect 17278 312771 18278 312873
rect 15678 312700 16678 312726
rect 17278 312700 18278 312726
rect 2848 312289 2874 312323
rect 19516 312209 19547 319133
rect 29952 317935 29955 323488
rect 30015 318754 30027 324477
rect 38946 323423 38954 323448
rect 38946 320213 38954 320239
rect 30015 318744 30721 318754
rect 30015 318728 30718 318744
rect 31823 316140 32061 316172
rect 31481 316120 31797 316138
rect 36071 315705 36098 316195
rect 31481 314920 31797 314932
rect 31481 314916 32061 314920
rect 31823 314882 32061 314916
rect 20809 312918 20821 312974
rect 14744 312035 19490 312183
rect 698110 295417 702856 295565
rect 696779 294626 696791 294682
rect 685539 292684 685777 292718
rect 685539 292680 686119 292684
rect 685803 292668 686119 292680
rect 681502 291405 681529 291895
rect 685803 291462 686119 291480
rect 685539 291428 685777 291460
rect 686882 288856 687585 288872
rect 686879 288846 687585 288856
rect 678646 287361 678654 287387
rect 678646 284152 678654 284177
rect 5137 283317 6021 283331
rect 5981 283307 6021 283317
rect 5995 281525 6021 283307
rect 15678 283064 16678 283219
rect 17278 283064 18278 283219
rect 687573 283123 687585 288846
rect 687645 284112 687648 289665
rect 698053 288467 698084 295391
rect 714726 295277 714752 295311
rect 699322 294874 700322 294900
rect 700922 294874 701922 294900
rect 699322 294727 700322 294829
rect 700922 294727 701922 294829
rect 707610 294301 708610 294441
rect 709211 294302 710211 294464
rect 687758 287389 687764 287837
rect 696817 287258 696821 288463
rect 687758 284317 687764 284791
rect 7389 282784 8389 282994
rect 8990 282784 9990 282994
rect 711579 282918 711595 295099
rect 714726 294043 714752 294077
rect 712409 282918 712431 290029
rect 15678 282739 16678 282894
rect 17278 282739 18278 282894
rect 7389 282222 8389 282263
rect 8990 282222 9990 282263
rect 707610 282137 708610 282178
rect 709211 282137 710211 282178
rect 699322 281506 700322 281661
rect 700922 281506 701922 281661
rect 5169 274371 5191 281482
rect 2848 270323 2874 270357
rect 6005 269301 6021 281482
rect 707610 281406 708610 281616
rect 709211 281406 710211 281616
rect 29836 279609 29842 280083
rect 20779 275937 20783 277142
rect 29836 276563 29842 277011
rect 7389 269936 8389 270098
rect 8990 269959 9990 270099
rect 15678 269571 16678 269673
rect 17278 269571 18278 269673
rect 15678 269500 16678 269526
rect 17278 269500 18278 269526
rect 2848 269089 2874 269123
rect 19516 269009 19547 275933
rect 29952 274735 29955 280288
rect 30015 275554 30027 281277
rect 699322 281181 700322 281336
rect 700922 281181 701922 281336
rect 711579 281093 711605 282875
rect 711579 281083 711619 281093
rect 711579 281069 712463 281083
rect 38946 280223 38954 280248
rect 38946 277013 38954 277039
rect 30015 275544 30721 275554
rect 30015 275528 30718 275544
rect 31823 272940 32061 272972
rect 31481 272920 31797 272938
rect 36071 272505 36098 272995
rect 31481 271720 31797 271732
rect 31481 271716 32061 271720
rect 31823 271682 32061 271716
rect 20809 269718 20821 269774
rect 14744 268835 19490 268983
rect 698110 250417 702856 250565
rect 696779 249626 696791 249682
rect 685539 247684 685777 247718
rect 685539 247680 686119 247684
rect 685803 247668 686119 247680
rect 681502 246405 681529 246895
rect 685803 246462 686119 246480
rect 685539 246428 685777 246460
rect 686882 243856 687585 243872
rect 686879 243846 687585 243856
rect 678646 242361 678654 242387
rect 5137 240117 6021 240131
rect 5981 240107 6021 240117
rect 5995 238325 6021 240107
rect 15678 239864 16678 240019
rect 17278 239864 18278 240019
rect 7389 239584 8389 239794
rect 8990 239584 9990 239794
rect 15678 239539 16678 239694
rect 17278 239539 18278 239694
rect 678646 239152 678654 239177
rect 7389 239022 8389 239063
rect 8990 239022 9990 239063
rect 5169 231171 5191 238282
rect 2848 227123 2874 227157
rect 6005 226101 6021 238282
rect 687573 238123 687585 243846
rect 687645 239112 687648 244665
rect 698053 243467 698084 250391
rect 714726 250277 714752 250311
rect 699322 249874 700322 249900
rect 700922 249874 701922 249900
rect 699322 249727 700322 249829
rect 700922 249727 701922 249829
rect 707610 249301 708610 249441
rect 709211 249302 710211 249464
rect 687758 242389 687764 242837
rect 696817 242258 696821 243463
rect 687758 239317 687764 239791
rect 29836 236409 29842 236883
rect 20779 232737 20783 233942
rect 29836 233363 29842 233811
rect 7389 226736 8389 226898
rect 8990 226759 9990 226899
rect 15678 226371 16678 226473
rect 17278 226371 18278 226473
rect 15678 226300 16678 226326
rect 17278 226300 18278 226326
rect 2848 225889 2874 225923
rect 19516 225809 19547 232733
rect 29952 231535 29955 237088
rect 30015 232354 30027 238077
rect 711579 237918 711595 250099
rect 714726 249043 714752 249077
rect 712409 237918 712431 245029
rect 707610 237137 708610 237178
rect 709211 237137 710211 237178
rect 38946 237023 38954 237048
rect 699322 236506 700322 236661
rect 700922 236506 701922 236661
rect 707610 236406 708610 236616
rect 709211 236406 710211 236616
rect 699322 236181 700322 236336
rect 700922 236181 701922 236336
rect 711579 236093 711605 237875
rect 711579 236083 711619 236093
rect 711579 236069 712463 236083
rect 38946 233813 38954 233839
rect 30015 232344 30721 232354
rect 30015 232328 30718 232344
rect 31823 229740 32061 229772
rect 31481 229720 31797 229738
rect 36071 229305 36098 229795
rect 31481 228520 31797 228532
rect 31481 228516 32061 228520
rect 31823 228482 32061 228516
rect 20809 226518 20821 226574
rect 14744 225635 19490 225783
rect 698110 205217 702856 205365
rect 696779 204426 696791 204482
rect 685539 202484 685777 202518
rect 685539 202480 686119 202484
rect 685803 202468 686119 202480
rect 681502 201205 681529 201695
rect 685803 201262 686119 201280
rect 685539 201228 685777 201260
rect 686882 198656 687585 198672
rect 686879 198646 687585 198656
rect 678646 197161 678654 197187
rect 5137 196917 6021 196931
rect 5981 196907 6021 196917
rect 5995 195125 6021 196907
rect 15678 196664 16678 196819
rect 17278 196664 18278 196819
rect 7389 196384 8389 196594
rect 8990 196384 9990 196594
rect 15678 196339 16678 196494
rect 17278 196339 18278 196494
rect 7389 195822 8389 195863
rect 8990 195822 9990 195863
rect 5169 187971 5191 195082
rect 2848 183923 2874 183957
rect 6005 182901 6021 195082
rect 29836 193209 29842 193683
rect 20779 189537 20783 190742
rect 29836 190163 29842 190611
rect 7389 183536 8389 183698
rect 8990 183559 9990 183699
rect 15678 183171 16678 183273
rect 17278 183171 18278 183273
rect 15678 183100 16678 183126
rect 17278 183100 18278 183126
rect 2848 182689 2874 182723
rect 19516 182609 19547 189533
rect 29952 188335 29955 193888
rect 30015 189154 30027 194877
rect 678646 193952 678654 193977
rect 38946 193823 38954 193848
rect 687573 192923 687585 198646
rect 687645 193912 687648 199465
rect 698053 198267 698084 205191
rect 714726 205077 714752 205111
rect 699322 204674 700322 204700
rect 700922 204674 701922 204700
rect 699322 204527 700322 204629
rect 700922 204527 701922 204629
rect 707610 204101 708610 204241
rect 709211 204102 710211 204264
rect 687758 197189 687764 197637
rect 696817 197058 696821 198263
rect 687758 194117 687764 194591
rect 711579 192718 711595 204899
rect 714726 203843 714752 203877
rect 712409 192718 712431 199829
rect 707610 191937 708610 191978
rect 709211 191937 710211 191978
rect 699322 191306 700322 191461
rect 700922 191306 701922 191461
rect 707610 191206 708610 191416
rect 709211 191206 710211 191416
rect 699322 190981 700322 191136
rect 700922 190981 701922 191136
rect 711579 190893 711605 192675
rect 711579 190883 711619 190893
rect 711579 190869 712463 190883
rect 38946 190613 38954 190639
rect 30015 189144 30721 189154
rect 30015 189128 30718 189144
rect 31823 186540 32061 186572
rect 31481 186520 31797 186538
rect 36071 186105 36098 186595
rect 31481 185320 31797 185332
rect 31481 185316 32061 185320
rect 31823 185282 32061 185316
rect 20809 183318 20821 183374
rect 14744 182435 19490 182583
rect 698110 160217 702856 160365
rect 696779 159426 696791 159482
rect 685539 157484 685777 157518
rect 685539 157480 686119 157484
rect 685803 157468 686119 157480
rect 681502 156205 681529 156695
rect 685803 156262 686119 156280
rect 685539 156228 685777 156260
rect 686882 153656 687585 153672
rect 686879 153646 687585 153656
rect 678646 152161 678654 152187
rect 678646 148952 678654 148977
rect 687573 147923 687585 153646
rect 687645 148912 687648 154465
rect 698053 153267 698084 160191
rect 714726 160077 714752 160111
rect 699322 159674 700322 159700
rect 700922 159674 701922 159700
rect 699322 159527 700322 159629
rect 700922 159527 701922 159629
rect 707610 159101 708610 159241
rect 709211 159102 710211 159264
rect 687758 152189 687764 152637
rect 696817 152058 696821 153263
rect 687758 149117 687764 149591
rect 711579 147718 711595 159899
rect 714726 158843 714752 158877
rect 712409 147718 712431 154829
rect 707610 146937 708610 146978
rect 709211 146937 710211 146978
rect 699322 146306 700322 146461
rect 700922 146306 701922 146461
rect 707610 146206 708610 146416
rect 709211 146206 710211 146416
rect 699322 145981 700322 146136
rect 700922 145981 701922 146136
rect 711579 145893 711605 147675
rect 711579 145883 711619 145893
rect 711579 145869 712463 145883
rect 698110 115017 702856 115165
rect 696779 114226 696791 114282
rect 685539 112284 685777 112318
rect 685539 112280 686119 112284
rect 685803 112268 686119 112280
rect 681502 111005 681529 111495
rect 685803 111062 686119 111080
rect 685539 111028 685777 111060
rect 686882 108456 687585 108472
rect 686879 108446 687585 108456
rect 678646 106961 678654 106987
rect 678646 103752 678654 103777
rect 687573 102723 687585 108446
rect 687645 103712 687648 109265
rect 698053 108067 698084 114991
rect 714726 114877 714752 114911
rect 699322 114474 700322 114500
rect 700922 114474 701922 114500
rect 699322 114327 700322 114429
rect 700922 114327 701922 114429
rect 707610 113901 708610 114041
rect 709211 113902 710211 114064
rect 687758 106989 687764 107437
rect 696817 106858 696821 108063
rect 687758 103917 687764 104391
rect 711579 102518 711595 114699
rect 714726 113643 714752 113677
rect 712409 102518 712431 109629
rect 707610 101737 708610 101778
rect 709211 101737 710211 101778
rect 699322 101106 700322 101261
rect 700922 101106 701922 101261
rect 707610 101006 708610 101216
rect 709211 101006 710211 101216
rect 699322 100781 700322 100936
rect 700922 100781 701922 100936
rect 711579 100693 711605 102475
rect 711579 100683 711619 100693
rect 711579 100669 712463 100683
rect 35930 75315 39318 75329
rect 35930 71355 39318 71413
rect 190152 38946 190177 38954
rect 193361 38946 193387 38954
rect 146187 38280 146453 38291
rect 144718 36866 144738 37390
rect 197405 36071 197895 36098
rect 248871 35930 248885 39318
rect 252787 35930 252845 39318
rect 298752 38946 298777 38954
rect 301961 38946 301987 38954
rect 353552 38946 353577 38954
rect 356761 38946 356787 38954
rect 408352 38946 408377 38954
rect 411561 38946 411587 38954
rect 463152 38946 463177 38954
rect 466361 38946 466387 38954
rect 517952 38946 517977 38954
rect 521161 38946 521187 38954
rect 306005 36071 306495 36098
rect 360805 36071 361295 36098
rect 415605 36071 416095 36098
rect 470405 36071 470895 36098
rect 525205 36071 525695 36098
rect 143407 35902 143463 35923
rect 143407 35793 143429 35902
rect 197428 31823 197460 32061
rect 198680 31823 198718 32061
rect 306028 31823 306060 32061
rect 307280 31823 307318 32061
rect 360828 31823 360860 32061
rect 362080 31823 362118 32061
rect 415628 31823 415660 32061
rect 416880 31823 416918 32061
rect 470428 31823 470460 32061
rect 471680 31823 471718 32061
rect 525228 31823 525260 32061
rect 526480 31823 526518 32061
rect 198680 31797 198684 31823
rect 307280 31797 307284 31823
rect 362080 31797 362084 31823
rect 416880 31797 416884 31823
rect 471680 31797 471684 31823
rect 526480 31797 526484 31823
rect 197462 31481 197480 31797
rect 198668 31481 198684 31797
rect 306062 31481 306080 31797
rect 307268 31481 307284 31797
rect 360862 31481 360880 31797
rect 362068 31481 362084 31797
rect 415662 31481 415680 31797
rect 416868 31481 416884 31797
rect 470462 31481 470480 31797
rect 471668 31481 471684 31797
rect 525262 31481 525280 31797
rect 526468 31481 526484 31797
rect 194846 30718 194856 30721
rect 303446 30718 303456 30721
rect 358246 30718 358256 30721
rect 413046 30718 413056 30721
rect 467846 30718 467856 30721
rect 522646 30718 522656 30721
rect 194846 30027 194872 30718
rect 303446 30027 303472 30718
rect 358246 30027 358272 30718
rect 413046 30027 413072 30718
rect 467846 30027 467872 30718
rect 522646 30027 522672 30718
rect 189123 30015 194872 30027
rect 297723 30015 303472 30027
rect 352523 30015 358272 30027
rect 407323 30015 413072 30027
rect 462123 30015 467872 30027
rect 516923 30015 522672 30027
rect 190112 29952 195665 29955
rect 298712 29952 304265 29955
rect 353512 29952 359065 29955
rect 408312 29952 413865 29955
rect 463112 29952 468665 29955
rect 517912 29952 523465 29955
rect 190317 29836 190791 29842
rect 193389 29836 193837 29842
rect 298917 29836 299391 29842
rect 301989 29836 302437 29842
rect 353717 29836 354191 29842
rect 356789 29836 357237 29842
rect 408517 29836 408991 29842
rect 411589 29836 412037 29842
rect 463317 29836 463791 29842
rect 466389 29836 466837 29842
rect 518117 29836 518591 29842
rect 521189 29836 521637 29842
rect 200626 20809 200682 20821
rect 309226 20809 309282 20821
rect 364026 20809 364082 20821
rect 418826 20809 418882 20821
rect 473626 20809 473682 20821
rect 528426 20809 528482 20821
rect 193258 20779 194463 20783
rect 301858 20779 303063 20783
rect 356658 20779 357863 20783
rect 411458 20779 412663 20783
rect 466258 20779 467463 20783
rect 521058 20779 522263 20783
rect 147509 19547 147573 19618
rect 194467 19516 201391 19547
rect 303067 19516 309991 19547
rect 357867 19516 364791 19547
rect 412667 19516 419591 19547
rect 467467 19516 474391 19547
rect 522267 19516 529191 19547
rect 133241 17478 133396 18478
rect 133566 17478 133721 18478
rect 146787 17478 146889 18478
rect 146934 17478 146960 18478
rect 187181 17278 187336 18278
rect 187506 17278 187661 18278
rect 200727 17278 200829 18278
rect 200874 17278 200900 18278
rect 133241 15878 133396 16878
rect 133566 15878 133721 16878
rect 146787 15878 146889 16878
rect 146934 15878 146960 16878
rect 187181 15678 187336 16678
rect 187506 15678 187661 16678
rect 200727 15678 200829 16678
rect 200874 15678 200900 16678
rect 201417 14744 201565 19490
rect 295781 17278 295936 18278
rect 296106 17278 296261 18278
rect 309327 17278 309429 18278
rect 309474 17278 309500 18278
rect 295781 15678 295936 16678
rect 296106 15678 296261 16678
rect 309327 15678 309429 16678
rect 309474 15678 309500 16678
rect 310017 14744 310165 19490
rect 350581 17278 350736 18278
rect 350906 17278 351061 18278
rect 364127 17278 364229 18278
rect 364274 17278 364300 18278
rect 350581 15678 350736 16678
rect 350906 15678 351061 16678
rect 364127 15678 364229 16678
rect 364274 15678 364300 16678
rect 364817 14744 364965 19490
rect 405381 17278 405536 18278
rect 405706 17278 405861 18278
rect 418927 17278 419029 18278
rect 419074 17278 419100 18278
rect 405381 15678 405536 16678
rect 405706 15678 405861 16678
rect 418927 15678 419029 16678
rect 419074 15678 419100 16678
rect 419617 14744 419765 19490
rect 460181 17278 460336 18278
rect 460506 17278 460661 18278
rect 473727 17278 473829 18278
rect 473874 17278 473900 18278
rect 460181 15678 460336 16678
rect 460506 15678 460661 16678
rect 473727 15678 473829 16678
rect 473874 15678 473900 16678
rect 474417 14744 474565 19490
rect 514981 17278 515136 18278
rect 515306 17278 515461 18278
rect 528527 17278 528629 18278
rect 528674 17278 528700 18278
rect 514981 15678 515136 16678
rect 515306 15678 515461 16678
rect 528527 15678 528629 16678
rect 528674 15678 528700 16678
rect 529217 14744 529365 19490
rect 133606 8990 133816 9990
rect 134337 8990 134378 9990
rect 146501 8990 146641 9990
rect 187406 8990 187616 9990
rect 188137 8990 188178 9990
rect 200301 8990 200441 9990
rect 296006 8990 296216 9990
rect 296737 8990 296778 9990
rect 308901 8990 309041 9990
rect 350806 8990 351016 9990
rect 351537 8990 351578 9990
rect 363701 8990 363841 9990
rect 405606 8990 405816 9990
rect 406337 8990 406378 9990
rect 418501 8990 418641 9990
rect 460406 8990 460616 9990
rect 461137 8990 461178 9990
rect 473301 8990 473441 9990
rect 515206 8990 515416 9990
rect 515937 8990 515978 9990
rect 528101 8990 528241 9990
rect 133606 7389 133816 8389
rect 134337 7389 134378 8389
rect 146502 7389 146664 8389
rect 187406 7389 187616 8389
rect 188137 7389 188178 8389
rect 200302 7389 200464 8389
rect 296006 7389 296216 8389
rect 296737 7389 296778 8389
rect 308902 7389 309064 8389
rect 350806 7389 351016 8389
rect 351537 7389 351578 8389
rect 363702 7389 363864 8389
rect 405606 7389 405816 8389
rect 406337 7389 406378 8389
rect 418502 7389 418664 8389
rect 460406 7389 460616 8389
rect 461137 7389 461178 8389
rect 473302 7389 473464 8389
rect 515206 7389 515416 8389
rect 515937 7389 515978 8389
rect 528102 7389 528264 8389
rect 187069 5995 188875 6021
rect 188918 6005 201099 6021
rect 295669 5995 297475 6021
rect 297518 6005 309699 6021
rect 350469 5995 352275 6021
rect 352318 6005 364499 6021
rect 405269 5995 407075 6021
rect 407118 6005 419299 6021
rect 460069 5995 461875 6021
rect 461918 6005 474099 6021
rect 514869 5995 516675 6021
rect 516718 6005 528899 6021
rect 187069 5981 187093 5995
rect 295669 5981 295693 5995
rect 350469 5981 350493 5995
rect 405269 5981 405293 5995
rect 460069 5981 460093 5995
rect 514869 5981 514893 5995
rect 187069 5137 187083 5981
rect 188918 5169 196029 5191
rect 295669 5137 295683 5981
rect 297518 5169 304629 5191
rect 350469 5137 350483 5981
rect 352318 5169 359429 5191
rect 405269 5137 405283 5981
rect 407118 5169 414229 5191
rect 460069 5137 460083 5981
rect 461918 5169 469029 5191
rect 514869 5137 514883 5981
rect 516718 5169 523829 5191
rect 200043 2848 200077 2874
rect 201277 2848 201311 2874
rect 308643 2848 308677 2874
rect 309877 2848 309911 2874
rect 363443 2848 363477 2874
rect 364677 2848 364711 2874
rect 418243 2848 418277 2874
rect 419477 2848 419511 2874
rect 473043 2848 473077 2874
rect 474277 2848 474311 2874
rect 527843 2848 527877 2874
rect 529077 2848 529111 2874
<< metal1 >>
rect 84010 995596 84016 995648
rect 84068 995636 84074 995648
rect 91738 995636 91744 995648
rect 84068 995608 91744 995636
rect 84068 995596 84074 995608
rect 91738 995596 91744 995608
rect 91796 995596 91802 995648
rect 238202 995596 238208 995648
rect 238260 995636 238266 995648
rect 245930 995636 245936 995648
rect 238260 995608 245936 995636
rect 238260 995596 238266 995608
rect 245930 995596 245936 995608
rect 245988 995596 245994 995648
rect 531958 995596 531964 995648
rect 532016 995636 532022 995648
rect 539686 995636 539692 995648
rect 532016 995608 539692 995636
rect 532016 995596 532022 995608
rect 539686 995596 539692 995608
rect 539744 995596 539750 995648
rect 135346 995460 135352 995512
rect 135404 995500 135410 995512
rect 143166 995500 143172 995512
rect 135404 995472 143172 995500
rect 135404 995460 135410 995472
rect 143166 995460 143172 995472
rect 143224 995460 143230 995512
rect 633802 995460 633808 995512
rect 633860 995500 633866 995512
rect 641530 995500 641536 995512
rect 633860 995472 641536 995500
rect 633860 995460 633866 995472
rect 641530 995460 641536 995472
rect 641588 995460 641594 995512
rect 289630 995256 289636 995308
rect 289688 995296 289694 995308
rect 297634 995296 297640 995308
rect 289688 995268 297640 995296
rect 289688 995256 289694 995268
rect 297634 995256 297640 995268
rect 297692 995256 297698 995308
rect 391474 995256 391480 995308
rect 391532 995296 391538 995308
rect 399478 995296 399484 995308
rect 391532 995268 399484 995296
rect 391532 995256 391538 995268
rect 399478 995256 399484 995268
rect 399536 995256 399542 995308
rect 480438 995256 480444 995308
rect 480496 995296 480502 995308
rect 488442 995296 488448 995308
rect 480496 995268 488448 995296
rect 480496 995256 480502 995268
rect 488442 995256 488448 995268
rect 488500 995256 488506 995308
rect 231854 995052 231860 995104
rect 231912 995092 231918 995104
rect 244182 995092 244188 995104
rect 231912 995064 244188 995092
rect 231912 995052 231918 995064
rect 244182 995052 244188 995064
rect 244240 995052 244246 995104
rect 463786 992264 463792 992316
rect 463844 992304 463850 992316
rect 475470 992304 475476 992316
rect 463844 992276 475476 992304
rect 463844 992264 463850 992276
rect 475470 992264 475476 992276
rect 475528 992304 475534 992316
rect 482922 992304 482928 992316
rect 475528 992276 482928 992304
rect 475528 992264 475534 992276
rect 482922 992264 482928 992276
rect 482980 992264 482986 992316
rect 141418 992060 141424 992112
rect 141476 992100 141482 992112
rect 154390 992100 154396 992112
rect 141476 992072 154396 992100
rect 141476 992060 141482 992072
rect 154390 992060 154396 992072
rect 154448 992060 154454 992112
rect 130286 990876 130292 990888
rect 130120 990848 130292 990876
rect 130120 990820 130148 990848
rect 130286 990836 130292 990848
rect 130344 990876 130350 990888
rect 130344 990848 130424 990876
rect 130344 990836 130350 990848
rect 79042 990768 79048 990820
rect 79100 990808 79106 990820
rect 110414 990808 110420 990820
rect 79100 990780 110420 990808
rect 79100 990768 79106 990780
rect 110414 990768 110420 990780
rect 110472 990768 110478 990820
rect 130102 990768 130108 990820
rect 130160 990768 130166 990820
rect 130396 990808 130424 990848
rect 419534 990836 419540 990888
rect 419592 990876 419598 990888
rect 438670 990876 438676 990888
rect 419592 990848 438676 990876
rect 419592 990836 419598 990848
rect 438670 990836 438676 990848
rect 438728 990836 438734 990888
rect 450262 990836 450268 990888
rect 450320 990876 450326 990888
rect 463602 990876 463608 990888
rect 450320 990848 463608 990876
rect 450320 990836 450326 990848
rect 463602 990836 463608 990848
rect 463660 990836 463666 990888
rect 143258 990808 143264 990820
rect 130396 990780 143264 990808
rect 143258 990768 143264 990780
rect 143316 990768 143322 990820
rect 173802 990768 173808 990820
rect 173860 990808 173866 990820
rect 179322 990808 179328 990820
rect 173860 990780 179328 990808
rect 173860 990768 173866 990780
rect 179322 990768 179328 990780
rect 179380 990768 179386 990820
rect 246942 990768 246948 990820
rect 247000 990808 247006 990820
rect 284662 990808 284668 990820
rect 247000 990780 284668 990808
rect 247000 990768 247006 990780
rect 284662 990768 284668 990780
rect 284720 990808 284726 990820
rect 286962 990808 286968 990820
rect 284720 990780 286968 990808
rect 284720 990768 284726 990780
rect 286962 990768 286968 990780
rect 287020 990768 287026 990820
rect 391750 990768 391756 990820
rect 391808 990808 391814 990820
rect 476114 990808 476120 990820
rect 391808 990780 476120 990808
rect 391808 990768 391814 990780
rect 476114 990768 476120 990780
rect 476172 990808 476178 990820
rect 527542 990808 527548 990820
rect 476172 990780 527548 990808
rect 476172 990768 476178 990780
rect 527542 990768 527548 990780
rect 527600 990808 527606 990820
rect 629294 990808 629300 990820
rect 527600 990780 629300 990808
rect 527600 990768 527606 990780
rect 629294 990768 629300 990780
rect 629352 990768 629358 990820
rect 187602 990700 187608 990752
rect 187660 990740 187666 990752
rect 187694 990740 187700 990752
rect 187660 990712 187700 990740
rect 187660 990700 187666 990712
rect 187694 990700 187700 990712
rect 187752 990700 187758 990752
rect 202874 990700 202880 990752
rect 202932 990740 202938 990752
rect 233050 990740 233056 990752
rect 202932 990712 233056 990740
rect 202932 990700 202938 990712
rect 233050 990700 233056 990712
rect 233108 990700 233114 990752
rect 244182 990700 244188 990752
rect 244240 990740 244246 990752
rect 295794 990740 295800 990752
rect 244240 990712 295800 990740
rect 244240 990700 244246 990712
rect 295794 990700 295800 990712
rect 295852 990740 295858 990752
rect 386322 990740 386328 990752
rect 295852 990712 386328 990740
rect 295852 990700 295858 990712
rect 386322 990700 386328 990712
rect 386380 990700 386386 990752
rect 482922 990700 482928 990752
rect 482980 990740 482986 990752
rect 526898 990740 526904 990752
rect 482980 990712 526904 990740
rect 482980 990700 482986 990712
rect 526898 990700 526904 990712
rect 526956 990740 526962 990752
rect 628650 990740 628656 990752
rect 526956 990712 628656 990740
rect 526956 990700 526962 990712
rect 628650 990700 628656 990712
rect 628708 990700 628714 990752
rect 79502 990632 79508 990684
rect 79560 990672 79566 990684
rect 79962 990672 79968 990684
rect 79560 990644 79968 990672
rect 79560 990632 79566 990644
rect 79962 990632 79968 990644
rect 80020 990672 80026 990684
rect 130930 990672 130936 990684
rect 80020 990644 130936 990672
rect 80020 990632 80026 990644
rect 130930 990632 130936 990644
rect 130988 990672 130994 990684
rect 182358 990672 182364 990684
rect 130988 990644 182364 990672
rect 130988 990632 130994 990644
rect 182358 990632 182364 990644
rect 182416 990672 182422 990684
rect 233694 990672 233700 990684
rect 182416 990644 233700 990672
rect 182416 990632 182422 990644
rect 233694 990632 233700 990644
rect 233752 990672 233758 990684
rect 285306 990672 285312 990684
rect 233752 990644 285312 990672
rect 233752 990632 233758 990644
rect 285306 990632 285312 990644
rect 285364 990672 285370 990684
rect 333514 990672 333520 990684
rect 285364 990644 333520 990672
rect 285364 990632 285370 990644
rect 333514 990632 333520 990644
rect 333572 990672 333578 990684
rect 387150 990672 387156 990684
rect 333572 990644 387156 990672
rect 333572 990632 333578 990644
rect 387150 990632 387156 990644
rect 387208 990672 387214 990684
rect 391750 990672 391756 990684
rect 387208 990644 391756 990672
rect 387208 990632 387214 990644
rect 391750 990632 391756 990644
rect 391808 990632 391814 990684
rect 391860 990644 405596 990672
rect 89990 990564 89996 990616
rect 90048 990604 90054 990616
rect 90048 990576 91140 990604
rect 90048 990564 90054 990576
rect 91112 990536 91140 990576
rect 110506 990564 110512 990616
rect 110564 990604 110570 990616
rect 130102 990604 130108 990616
rect 110564 990576 130108 990604
rect 110564 990564 110570 990576
rect 130102 990564 130108 990576
rect 130160 990564 130166 990616
rect 179322 990564 179328 990616
rect 179380 990604 179386 990616
rect 181714 990604 181720 990616
rect 179380 990576 181720 990604
rect 179380 990564 179386 990576
rect 181714 990564 181720 990576
rect 181772 990564 181778 990616
rect 186682 990564 186688 990616
rect 186740 990604 186746 990616
rect 194686 990604 194692 990616
rect 186740 990576 194692 990604
rect 186740 990564 186746 990576
rect 194686 990564 194692 990576
rect 194744 990564 194750 990616
rect 386506 990604 386512 990616
rect 386419 990576 386512 990604
rect 386506 990564 386512 990576
rect 386564 990604 386570 990616
rect 391860 990604 391888 990644
rect 386564 990576 391888 990604
rect 386564 990564 386570 990576
rect 91112 990508 110368 990536
rect 110340 990468 110368 990508
rect 164142 990496 164148 990548
rect 164200 990536 164206 990548
rect 192846 990536 192852 990548
rect 164200 990508 192852 990536
rect 164200 990496 164206 990508
rect 192846 990496 192852 990508
rect 192904 990536 192910 990548
rect 193214 990536 193220 990548
rect 192904 990508 193220 990536
rect 192904 990496 192910 990508
rect 193214 990496 193220 990508
rect 193272 990496 193278 990548
rect 212442 990496 212448 990548
rect 212500 990536 212506 990548
rect 231854 990536 231860 990548
rect 212500 990508 231860 990536
rect 212500 990496 212506 990508
rect 231854 990496 231860 990508
rect 231912 990496 231918 990548
rect 286962 990496 286968 990548
rect 287020 990536 287026 990548
rect 386524 990536 386552 990564
rect 287020 990508 386552 990536
rect 405568 990536 405596 990644
rect 596082 990632 596088 990684
rect 596140 990672 596146 990684
rect 596140 990644 598980 990672
rect 596140 990632 596146 990644
rect 419534 990604 419540 990616
rect 405752 990576 419540 990604
rect 405752 990536 405780 990576
rect 419534 990564 419540 990576
rect 419592 990564 419598 990616
rect 438762 990564 438768 990616
rect 438820 990604 438826 990616
rect 450262 990604 450268 990616
rect 438820 990576 450268 990604
rect 438820 990564 438826 990576
rect 450262 990564 450268 990576
rect 450320 990564 450326 990616
rect 469306 990564 469312 990616
rect 469364 990604 469370 990616
rect 576854 990604 576860 990616
rect 469364 990576 483060 990604
rect 469364 990564 469370 990576
rect 483032 990548 483060 990576
rect 565740 990576 576860 990604
rect 469030 990536 469036 990548
rect 405568 990508 405780 990536
rect 449820 990508 469036 990536
rect 287020 990496 287026 990508
rect 141326 990468 141332 990480
rect 110340 990440 141332 990468
rect 141326 990428 141332 990440
rect 141384 990428 141390 990480
rect 143258 990428 143264 990480
rect 143316 990468 143322 990480
rect 160094 990468 160100 990480
rect 143316 990440 160100 990468
rect 143316 990428 143322 990440
rect 160094 990428 160100 990440
rect 160152 990428 160158 990480
rect 181714 990428 181720 990480
rect 181772 990468 181778 990480
rect 187602 990468 187608 990480
rect 181772 990440 187608 990468
rect 181772 990428 181778 990440
rect 187602 990428 187608 990440
rect 187660 990428 187666 990480
rect 187694 990428 187700 990480
rect 187752 990468 187758 990480
rect 202874 990468 202880 990480
rect 187752 990440 202880 990468
rect 187752 990428 187758 990440
rect 202874 990428 202880 990440
rect 202932 990428 202938 990480
rect 233050 990428 233056 990480
rect 233108 990468 233114 990480
rect 246942 990468 246948 990480
rect 233108 990440 246948 990468
rect 233108 990428 233114 990440
rect 246942 990428 246948 990440
rect 247000 990428 247006 990480
rect 449820 990468 449848 990508
rect 469030 990496 469036 990508
rect 469088 990496 469094 990548
rect 483014 990496 483020 990548
rect 483072 990496 483078 990548
rect 560202 990496 560208 990548
rect 560260 990536 560266 990548
rect 565740 990536 565768 990576
rect 576854 990564 576860 990576
rect 576912 990564 576918 990616
rect 560260 990508 565768 990536
rect 598952 990536 598980 990644
rect 623682 990604 623688 990616
rect 604564 990576 623688 990604
rect 604564 990536 604592 990576
rect 623682 990564 623688 990576
rect 623740 990564 623746 990616
rect 598952 990508 604592 990536
rect 560260 990496 560266 990508
rect 623866 990496 623872 990548
rect 623924 990536 623930 990548
rect 639782 990536 639788 990548
rect 623924 990508 639788 990536
rect 623924 990496 623930 990508
rect 639782 990496 639788 990508
rect 639840 990496 639846 990548
rect 540974 990468 540980 990480
rect 430592 990440 449848 990468
rect 540900 990440 540980 990468
rect 154390 990360 154396 990412
rect 154448 990400 154454 990412
rect 154574 990400 154580 990412
rect 154448 990372 154580 990400
rect 154448 990360 154454 990372
rect 154574 990360 154580 990372
rect 154632 990360 154638 990412
rect 386322 990360 386328 990412
rect 386380 990400 386386 990412
rect 397638 990400 397644 990412
rect 386380 990372 397644 990400
rect 386380 990360 386386 990372
rect 397638 990360 397644 990372
rect 397696 990360 397702 990412
rect 424962 990360 424968 990412
rect 425020 990400 425026 990412
rect 430592 990400 430620 990440
rect 540900 990412 540928 990440
rect 540974 990428 540980 990440
rect 541032 990428 541038 990480
rect 425020 990372 430620 990400
rect 425020 990360 425026 990372
rect 483014 990360 483020 990412
rect 483072 990400 483078 990412
rect 486602 990400 486608 990412
rect 483072 990372 486608 990400
rect 483072 990360 483078 990372
rect 486602 990360 486608 990372
rect 486660 990400 486666 990412
rect 521654 990400 521660 990412
rect 486660 990372 502288 990400
rect 486660 990360 486666 990372
rect 502260 990332 502288 990372
rect 511920 990372 521660 990400
rect 507762 990332 507768 990344
rect 502260 990304 507768 990332
rect 507762 990292 507768 990304
rect 507820 990292 507826 990344
rect 507854 990292 507860 990344
rect 507912 990332 507918 990344
rect 511920 990332 511948 990372
rect 521654 990360 521660 990372
rect 521712 990360 521718 990412
rect 540882 990360 540888 990412
rect 540940 990360 540946 990412
rect 507912 990304 511948 990332
rect 507912 990292 507918 990304
rect 154574 990224 154580 990276
rect 154632 990264 154638 990276
rect 164142 990264 164148 990276
rect 154632 990236 164148 990264
rect 154632 990224 154638 990236
rect 164142 990224 164148 990236
rect 164200 990224 164206 990276
rect 397638 990224 397644 990276
rect 397696 990264 397702 990276
rect 405734 990264 405740 990276
rect 397696 990236 405740 990264
rect 397696 990224 397702 990236
rect 405734 990224 405740 990236
rect 405792 990224 405798 990276
rect 521654 990224 521660 990276
rect 521712 990264 521718 990276
rect 537846 990264 537852 990276
rect 521712 990236 537852 990264
rect 521712 990224 521718 990236
rect 537846 990224 537852 990236
rect 537904 990264 537910 990276
rect 540882 990264 540888 990276
rect 537904 990236 540888 990264
rect 537904 990224 537910 990236
rect 540882 990224 540888 990236
rect 540940 990224 540946 990276
rect 42242 990156 42248 990208
rect 42300 990196 42306 990208
rect 79962 990196 79968 990208
rect 42300 990168 79968 990196
rect 42300 990156 42306 990168
rect 79962 990156 79968 990168
rect 80020 990156 80026 990208
rect 639782 990156 639788 990208
rect 639840 990196 639846 990208
rect 673638 990196 673644 990208
rect 639840 990168 673644 990196
rect 639840 990156 639846 990168
rect 673638 990156 673644 990168
rect 673696 990156 673702 990208
rect 42426 990088 42432 990140
rect 42484 990128 42490 990140
rect 79042 990128 79048 990140
rect 42484 990100 79048 990128
rect 42484 990088 42490 990100
rect 79042 990088 79048 990100
rect 79100 990088 79106 990140
rect 89990 990088 89996 990140
rect 90048 990088 90054 990140
rect 405734 990088 405740 990140
rect 405792 990128 405798 990140
rect 424962 990128 424968 990140
rect 405792 990100 424968 990128
rect 405792 990088 405798 990100
rect 424962 990088 424968 990100
rect 425020 990088 425026 990140
rect 628650 990088 628656 990140
rect 628708 990088 628714 990140
rect 629294 990088 629300 990140
rect 629352 990128 629358 990140
rect 673546 990128 673552 990140
rect 629352 990100 673552 990128
rect 629352 990088 629358 990100
rect 673546 990088 673552 990100
rect 673604 990088 673610 990140
rect 42518 990020 42524 990072
rect 42576 990060 42582 990072
rect 90008 990060 90036 990088
rect 42576 990032 90036 990060
rect 628668 990060 628696 990088
rect 673454 990060 673460 990072
rect 628668 990032 673460 990060
rect 42576 990020 42582 990032
rect 673454 990020 673460 990032
rect 673512 990020 673518 990072
rect 41782 969348 41788 969400
rect 41840 969388 41846 969400
rect 42334 969388 42340 969400
rect 41840 969360 42340 969388
rect 41840 969348 41846 969360
rect 42334 969348 42340 969360
rect 42392 969348 42398 969400
rect 41782 968464 41788 968516
rect 41840 968504 41846 968516
rect 42518 968504 42524 968516
rect 41840 968476 42524 968504
rect 41840 968464 41846 968476
rect 42518 968464 42524 968476
rect 42576 968464 42582 968516
rect 673454 965268 673460 965320
rect 673512 965308 673518 965320
rect 675386 965308 675392 965320
rect 673512 965280 675392 965308
rect 673512 965268 673518 965280
rect 675386 965268 675392 965280
rect 675444 965268 675450 965320
rect 673546 964724 673552 964776
rect 673604 964764 673610 964776
rect 675386 964764 675392 964776
rect 673604 964736 675392 964764
rect 673604 964724 673610 964736
rect 675386 964724 675392 964736
rect 675444 964724 675450 964776
rect 41782 962412 41788 962464
rect 41840 962452 41846 962464
rect 42334 962452 42340 962464
rect 41840 962424 42340 962452
rect 41840 962412 41846 962424
rect 42334 962412 42340 962424
rect 42392 962412 42398 962464
rect 41782 956428 41788 956480
rect 41840 956468 41846 956480
rect 42426 956468 42432 956480
rect 41840 956440 42432 956468
rect 41840 956428 41846 956440
rect 42426 956428 42432 956440
rect 42484 956428 42490 956480
rect 673638 953300 673644 953352
rect 673696 953340 673702 953352
rect 675386 953340 675392 953352
rect 673696 953312 675392 953340
rect 673696 953300 673702 953312
rect 675386 953300 675392 953312
rect 675444 953300 675450 953352
rect 44266 930112 44272 930164
rect 44324 930152 44330 930164
rect 45462 930152 45468 930164
rect 44324 930124 45468 930152
rect 44324 930112 44330 930124
rect 45462 930112 45468 930124
rect 45520 930112 45526 930164
rect 39666 922904 39672 922956
rect 39724 922944 39730 922956
rect 44266 922944 44272 922956
rect 39724 922916 44272 922944
rect 39724 922904 39730 922916
rect 44266 922904 44272 922916
rect 44324 922904 44330 922956
rect 39850 914676 39856 914728
rect 39908 914716 39914 914728
rect 41414 914716 41420 914728
rect 39908 914688 41420 914716
rect 39908 914676 39914 914688
rect 41414 914676 41420 914688
rect 41472 914716 41478 914728
rect 42242 914716 42248 914728
rect 41472 914688 42248 914716
rect 41472 914676 41478 914688
rect 42242 914676 42248 914688
rect 42300 914676 42306 914728
rect 673546 910732 673552 910784
rect 673604 910772 673610 910784
rect 677778 910772 677784 910784
rect 673604 910744 677784 910772
rect 673604 910732 673610 910744
rect 677778 910732 677784 910744
rect 677836 910732 677842 910784
rect 673178 908012 673184 908064
rect 673236 908052 673242 908064
rect 673454 908052 673460 908064
rect 673236 908024 673460 908052
rect 673236 908012 673242 908024
rect 673454 908012 673460 908024
rect 673512 908012 673518 908064
rect 673178 888768 673184 888820
rect 673236 888808 673242 888820
rect 673454 888808 673460 888820
rect 673236 888780 673460 888808
rect 673236 888768 673242 888780
rect 673454 888768 673460 888780
rect 673512 888768 673518 888820
rect 39850 879792 39856 879844
rect 39908 879832 39914 879844
rect 40126 879832 40132 879844
rect 39908 879804 40132 879832
rect 39908 879792 39914 879804
rect 40126 879792 40132 879804
rect 40184 879832 40190 879844
rect 44174 879832 44180 879844
rect 40184 879804 44180 879832
rect 40184 879792 40190 879804
rect 44174 879792 44180 879804
rect 44232 879832 44238 879844
rect 45830 879832 45836 879844
rect 44232 879804 45836 879832
rect 44232 879792 44238 879804
rect 45830 879792 45836 879804
rect 45888 879792 45894 879844
rect 41414 875576 41420 875628
rect 41472 875616 41478 875628
rect 42242 875616 42248 875628
rect 41472 875588 42248 875616
rect 41472 875576 41478 875588
rect 42242 875576 42248 875588
rect 42300 875576 42306 875628
rect 673546 875508 673552 875560
rect 673604 875548 673610 875560
rect 675386 875548 675392 875560
rect 673604 875520 675392 875548
rect 673604 875508 673610 875520
rect 675386 875508 675392 875520
rect 675444 875508 675450 875560
rect 673638 875032 673644 875084
rect 673696 875032 673702 875084
rect 673656 874948 673684 875032
rect 673638 874896 673644 874948
rect 673696 874896 673702 874948
rect 673730 869388 673736 869440
rect 673788 869428 673794 869440
rect 675202 869428 675208 869440
rect 673788 869400 675208 869428
rect 673788 869388 673794 869400
rect 675202 869388 675208 869400
rect 675260 869388 675266 869440
rect 673638 864968 673644 865020
rect 673696 865008 673702 865020
rect 673822 865008 673828 865020
rect 673696 864980 673828 865008
rect 673696 864968 673702 864980
rect 673822 864968 673828 864980
rect 673880 865008 673886 865020
rect 675386 865008 675392 865020
rect 673880 864980 675392 865008
rect 673880 864968 673886 864980
rect 675386 864968 675392 864980
rect 675444 864968 675450 865020
rect 673546 836272 673552 836324
rect 673604 836312 673610 836324
rect 673604 836284 673684 836312
rect 673604 836272 673610 836284
rect 673656 836256 673684 836284
rect 673638 836204 673644 836256
rect 673696 836204 673702 836256
rect 673546 830764 673552 830816
rect 673604 830804 673610 830816
rect 673638 830804 673644 830816
rect 673604 830776 673644 830804
rect 673604 830764 673610 830776
rect 673638 830764 673644 830776
rect 673696 830764 673702 830816
rect 673546 821040 673552 821092
rect 673604 821080 673610 821092
rect 674098 821080 674104 821092
rect 673604 821052 674104 821080
rect 673604 821040 673610 821052
rect 674098 821040 674104 821052
rect 674156 821040 674162 821092
rect 42242 807304 42248 807356
rect 42300 807344 42306 807356
rect 42702 807344 42708 807356
rect 42300 807316 42708 807344
rect 42300 807304 42306 807316
rect 42702 807304 42708 807316
rect 42760 807304 42766 807356
rect 44542 805944 44548 805996
rect 44600 805984 44606 805996
rect 44726 805984 44732 805996
rect 44600 805956 44732 805984
rect 44600 805944 44606 805956
rect 44726 805944 44732 805956
rect 44784 805944 44790 805996
rect 41782 798328 41788 798380
rect 41840 798368 41846 798380
rect 42518 798368 42524 798380
rect 41840 798340 42524 798368
rect 41840 798328 41846 798340
rect 42518 798328 42524 798340
rect 42576 798328 42582 798380
rect 674098 797580 674104 797632
rect 674156 797620 674162 797632
rect 675294 797620 675300 797632
rect 674156 797592 675300 797620
rect 674156 797580 674162 797592
rect 675294 797580 675300 797592
rect 675352 797580 675358 797632
rect 41782 787856 41788 787908
rect 41840 787896 41846 787908
rect 42426 787896 42432 787908
rect 41840 787868 42432 787896
rect 41840 787856 41846 787868
rect 42426 787856 42432 787868
rect 42484 787896 42490 787908
rect 42702 787896 42708 787908
rect 42484 787868 42708 787896
rect 42484 787856 42490 787868
rect 42702 787856 42708 787868
rect 42760 787856 42766 787908
rect 42242 787176 42248 787228
rect 42300 787216 42306 787228
rect 42610 787216 42616 787228
rect 42300 787188 42616 787216
rect 42300 787176 42306 787188
rect 42610 787176 42616 787188
rect 42668 787176 42674 787228
rect 674006 786428 674012 786480
rect 674064 786468 674070 786480
rect 675294 786468 675300 786480
rect 674064 786440 675300 786468
rect 674064 786428 674070 786440
rect 675294 786428 675300 786440
rect 675352 786428 675358 786480
rect 673638 785272 673644 785324
rect 673696 785312 673702 785324
rect 675386 785312 675392 785324
rect 673696 785284 675392 785312
rect 673696 785272 673702 785284
rect 675386 785272 675392 785284
rect 675444 785272 675450 785324
rect 672994 778336 673000 778388
rect 673052 778336 673058 778388
rect 673012 778240 673040 778336
rect 673086 778240 673092 778252
rect 673012 778212 673092 778240
rect 673086 778200 673092 778212
rect 673144 778200 673150 778252
rect 673454 774868 673460 774920
rect 673512 774908 673518 774920
rect 673822 774908 673828 774920
rect 673512 774880 673828 774908
rect 673512 774868 673518 774880
rect 673822 774868 673828 774880
rect 673880 774908 673886 774920
rect 675386 774908 675392 774920
rect 673880 774880 675392 774908
rect 673880 774868 673886 774880
rect 675386 774868 675392 774880
rect 675444 774868 675450 774920
rect 672810 772760 672816 772812
rect 672868 772800 672874 772812
rect 673086 772800 673092 772812
rect 672868 772772 673092 772800
rect 672868 772760 672874 772772
rect 673086 772760 673092 772772
rect 673144 772760 673150 772812
rect 42518 768612 42524 768664
rect 42576 768652 42582 768664
rect 42702 768652 42708 768664
rect 42576 768624 42708 768652
rect 42576 768612 42582 768624
rect 42702 768612 42708 768624
rect 42760 768612 42766 768664
rect 673546 768612 673552 768664
rect 673604 768652 673610 768664
rect 674006 768652 674012 768664
rect 673604 768624 674012 768652
rect 673604 768612 673610 768624
rect 674006 768612 674012 768624
rect 674064 768612 674070 768664
rect 41782 754468 41788 754520
rect 41840 754508 41846 754520
rect 42518 754508 42524 754520
rect 41840 754480 42524 754508
rect 41840 754468 41846 754480
rect 42518 754468 42524 754480
rect 42576 754508 42582 754520
rect 42702 754508 42708 754520
rect 42576 754480 42708 754508
rect 42576 754468 42582 754480
rect 42702 754468 42708 754480
rect 42760 754468 42766 754520
rect 41782 744404 41788 744456
rect 41840 744444 41846 744456
rect 42610 744444 42616 744456
rect 41840 744416 42616 744444
rect 41840 744404 41846 744416
rect 42610 744404 42616 744416
rect 42668 744404 42674 744456
rect 673546 741888 673552 741940
rect 673604 741928 673610 741940
rect 674190 741928 674196 741940
rect 673604 741900 674196 741928
rect 673604 741888 673610 741900
rect 674190 741888 674196 741900
rect 674248 741928 674254 741940
rect 675386 741928 675392 741940
rect 674248 741900 675392 741928
rect 674248 741888 674254 741900
rect 675386 741888 675392 741900
rect 675444 741888 675450 741940
rect 673638 741344 673644 741396
rect 673696 741384 673702 741396
rect 675386 741384 675392 741396
rect 673696 741356 675392 741384
rect 673696 741344 673702 741356
rect 675386 741344 675392 741356
rect 675444 741344 675450 741396
rect 672994 739712 673000 739764
rect 673052 739712 673058 739764
rect 673012 739616 673040 739712
rect 673178 739616 673184 739628
rect 673012 739588 673184 739616
rect 673178 739576 673184 739588
rect 673236 739576 673242 739628
rect 673454 730124 673460 730176
rect 673512 730164 673518 730176
rect 675386 730164 675392 730176
rect 673512 730136 675392 730164
rect 673512 730124 673518 730136
rect 675386 730124 675392 730136
rect 675444 730124 675450 730176
rect 673822 729988 673828 730040
rect 673880 730028 673886 730040
rect 675110 730028 675116 730040
rect 673880 730000 675116 730028
rect 673880 729988 673886 730000
rect 675110 729988 675116 730000
rect 675168 729988 675174 730040
rect 674006 720400 674012 720452
rect 674064 720440 674070 720452
rect 674190 720440 674196 720452
rect 674064 720412 674196 720440
rect 674064 720400 674070 720412
rect 674190 720400 674196 720412
rect 674248 720400 674254 720452
rect 41782 711288 41788 711340
rect 41840 711328 41846 711340
rect 42518 711328 42524 711340
rect 41840 711300 42524 711328
rect 41840 711288 41846 711300
rect 42518 711288 42524 711300
rect 42576 711288 42582 711340
rect 674006 710676 674012 710728
rect 674064 710716 674070 710728
rect 675294 710716 675300 710728
rect 674064 710688 675300 710716
rect 674064 710676 674070 710688
rect 675294 710676 675300 710688
rect 675352 710676 675358 710728
rect 42242 700952 42248 701004
rect 42300 700992 42306 701004
rect 42518 700992 42524 701004
rect 42300 700964 42524 700992
rect 42300 700952 42306 700964
rect 42518 700952 42524 700964
rect 42576 700952 42582 701004
rect 41782 700816 41788 700868
rect 41840 700856 41846 700868
rect 42610 700856 42616 700868
rect 41840 700828 42616 700856
rect 41840 700816 41846 700828
rect 42610 700816 42616 700828
rect 42668 700816 42674 700868
rect 673638 695920 673644 695972
rect 673696 695960 673702 695972
rect 675386 695960 675392 695972
rect 673696 695932 675392 695960
rect 673696 695920 673702 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 673086 695512 673092 695564
rect 673144 695552 673150 695564
rect 673178 695552 673184 695564
rect 673144 695524 673184 695552
rect 673144 695512 673150 695524
rect 673178 695512 673184 695524
rect 673236 695512 673242 695564
rect 44634 695444 44640 695496
rect 44692 695484 44698 695496
rect 44910 695484 44916 695496
rect 44692 695456 44916 695484
rect 44692 695444 44698 695456
rect 44910 695444 44916 695456
rect 44968 695444 44974 695496
rect 673546 695308 673552 695360
rect 673604 695348 673610 695360
rect 673822 695348 673828 695360
rect 673604 695320 673828 695348
rect 673604 695308 673610 695320
rect 673822 695308 673828 695320
rect 673880 695348 673886 695360
rect 675386 695348 675392 695360
rect 673880 695320 675392 695348
rect 673880 695308 673886 695320
rect 675386 695308 675392 695320
rect 675444 695308 675450 695360
rect 44726 676200 44732 676252
rect 44784 676240 44790 676252
rect 44910 676240 44916 676252
rect 44784 676212 44916 676240
rect 44784 676200 44790 676212
rect 44910 676200 44916 676212
rect 44968 676200 44974 676252
rect 42334 669168 42340 669180
rect 41800 669140 42340 669168
rect 41800 669112 41828 669140
rect 42334 669128 42340 669140
rect 42392 669128 42398 669180
rect 41782 669060 41788 669112
rect 41840 669060 41846 669112
rect 673178 662464 673184 662516
rect 673236 662464 673242 662516
rect 44542 662396 44548 662448
rect 44600 662436 44606 662448
rect 44726 662436 44732 662448
rect 44600 662408 44732 662436
rect 44600 662396 44606 662408
rect 44726 662396 44732 662408
rect 44784 662396 44790 662448
rect 673196 662380 673224 662464
rect 673178 662328 673184 662380
rect 673236 662328 673242 662380
rect 41782 657636 41788 657688
rect 41840 657676 41846 657688
rect 42518 657676 42524 657688
rect 41840 657648 42524 657676
rect 41840 657636 41846 657648
rect 42518 657636 42524 657648
rect 42576 657636 42582 657688
rect 41782 657092 41788 657144
rect 41840 657132 41846 657144
rect 42334 657132 42340 657144
rect 41840 657104 42340 657132
rect 41840 657092 41846 657104
rect 42334 657092 42340 657104
rect 42392 657132 42398 657144
rect 42610 657132 42616 657144
rect 42392 657104 42616 657132
rect 42392 657092 42398 657104
rect 42610 657092 42616 657104
rect 42668 657092 42674 657144
rect 44634 656820 44640 656872
rect 44692 656860 44698 656872
rect 44818 656860 44824 656872
rect 44692 656832 44824 656860
rect 44692 656820 44698 656832
rect 44818 656820 44824 656832
rect 44876 656820 44882 656872
rect 673638 651720 673644 651772
rect 673696 651760 673702 651772
rect 675386 651760 675392 651772
rect 673696 651732 675392 651760
rect 673696 651720 673702 651732
rect 675386 651720 675392 651732
rect 675444 651720 675450 651772
rect 673546 651108 673552 651160
rect 673604 651148 673610 651160
rect 675386 651148 675392 651160
rect 673604 651120 675392 651148
rect 673604 651108 673610 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 673454 639684 673460 639736
rect 673512 639724 673518 639736
rect 675386 639724 675392 639736
rect 673512 639696 675392 639724
rect 673512 639684 673518 639696
rect 675386 639684 675392 639696
rect 675444 639684 675450 639736
rect 672810 637508 672816 637560
rect 672868 637548 672874 637560
rect 673086 637548 673092 637560
rect 672868 637520 673092 637548
rect 672868 637508 672874 637520
rect 673086 637508 673092 637520
rect 673144 637508 673150 637560
rect 42518 633496 42524 633548
rect 42576 633496 42582 633548
rect 42536 633344 42564 633496
rect 42518 633292 42524 633344
rect 42576 633292 42582 633344
rect 42334 633224 42340 633276
rect 42392 633264 42398 633276
rect 42610 633264 42616 633276
rect 42392 633236 42616 633264
rect 42392 633224 42398 633236
rect 42610 633224 42616 633236
rect 42668 633224 42674 633276
rect 41782 625880 41788 625932
rect 41840 625920 41846 625932
rect 42426 625920 42432 625932
rect 41840 625892 42432 625920
rect 41840 625880 41846 625892
rect 42426 625880 42432 625892
rect 42484 625880 42490 625932
rect 672810 618264 672816 618316
rect 672868 618304 672874 618316
rect 672994 618304 673000 618316
rect 672868 618276 673000 618304
rect 672868 618264 672874 618276
rect 672994 618264 673000 618276
rect 673052 618264 673058 618316
rect 41874 614456 41880 614508
rect 41932 614496 41938 614508
rect 42242 614496 42248 614508
rect 41932 614468 42248 614496
rect 41932 614456 41938 614468
rect 42242 614456 42248 614468
rect 42300 614496 42306 614508
rect 42610 614496 42616 614508
rect 42300 614468 42616 614496
rect 42300 614456 42306 614468
rect 42610 614456 42616 614468
rect 42668 614456 42674 614508
rect 41782 614388 41788 614440
rect 41840 614428 41846 614440
rect 42518 614428 42524 614440
rect 41840 614400 42524 614428
rect 41840 614388 41846 614400
rect 42518 614388 42524 614400
rect 42576 614388 42582 614440
rect 673638 606704 673644 606756
rect 673696 606744 673702 606756
rect 675386 606744 675392 606756
rect 673696 606716 675392 606744
rect 673696 606704 673702 606716
rect 675386 606704 675392 606716
rect 675444 606704 675450 606756
rect 673546 605616 673552 605668
rect 673604 605656 673610 605668
rect 675294 605656 675300 605668
rect 673604 605628 675300 605656
rect 673604 605616 673610 605628
rect 675294 605616 675300 605628
rect 675352 605616 675358 605668
rect 44634 604528 44640 604580
rect 44692 604528 44698 604580
rect 44652 604444 44680 604528
rect 44634 604392 44640 604444
rect 44692 604392 44698 604444
rect 673546 604392 673552 604444
rect 673604 604432 673610 604444
rect 673822 604432 673828 604444
rect 673604 604404 673828 604432
rect 673604 604392 673610 604404
rect 673822 604392 673828 604404
rect 673880 604392 673886 604444
rect 672810 598952 672816 599004
rect 672868 598992 672874 599004
rect 673086 598992 673092 599004
rect 672868 598964 673092 598992
rect 672868 598952 672874 598964
rect 673086 598952 673092 598964
rect 673144 598952 673150 599004
rect 673454 594872 673460 594924
rect 673512 594912 673518 594924
rect 675386 594912 675392 594924
rect 673512 594884 675392 594912
rect 673512 594872 673518 594884
rect 675386 594872 675392 594884
rect 675444 594872 675450 594924
rect 673086 585188 673092 585200
rect 673012 585160 673092 585188
rect 673012 585132 673040 585160
rect 673086 585148 673092 585160
rect 673144 585148 673150 585200
rect 672994 585080 673000 585132
rect 673052 585080 673058 585132
rect 42242 584196 42248 584248
rect 42300 584236 42306 584248
rect 42610 584236 42616 584248
rect 42300 584208 42616 584236
rect 42300 584196 42306 584208
rect 42610 584196 42616 584208
rect 42668 584196 42674 584248
rect 41782 581680 41788 581732
rect 41840 581720 41846 581732
rect 42426 581720 42432 581732
rect 41840 581692 42432 581720
rect 41840 581680 41846 581692
rect 42426 581680 42432 581692
rect 42484 581680 42490 581732
rect 41782 572228 41788 572280
rect 41840 572268 41846 572280
rect 42242 572268 42248 572280
rect 41840 572240 42248 572268
rect 41840 572228 41846 572240
rect 42242 572228 42248 572240
rect 42300 572268 42306 572280
rect 42518 572268 42524 572280
rect 42300 572240 42524 572268
rect 42300 572228 42306 572240
rect 42518 572228 42524 572240
rect 42576 572228 42582 572280
rect 41782 571616 41788 571668
rect 41840 571656 41846 571668
rect 42610 571656 42616 571668
rect 41840 571628 42616 571656
rect 41840 571616 41846 571628
rect 42610 571616 42616 571628
rect 42668 571616 42674 571668
rect 672810 569916 672816 569968
rect 672868 569956 672874 569968
rect 672994 569956 673000 569968
rect 672868 569928 673000 569956
rect 672868 569916 672874 569928
rect 672994 569916 673000 569928
rect 673052 569916 673058 569968
rect 673546 565836 673552 565888
rect 673604 565876 673610 565888
rect 673914 565876 673920 565888
rect 673604 565848 673920 565876
rect 673604 565836 673610 565848
rect 673914 565836 673920 565848
rect 673972 565836 673978 565888
rect 673638 561484 673644 561536
rect 673696 561524 673702 561536
rect 675386 561524 675392 561536
rect 673696 561496 675392 561524
rect 673696 561484 673702 561496
rect 675386 561484 675392 561496
rect 675444 561484 675450 561536
rect 672810 560260 672816 560312
rect 672868 560300 672874 560312
rect 672994 560300 673000 560312
rect 672868 560272 673000 560300
rect 672868 560260 672874 560272
rect 672994 560260 673000 560272
rect 673052 560260 673058 560312
rect 673546 559920 673552 559972
rect 673604 559960 673610 559972
rect 673914 559960 673920 559972
rect 673604 559932 673920 559960
rect 673604 559920 673610 559932
rect 673914 559920 673920 559932
rect 673972 559960 673978 559972
rect 675386 559960 675392 559972
rect 673972 559932 675392 559960
rect 673972 559920 673978 559932
rect 675386 559920 675392 559932
rect 675444 559920 675450 559972
rect 673454 550468 673460 550520
rect 673512 550508 673518 550520
rect 675386 550508 675392 550520
rect 673512 550480 675392 550508
rect 673512 550468 673518 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 672994 546524 673000 546576
rect 673052 546564 673058 546576
rect 673052 546536 673132 546564
rect 673052 546524 673058 546536
rect 673104 546372 673132 546536
rect 673086 546320 673092 546372
rect 673144 546320 673150 546372
rect 44726 540948 44732 541000
rect 44784 540988 44790 541000
rect 44910 540988 44916 541000
rect 44784 540960 44916 540988
rect 44784 540948 44790 540960
rect 44910 540948 44916 540960
rect 44968 540948 44974 541000
rect 41782 538500 41788 538552
rect 41840 538540 41846 538552
rect 42426 538540 42432 538552
rect 41840 538512 42432 538540
rect 41840 538500 41846 538512
rect 42426 538500 42432 538512
rect 42484 538500 42490 538552
rect 41782 528436 41788 528488
rect 41840 528476 41846 528488
rect 42426 528476 42432 528488
rect 41840 528448 42432 528476
rect 41840 528436 41846 528448
rect 42426 528436 42432 528448
rect 42484 528476 42490 528488
rect 42610 528476 42616 528488
rect 42484 528448 42616 528476
rect 42484 528436 42490 528448
rect 42610 528436 42616 528448
rect 42668 528436 42674 528488
rect 673086 527144 673092 527196
rect 673144 527144 673150 527196
rect 673104 527048 673132 527144
rect 673178 527048 673184 527060
rect 673104 527020 673184 527048
rect 673178 527008 673184 527020
rect 673236 527008 673242 527060
rect 673730 522928 673736 522980
rect 673788 522968 673794 522980
rect 673914 522968 673920 522980
rect 673788 522940 673920 522968
rect 673788 522928 673794 522940
rect 673914 522928 673920 522940
rect 673972 522928 673978 522980
rect 673178 521568 673184 521620
rect 673236 521608 673242 521620
rect 676122 521608 676128 521620
rect 673236 521580 676128 521608
rect 673236 521568 673242 521580
rect 676122 521568 676128 521580
rect 676180 521568 676186 521620
rect 44542 496816 44548 496868
rect 44600 496856 44606 496868
rect 44726 496856 44732 496868
rect 44600 496828 44732 496856
rect 44600 496816 44606 496828
rect 44726 496816 44732 496828
rect 44784 496816 44790 496868
rect 673730 463632 673736 463684
rect 673788 463672 673794 463684
rect 677686 463672 677692 463684
rect 673788 463644 677692 463672
rect 673788 463632 673794 463644
rect 677686 463632 677692 463644
rect 677744 463632 677750 463684
rect 39390 458192 39396 458244
rect 39448 458232 39454 458244
rect 44266 458232 44272 458244
rect 39448 458204 44272 458232
rect 39448 458192 39454 458204
rect 44266 458192 44272 458204
rect 44324 458192 44330 458244
rect 672994 449896 673000 449948
rect 673052 449936 673058 449948
rect 673362 449936 673368 449948
rect 673052 449908 673368 449936
rect 673052 449896 673058 449908
rect 673362 449896 673368 449908
rect 673420 449896 673426 449948
rect 39850 448264 39856 448316
rect 39908 448304 39914 448316
rect 42242 448304 42248 448316
rect 39908 448276 42248 448304
rect 39908 448264 39914 448276
rect 42242 448264 42248 448276
rect 42300 448264 42306 448316
rect 676214 440172 676220 440224
rect 676272 440212 676278 440224
rect 677686 440212 677692 440224
rect 676272 440184 677692 440212
rect 676272 440172 676278 440184
rect 677686 440172 677692 440184
rect 677744 440172 677750 440224
rect 42242 413380 42248 413432
rect 42300 413420 42306 413432
rect 42610 413420 42616 413432
rect 42300 413392 42616 413420
rect 42300 413380 42306 413392
rect 42610 413380 42616 413392
rect 42668 413380 42674 413432
rect 672810 412496 672816 412548
rect 672868 412536 672874 412548
rect 676214 412536 676220 412548
rect 672868 412508 676220 412536
rect 672868 412496 672874 412508
rect 676214 412496 676220 412508
rect 676272 412496 676278 412548
rect 41782 410932 41788 410984
rect 41840 410972 41846 410984
rect 42518 410972 42524 410984
rect 41840 410944 42524 410972
rect 41840 410932 41846 410944
rect 42518 410932 42524 410944
rect 42576 410932 42582 410984
rect 672534 405628 672540 405680
rect 672592 405668 672598 405680
rect 672718 405668 672724 405680
rect 672592 405640 672724 405668
rect 672592 405628 672598 405640
rect 672718 405628 672724 405640
rect 672776 405628 672782 405680
rect 673454 401548 673460 401600
rect 673512 401588 673518 401600
rect 675294 401588 675300 401600
rect 673512 401560 675300 401588
rect 673512 401548 673518 401560
rect 675294 401548 675300 401560
rect 675352 401548 675358 401600
rect 41782 401480 41788 401532
rect 41840 401520 41846 401532
rect 42242 401520 42248 401532
rect 41840 401492 42248 401520
rect 41840 401480 41846 401492
rect 42242 401480 42248 401492
rect 42300 401520 42306 401532
rect 42610 401520 42616 401532
rect 42300 401492 42616 401520
rect 42300 401480 42306 401492
rect 42610 401480 42616 401492
rect 42668 401480 42674 401532
rect 41966 400120 41972 400172
rect 42024 400160 42030 400172
rect 42426 400160 42432 400172
rect 42024 400132 42432 400160
rect 42024 400120 42030 400132
rect 42426 400120 42432 400132
rect 42484 400120 42490 400172
rect 672534 386384 672540 386436
rect 672592 386424 672598 386436
rect 672810 386424 672816 386436
rect 672592 386396 672816 386424
rect 672592 386384 672598 386396
rect 672810 386384 672816 386396
rect 672868 386384 672874 386436
rect 673546 384004 673552 384056
rect 673604 384044 673610 384056
rect 675386 384044 675392 384056
rect 673604 384016 675392 384044
rect 673604 384004 673610 384016
rect 675386 384004 675392 384016
rect 675444 384004 675450 384056
rect 673638 382712 673644 382764
rect 673696 382752 673702 382764
rect 675386 382752 675392 382764
rect 673696 382724 675392 382752
rect 673696 382712 673702 382724
rect 675386 382712 675392 382724
rect 675444 382712 675450 382764
rect 42334 380876 42340 380928
rect 42392 380916 42398 380928
rect 42610 380916 42616 380928
rect 42392 380888 42616 380916
rect 42392 380876 42398 380888
rect 42610 380876 42616 380888
rect 42668 380876 42674 380928
rect 673822 372308 673828 372360
rect 673880 372348 673886 372360
rect 675386 372348 675392 372360
rect 673880 372320 675392 372348
rect 673880 372308 673886 372320
rect 675386 372308 675392 372320
rect 675444 372308 675450 372360
rect 41782 368636 41788 368688
rect 41840 368676 41846 368688
rect 42518 368676 42524 368688
rect 41840 368648 42524 368676
rect 41840 368636 41846 368648
rect 42518 368636 42524 368648
rect 42576 368636 42582 368688
rect 42518 367004 42524 367056
rect 42576 367004 42582 367056
rect 42536 366976 42564 367004
rect 42794 366976 42800 366988
rect 42536 366948 42800 366976
rect 42794 366936 42800 366948
rect 42852 366936 42858 366988
rect 41782 357484 41788 357536
rect 41840 357524 41846 357536
rect 42334 357524 42340 357536
rect 41840 357496 42340 357524
rect 41840 357484 41846 357496
rect 42334 357484 42340 357496
rect 42392 357524 42398 357536
rect 42610 357524 42616 357536
rect 42392 357496 42616 357524
rect 42392 357484 42398 357496
rect 42610 357484 42616 357496
rect 42668 357484 42674 357536
rect 41782 356668 41788 356720
rect 41840 356708 41846 356720
rect 42426 356708 42432 356720
rect 41840 356680 42432 356708
rect 41840 356668 41846 356680
rect 42426 356668 42432 356680
rect 42484 356668 42490 356720
rect 672626 353376 672632 353388
rect 672552 353348 672632 353376
rect 672552 353252 672580 353348
rect 672626 353336 672632 353348
rect 672684 353336 672690 353388
rect 672534 353200 672540 353252
rect 672592 353200 672598 353252
rect 42702 347692 42708 347744
rect 42760 347732 42766 347744
rect 42886 347732 42892 347744
rect 42760 347704 42892 347732
rect 42760 347692 42766 347704
rect 42886 347692 42892 347704
rect 42944 347692 42950 347744
rect 672534 347692 672540 347744
rect 672592 347732 672598 347744
rect 672718 347732 672724 347744
rect 672592 347704 672724 347732
rect 672592 347692 672598 347704
rect 672718 347692 672724 347704
rect 672776 347692 672782 347744
rect 673638 338512 673644 338564
rect 673696 338552 673702 338564
rect 675386 338552 675392 338564
rect 673696 338524 675392 338552
rect 673696 338512 673702 338524
rect 675386 338512 675392 338524
rect 675444 338512 675450 338564
rect 42334 334636 42340 334688
rect 42392 334676 42398 334688
rect 42610 334676 42616 334688
rect 42392 334648 42616 334676
rect 42392 334636 42398 334648
rect 42610 334636 42616 334648
rect 42668 334636 42674 334688
rect 42610 328448 42616 328500
rect 42668 328488 42674 328500
rect 42886 328488 42892 328500
rect 42668 328460 42892 328488
rect 42668 328448 42674 328460
rect 42886 328448 42892 328460
rect 42944 328448 42950 328500
rect 672442 328448 672448 328500
rect 672500 328488 672506 328500
rect 672718 328488 672724 328500
rect 672500 328460 672724 328488
rect 672500 328448 672506 328460
rect 672718 328448 672724 328460
rect 672776 328448 672782 328500
rect 673822 327088 673828 327140
rect 673880 327128 673886 327140
rect 675386 327128 675392 327140
rect 673880 327100 675392 327128
rect 673880 327088 673886 327100
rect 675386 327088 675392 327100
rect 675444 327088 675450 327140
rect 41782 324504 41788 324556
rect 41840 324544 41846 324556
rect 41840 324516 42564 324544
rect 41840 324504 41846 324516
rect 42536 324488 42564 324516
rect 42518 324436 42524 324488
rect 42576 324436 42582 324488
rect 42334 314576 42340 314628
rect 42392 314576 42398 314628
rect 42352 314548 42380 314576
rect 42610 314548 42616 314560
rect 41800 314520 42616 314548
rect 41800 314492 41828 314520
rect 42610 314508 42616 314520
rect 42668 314508 42674 314560
rect 41782 314440 41788 314492
rect 41840 314440 41846 314492
rect 42518 314440 42524 314492
rect 42576 314480 42582 314492
rect 42794 314480 42800 314492
rect 42576 314452 42800 314480
rect 42576 314440 42582 314452
rect 42794 314440 42800 314452
rect 42852 314440 42858 314492
rect 41782 313760 41788 313812
rect 41840 313800 41846 313812
rect 42426 313800 42432 313812
rect 41840 313772 42432 313800
rect 41840 313760 41846 313772
rect 42426 313760 42432 313772
rect 42484 313760 42490 313812
rect 672534 309068 672540 309120
rect 672592 309108 672598 309120
rect 672810 309108 672816 309120
rect 672592 309080 672816 309108
rect 672592 309068 672598 309080
rect 672810 309068 672816 309080
rect 672868 309068 672874 309120
rect 42426 307912 42432 307964
rect 42484 307952 42490 307964
rect 42702 307952 42708 307964
rect 42484 307924 42708 307952
rect 42484 307912 42490 307924
rect 42702 307912 42708 307924
rect 42760 307912 42766 307964
rect 673454 304920 673460 304972
rect 673512 304960 673518 304972
rect 673822 304960 673828 304972
rect 673512 304932 673828 304960
rect 673512 304920 673518 304932
rect 673822 304920 673828 304932
rect 673880 304920 673886 304972
rect 42610 295332 42616 295384
rect 42668 295372 42674 295384
rect 42794 295372 42800 295384
rect 42668 295344 42800 295372
rect 42668 295332 42674 295344
rect 42794 295332 42800 295344
rect 42852 295332 42858 295384
rect 673638 293496 673644 293548
rect 673696 293536 673702 293548
rect 675018 293536 675024 293548
rect 673696 293508 675024 293536
rect 673696 293496 673702 293508
rect 675018 293496 675024 293508
rect 675076 293496 675082 293548
rect 673822 293156 673828 293208
rect 673880 293196 673886 293208
rect 675386 293196 675392 293208
rect 673880 293168 675392 293196
rect 673880 293156 673886 293168
rect 675386 293156 675392 293168
rect 675444 293156 675450 293208
rect 672626 289824 672632 289876
rect 672684 289864 672690 289876
rect 672810 289864 672816 289876
rect 672684 289836 672816 289864
rect 672684 289824 672690 289836
rect 672810 289824 672816 289836
rect 672868 289824 672874 289876
rect 673454 283024 673460 283076
rect 673512 283064 673518 283076
rect 674926 283064 674932 283076
rect 673512 283036 674932 283064
rect 673512 283024 673518 283036
rect 674926 283024 674932 283036
rect 674984 283064 674990 283076
rect 675386 283064 675392 283076
rect 674984 283036 675392 283064
rect 674984 283024 674990 283036
rect 675386 283024 675392 283036
rect 675444 283024 675450 283076
rect 41782 282276 41788 282328
rect 41840 282316 41846 282328
rect 42426 282316 42432 282328
rect 41840 282288 42432 282316
rect 41840 282276 41846 282288
rect 42426 282276 42432 282288
rect 42484 282316 42490 282328
rect 42610 282316 42616 282328
rect 42484 282288 42616 282316
rect 42484 282276 42490 282288
rect 42610 282276 42616 282288
rect 42668 282276 42674 282328
rect 42702 282208 42708 282260
rect 42760 282208 42766 282260
rect 42720 282056 42748 282208
rect 42702 282004 42708 282056
rect 42760 282004 42766 282056
rect 673914 276020 673920 276072
rect 673972 276060 673978 276072
rect 675202 276060 675208 276072
rect 673972 276032 675208 276060
rect 673972 276020 673978 276032
rect 675202 276020 675208 276032
rect 675260 276020 675266 276072
rect 42518 275952 42524 276004
rect 42576 275992 42582 276004
rect 42794 275992 42800 276004
rect 42576 275964 42800 275992
rect 42576 275952 42582 275964
rect 42794 275952 42800 275964
rect 42852 275952 42858 276004
rect 41782 270784 41788 270836
rect 41840 270824 41846 270836
rect 42518 270824 42524 270836
rect 41840 270796 42524 270824
rect 41840 270784 41846 270796
rect 42518 270784 42524 270796
rect 42576 270784 42582 270836
rect 41782 270240 41788 270292
rect 41840 270280 41846 270292
rect 42334 270280 42340 270292
rect 41840 270252 42340 270280
rect 41840 270240 41846 270252
rect 42334 270240 42340 270252
rect 42392 270280 42398 270292
rect 42702 270280 42708 270292
rect 42392 270252 42708 270280
rect 42392 270240 42398 270252
rect 42702 270240 42708 270252
rect 42760 270240 42766 270292
rect 673730 266296 673736 266348
rect 673788 266336 673794 266348
rect 674926 266336 674932 266348
rect 673788 266308 674932 266336
rect 673788 266296 673794 266308
rect 674926 266296 674932 266308
rect 674984 266296 674990 266348
rect 673822 248140 673828 248192
rect 673880 248180 673886 248192
rect 675386 248180 675392 248192
rect 673880 248152 675392 248180
rect 673880 248140 673886 248152
rect 675386 248140 675392 248152
rect 675444 248140 675450 248192
rect 673638 247460 673644 247512
rect 673696 247500 673702 247512
rect 673914 247500 673920 247512
rect 673696 247472 673920 247500
rect 673696 247460 673702 247472
rect 673914 247460 673920 247472
rect 673972 247500 673978 247512
rect 675386 247500 675392 247512
rect 673972 247472 675392 247500
rect 673972 247460 673978 247472
rect 675386 247460 675392 247472
rect 675444 247460 675450 247512
rect 42334 246984 42340 247036
rect 42392 247024 42398 247036
rect 42702 247024 42708 247036
rect 42392 246996 42708 247024
rect 42392 246984 42398 246996
rect 42702 246984 42708 246996
rect 42760 246984 42766 247036
rect 41782 239028 41788 239080
rect 41840 239068 41846 239080
rect 42426 239068 42432 239080
rect 41840 239040 42432 239068
rect 41840 239028 41846 239040
rect 42426 239028 42432 239040
rect 42484 239068 42490 239080
rect 42610 239068 42616 239080
rect 42484 239040 42616 239068
rect 42484 239028 42490 239040
rect 42610 239028 42616 239040
rect 42668 239028 42674 239080
rect 673730 237668 673736 237720
rect 673788 237708 673794 237720
rect 675386 237708 675392 237720
rect 673788 237680 675392 237708
rect 673788 237668 673794 237680
rect 675386 237668 675392 237680
rect 675444 237668 675450 237720
rect 41782 228624 41788 228676
rect 41840 228664 41846 228676
rect 42518 228664 42524 228676
rect 41840 228636 42524 228664
rect 41840 228624 41846 228636
rect 42518 228624 42524 228636
rect 42576 228624 42582 228676
rect 41782 228012 41788 228064
rect 41840 228052 41846 228064
rect 42426 228052 42432 228064
rect 41840 228024 42432 228052
rect 41840 228012 41846 228024
rect 42426 228012 42432 228024
rect 42484 228052 42490 228064
rect 42702 228052 42708 228064
rect 42484 228024 42708 228052
rect 42484 228012 42490 228024
rect 42702 228012 42708 228024
rect 42760 228012 42766 228064
rect 42242 227876 42248 227928
rect 42300 227916 42306 227928
rect 42518 227916 42524 227928
rect 42300 227888 42524 227916
rect 42300 227876 42306 227888
rect 42518 227876 42524 227888
rect 42576 227876 42582 227928
rect 672718 212508 672724 212560
rect 672776 212548 672782 212560
rect 672902 212548 672908 212560
rect 672776 212520 672908 212548
rect 672776 212508 672782 212520
rect 672902 212508 672908 212520
rect 672960 212508 672966 212560
rect 673546 203872 673552 203924
rect 673604 203912 673610 203924
rect 673822 203912 673828 203924
rect 673604 203884 673828 203912
rect 673604 203872 673610 203884
rect 673822 203872 673828 203884
rect 673880 203912 673886 203924
rect 675386 203912 675392 203924
rect 673880 203884 675392 203912
rect 673880 203872 673886 203884
rect 675386 203872 675392 203884
rect 675444 203872 675450 203924
rect 673454 203328 673460 203380
rect 673512 203368 673518 203380
rect 673638 203368 673644 203380
rect 673512 203340 673644 203368
rect 673512 203328 673518 203340
rect 673638 203328 673644 203340
rect 673696 203368 673702 203380
rect 675386 203368 675392 203380
rect 673696 203340 675392 203368
rect 673696 203328 673702 203340
rect 675386 203328 675392 203340
rect 675444 203328 675450 203380
rect 672534 198704 672540 198756
rect 672592 198744 672598 198756
rect 672718 198744 672724 198756
rect 672592 198716 672724 198744
rect 672592 198704 672598 198716
rect 672718 198704 672724 198716
rect 672776 198704 672782 198756
rect 41782 196732 41788 196784
rect 41840 196772 41846 196784
rect 42334 196772 42340 196784
rect 41840 196744 42340 196772
rect 41840 196732 41846 196744
rect 42334 196732 42340 196744
rect 42392 196732 42398 196784
rect 41782 195848 41788 195900
rect 41840 195888 41846 195900
rect 42610 195888 42616 195900
rect 41840 195860 42616 195888
rect 41840 195848 41846 195860
rect 42610 195848 42616 195860
rect 42668 195888 42674 195900
rect 44634 195888 44640 195900
rect 42668 195860 44640 195888
rect 42668 195848 42674 195860
rect 44634 195848 44640 195860
rect 44692 195848 44698 195900
rect 673730 191972 673736 192024
rect 673788 192012 673794 192024
rect 674006 192012 674012 192024
rect 673788 191984 674012 192012
rect 673788 191972 673794 191984
rect 674006 191972 674012 191984
rect 674064 191972 674070 192024
rect 41782 189796 41788 189848
rect 41840 189836 41846 189848
rect 42334 189836 42340 189848
rect 41840 189808 42340 189836
rect 41840 189796 41846 189808
rect 42334 189796 42340 189808
rect 42392 189796 42398 189848
rect 42242 184220 42248 184272
rect 42300 184260 42306 184272
rect 42426 184260 42432 184272
rect 42300 184232 42432 184260
rect 42300 184220 42306 184232
rect 42426 184220 42432 184232
rect 42484 184220 42490 184272
rect 44450 173884 44456 173936
rect 44508 173924 44514 173936
rect 44726 173924 44732 173936
rect 44508 173896 44732 173924
rect 44508 173884 44514 173896
rect 44726 173884 44732 173896
rect 44784 173884 44790 173936
rect 672718 173884 672724 173936
rect 672776 173924 672782 173936
rect 672902 173924 672908 173936
rect 672776 173896 672908 173924
rect 672776 173884 672782 173896
rect 672902 173884 672908 173896
rect 672960 173884 672966 173936
rect 673822 173884 673828 173936
rect 673880 173924 673886 173936
rect 674006 173924 674012 173936
rect 673880 173896 674012 173924
rect 673880 173884 673886 173896
rect 674006 173884 674012 173896
rect 674064 173884 674070 173936
rect 44726 160188 44732 160200
rect 44652 160160 44732 160188
rect 44652 160064 44680 160160
rect 44726 160148 44732 160160
rect 44784 160148 44790 160200
rect 672534 160080 672540 160132
rect 672592 160120 672598 160132
rect 672718 160120 672724 160132
rect 672592 160092 672724 160120
rect 672592 160080 672598 160092
rect 672718 160080 672724 160092
rect 672776 160080 672782 160132
rect 673638 160080 673644 160132
rect 673696 160120 673702 160132
rect 673822 160120 673828 160132
rect 673696 160092 673828 160120
rect 673696 160080 673702 160092
rect 673822 160080 673828 160092
rect 673880 160080 673886 160132
rect 44634 160012 44640 160064
rect 44692 160012 44698 160064
rect 673546 158312 673552 158364
rect 673604 158352 673610 158364
rect 675386 158352 675392 158364
rect 673604 158324 675392 158352
rect 673604 158312 673610 158324
rect 675386 158312 675392 158324
rect 675444 158312 675450 158364
rect 673454 157292 673460 157344
rect 673512 157332 673518 157344
rect 675386 157332 675392 157344
rect 673512 157304 675392 157332
rect 673512 157292 673518 157304
rect 675386 157292 675392 157304
rect 675444 157292 675450 157344
rect 44634 154504 44640 154556
rect 44692 154544 44698 154556
rect 44726 154544 44732 154556
rect 44692 154516 44732 154544
rect 44692 154504 44698 154516
rect 44726 154504 44732 154516
rect 44784 154504 44790 154556
rect 673638 147840 673644 147892
rect 673696 147880 673702 147892
rect 674006 147880 674012 147892
rect 673696 147852 674012 147880
rect 673696 147840 673702 147852
rect 674006 147840 674012 147852
rect 674064 147880 674070 147892
rect 675386 147880 675392 147892
rect 674064 147852 675392 147880
rect 674064 147840 674070 147852
rect 675386 147840 675392 147852
rect 675444 147840 675450 147892
rect 44726 140808 44732 140820
rect 44652 140780 44732 140808
rect 44652 140752 44680 140780
rect 44726 140768 44732 140780
rect 44784 140768 44790 140820
rect 44634 140700 44640 140752
rect 44692 140700 44698 140752
rect 44726 121564 44732 121576
rect 44652 121536 44732 121564
rect 44652 121440 44680 121536
rect 44726 121524 44732 121536
rect 44784 121524 44790 121576
rect 44634 121388 44640 121440
rect 44692 121388 44698 121440
rect 672718 115880 672724 115932
rect 672776 115920 672782 115932
rect 672810 115920 672816 115932
rect 672776 115892 672816 115920
rect 672776 115880 672782 115892
rect 672810 115880 672816 115892
rect 672868 115880 672874 115932
rect 673546 112752 673552 112804
rect 673604 112792 673610 112804
rect 675386 112792 675392 112804
rect 673604 112764 675392 112792
rect 673604 112752 673610 112764
rect 675386 112752 675392 112764
rect 675444 112752 675450 112804
rect 673454 112072 673460 112124
rect 673512 112112 673518 112124
rect 675386 112112 675392 112124
rect 673512 112084 675392 112112
rect 673512 112072 673518 112084
rect 675386 112072 675392 112084
rect 675444 112072 675450 112124
rect 672810 102184 672816 102196
rect 672736 102156 672816 102184
rect 672736 102128 672764 102156
rect 672810 102144 672816 102156
rect 672868 102144 672874 102196
rect 673638 102144 673644 102196
rect 673696 102184 673702 102196
rect 673822 102184 673828 102196
rect 673696 102156 673828 102184
rect 673696 102144 673702 102156
rect 673822 102144 673828 102156
rect 673880 102144 673886 102196
rect 672718 102076 672724 102128
rect 672776 102076 672782 102128
rect 673638 102008 673644 102060
rect 673696 102048 673702 102060
rect 675386 102048 675392 102060
rect 673696 102020 675392 102048
rect 673696 102008 673702 102020
rect 675386 102008 675392 102020
rect 675444 102008 675450 102060
rect 44266 96568 44272 96620
rect 44324 96608 44330 96620
rect 44542 96608 44548 96620
rect 44324 96580 44548 96608
rect 44324 96568 44330 96580
rect 44542 96568 44548 96580
rect 44600 96568 44606 96620
rect 672810 82900 672816 82952
rect 672868 82900 672874 82952
rect 672828 82748 672856 82900
rect 672810 82696 672816 82748
rect 672868 82696 672874 82748
rect 44266 77256 44272 77308
rect 44324 77296 44330 77308
rect 44358 77296 44364 77308
rect 44324 77268 44364 77296
rect 44324 77256 44330 77268
rect 44358 77256 44364 77268
rect 44416 77256 44422 77308
rect 39666 75216 39672 75268
rect 39724 75216 39730 75268
rect 39684 74996 39712 75216
rect 39666 74944 39672 74996
rect 39724 74944 39730 74996
rect 39574 67940 39580 67992
rect 39632 67980 39638 67992
rect 41414 67980 41420 67992
rect 39632 67952 41420 67980
rect 39632 67940 39638 67952
rect 41414 67940 41420 67952
rect 41472 67940 41478 67992
rect 41414 64608 41420 64660
rect 41472 64648 41478 64660
rect 42702 64648 42708 64660
rect 41472 64620 42708 64648
rect 41472 64608 41478 64620
rect 42702 64608 42708 64620
rect 42760 64608 42766 64660
rect 39666 52368 39672 52420
rect 39724 52408 39730 52420
rect 39850 52408 39856 52420
rect 39724 52380 39856 52408
rect 39724 52368 39730 52380
rect 39850 52368 39856 52380
rect 39908 52368 39914 52420
rect 45462 47880 45468 47932
rect 45520 47920 45526 47932
rect 179414 47920 179420 47932
rect 45520 47892 179420 47920
rect 45520 47880 45526 47892
rect 179414 47880 179420 47892
rect 179472 47880 179478 47932
rect 518802 47880 518808 47932
rect 518860 47920 518866 47932
rect 673638 47920 673644 47932
rect 518860 47892 673644 47920
rect 518860 47880 518866 47892
rect 673638 47880 673644 47892
rect 673696 47880 673702 47932
rect 39850 47812 39856 47864
rect 39908 47852 39914 47864
rect 189166 47852 189172 47864
rect 39908 47824 189172 47852
rect 39908 47812 39914 47824
rect 189166 47812 189172 47824
rect 189224 47812 189230 47864
rect 527450 47812 527456 47864
rect 527508 47852 527514 47864
rect 673546 47852 673552 47864
rect 527508 47824 673552 47852
rect 527508 47812 527514 47824
rect 673546 47812 673552 47824
rect 673604 47812 673610 47864
rect 45554 47744 45560 47796
rect 45612 47784 45618 47796
rect 149054 47784 149060 47796
rect 45612 47756 149060 47784
rect 45612 47744 45618 47756
rect 149054 47744 149060 47756
rect 149112 47744 149118 47796
rect 528646 47744 528652 47796
rect 528704 47784 528710 47796
rect 672810 47784 672816 47796
rect 528704 47756 672816 47784
rect 528704 47744 528710 47756
rect 672810 47744 672816 47756
rect 672868 47744 672874 47796
rect 39758 47676 39764 47728
rect 39816 47716 39822 47728
rect 86310 47716 86316 47728
rect 39816 47688 86316 47716
rect 39816 47676 39822 47688
rect 86310 47676 86316 47688
rect 86368 47676 86374 47728
rect 212534 47648 212540 47660
rect 198936 47620 212540 47648
rect 195974 47580 195980 47592
rect 193232 47552 195980 47580
rect 179414 47472 179420 47524
rect 179472 47512 179478 47524
rect 193232 47512 193260 47552
rect 195974 47540 195980 47552
rect 196032 47580 196038 47592
rect 198642 47580 198648 47592
rect 196032 47552 198648 47580
rect 196032 47540 196038 47552
rect 198642 47540 198648 47552
rect 198700 47540 198706 47592
rect 198734 47540 198740 47592
rect 198792 47580 198798 47592
rect 198936 47580 198964 47620
rect 212534 47608 212540 47620
rect 212592 47608 212598 47660
rect 270494 47608 270500 47660
rect 270552 47608 270558 47660
rect 270512 47580 270540 47608
rect 198792 47552 198964 47580
rect 270420 47552 270540 47580
rect 198792 47540 198798 47552
rect 270420 47524 270448 47552
rect 303614 47540 303620 47592
rect 303672 47580 303678 47592
rect 304534 47580 304540 47592
rect 303672 47552 304540 47580
rect 303672 47540 303678 47552
rect 304534 47540 304540 47552
rect 304592 47580 304598 47592
rect 359366 47580 359372 47592
rect 304592 47552 359372 47580
rect 304592 47540 304598 47552
rect 359366 47540 359372 47552
rect 359424 47580 359430 47592
rect 361482 47580 361488 47592
rect 359424 47552 361488 47580
rect 359424 47540 359430 47552
rect 361482 47540 361488 47552
rect 361540 47540 361546 47592
rect 179472 47484 193260 47512
rect 179472 47472 179478 47484
rect 231762 47472 231768 47524
rect 231820 47512 231826 47524
rect 251174 47512 251180 47524
rect 231820 47484 231992 47512
rect 231820 47472 231826 47484
rect 231964 47444 231992 47484
rect 237392 47484 251180 47512
rect 237392 47444 237420 47484
rect 251174 47472 251180 47484
rect 251232 47472 251238 47524
rect 270402 47472 270408 47524
rect 270460 47472 270466 47524
rect 416774 47512 416780 47524
rect 400232 47484 416780 47512
rect 231964 47416 237420 47444
rect 289722 47404 289728 47456
rect 289780 47444 289786 47456
rect 289780 47416 295288 47444
rect 289780 47404 289786 47416
rect 86310 47336 86316 47388
rect 86368 47376 86374 47388
rect 199010 47376 199016 47388
rect 86368 47348 199016 47376
rect 86368 47336 86374 47348
rect 199010 47336 199016 47348
rect 199068 47376 199074 47388
rect 201402 47376 201408 47388
rect 199068 47348 201408 47376
rect 199068 47336 199074 47348
rect 201402 47336 201408 47348
rect 201460 47336 201466 47388
rect 251174 47336 251180 47388
rect 251232 47376 251238 47388
rect 270402 47376 270408 47388
rect 251232 47348 270408 47376
rect 251232 47336 251238 47348
rect 270402 47336 270408 47348
rect 270460 47336 270466 47388
rect 295260 47376 295288 47416
rect 364150 47404 364156 47456
rect 364208 47444 364214 47456
rect 400232 47444 400260 47484
rect 416774 47472 416780 47484
rect 416832 47472 416838 47524
rect 364208 47416 400260 47444
rect 364208 47404 364214 47416
rect 303614 47376 303620 47388
rect 295260 47348 303620 47376
rect 303614 47336 303620 47348
rect 303672 47336 303678 47388
rect 361482 47336 361488 47388
rect 361540 47376 361546 47388
rect 414198 47376 414204 47388
rect 361540 47348 414204 47376
rect 361540 47336 361546 47348
rect 414198 47336 414204 47348
rect 414256 47376 414262 47388
rect 417970 47376 417976 47388
rect 414256 47348 417976 47376
rect 414256 47336 414262 47348
rect 417970 47336 417976 47348
rect 418028 47336 418034 47388
rect 418062 47336 418068 47388
rect 418120 47376 418126 47388
rect 471974 47376 471980 47388
rect 418120 47348 471980 47376
rect 418120 47336 418126 47348
rect 471974 47336 471980 47348
rect 472032 47376 472038 47388
rect 526806 47376 526812 47388
rect 472032 47348 526812 47376
rect 472032 47336 472038 47348
rect 526806 47336 526812 47348
rect 526864 47336 526870 47388
rect 199654 47268 199660 47320
rect 199712 47308 199718 47320
rect 199712 47280 276060 47308
rect 199712 47268 199718 47280
rect 217962 47200 217968 47252
rect 218020 47240 218026 47252
rect 240134 47240 240140 47252
rect 218020 47212 240140 47240
rect 218020 47200 218026 47212
rect 240134 47200 240140 47212
rect 240192 47200 240198 47252
rect 276032 47240 276060 47280
rect 285582 47268 285588 47320
rect 285640 47308 285646 47320
rect 307570 47308 307576 47320
rect 285640 47280 307576 47308
rect 285640 47268 285646 47280
rect 307570 47268 307576 47280
rect 307628 47308 307634 47320
rect 362402 47308 362408 47320
rect 307628 47280 362408 47308
rect 307628 47268 307634 47280
rect 362402 47268 362408 47280
rect 362460 47308 362466 47320
rect 364150 47308 364156 47320
rect 362460 47280 364156 47308
rect 362460 47268 362466 47280
rect 364150 47268 364156 47280
rect 364208 47268 364214 47320
rect 406746 47268 406752 47320
rect 406804 47308 406810 47320
rect 461486 47308 461492 47320
rect 406804 47280 461492 47308
rect 406804 47268 406810 47280
rect 461486 47268 461492 47280
rect 461544 47308 461550 47320
rect 516318 47308 516324 47320
rect 461544 47280 516324 47308
rect 461544 47268 461550 47280
rect 516318 47268 516324 47280
rect 516376 47308 516382 47320
rect 518802 47308 518808 47320
rect 516376 47280 518808 47308
rect 516376 47268 516382 47280
rect 518802 47268 518808 47280
rect 518860 47268 518866 47320
rect 276032 47212 285720 47240
rect 200850 47132 200856 47184
rect 200908 47172 200914 47184
rect 242894 47172 242900 47184
rect 200908 47144 242900 47172
rect 200908 47132 200914 47144
rect 242894 47132 242900 47144
rect 242952 47132 242958 47184
rect 149054 47064 149060 47116
rect 149112 47104 149118 47116
rect 154574 47104 154580 47116
rect 149112 47076 154580 47104
rect 149112 47064 149118 47076
rect 154574 47064 154580 47076
rect 154632 47064 154638 47116
rect 188522 47104 188528 47116
rect 186608 47076 188528 47104
rect 173802 46996 173808 47048
rect 173860 47036 173866 47048
rect 173860 47008 179368 47036
rect 173860 46996 173866 47008
rect 179340 46968 179368 47008
rect 186608 46968 186636 47076
rect 188522 47064 188528 47076
rect 188580 47104 188586 47116
rect 192846 47104 192852 47116
rect 188580 47076 192852 47104
rect 188580 47064 188586 47076
rect 192846 47064 192852 47076
rect 192904 47104 192910 47116
rect 192904 47076 198688 47104
rect 192904 47064 192910 47076
rect 179340 46940 186636 46968
rect 186682 46928 186688 46980
rect 186740 46968 186746 46980
rect 194686 46968 194692 46980
rect 186740 46940 194692 46968
rect 186740 46928 186746 46940
rect 194686 46928 194692 46940
rect 194744 46928 194750 46980
rect 198660 46968 198688 47076
rect 201402 47064 201408 47116
rect 201460 47104 201466 47116
rect 247402 47104 247408 47116
rect 201460 47076 247408 47104
rect 201460 47064 201466 47076
rect 247402 47064 247408 47076
rect 247460 47104 247466 47116
rect 285582 47104 285588 47116
rect 247460 47076 285588 47104
rect 247460 47064 247466 47076
rect 285582 47064 285588 47076
rect 285640 47064 285646 47116
rect 285692 47104 285720 47212
rect 309410 47200 309416 47252
rect 309468 47240 309474 47252
rect 352558 47240 352564 47252
rect 309468 47212 352564 47240
rect 309468 47200 309474 47212
rect 352558 47200 352564 47212
rect 352616 47200 352622 47252
rect 364242 47200 364248 47252
rect 364300 47240 364306 47252
rect 407390 47240 407396 47252
rect 364300 47212 407396 47240
rect 364300 47200 364306 47212
rect 407390 47200 407396 47212
rect 407448 47200 407454 47252
rect 416774 47200 416780 47252
rect 416832 47240 416838 47252
rect 417234 47240 417240 47252
rect 416832 47212 417240 47240
rect 416832 47200 416838 47212
rect 417234 47200 417240 47212
rect 417292 47240 417298 47252
rect 418062 47240 418068 47252
rect 417292 47212 418068 47240
rect 417292 47200 417298 47212
rect 418062 47200 418068 47212
rect 418120 47200 418126 47252
rect 419074 47200 419080 47252
rect 419132 47240 419138 47252
rect 462130 47240 462136 47252
rect 419132 47212 462136 47240
rect 419132 47200 419138 47212
rect 462130 47200 462136 47212
rect 462188 47200 462194 47252
rect 473814 47200 473820 47252
rect 473872 47240 473878 47252
rect 516962 47240 516968 47252
rect 473872 47212 516968 47240
rect 473872 47200 473878 47212
rect 516962 47200 516968 47212
rect 517020 47200 517026 47252
rect 299474 47132 299480 47184
rect 299532 47172 299538 47184
rect 305730 47172 305736 47184
rect 299532 47144 305736 47172
rect 299532 47132 299538 47144
rect 305730 47132 305736 47144
rect 305788 47172 305794 47184
rect 351914 47172 351920 47184
rect 305788 47144 351920 47172
rect 305788 47132 305794 47144
rect 351914 47132 351920 47144
rect 351972 47132 351978 47184
rect 360562 47132 360568 47184
rect 360620 47172 360626 47184
rect 406746 47172 406752 47184
rect 360620 47144 406752 47172
rect 360620 47132 360626 47144
rect 406746 47132 406752 47144
rect 406804 47132 406810 47184
rect 468294 47172 468300 47184
rect 417896 47144 468300 47172
rect 417896 47116 417924 47144
rect 468294 47132 468300 47144
rect 468352 47172 468358 47184
rect 527450 47172 527456 47184
rect 468352 47144 527456 47172
rect 468352 47132 468358 47144
rect 527450 47132 527456 47144
rect 527508 47132 527514 47184
rect 303890 47104 303896 47116
rect 285692 47076 303896 47104
rect 303890 47064 303896 47076
rect 303948 47104 303954 47116
rect 308214 47104 308220 47116
rect 303948 47076 308220 47104
rect 303948 47064 303954 47076
rect 308214 47064 308220 47076
rect 308272 47104 308278 47116
rect 358722 47104 358728 47116
rect 308272 47076 358728 47104
rect 308272 47064 308278 47076
rect 358722 47064 358728 47076
rect 358780 47104 358786 47116
rect 363046 47104 363052 47116
rect 358780 47076 363052 47104
rect 358780 47064 358786 47076
rect 363046 47064 363052 47076
rect 363104 47104 363110 47116
rect 413554 47104 413560 47116
rect 363104 47076 413560 47104
rect 363104 47064 363110 47076
rect 413554 47064 413560 47076
rect 413612 47104 413618 47116
rect 417878 47104 417884 47116
rect 413612 47076 417884 47104
rect 413612 47064 413618 47076
rect 417878 47064 417884 47076
rect 417936 47064 417942 47116
rect 417970 47064 417976 47116
rect 418028 47104 418034 47116
rect 468938 47104 468944 47116
rect 418028 47076 468944 47104
rect 418028 47064 418034 47076
rect 468938 47064 468944 47076
rect 468996 47104 469002 47116
rect 523770 47104 523776 47116
rect 468996 47076 523776 47104
rect 468996 47064 469002 47076
rect 523770 47064 523776 47076
rect 523828 47104 523834 47116
rect 569126 47104 569132 47116
rect 523828 47076 569132 47104
rect 523828 47064 523834 47076
rect 569126 47064 569132 47076
rect 569184 47064 569190 47116
rect 201586 47036 201592 47048
rect 198752 47008 201592 47036
rect 198752 46968 198780 47008
rect 201586 46996 201592 47008
rect 201644 47036 201650 47048
rect 217962 47036 217968 47048
rect 201644 47008 217968 47036
rect 201644 46996 201650 47008
rect 217962 46996 217968 47008
rect 218020 46996 218026 47048
rect 198660 46940 198780 46968
rect 514478 46928 514484 46980
rect 514536 46968 514542 46980
rect 522482 46968 522488 46980
rect 514536 46940 522488 46968
rect 514536 46928 514542 46940
rect 522482 46928 522488 46940
rect 522540 46928 522546 46980
rect 526806 46928 526812 46980
rect 526864 46968 526870 46980
rect 634814 46968 634820 46980
rect 526864 46940 634820 46968
rect 526864 46928 526870 46940
rect 634814 46928 634820 46940
rect 634872 46928 634878 46980
rect 42242 45636 42248 45688
rect 42300 45676 42306 45688
rect 145098 45676 145104 45688
rect 42300 45648 145104 45676
rect 42300 45636 42306 45648
rect 145098 45636 145104 45648
rect 145156 45636 145162 45688
rect 42702 45568 42708 45620
rect 42760 45608 42766 45620
rect 140958 45608 140964 45620
rect 42760 45580 140964 45608
rect 42760 45568 42766 45580
rect 140958 45568 140964 45580
rect 141016 45568 141022 45620
rect 242894 45500 242900 45552
rect 242952 45540 242958 45552
rect 297726 45540 297732 45552
rect 242952 45512 297732 45540
rect 242952 45500 242958 45512
rect 297726 45500 297732 45512
rect 297784 45500 297790 45552
rect 579154 45500 579160 45552
rect 579212 45540 579218 45552
rect 673454 45540 673460 45552
rect 579212 45512 673460 45540
rect 579212 45500 579218 45512
rect 673454 45500 673460 45512
rect 673512 45500 673518 45552
rect 145098 44208 145104 44260
rect 145156 44248 145162 44260
rect 195330 44248 195336 44260
rect 145156 44220 195336 44248
rect 145156 44208 145162 44220
rect 195330 44208 195336 44220
rect 195388 44208 195394 44260
rect 140958 44140 140964 44192
rect 141016 44180 141022 44192
rect 254026 44180 254032 44192
rect 141016 44152 254032 44180
rect 141016 44140 141022 44152
rect 254026 44140 254032 44152
rect 254084 44180 254090 44192
rect 569218 44180 569224 44192
rect 254084 44152 569224 44180
rect 254084 44140 254090 44152
rect 569218 44140 569224 44152
rect 569276 44140 569282 44192
rect 299474 42004 299480 42016
rect 296916 41976 299480 42004
rect 296916 41948 296944 41976
rect 299474 41964 299480 41976
rect 299532 41964 299538 42016
rect 302234 41964 302240 42016
rect 302292 42004 302298 42016
rect 304994 42004 305000 42016
rect 302292 41976 305000 42004
rect 302292 41964 302298 41976
rect 304994 41964 305000 41976
rect 305052 41964 305058 42016
rect 411530 42004 411536 42016
rect 410260 41976 411536 42004
rect 410260 41948 410288 41976
rect 411530 41964 411536 41976
rect 411588 42004 411594 42016
rect 414566 42004 414572 42016
rect 411588 41976 414572 42004
rect 411588 41964 411594 41976
rect 414566 41964 414572 41976
rect 414624 42004 414630 42016
rect 415854 42004 415860 42016
rect 414624 41976 415860 42004
rect 414624 41964 414630 41976
rect 415854 41964 415860 41976
rect 415912 42004 415918 42016
rect 418246 42004 418252 42016
rect 415912 41976 418252 42004
rect 415912 41964 415918 41976
rect 418246 41964 418252 41976
rect 418304 41964 418310 42016
rect 466362 42004 466368 42016
rect 465092 41976 466368 42004
rect 465092 41948 465120 41976
rect 466362 41964 466368 41976
rect 466420 42004 466426 42016
rect 469398 42004 469404 42016
rect 466420 41976 469404 42004
rect 466420 41964 466426 41976
rect 469398 41964 469404 41976
rect 469456 42004 469462 42016
rect 470686 42004 470692 42016
rect 469456 41976 470692 42004
rect 469456 41964 469462 41976
rect 470686 41964 470692 41976
rect 470744 42004 470750 42016
rect 473078 42004 473084 42016
rect 470744 41976 473084 42004
rect 470744 41964 470750 41976
rect 473078 41964 473084 41976
rect 473136 41964 473142 42016
rect 296898 41936 296904 41948
rect 295352 41908 296904 41936
rect 189258 41828 189264 41880
rect 189316 41868 189322 41880
rect 191098 41868 191104 41880
rect 189316 41840 191104 41868
rect 189316 41828 189322 41840
rect 191098 41828 191104 41840
rect 191156 41868 191162 41880
rect 192294 41868 192300 41880
rect 191156 41840 192300 41868
rect 191156 41828 191162 41840
rect 192294 41828 192300 41840
rect 192352 41868 192358 41880
rect 192352 41840 193628 41868
rect 192352 41828 192358 41840
rect 193600 41812 193628 41840
rect 195422 41828 195428 41880
rect 195480 41868 195486 41880
rect 199562 41868 199568 41880
rect 195480 41840 199568 41868
rect 195480 41828 195486 41840
rect 199562 41828 199568 41840
rect 199620 41828 199626 41880
rect 193582 41760 193588 41812
rect 193640 41800 193646 41812
rect 196434 41800 196440 41812
rect 193640 41772 196440 41800
rect 193640 41760 193646 41772
rect 196434 41760 196440 41772
rect 196492 41760 196498 41812
rect 198458 41760 198464 41812
rect 198516 41800 198522 41812
rect 200114 41800 200120 41812
rect 198516 41772 200120 41800
rect 198516 41760 198522 41772
rect 200114 41760 200120 41772
rect 200172 41760 200178 41812
rect 253934 41556 253940 41608
rect 253992 41596 253998 41608
rect 253992 41568 256740 41596
rect 253992 41556 253998 41568
rect 256712 41528 256740 41568
rect 256712 41500 275968 41528
rect 275940 41460 275968 41500
rect 295352 41460 295380 41908
rect 296898 41896 296904 41908
rect 296956 41896 296962 41948
rect 352650 41896 352656 41948
rect 352708 41936 352714 41948
rect 355502 41936 355508 41948
rect 352708 41908 355508 41936
rect 352708 41896 352714 41908
rect 355502 41896 355508 41908
rect 355560 41896 355566 41948
rect 356974 41896 356980 41948
rect 357032 41936 357038 41948
rect 359826 41936 359832 41948
rect 357032 41908 359832 41936
rect 357032 41896 357038 41908
rect 359826 41896 359832 41908
rect 359884 41936 359890 41948
rect 361114 41936 361120 41948
rect 359884 41908 361120 41936
rect 359884 41896 359890 41908
rect 361114 41896 361120 41908
rect 361172 41896 361178 41948
rect 407482 41896 407488 41948
rect 407540 41936 407546 41948
rect 410242 41936 410248 41948
rect 407540 41908 410248 41936
rect 407540 41896 407546 41908
rect 410242 41896 410248 41908
rect 410300 41896 410306 41948
rect 411162 41896 411168 41948
rect 411220 41936 411226 41948
rect 411220 41908 415624 41936
rect 411220 41896 411226 41908
rect 297910 41828 297916 41880
rect 297968 41868 297974 41880
rect 300670 41868 300676 41880
rect 297968 41840 300676 41868
rect 297968 41828 297974 41840
rect 300670 41828 300676 41840
rect 300728 41828 300734 41880
rect 352006 41828 352012 41880
rect 352064 41868 352070 41880
rect 354306 41868 354312 41880
rect 352064 41840 354312 41868
rect 352064 41828 352070 41840
rect 354306 41828 354312 41840
rect 354364 41868 354370 41880
rect 360470 41868 360476 41880
rect 354364 41840 360476 41868
rect 354364 41828 354370 41840
rect 360470 41828 360476 41840
rect 360528 41828 360534 41880
rect 295426 41760 295432 41812
rect 295484 41800 295490 41812
rect 303154 41800 303160 41812
rect 295484 41772 303160 41800
rect 295484 41760 295490 41772
rect 303154 41760 303160 41772
rect 303212 41760 303218 41812
rect 305270 41760 305276 41812
rect 305328 41800 305334 41812
rect 306558 41800 306564 41812
rect 305328 41772 306564 41800
rect 305328 41760 305334 41772
rect 306558 41760 306564 41772
rect 306616 41800 306622 41812
rect 308674 41800 308680 41812
rect 306616 41772 308680 41800
rect 306616 41760 306622 41772
rect 308674 41760 308680 41772
rect 308732 41760 308738 41812
rect 350166 41760 350172 41812
rect 350224 41800 350230 41812
rect 357986 41800 357992 41812
rect 350224 41772 357992 41800
rect 350224 41760 350230 41772
rect 357986 41760 357992 41772
rect 358044 41760 358050 41812
rect 361132 41800 361160 41896
rect 409322 41828 409328 41880
rect 409380 41868 409386 41880
rect 412358 41868 412364 41880
rect 409380 41840 412364 41868
rect 409380 41828 409386 41840
rect 412358 41828 412364 41840
rect 412416 41868 412422 41880
rect 415486 41868 415492 41880
rect 412416 41840 415492 41868
rect 412416 41828 412422 41840
rect 415486 41828 415492 41840
rect 415544 41828 415550 41880
rect 415596 41868 415624 41908
rect 462314 41896 462320 41948
rect 462372 41936 462378 41948
rect 465074 41936 465080 41948
rect 462372 41908 465080 41936
rect 462372 41896 462378 41908
rect 465074 41896 465080 41908
rect 465132 41896 465138 41948
rect 465994 41896 466000 41948
rect 466052 41936 466058 41948
rect 474366 41936 474372 41948
rect 466052 41908 474372 41936
rect 466052 41896 466058 41908
rect 474366 41896 474372 41908
rect 474424 41896 474430 41948
rect 523218 41896 523224 41948
rect 523276 41936 523282 41948
rect 527358 41936 527364 41948
rect 523276 41908 527364 41936
rect 523276 41896 523282 41908
rect 527358 41896 527364 41908
rect 527416 41896 527422 41948
rect 419534 41868 419540 41880
rect 415596 41840 419540 41868
rect 419534 41828 419540 41840
rect 419592 41828 419598 41880
rect 459830 41828 459836 41880
rect 459888 41868 459894 41880
rect 467558 41868 467564 41880
rect 459888 41840 467564 41868
rect 459888 41828 459894 41840
rect 467558 41828 467564 41840
rect 467616 41828 467622 41880
rect 468478 41828 468484 41880
rect 468536 41868 468542 41880
rect 472526 41868 472532 41880
rect 468536 41840 472532 41868
rect 468536 41828 468542 41840
rect 472526 41828 472532 41840
rect 472584 41828 472590 41880
rect 518894 41828 518900 41880
rect 518952 41868 518958 41880
rect 524874 41868 524880 41880
rect 518952 41840 524880 41868
rect 518952 41828 518958 41840
rect 524874 41828 524880 41840
rect 524932 41828 524938 41880
rect 363506 41800 363512 41812
rect 361132 41772 363512 41800
rect 363506 41760 363512 41772
rect 363564 41760 363570 41812
rect 404998 41760 405004 41812
rect 405056 41800 405062 41812
rect 412726 41800 412732 41812
rect 405056 41772 412732 41800
rect 405056 41760 405062 41772
rect 412726 41760 412732 41772
rect 412784 41760 412790 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
rect 517054 41760 517060 41812
rect 517112 41800 517118 41812
rect 520090 41800 520096 41812
rect 517112 41772 520096 41800
rect 517112 41760 517118 41772
rect 520090 41760 520096 41772
rect 520148 41800 520154 41812
rect 521378 41800 521384 41812
rect 520148 41772 521384 41800
rect 520148 41760 520154 41772
rect 521378 41760 521384 41772
rect 521436 41800 521442 41812
rect 524414 41800 524420 41812
rect 521436 41772 524420 41800
rect 521436 41760 521442 41772
rect 524414 41760 524420 41772
rect 524472 41800 524478 41812
rect 525702 41800 525708 41812
rect 524472 41772 525708 41800
rect 524472 41760 524478 41772
rect 525702 41760 525708 41772
rect 525760 41800 525766 41812
rect 527910 41800 527916 41812
rect 525760 41772 527916 41800
rect 525760 41760 525766 41772
rect 527910 41760 527916 41772
rect 527968 41760 527974 41812
rect 275940 41432 295380 41460
rect 133092 40196 133098 40248
rect 133150 40236 133156 40248
rect 143810 40236 143816 40248
rect 133150 40208 143816 40236
rect 133150 40196 133156 40208
rect 143810 40196 143816 40208
rect 143868 40196 143874 40248
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143066 40100 143072 40112
rect 141048 40072 143072 40100
rect 141048 40060 141054 40072
rect 142586 39950 142614 40072
rect 143066 40060 143072 40072
rect 143124 40100 143130 40112
rect 143350 40100 143356 40112
rect 143124 40072 143356 40100
rect 143124 40060 143130 40072
rect 143350 40060 143356 40072
rect 143408 40100 143414 40112
rect 143408 40072 144684 40100
rect 143408 40060 143414 40072
rect 144656 39984 144684 40072
rect 252094 39652 252100 39704
rect 252152 39692 252158 39704
rect 254026 39692 254032 39704
rect 252152 39664 254032 39692
rect 252152 39652 252158 39664
rect 254026 39652 254032 39664
rect 254084 39652 254090 39704
<< via1 >>
rect 84016 995596 84068 995648
rect 91744 995596 91796 995648
rect 238208 995596 238260 995648
rect 245936 995596 245988 995648
rect 531964 995596 532016 995648
rect 539692 995596 539744 995648
rect 135352 995460 135404 995512
rect 143172 995460 143224 995512
rect 633808 995460 633860 995512
rect 641536 995460 641588 995512
rect 289636 995256 289688 995308
rect 297640 995256 297692 995308
rect 391480 995256 391532 995308
rect 399484 995256 399536 995308
rect 480444 995256 480496 995308
rect 488448 995256 488500 995308
rect 231860 995052 231912 995104
rect 244188 995052 244240 995104
rect 463792 992264 463844 992316
rect 475476 992264 475528 992316
rect 482928 992264 482980 992316
rect 141424 992060 141476 992112
rect 154396 992060 154448 992112
rect 130292 990836 130344 990888
rect 79048 990768 79100 990820
rect 110420 990768 110472 990820
rect 130108 990768 130160 990820
rect 419540 990836 419592 990888
rect 438676 990836 438728 990888
rect 450268 990836 450320 990888
rect 463608 990836 463660 990888
rect 143264 990768 143316 990820
rect 173808 990768 173860 990820
rect 179328 990768 179380 990820
rect 246948 990768 247000 990820
rect 284668 990768 284720 990820
rect 286968 990768 287020 990820
rect 391756 990768 391808 990820
rect 476120 990768 476172 990820
rect 527548 990768 527600 990820
rect 629300 990768 629352 990820
rect 187608 990700 187660 990752
rect 187700 990700 187752 990752
rect 202880 990700 202932 990752
rect 233056 990700 233108 990752
rect 244188 990700 244240 990752
rect 295800 990700 295852 990752
rect 386328 990700 386380 990752
rect 482928 990700 482980 990752
rect 526904 990700 526956 990752
rect 628656 990700 628708 990752
rect 79508 990632 79560 990684
rect 79968 990632 80020 990684
rect 130936 990632 130988 990684
rect 182364 990632 182416 990684
rect 233700 990632 233752 990684
rect 285312 990632 285364 990684
rect 333520 990632 333572 990684
rect 387156 990632 387208 990684
rect 391756 990632 391808 990684
rect 89996 990564 90048 990616
rect 110512 990564 110564 990616
rect 130108 990564 130160 990616
rect 179328 990564 179380 990616
rect 181720 990564 181772 990616
rect 186688 990564 186740 990616
rect 194692 990564 194744 990616
rect 386512 990564 386564 990616
rect 164148 990496 164200 990548
rect 192852 990496 192904 990548
rect 193220 990496 193272 990548
rect 212448 990496 212500 990548
rect 231860 990496 231912 990548
rect 286968 990496 287020 990548
rect 596088 990632 596140 990684
rect 419540 990564 419592 990616
rect 438768 990564 438820 990616
rect 450268 990564 450320 990616
rect 469312 990564 469364 990616
rect 141332 990428 141384 990480
rect 143264 990428 143316 990480
rect 160100 990428 160152 990480
rect 181720 990428 181772 990480
rect 187608 990428 187660 990480
rect 187700 990428 187752 990480
rect 202880 990428 202932 990480
rect 233056 990428 233108 990480
rect 246948 990428 247000 990480
rect 469036 990496 469088 990548
rect 483020 990496 483072 990548
rect 560208 990496 560260 990548
rect 576860 990564 576912 990616
rect 623688 990564 623740 990616
rect 623872 990496 623924 990548
rect 639788 990496 639840 990548
rect 154396 990360 154448 990412
rect 154580 990360 154632 990412
rect 386328 990360 386380 990412
rect 397644 990360 397696 990412
rect 424968 990360 425020 990412
rect 540980 990428 541032 990480
rect 483020 990360 483072 990412
rect 486608 990360 486660 990412
rect 507768 990292 507820 990344
rect 507860 990292 507912 990344
rect 521660 990360 521712 990412
rect 540888 990360 540940 990412
rect 154580 990224 154632 990276
rect 164148 990224 164200 990276
rect 397644 990224 397696 990276
rect 405740 990224 405792 990276
rect 521660 990224 521712 990276
rect 537852 990224 537904 990276
rect 540888 990224 540940 990276
rect 42248 990156 42300 990208
rect 79968 990156 80020 990208
rect 639788 990156 639840 990208
rect 673644 990156 673696 990208
rect 42432 990088 42484 990140
rect 79048 990088 79100 990140
rect 89996 990088 90048 990140
rect 405740 990088 405792 990140
rect 424968 990088 425020 990140
rect 628656 990088 628708 990140
rect 629300 990088 629352 990140
rect 673552 990088 673604 990140
rect 42524 990020 42576 990072
rect 673460 990020 673512 990072
rect 41788 969348 41840 969400
rect 42340 969348 42392 969400
rect 41788 968464 41840 968516
rect 42524 968464 42576 968516
rect 673460 965268 673512 965320
rect 675392 965268 675444 965320
rect 673552 964724 673604 964776
rect 675392 964724 675444 964776
rect 41788 962412 41840 962464
rect 42340 962412 42392 962464
rect 41788 956428 41840 956480
rect 42432 956428 42484 956480
rect 673644 953300 673696 953352
rect 675392 953300 675444 953352
rect 44272 930112 44324 930164
rect 45468 930112 45520 930164
rect 39672 922904 39724 922956
rect 44272 922904 44324 922956
rect 39856 914676 39908 914728
rect 41420 914676 41472 914728
rect 42248 914676 42300 914728
rect 673552 910732 673604 910784
rect 677784 910732 677836 910784
rect 673184 908012 673236 908064
rect 673460 908012 673512 908064
rect 673184 888768 673236 888820
rect 673460 888768 673512 888820
rect 39856 879792 39908 879844
rect 40132 879792 40184 879844
rect 44180 879792 44232 879844
rect 45836 879792 45888 879844
rect 41420 875576 41472 875628
rect 42248 875576 42300 875628
rect 673552 875508 673604 875560
rect 675392 875508 675444 875560
rect 673644 875032 673696 875084
rect 673644 874896 673696 874948
rect 673736 869388 673788 869440
rect 675208 869388 675260 869440
rect 673644 864968 673696 865020
rect 673828 864968 673880 865020
rect 675392 864968 675444 865020
rect 673552 836272 673604 836324
rect 673644 836204 673696 836256
rect 673552 830764 673604 830816
rect 673644 830764 673696 830816
rect 673552 821040 673604 821092
rect 674104 821040 674156 821092
rect 42248 807304 42300 807356
rect 42708 807304 42760 807356
rect 44548 805944 44600 805996
rect 44732 805944 44784 805996
rect 41788 798328 41840 798380
rect 42524 798328 42576 798380
rect 674104 797580 674156 797632
rect 675300 797580 675352 797632
rect 41788 787856 41840 787908
rect 42432 787856 42484 787908
rect 42708 787856 42760 787908
rect 42248 787176 42300 787228
rect 42616 787176 42668 787228
rect 674012 786428 674064 786480
rect 675300 786428 675352 786480
rect 673644 785272 673696 785324
rect 675392 785272 675444 785324
rect 673000 778336 673052 778388
rect 673092 778200 673144 778252
rect 673460 774868 673512 774920
rect 673828 774868 673880 774920
rect 675392 774868 675444 774920
rect 672816 772760 672868 772812
rect 673092 772760 673144 772812
rect 42524 768612 42576 768664
rect 42708 768612 42760 768664
rect 673552 768612 673604 768664
rect 674012 768612 674064 768664
rect 41788 754468 41840 754520
rect 42524 754468 42576 754520
rect 42708 754468 42760 754520
rect 41788 744404 41840 744456
rect 42616 744404 42668 744456
rect 673552 741888 673604 741940
rect 674196 741888 674248 741940
rect 675392 741888 675444 741940
rect 673644 741344 673696 741396
rect 675392 741344 675444 741396
rect 673000 739712 673052 739764
rect 673184 739576 673236 739628
rect 673460 730124 673512 730176
rect 675392 730124 675444 730176
rect 673828 729988 673880 730040
rect 675116 729988 675168 730040
rect 674012 720400 674064 720452
rect 674196 720400 674248 720452
rect 41788 711288 41840 711340
rect 42524 711288 42576 711340
rect 674012 710676 674064 710728
rect 675300 710676 675352 710728
rect 42248 700952 42300 701004
rect 42524 700952 42576 701004
rect 41788 700816 41840 700868
rect 42616 700816 42668 700868
rect 673644 695920 673696 695972
rect 675392 695920 675444 695972
rect 673092 695512 673144 695564
rect 673184 695512 673236 695564
rect 44640 695444 44692 695496
rect 44916 695444 44968 695496
rect 673552 695308 673604 695360
rect 673828 695308 673880 695360
rect 675392 695308 675444 695360
rect 44732 676200 44784 676252
rect 44916 676200 44968 676252
rect 42340 669128 42392 669180
rect 41788 669060 41840 669112
rect 673184 662464 673236 662516
rect 44548 662396 44600 662448
rect 44732 662396 44784 662448
rect 673184 662328 673236 662380
rect 41788 657636 41840 657688
rect 42524 657636 42576 657688
rect 41788 657092 41840 657144
rect 42340 657092 42392 657144
rect 42616 657092 42668 657144
rect 44640 656820 44692 656872
rect 44824 656820 44876 656872
rect 673644 651720 673696 651772
rect 675392 651720 675444 651772
rect 673552 651108 673604 651160
rect 675392 651108 675444 651160
rect 673460 639684 673512 639736
rect 675392 639684 675444 639736
rect 672816 637508 672868 637560
rect 673092 637508 673144 637560
rect 42524 633496 42576 633548
rect 42524 633292 42576 633344
rect 42340 633224 42392 633276
rect 42616 633224 42668 633276
rect 41788 625880 41840 625932
rect 42432 625880 42484 625932
rect 672816 618264 672868 618316
rect 673000 618264 673052 618316
rect 41880 614456 41932 614508
rect 42248 614456 42300 614508
rect 42616 614456 42668 614508
rect 41788 614388 41840 614440
rect 42524 614388 42576 614440
rect 673644 606704 673696 606756
rect 675392 606704 675444 606756
rect 673552 605616 673604 605668
rect 675300 605616 675352 605668
rect 44640 604528 44692 604580
rect 44640 604392 44692 604444
rect 673552 604392 673604 604444
rect 673828 604392 673880 604444
rect 672816 598952 672868 599004
rect 673092 598952 673144 599004
rect 673460 594872 673512 594924
rect 675392 594872 675444 594924
rect 673092 585148 673144 585200
rect 673000 585080 673052 585132
rect 42248 584196 42300 584248
rect 42616 584196 42668 584248
rect 41788 581680 41840 581732
rect 42432 581680 42484 581732
rect 41788 572228 41840 572280
rect 42248 572228 42300 572280
rect 42524 572228 42576 572280
rect 41788 571616 41840 571668
rect 42616 571616 42668 571668
rect 672816 569916 672868 569968
rect 673000 569916 673052 569968
rect 673552 565836 673604 565888
rect 673920 565836 673972 565888
rect 673644 561484 673696 561536
rect 675392 561484 675444 561536
rect 672816 560260 672868 560312
rect 673000 560260 673052 560312
rect 673552 559920 673604 559972
rect 673920 559920 673972 559972
rect 675392 559920 675444 559972
rect 673460 550468 673512 550520
rect 675392 550468 675444 550520
rect 673000 546524 673052 546576
rect 673092 546320 673144 546372
rect 44732 540948 44784 541000
rect 44916 540948 44968 541000
rect 41788 538500 41840 538552
rect 42432 538500 42484 538552
rect 41788 528436 41840 528488
rect 42432 528436 42484 528488
rect 42616 528436 42668 528488
rect 673092 527144 673144 527196
rect 673184 527008 673236 527060
rect 673736 522928 673788 522980
rect 673920 522928 673972 522980
rect 673184 521568 673236 521620
rect 676128 521568 676180 521620
rect 44548 496816 44600 496868
rect 44732 496816 44784 496868
rect 673736 463632 673788 463684
rect 677692 463632 677744 463684
rect 39396 458192 39448 458244
rect 44272 458192 44324 458244
rect 673000 449896 673052 449948
rect 673368 449896 673420 449948
rect 39856 448264 39908 448316
rect 42248 448264 42300 448316
rect 676220 440172 676272 440224
rect 677692 440172 677744 440224
rect 42248 413380 42300 413432
rect 42616 413380 42668 413432
rect 672816 412496 672868 412548
rect 676220 412496 676272 412548
rect 41788 410932 41840 410984
rect 42524 410932 42576 410984
rect 672540 405628 672592 405680
rect 672724 405628 672776 405680
rect 673460 401548 673512 401600
rect 675300 401548 675352 401600
rect 41788 401480 41840 401532
rect 42248 401480 42300 401532
rect 42616 401480 42668 401532
rect 41972 400120 42024 400172
rect 42432 400120 42484 400172
rect 672540 386384 672592 386436
rect 672816 386384 672868 386436
rect 673552 384004 673604 384056
rect 675392 384004 675444 384056
rect 673644 382712 673696 382764
rect 675392 382712 675444 382764
rect 42340 380876 42392 380928
rect 42616 380876 42668 380928
rect 673828 372308 673880 372360
rect 675392 372308 675444 372360
rect 41788 368636 41840 368688
rect 42524 368636 42576 368688
rect 42524 367004 42576 367056
rect 42800 366936 42852 366988
rect 41788 357484 41840 357536
rect 42340 357484 42392 357536
rect 42616 357484 42668 357536
rect 41788 356668 41840 356720
rect 42432 356668 42484 356720
rect 672632 353336 672684 353388
rect 672540 353200 672592 353252
rect 42708 347692 42760 347744
rect 42892 347692 42944 347744
rect 672540 347692 672592 347744
rect 672724 347692 672776 347744
rect 673644 338512 673696 338564
rect 675392 338512 675444 338564
rect 42340 334636 42392 334688
rect 42616 334636 42668 334688
rect 42616 328448 42668 328500
rect 42892 328448 42944 328500
rect 672448 328448 672500 328500
rect 672724 328448 672776 328500
rect 673828 327088 673880 327140
rect 675392 327088 675444 327140
rect 41788 324504 41840 324556
rect 42524 324436 42576 324488
rect 42340 314576 42392 314628
rect 42616 314508 42668 314560
rect 41788 314440 41840 314492
rect 42524 314440 42576 314492
rect 42800 314440 42852 314492
rect 41788 313760 41840 313812
rect 42432 313760 42484 313812
rect 672540 309068 672592 309120
rect 672816 309068 672868 309120
rect 42432 307912 42484 307964
rect 42708 307912 42760 307964
rect 673460 304920 673512 304972
rect 673828 304920 673880 304972
rect 42616 295332 42668 295384
rect 42800 295332 42852 295384
rect 673644 293496 673696 293548
rect 675024 293496 675076 293548
rect 673828 293156 673880 293208
rect 675392 293156 675444 293208
rect 672632 289824 672684 289876
rect 672816 289824 672868 289876
rect 673460 283024 673512 283076
rect 674932 283024 674984 283076
rect 675392 283024 675444 283076
rect 41788 282276 41840 282328
rect 42432 282276 42484 282328
rect 42616 282276 42668 282328
rect 42708 282208 42760 282260
rect 42708 282004 42760 282056
rect 673920 276020 673972 276072
rect 675208 276020 675260 276072
rect 42524 275952 42576 276004
rect 42800 275952 42852 276004
rect 41788 270784 41840 270836
rect 42524 270784 42576 270836
rect 41788 270240 41840 270292
rect 42340 270240 42392 270292
rect 42708 270240 42760 270292
rect 673736 266296 673788 266348
rect 674932 266296 674984 266348
rect 673828 248140 673880 248192
rect 675392 248140 675444 248192
rect 673644 247460 673696 247512
rect 673920 247460 673972 247512
rect 675392 247460 675444 247512
rect 42340 246984 42392 247036
rect 42708 246984 42760 247036
rect 41788 239028 41840 239080
rect 42432 239028 42484 239080
rect 42616 239028 42668 239080
rect 673736 237668 673788 237720
rect 675392 237668 675444 237720
rect 41788 228624 41840 228676
rect 42524 228624 42576 228676
rect 41788 228012 41840 228064
rect 42432 228012 42484 228064
rect 42708 228012 42760 228064
rect 42248 227876 42300 227928
rect 42524 227876 42576 227928
rect 672724 212508 672776 212560
rect 672908 212508 672960 212560
rect 673552 203872 673604 203924
rect 673828 203872 673880 203924
rect 675392 203872 675444 203924
rect 673460 203328 673512 203380
rect 673644 203328 673696 203380
rect 675392 203328 675444 203380
rect 672540 198704 672592 198756
rect 672724 198704 672776 198756
rect 41788 196732 41840 196784
rect 42340 196732 42392 196784
rect 41788 195848 41840 195900
rect 42616 195848 42668 195900
rect 44640 195848 44692 195900
rect 673736 191972 673788 192024
rect 674012 191972 674064 192024
rect 41788 189796 41840 189848
rect 42340 189796 42392 189848
rect 42248 184220 42300 184272
rect 42432 184220 42484 184272
rect 44456 173884 44508 173936
rect 44732 173884 44784 173936
rect 672724 173884 672776 173936
rect 672908 173884 672960 173936
rect 673828 173884 673880 173936
rect 674012 173884 674064 173936
rect 44732 160148 44784 160200
rect 672540 160080 672592 160132
rect 672724 160080 672776 160132
rect 673644 160080 673696 160132
rect 673828 160080 673880 160132
rect 44640 160012 44692 160064
rect 673552 158312 673604 158364
rect 675392 158312 675444 158364
rect 673460 157292 673512 157344
rect 675392 157292 675444 157344
rect 44640 154504 44692 154556
rect 44732 154504 44784 154556
rect 673644 147840 673696 147892
rect 674012 147840 674064 147892
rect 675392 147840 675444 147892
rect 44732 140768 44784 140820
rect 44640 140700 44692 140752
rect 44732 121524 44784 121576
rect 44640 121388 44692 121440
rect 672724 115880 672776 115932
rect 672816 115880 672868 115932
rect 673552 112752 673604 112804
rect 675392 112752 675444 112804
rect 673460 112072 673512 112124
rect 675392 112072 675444 112124
rect 672816 102144 672868 102196
rect 673644 102144 673696 102196
rect 673828 102144 673880 102196
rect 672724 102076 672776 102128
rect 673644 102008 673696 102060
rect 675392 102008 675444 102060
rect 44272 96568 44324 96620
rect 44548 96568 44600 96620
rect 672816 82900 672868 82952
rect 672816 82696 672868 82748
rect 44272 77256 44324 77308
rect 44364 77256 44416 77308
rect 39672 75216 39724 75268
rect 39672 74944 39724 74996
rect 39580 67940 39632 67992
rect 41420 67940 41472 67992
rect 41420 64608 41472 64660
rect 42708 64608 42760 64660
rect 39672 52368 39724 52420
rect 39856 52368 39908 52420
rect 45468 47880 45520 47932
rect 179420 47880 179472 47932
rect 518808 47880 518860 47932
rect 673644 47880 673696 47932
rect 39856 47812 39908 47864
rect 189172 47812 189224 47864
rect 527456 47812 527508 47864
rect 673552 47812 673604 47864
rect 45560 47744 45612 47796
rect 149060 47744 149112 47796
rect 528652 47744 528704 47796
rect 672816 47744 672868 47796
rect 39764 47676 39816 47728
rect 86316 47676 86368 47728
rect 179420 47472 179472 47524
rect 195980 47540 196032 47592
rect 198648 47540 198700 47592
rect 198740 47540 198792 47592
rect 212540 47608 212592 47660
rect 270500 47608 270552 47660
rect 303620 47540 303672 47592
rect 304540 47540 304592 47592
rect 359372 47540 359424 47592
rect 361488 47540 361540 47592
rect 231768 47472 231820 47524
rect 251180 47472 251232 47524
rect 270408 47472 270460 47524
rect 289728 47404 289780 47456
rect 86316 47336 86368 47388
rect 199016 47336 199068 47388
rect 201408 47336 201460 47388
rect 251180 47336 251232 47388
rect 270408 47336 270460 47388
rect 364156 47404 364208 47456
rect 416780 47472 416832 47524
rect 303620 47336 303672 47388
rect 361488 47336 361540 47388
rect 414204 47336 414256 47388
rect 417976 47336 418028 47388
rect 418068 47336 418120 47388
rect 471980 47336 472032 47388
rect 526812 47336 526864 47388
rect 199660 47268 199712 47320
rect 217968 47200 218020 47252
rect 240140 47200 240192 47252
rect 285588 47268 285640 47320
rect 307576 47268 307628 47320
rect 362408 47268 362460 47320
rect 364156 47268 364208 47320
rect 406752 47268 406804 47320
rect 461492 47268 461544 47320
rect 516324 47268 516376 47320
rect 518808 47268 518860 47320
rect 200856 47132 200908 47184
rect 242900 47132 242952 47184
rect 149060 47064 149112 47116
rect 154580 47064 154632 47116
rect 173808 46996 173860 47048
rect 188528 47064 188580 47116
rect 192852 47064 192904 47116
rect 186688 46928 186740 46980
rect 194692 46928 194744 46980
rect 201408 47064 201460 47116
rect 247408 47064 247460 47116
rect 285588 47064 285640 47116
rect 309416 47200 309468 47252
rect 352564 47200 352616 47252
rect 364248 47200 364300 47252
rect 407396 47200 407448 47252
rect 416780 47200 416832 47252
rect 417240 47200 417292 47252
rect 418068 47200 418120 47252
rect 419080 47200 419132 47252
rect 462136 47200 462188 47252
rect 473820 47200 473872 47252
rect 516968 47200 517020 47252
rect 299480 47132 299532 47184
rect 305736 47132 305788 47184
rect 351920 47132 351972 47184
rect 360568 47132 360620 47184
rect 406752 47132 406804 47184
rect 468300 47132 468352 47184
rect 527456 47132 527508 47184
rect 303896 47064 303948 47116
rect 308220 47064 308272 47116
rect 358728 47064 358780 47116
rect 363052 47064 363104 47116
rect 413560 47064 413612 47116
rect 417884 47064 417936 47116
rect 417976 47064 418028 47116
rect 468944 47064 468996 47116
rect 523776 47064 523828 47116
rect 569132 47064 569184 47116
rect 201592 46996 201644 47048
rect 217968 46996 218020 47048
rect 514484 46928 514536 46980
rect 522488 46928 522540 46980
rect 526812 46928 526864 46980
rect 634820 46928 634872 46980
rect 42248 45636 42300 45688
rect 145104 45636 145156 45688
rect 42708 45568 42760 45620
rect 140964 45568 141016 45620
rect 242900 45500 242952 45552
rect 297732 45500 297784 45552
rect 579160 45500 579212 45552
rect 673460 45500 673512 45552
rect 145104 44208 145156 44260
rect 195336 44208 195388 44260
rect 140964 44140 141016 44192
rect 254032 44140 254084 44192
rect 569224 44140 569276 44192
rect 299480 41964 299532 42016
rect 302240 41964 302292 42016
rect 305000 41964 305052 42016
rect 411536 41964 411588 42016
rect 414572 41964 414624 42016
rect 415860 41964 415912 42016
rect 418252 41964 418304 42016
rect 466368 41964 466420 42016
rect 469404 41964 469456 42016
rect 470692 41964 470744 42016
rect 473084 41964 473136 42016
rect 189264 41828 189316 41880
rect 191104 41828 191156 41880
rect 192300 41828 192352 41880
rect 195428 41828 195480 41880
rect 199568 41828 199620 41880
rect 193588 41760 193640 41812
rect 196440 41760 196492 41812
rect 198464 41760 198516 41812
rect 200120 41760 200172 41812
rect 253940 41556 253992 41608
rect 296904 41896 296956 41948
rect 352656 41896 352708 41948
rect 355508 41896 355560 41948
rect 356980 41896 357032 41948
rect 359832 41896 359884 41948
rect 361120 41896 361172 41948
rect 407488 41896 407540 41948
rect 410248 41896 410300 41948
rect 411168 41896 411220 41948
rect 297916 41828 297968 41880
rect 300676 41828 300728 41880
rect 352012 41828 352064 41880
rect 354312 41828 354364 41880
rect 360476 41828 360528 41880
rect 295432 41760 295484 41812
rect 303160 41760 303212 41812
rect 305276 41760 305328 41812
rect 306564 41760 306616 41812
rect 308680 41760 308732 41812
rect 350172 41760 350224 41812
rect 357992 41760 358044 41812
rect 409328 41828 409380 41880
rect 412364 41828 412416 41880
rect 415492 41828 415544 41880
rect 462320 41896 462372 41948
rect 465080 41896 465132 41948
rect 466000 41896 466052 41948
rect 474372 41896 474424 41948
rect 523224 41896 523276 41948
rect 527364 41896 527416 41948
rect 419540 41828 419592 41880
rect 459836 41828 459888 41880
rect 467564 41828 467616 41880
rect 468484 41828 468536 41880
rect 472532 41828 472584 41880
rect 518900 41828 518952 41880
rect 524880 41828 524932 41880
rect 363512 41760 363564 41812
rect 405004 41760 405056 41812
rect 412732 41760 412784 41812
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
rect 517060 41760 517112 41812
rect 520096 41760 520148 41812
rect 521384 41760 521436 41812
rect 524420 41760 524472 41812
rect 525708 41760 525760 41812
rect 527916 41760 527968 41812
rect 133098 40196 133150 40248
rect 143816 40196 143868 40248
rect 140996 40060 141048 40112
rect 143072 40060 143124 40112
rect 143356 40060 143408 40112
rect 252100 39652 252152 39704
rect 254032 39652 254084 39704
<< metal2 >>
rect 333518 997656 333574 997665
rect 333518 997591 333574 997600
rect 45926 996568 45982 996577
rect 45926 996503 45982 996512
rect 42248 990208 42300 990214
rect 42248 990150 42300 990156
rect 45466 990176 45522 990185
rect 41722 969870 41828 969898
rect 41800 969406 41828 969870
rect 41788 969400 41840 969406
rect 41788 969342 41840 969348
rect 41713 969217 42193 969273
rect 41788 968516 41840 968522
rect 41788 968458 41840 968464
rect 41800 968063 41828 968458
rect 41722 968035 41828 968063
rect 41713 967377 42193 967433
rect 41713 965537 42193 965593
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 41713 963053 42193 963109
rect 41713 962501 42193 962557
rect 41788 962464 41840 962470
rect 41788 962406 41840 962412
rect 41800 961874 41828 962406
rect 41722 961846 41828 961874
rect 41713 961213 42193 961269
rect 41713 960569 42193 960625
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 41713 958729 42193 958785
rect 41713 958177 42193 958233
rect 41722 957547 41920 957575
rect 41892 957386 41920 957547
rect 42260 957386 42288 990150
rect 42432 990140 42484 990146
rect 45466 990111 45522 990120
rect 42432 990082 42484 990088
rect 42340 969400 42392 969406
rect 42340 969342 42392 969348
rect 42352 962470 42380 969342
rect 42340 962464 42392 962470
rect 42340 962406 42392 962412
rect 41892 957358 42288 957386
rect 41722 956903 41828 956931
rect 41800 956486 41828 956903
rect 41788 956480 41840 956486
rect 41788 956422 41840 956428
rect 41713 956337 42193 956393
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 39330 922962 39712 922978
rect 39330 922956 39724 922962
rect 39330 922950 39672 922956
rect 39672 922898 39724 922904
rect 39567 919006 39896 919034
rect 39868 914734 39896 919006
rect 42260 914734 42288 957358
rect 42444 956486 42472 990082
rect 42524 990072 42576 990078
rect 42524 990014 42576 990020
rect 42536 968522 42564 990014
rect 42524 968516 42576 968522
rect 42524 968458 42576 968464
rect 42432 956480 42484 956486
rect 42432 956422 42484 956428
rect 39856 914728 39908 914734
rect 39856 914670 39908 914676
rect 41420 914728 41472 914734
rect 41420 914670 41472 914676
rect 42248 914728 42300 914734
rect 42248 914670 42300 914676
rect 39330 912206 39712 912234
rect 39684 908177 39712 912206
rect 39670 908168 39726 908177
rect 39670 908103 39726 908112
rect 40406 908032 40462 908041
rect 40406 907967 40462 907976
rect 40420 889001 40448 907967
rect 40406 888992 40462 889001
rect 40406 888927 40462 888936
rect 40130 880016 40186 880025
rect 39606 879974 39896 880002
rect 39868 879850 39896 879974
rect 40130 879951 40186 879960
rect 40144 879850 40172 879951
rect 39856 879844 39908 879850
rect 39856 879786 39908 879792
rect 40132 879844 40184 879850
rect 40132 879786 40184 879792
rect 41432 875634 41460 914670
rect 41420 875628 41472 875634
rect 41420 875570 41472 875576
rect 42248 875628 42300 875634
rect 42248 875570 42300 875576
rect 41432 875129 41460 875570
rect 41418 875120 41474 875129
rect 41418 875055 41474 875064
rect 39854 837584 39910 837593
rect 39854 837519 39910 837528
rect 39868 832697 39896 837519
rect 39854 832688 39910 832697
rect 39854 832623 39910 832632
rect 39606 827750 39712 827778
rect 39684 827529 39712 827750
rect 39670 827520 39726 827529
rect 39670 827455 39726 827464
rect 42260 807362 42288 875570
rect 42248 807356 42300 807362
rect 42248 807298 42300 807304
rect 41722 800075 41828 800103
rect 41800 799898 41828 800075
rect 41800 799870 42288 799898
rect 41713 799417 42193 799473
rect 41788 798380 41840 798386
rect 41788 798322 41840 798328
rect 41800 798266 41828 798322
rect 41722 798238 41828 798266
rect 41713 797577 42193 797633
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 42260 792282 42288 799870
rect 41800 792254 42288 792282
rect 41800 792099 41828 792254
rect 41722 792071 41828 792099
rect 41713 791413 42193 791469
rect 41713 790769 42193 790825
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 42444 788066 42472 956422
rect 42536 798386 42564 968458
rect 45480 930170 45508 990111
rect 44272 930164 44324 930170
rect 44272 930106 44324 930112
rect 45468 930164 45520 930170
rect 45468 930106 45520 930112
rect 44284 922962 44312 930106
rect 44272 922956 44324 922962
rect 44272 922898 44324 922904
rect 44180 879844 44232 879850
rect 44180 879786 44232 879792
rect 42708 807356 42760 807362
rect 42708 807298 42760 807304
rect 42524 798380 42576 798386
rect 42524 798322 42576 798328
rect 42260 788038 42472 788066
rect 41788 787908 41840 787914
rect 41788 787850 41840 787856
rect 41800 787794 41828 787850
rect 41722 787766 41828 787794
rect 42260 787250 42288 788038
rect 42432 787908 42484 787914
rect 42432 787850 42484 787856
rect 41800 787234 42288 787250
rect 41800 787228 42300 787234
rect 41800 787222 42248 787228
rect 41800 787114 41828 787222
rect 42248 787170 42300 787176
rect 42260 787139 42288 787170
rect 41722 787086 41828 787114
rect 42444 786978 42472 787850
rect 42260 786950 42472 786978
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 42260 757058 42288 786950
rect 42536 768670 42564 798322
rect 42720 787914 42748 807298
rect 42708 787908 42760 787914
rect 42708 787850 42760 787856
rect 42616 787228 42668 787234
rect 42616 787170 42668 787176
rect 42524 768664 42576 768670
rect 42524 768606 42576 768612
rect 42260 757030 42380 757058
rect 41722 756894 42288 756922
rect 41713 756217 42193 756273
rect 41722 755035 41828 755063
rect 41800 754526 41828 755035
rect 41788 754520 41840 754526
rect 41788 754462 41840 754468
rect 41713 754377 42193 754433
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 42260 749034 42288 756894
rect 41800 749006 42288 749034
rect 41800 748898 41828 749006
rect 41722 748870 41828 748898
rect 41713 748213 42193 748269
rect 41713 747569 42193 747625
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 42352 744682 42380 757030
rect 42524 754520 42576 754526
rect 42524 754462 42576 754468
rect 41800 744654 42380 744682
rect 41800 744575 41828 744654
rect 41722 744547 41828 744575
rect 41788 744456 41840 744462
rect 41788 744398 41840 744404
rect 41800 743931 41828 744398
rect 41722 743903 41828 743931
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 42260 713810 42288 744654
rect 42536 744546 42564 754462
rect 42352 744518 42564 744546
rect 42352 713946 42380 744518
rect 42628 744462 42656 787170
rect 42708 768664 42760 768670
rect 42708 768606 42760 768612
rect 42720 754526 42748 768606
rect 42708 754520 42760 754526
rect 42708 754462 42760 754468
rect 42616 744456 42668 744462
rect 42616 744398 42668 744404
rect 42352 713918 42564 713946
rect 42260 713782 42380 713810
rect 41722 713675 42288 713703
rect 41713 713017 42193 713073
rect 41722 711835 41828 711863
rect 41800 711346 41828 711835
rect 41788 711340 41840 711346
rect 41788 711282 41840 711288
rect 41713 711177 42193 711233
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 42260 705786 42288 713675
rect 41800 705758 42288 705786
rect 41800 705699 41828 705758
rect 42352 705699 42380 713782
rect 42536 711346 42564 713918
rect 42524 711340 42576 711346
rect 42524 711282 42576 711288
rect 41722 705671 41828 705699
rect 42260 705671 42380 705699
rect 41713 705013 42193 705069
rect 41713 704369 42193 704425
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 42260 701375 42288 705671
rect 42536 705514 42564 711282
rect 41722 701347 42288 701375
rect 42260 701010 42288 701347
rect 42352 705486 42564 705514
rect 42248 701004 42300 701010
rect 42248 700946 42300 700952
rect 41788 700868 41840 700874
rect 41788 700810 41840 700816
rect 41800 700754 41828 700810
rect 41722 700726 41828 700754
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41722 670475 42288 670503
rect 41713 669817 42193 669873
rect 41788 669112 41840 669118
rect 41788 669054 41840 669060
rect 41800 668658 41828 669054
rect 41722 668630 41828 668658
rect 41713 667977 42193 668033
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 42260 662538 42288 670475
rect 42352 669186 42380 705486
rect 42524 701004 42576 701010
rect 42524 700946 42576 700952
rect 42340 669180 42392 669186
rect 42340 669122 42392 669128
rect 41708 662510 42288 662538
rect 41708 662485 41736 662510
rect 42352 662499 42380 669122
rect 42352 662471 42472 662499
rect 41713 661813 42193 661869
rect 41713 661169 42193 661225
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41722 658158 41828 658186
rect 41800 657694 41828 658158
rect 41788 657688 41840 657694
rect 41788 657630 41840 657636
rect 41722 657478 41828 657506
rect 41800 657150 41828 657478
rect 41788 657144 41840 657150
rect 41788 657086 41840 657092
rect 42340 657144 42392 657150
rect 42340 657086 42392 657092
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 42352 633282 42380 657086
rect 42340 633276 42392 633282
rect 42340 633218 42392 633224
rect 41722 627286 42288 627314
rect 41713 626617 42193 626673
rect 41788 625932 41840 625938
rect 41788 625874 41840 625880
rect 41800 625463 41828 625874
rect 41722 625435 41828 625463
rect 41713 624777 42193 624833
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42260 619426 42288 627286
rect 42444 625938 42472 662471
rect 42536 657694 42564 700946
rect 42628 700874 42656 744398
rect 42616 700868 42668 700874
rect 42616 700810 42668 700816
rect 42524 657688 42576 657694
rect 42524 657630 42576 657636
rect 42536 633554 42564 657630
rect 42628 657150 42656 700810
rect 42616 657144 42668 657150
rect 42616 657086 42668 657092
rect 42524 633548 42576 633554
rect 42524 633490 42576 633496
rect 42524 633344 42576 633350
rect 42524 633286 42576 633292
rect 42432 625932 42484 625938
rect 42432 625874 42484 625880
rect 41800 619398 42288 619426
rect 41800 619290 41828 619398
rect 41722 619262 41828 619290
rect 41713 618613 42193 618669
rect 41713 617969 42193 618025
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41722 614947 41828 614975
rect 41800 614446 41828 614947
rect 41880 614508 41932 614514
rect 41880 614450 41932 614456
rect 42248 614508 42300 614514
rect 42248 614450 42300 614456
rect 41788 614440 41840 614446
rect 41788 614382 41840 614388
rect 41892 614331 41920 614450
rect 41722 614303 41920 614331
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 42260 584254 42288 614450
rect 42248 584248 42300 584254
rect 42248 584190 42300 584196
rect 41722 584075 42288 584103
rect 41713 583417 42193 583473
rect 41722 582235 41828 582263
rect 41800 581738 41828 582235
rect 41788 581732 41840 581738
rect 41788 581674 41840 581680
rect 41713 581577 42193 581633
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 42260 576178 42288 584075
rect 42444 581738 42472 625874
rect 42536 614446 42564 633286
rect 42616 633276 42668 633282
rect 42616 633218 42668 633224
rect 42628 614514 42656 633218
rect 42616 614508 42668 614514
rect 42616 614450 42668 614456
rect 42524 614440 42576 614446
rect 42524 614382 42576 614388
rect 42432 581732 42484 581738
rect 42432 581674 42484 581680
rect 41892 576150 42288 576178
rect 41892 576099 41920 576150
rect 41722 576071 41920 576099
rect 41713 575413 42193 575469
rect 41713 574769 42193 574825
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41788 572280 41840 572286
rect 41788 572222 41840 572228
rect 42248 572280 42300 572286
rect 42248 572222 42300 572228
rect 41800 571775 41828 572222
rect 41722 571747 41828 571775
rect 41788 571668 41840 571674
rect 41788 571610 41840 571616
rect 41800 571146 41828 571610
rect 41722 571118 41828 571146
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 42260 541090 42288 572222
rect 42260 541062 42380 541090
rect 41722 540875 42288 540903
rect 41713 540217 42193 540273
rect 41722 539022 41828 539050
rect 41800 538558 41828 539022
rect 41788 538552 41840 538558
rect 41788 538494 41840 538500
rect 41713 538377 42193 538433
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 42260 532930 42288 540875
rect 41708 532902 42288 532930
rect 41708 532885 41736 532902
rect 41713 532213 42193 532269
rect 41713 531569 42193 531625
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 42352 528850 42380 541062
rect 42444 538558 42472 581674
rect 42536 572286 42564 614382
rect 42616 584248 42668 584254
rect 42616 584190 42668 584196
rect 42524 572280 42576 572286
rect 42524 572222 42576 572228
rect 42628 571674 42656 584190
rect 42616 571668 42668 571674
rect 42616 571610 42668 571616
rect 42432 538552 42484 538558
rect 42484 538500 42564 538506
rect 42432 538494 42564 538500
rect 42444 538478 42564 538494
rect 41892 528822 42380 528850
rect 41892 528578 41920 528822
rect 41722 528550 41920 528578
rect 41788 528488 41840 528494
rect 41788 528430 41840 528436
rect 41800 527931 41828 528430
rect 41722 527903 41828 527931
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 39606 493190 39804 493218
rect 39776 492969 39804 493190
rect 39762 492960 39818 492969
rect 39762 492895 39818 492904
rect 39396 458244 39448 458250
rect 39396 458186 39448 458192
rect 39408 451874 39436 458186
rect 39946 455424 40002 455433
rect 39946 455359 40002 455368
rect 39670 451888 39726 451897
rect 39330 451846 39670 451874
rect 39670 451823 39726 451832
rect 39856 448316 39908 448322
rect 39856 448258 39908 448264
rect 39868 447794 39896 448258
rect 39567 447766 39896 447794
rect 39670 441008 39726 441017
rect 39330 440966 39670 440994
rect 39960 440994 39988 455359
rect 42260 448322 42288 528822
rect 42432 528488 42484 528494
rect 42432 528430 42484 528436
rect 42248 448316 42300 448322
rect 42248 448258 42300 448264
rect 39726 440966 39988 440994
rect 39670 440943 39726 440952
rect 42260 413438 42288 448258
rect 42248 413432 42300 413438
rect 42248 413374 42300 413380
rect 41722 413275 42288 413303
rect 41713 412617 42193 412673
rect 41722 411454 41828 411482
rect 41800 410990 41828 411454
rect 41788 410984 41840 410990
rect 41788 410926 41840 410932
rect 41713 410777 42193 410833
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 42260 405299 42288 413275
rect 41722 405271 42288 405299
rect 41713 404613 42193 404669
rect 41713 403969 42193 404025
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41788 401532 41840 401538
rect 41788 401474 41840 401480
rect 42248 401532 42300 401538
rect 42248 401474 42300 401480
rect 41800 400975 41828 401474
rect 41722 400947 41828 400975
rect 41722 400302 42012 400330
rect 41984 400178 42012 400302
rect 42260 400217 42288 401474
rect 42246 400208 42302 400217
rect 41972 400172 42024 400178
rect 42444 400178 42472 528430
rect 42536 410990 42564 538478
rect 42628 528494 42656 571610
rect 42616 528488 42668 528494
rect 42616 528430 42668 528436
rect 42616 413432 42668 413438
rect 42616 413374 42668 413380
rect 42524 410984 42576 410990
rect 42524 410926 42576 410932
rect 42246 400143 42302 400152
rect 42432 400172 42484 400178
rect 41972 400114 42024 400120
rect 42432 400114 42484 400120
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 42340 380928 42392 380934
rect 42340 380870 42392 380876
rect 41722 370075 42288 370103
rect 41713 369417 42193 369473
rect 41788 368688 41840 368694
rect 41788 368630 41840 368636
rect 41800 368263 41828 368630
rect 41722 368235 41828 368263
rect 41713 367577 42193 367633
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 42260 362250 42288 370075
rect 41892 362222 42288 362250
rect 41892 362114 41920 362222
rect 41722 362086 41920 362114
rect 41713 361413 42193 361469
rect 41713 360769 42193 360825
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41722 357734 41828 357762
rect 41800 357542 41828 357734
rect 42352 357542 42380 380870
rect 41788 357536 41840 357542
rect 41788 357478 41840 357484
rect 42340 357536 42392 357542
rect 42340 357478 42392 357484
rect 41722 357103 41828 357131
rect 41800 356726 41828 357103
rect 42444 356726 42472 400114
rect 42536 368694 42564 410926
rect 42628 401538 42656 413374
rect 42616 401532 42668 401538
rect 42616 401474 42668 401480
rect 42614 400208 42670 400217
rect 42614 400143 42670 400152
rect 42628 380934 42656 400143
rect 42616 380928 42668 380934
rect 42616 380870 42668 380876
rect 42524 368688 42576 368694
rect 42524 368630 42576 368636
rect 42536 367062 42564 368630
rect 42524 367056 42576 367062
rect 42524 366998 42576 367004
rect 42800 366988 42852 366994
rect 42800 366930 42852 366936
rect 42616 357536 42668 357542
rect 42616 357478 42668 357484
rect 41788 356720 41840 356726
rect 41788 356662 41840 356668
rect 42432 356720 42484 356726
rect 42432 356662 42484 356668
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 42340 334688 42392 334694
rect 42340 334630 42392 334636
rect 41722 326862 42288 326890
rect 41713 326217 42193 326273
rect 41722 325035 41828 325063
rect 41800 324562 41828 325035
rect 41788 324556 41840 324562
rect 41788 324498 41840 324504
rect 41713 324377 42193 324433
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 42260 318899 42288 326862
rect 41722 318871 42288 318899
rect 41713 318213 42193 318269
rect 41713 317569 42193 317625
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 42352 314634 42380 334630
rect 42340 314628 42392 314634
rect 41722 314547 41828 314575
rect 42340 314570 42392 314576
rect 41800 314498 41828 314547
rect 41788 314492 41840 314498
rect 41788 314434 41840 314440
rect 41722 313903 41828 313931
rect 41800 313818 41828 313903
rect 42444 313818 42472 356662
rect 42628 334694 42656 357478
rect 42812 347834 42840 366930
rect 42720 347806 42840 347834
rect 42720 347750 42748 347806
rect 42708 347744 42760 347750
rect 42708 347686 42760 347692
rect 42892 347744 42944 347750
rect 42892 347686 42944 347692
rect 42616 334688 42668 334694
rect 42616 334630 42668 334636
rect 42904 328506 42932 347686
rect 42616 328500 42668 328506
rect 42616 328442 42668 328448
rect 42892 328500 42944 328506
rect 42892 328442 42944 328448
rect 42524 324488 42576 324494
rect 42628 324442 42656 328442
rect 42576 324436 42656 324442
rect 42524 324430 42656 324436
rect 42536 324414 42656 324430
rect 42536 314498 42564 324414
rect 42616 314560 42668 314566
rect 42616 314502 42668 314508
rect 42524 314492 42576 314498
rect 42524 314434 42576 314440
rect 41788 313812 41840 313818
rect 41788 313754 41840 313760
rect 42432 313812 42484 313818
rect 42432 313754 42484 313760
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 42444 307970 42472 313754
rect 42432 307964 42484 307970
rect 42432 307906 42484 307912
rect 42628 295474 42656 314502
rect 42800 314492 42852 314498
rect 42800 314434 42852 314440
rect 42708 307964 42760 307970
rect 42708 307906 42760 307912
rect 42536 295446 42656 295474
rect 41722 283675 41920 283703
rect 41892 283234 41920 283675
rect 41892 283206 42288 283234
rect 41713 283017 42193 283073
rect 41788 282328 41840 282334
rect 41788 282270 41840 282276
rect 41800 281874 41828 282270
rect 41722 281846 41828 281874
rect 41713 281177 42193 281233
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41722 275671 41828 275699
rect 41800 275618 41828 275671
rect 42260 275618 42288 283206
rect 42432 282328 42484 282334
rect 42432 282270 42484 282276
rect 41800 275590 42288 275618
rect 41713 275013 42193 275069
rect 41713 274369 42193 274425
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41722 271374 41828 271402
rect 41800 270842 41828 271374
rect 41788 270836 41840 270842
rect 41788 270778 41840 270784
rect 41722 270694 41828 270722
rect 41800 270298 41828 270694
rect 41788 270292 41840 270298
rect 41788 270234 41840 270240
rect 42340 270292 42392 270298
rect 42340 270234 42392 270240
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 42352 247042 42380 270234
rect 42340 247036 42392 247042
rect 42340 246978 42392 246984
rect 41722 240502 42288 240530
rect 41713 239817 42193 239873
rect 41788 239080 41840 239086
rect 41788 239022 41840 239028
rect 41800 238663 41828 239022
rect 41722 238635 41828 238663
rect 41713 237977 42193 238033
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 42260 232642 42288 240502
rect 42444 239086 42472 282270
rect 42536 282146 42564 295446
rect 42616 295384 42668 295390
rect 42616 295326 42668 295332
rect 42628 282334 42656 295326
rect 42616 282328 42668 282334
rect 42616 282270 42668 282276
rect 42720 282266 42748 307906
rect 42812 295390 42840 314434
rect 42800 295384 42852 295390
rect 42800 295326 42852 295332
rect 42708 282260 42760 282266
rect 42708 282202 42760 282208
rect 42536 282118 42840 282146
rect 42708 282056 42760 282062
rect 42708 281998 42760 282004
rect 42524 276004 42576 276010
rect 42524 275946 42576 275952
rect 42536 270842 42564 275946
rect 42524 270836 42576 270842
rect 42524 270778 42576 270784
rect 42432 239080 42484 239086
rect 42432 239022 42484 239028
rect 41892 232614 42288 232642
rect 41892 232506 41920 232614
rect 41722 232478 41920 232506
rect 41713 231813 42193 231869
rect 41713 231169 42193 231225
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 42536 228682 42564 270778
rect 42720 270298 42748 281998
rect 42812 276010 42840 282118
rect 42800 276004 42852 276010
rect 42800 275946 42852 275952
rect 42708 270292 42760 270298
rect 42708 270234 42760 270240
rect 42708 247036 42760 247042
rect 42708 246978 42760 246984
rect 42616 239080 42668 239086
rect 42616 239022 42668 239028
rect 41788 228676 41840 228682
rect 41788 228618 41840 228624
rect 42524 228676 42576 228682
rect 42524 228618 42576 228624
rect 41800 228154 41828 228618
rect 41722 228126 41828 228154
rect 41788 228064 41840 228070
rect 41788 228006 41840 228012
rect 42432 228064 42484 228070
rect 42432 228006 42484 228012
rect 41800 227531 41828 228006
rect 42248 227928 42300 227934
rect 42248 227870 42300 227876
rect 41722 227503 41828 227531
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41722 197254 41828 197282
rect 41800 196790 41828 197254
rect 41788 196784 41840 196790
rect 41788 196726 41840 196732
rect 41713 196617 42193 196673
rect 41788 195900 41840 195906
rect 41788 195842 41840 195848
rect 41800 195463 41828 195842
rect 41722 195435 41828 195463
rect 41713 194777 42193 194833
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41788 189848 41840 189854
rect 41788 189790 41840 189796
rect 41800 189299 41828 189790
rect 41722 189271 41828 189299
rect 41713 188613 42193 188669
rect 41713 187969 42193 188025
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41722 184947 41828 184975
rect 41800 184498 41828 184947
rect 42260 184498 42288 227870
rect 42340 196784 42392 196790
rect 42340 196726 42392 196732
rect 42352 189854 42380 196726
rect 42340 189848 42392 189854
rect 42340 189790 42392 189796
rect 41800 184470 42380 184498
rect 41722 184303 41920 184331
rect 41892 184226 41920 184303
rect 42260 184278 42288 184309
rect 42248 184272 42300 184278
rect 41892 184220 42248 184226
rect 41892 184214 42300 184220
rect 41892 184198 42288 184214
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 39606 120278 39804 120306
rect 39776 120193 39804 120278
rect 39762 120184 39818 120193
rect 39762 120119 39818 120128
rect 41418 115968 41474 115977
rect 41418 115903 41474 115912
rect 39394 84280 39450 84289
rect 39394 84215 39450 84224
rect 39408 79098 39436 84215
rect 39316 79070 39528 79098
rect 39316 78948 39344 79070
rect 39500 78962 39528 79070
rect 39500 78934 39712 78962
rect 39684 75274 39712 78934
rect 39672 75268 39724 75274
rect 39672 75210 39724 75216
rect 39592 75126 39804 75154
rect 39592 75018 39620 75126
rect 39567 74990 39620 75018
rect 39672 74996 39724 75002
rect 39672 74938 39724 74944
rect 39330 68190 39620 68218
rect 39592 67998 39620 68190
rect 39580 67992 39632 67998
rect 39580 67934 39632 67940
rect 39684 52426 39712 74938
rect 39672 52420 39724 52426
rect 39672 52362 39724 52368
rect 39776 47734 39804 75126
rect 41432 67998 41460 115903
rect 41420 67992 41472 67998
rect 41420 67934 41472 67940
rect 41432 64666 41460 67934
rect 41420 64660 41472 64666
rect 41420 64602 41472 64608
rect 39856 52420 39908 52426
rect 39856 52362 39908 52368
rect 39868 47870 39896 52362
rect 39856 47864 39908 47870
rect 39856 47806 39908 47812
rect 39764 47728 39816 47734
rect 39764 47670 39816 47676
rect 42260 45694 42288 184198
rect 42352 115977 42380 184470
rect 42444 184278 42472 228006
rect 42536 227934 42564 228618
rect 42524 227928 42576 227934
rect 42524 227870 42576 227876
rect 42628 195906 42656 239022
rect 42720 228070 42748 246978
rect 42708 228064 42760 228070
rect 42708 228006 42760 228012
rect 42616 195900 42668 195906
rect 42616 195842 42668 195848
rect 42432 184272 42484 184278
rect 42432 184214 42484 184220
rect 44192 120193 44220 879786
rect 44284 458250 44312 922898
rect 44362 917280 44418 917289
rect 44362 917215 44418 917224
rect 44272 458244 44324 458250
rect 44272 458186 44324 458192
rect 44376 448633 44404 917215
rect 45940 879866 45968 996503
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 78876 992202 78904 995452
rect 78876 992174 79088 992202
rect 79060 990826 79088 992174
rect 79048 990820 79100 990826
rect 79048 990762 79100 990768
rect 79060 990146 79088 990762
rect 79520 990690 79548 995452
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 82569 995407 82625 995887
rect 83213 995407 83269 995887
rect 83885 995654 84056 995661
rect 83885 995648 84068 995654
rect 83885 995633 84016 995648
rect 84016 995590 84068 995596
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 89377 995407 89433 995887
rect 79508 990684 79560 990690
rect 79508 990626 79560 990632
rect 79968 990684 80020 990690
rect 79968 990626 80020 990632
rect 79980 990214 80008 990626
rect 90008 990622 90036 995452
rect 91217 995407 91273 995887
rect 91744 995648 91796 995654
rect 91744 995590 91796 995596
rect 91756 995466 91784 995590
rect 91756 995438 91862 995466
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 130304 990894 130332 995452
rect 130292 990888 130344 990894
rect 130292 990830 130344 990836
rect 110420 990820 110472 990826
rect 110420 990762 110472 990768
rect 130108 990820 130160 990826
rect 130108 990762 130160 990768
rect 110432 990706 110460 990762
rect 110432 990678 110552 990706
rect 110524 990622 110552 990678
rect 130120 990622 130148 990762
rect 130948 990690 130976 995452
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 133969 995407 134025 995887
rect 134613 995407 134669 995887
rect 135352 995512 135404 995518
rect 135286 995460 135352 995466
rect 135286 995454 135404 995460
rect 135286 995438 135392 995454
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140777 995407 140833 995887
rect 141436 992118 141464 995452
rect 142617 995407 142673 995887
rect 143172 995512 143224 995518
rect 143224 995460 143290 995466
rect 143172 995454 143290 995460
rect 143184 995438 143290 995454
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 181717 995438 181760 995466
rect 182361 995438 182404 995466
rect 141424 992112 141476 992118
rect 141424 992054 141476 992060
rect 154396 992112 154448 992118
rect 154396 992054 154448 992060
rect 141436 990978 141464 992054
rect 141344 990950 141464 990978
rect 130936 990684 130988 990690
rect 130936 990626 130988 990632
rect 89996 990616 90048 990622
rect 89996 990558 90048 990564
rect 110512 990616 110564 990622
rect 110512 990558 110564 990564
rect 130108 990616 130160 990622
rect 130108 990558 130160 990564
rect 79968 990208 80020 990214
rect 79968 990150 80020 990156
rect 90008 990146 90036 990558
rect 141344 990486 141372 990950
rect 143264 990820 143316 990826
rect 143264 990762 143316 990768
rect 143276 990486 143304 990762
rect 141332 990480 141384 990486
rect 141332 990422 141384 990428
rect 143264 990480 143316 990486
rect 143264 990422 143316 990428
rect 154408 990418 154436 992054
rect 173808 990820 173860 990826
rect 173808 990762 173860 990768
rect 179328 990820 179380 990826
rect 179328 990762 179380 990768
rect 173820 990729 173848 990762
rect 160098 990720 160154 990729
rect 160098 990655 160154 990664
rect 173806 990720 173862 990729
rect 173806 990655 173862 990664
rect 160112 990486 160140 990655
rect 179340 990622 179368 990762
rect 181732 990622 181760 995438
rect 182376 990690 182404 995438
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 185369 995407 185425 995887
rect 186013 995407 186069 995887
rect 186685 995438 186728 995466
rect 182364 990684 182416 990690
rect 182364 990626 182416 990632
rect 186700 990622 186728 995438
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 192177 995407 192233 995887
rect 192849 995438 192892 995466
rect 187608 990752 187660 990758
rect 187608 990694 187660 990700
rect 187700 990752 187752 990758
rect 187700 990694 187752 990700
rect 179328 990616 179380 990622
rect 179328 990558 179380 990564
rect 181720 990616 181772 990622
rect 181720 990558 181772 990564
rect 186688 990616 186740 990622
rect 186688 990558 186740 990564
rect 164148 990548 164200 990554
rect 164148 990490 164200 990496
rect 160100 990480 160152 990486
rect 160100 990422 160152 990428
rect 154396 990412 154448 990418
rect 154396 990354 154448 990360
rect 154580 990412 154632 990418
rect 154580 990354 154632 990360
rect 154592 990282 154620 990354
rect 164160 990282 164188 990490
rect 181732 990486 181760 990558
rect 187620 990486 187648 990694
rect 187712 990486 187740 990694
rect 192864 990554 192892 995438
rect 194017 995407 194073 995887
rect 194689 995438 194732 995466
rect 194704 990622 194732 995438
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 233068 995438 233117 995466
rect 233712 995438 233761 995466
rect 231860 995104 231912 995110
rect 231860 995046 231912 995052
rect 202880 990752 202932 990758
rect 202880 990694 202932 990700
rect 194692 990616 194744 990622
rect 193218 990584 193274 990593
rect 192852 990548 192904 990554
rect 194692 990558 194744 990564
rect 193218 990519 193220 990528
rect 192852 990490 192904 990496
rect 193272 990519 193274 990528
rect 193220 990490 193272 990496
rect 202892 990486 202920 990694
rect 212446 990584 212502 990593
rect 231872 990554 231900 995046
rect 233068 990758 233096 995438
rect 233056 990752 233108 990758
rect 233056 990694 233108 990700
rect 212446 990519 212448 990528
rect 212500 990519 212502 990528
rect 231860 990548 231912 990554
rect 212448 990490 212500 990496
rect 231860 990490 231912 990496
rect 233068 990486 233096 990694
rect 233712 990690 233740 995438
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 236769 995407 236825 995887
rect 237413 995407 237469 995887
rect 238208 995648 238260 995654
rect 238208 995590 238260 995596
rect 238220 995466 238248 995590
rect 238085 995438 238248 995466
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 243577 995407 243633 995887
rect 244200 995438 244249 995466
rect 244200 995110 244228 995438
rect 245417 995407 245473 995887
rect 245936 995648 245988 995654
rect 245936 995590 245988 995596
rect 245948 995466 245976 995590
rect 245948 995438 246089 995466
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 244188 995104 244240 995110
rect 244188 995046 244240 995052
rect 244200 990758 244228 995046
rect 284680 990826 284708 995452
rect 246948 990820 247000 990826
rect 246948 990762 247000 990768
rect 284668 990820 284720 990826
rect 284668 990762 284720 990768
rect 244188 990752 244240 990758
rect 244188 990694 244240 990700
rect 233700 990684 233752 990690
rect 233700 990626 233752 990632
rect 246960 990486 246988 990762
rect 285324 990690 285352 995452
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 288369 995407 288425 995887
rect 289013 995407 289069 995887
rect 289648 995314 289676 995452
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 295177 995407 295233 995887
rect 289636 995308 289688 995314
rect 289636 995250 289688 995256
rect 286968 990820 287020 990826
rect 286968 990762 287020 990768
rect 285312 990684 285364 990690
rect 285312 990626 285364 990632
rect 286980 990554 287008 990762
rect 295812 990758 295840 995452
rect 297017 995407 297073 995887
rect 297652 995314 297680 995452
rect 297640 995308 297692 995314
rect 297640 995250 297692 995256
rect 295800 990752 295852 990758
rect 295800 990694 295852 990700
rect 333532 990690 333560 997591
rect 585704 996441 585732 997628
rect 672630 996568 672686 996577
rect 672630 996503 672686 996512
rect 585690 996432 585746 996441
rect 585690 996367 585746 996376
rect 672446 996432 672502 996441
rect 672446 996367 672502 996376
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 386328 990752 386380 990758
rect 386328 990694 386380 990700
rect 333520 990684 333572 990690
rect 333520 990626 333572 990632
rect 286968 990548 287020 990554
rect 286968 990490 287020 990496
rect 181720 990480 181772 990486
rect 181720 990422 181772 990428
rect 187608 990480 187660 990486
rect 187608 990422 187660 990428
rect 187700 990480 187752 990486
rect 187700 990422 187752 990428
rect 202880 990480 202932 990486
rect 202880 990422 202932 990428
rect 233056 990480 233108 990486
rect 233056 990422 233108 990428
rect 246948 990480 247000 990486
rect 246948 990422 247000 990428
rect 386340 990418 386368 990694
rect 386524 990622 386552 995452
rect 387168 990690 387196 995452
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 390169 995407 390225 995887
rect 390813 995407 390869 995887
rect 391492 995314 391520 995452
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396977 995407 397033 995887
rect 391480 995308 391532 995314
rect 391480 995250 391532 995256
rect 391756 990820 391808 990826
rect 391756 990762 391808 990768
rect 391768 990690 391796 990762
rect 387156 990684 387208 990690
rect 387156 990626 387208 990632
rect 391756 990684 391808 990690
rect 391756 990626 391808 990632
rect 386512 990616 386564 990622
rect 386512 990558 386564 990564
rect 397656 990418 397684 995452
rect 398817 995407 398873 995887
rect 399496 995314 399524 995452
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 399484 995308 399536 995314
rect 399484 995250 399536 995256
rect 475488 992322 475516 995452
rect 463792 992316 463844 992322
rect 463792 992258 463844 992264
rect 475476 992316 475528 992322
rect 475476 992258 475528 992264
rect 419540 990888 419592 990894
rect 419540 990830 419592 990836
rect 438676 990888 438728 990894
rect 438676 990830 438728 990836
rect 450268 990888 450320 990894
rect 450268 990830 450320 990836
rect 463608 990888 463660 990894
rect 463804 990842 463832 992258
rect 463660 990836 463832 990842
rect 463608 990830 463832 990836
rect 419552 990622 419580 990830
rect 419540 990616 419592 990622
rect 419540 990558 419592 990564
rect 438688 990570 438716 990830
rect 450280 990622 450308 990830
rect 463620 990814 463832 990830
rect 476132 990826 476160 995452
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 479169 995407 479225 995887
rect 479813 995407 479869 995887
rect 480456 995314 480484 995452
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485977 995407 486033 995887
rect 480444 995308 480496 995314
rect 480444 995250 480496 995256
rect 482928 992316 482980 992322
rect 482928 992258 482980 992264
rect 476120 990820 476172 990826
rect 476120 990762 476172 990768
rect 482940 990758 482968 992258
rect 482928 990752 482980 990758
rect 482928 990694 482980 990700
rect 438768 990616 438820 990622
rect 438688 990564 438768 990570
rect 438688 990558 438820 990564
rect 450268 990616 450320 990622
rect 469312 990616 469364 990622
rect 450268 990558 450320 990564
rect 469048 990564 469312 990570
rect 469048 990558 469364 990564
rect 438688 990542 438808 990558
rect 469048 990554 469352 990558
rect 469036 990548 469352 990554
rect 469088 990542 469352 990548
rect 483020 990548 483072 990554
rect 469036 990490 469088 990496
rect 483020 990490 483072 990496
rect 483032 990418 483060 990490
rect 486620 990418 486648 995452
rect 487817 995407 487873 995887
rect 488460 995314 488488 995452
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 488448 995308 488500 995314
rect 488448 995250 488500 995256
rect 526916 990758 526944 995452
rect 527560 990826 527588 995452
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 530569 995407 530625 995887
rect 531213 995407 531269 995887
rect 531964 995648 532016 995654
rect 531964 995590 532016 995596
rect 531976 995466 532004 995590
rect 531898 995438 532004 995466
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 537377 995407 537433 995887
rect 537850 995480 537906 995489
rect 537850 995415 537906 995424
rect 538034 995480 538090 995489
rect 538034 995415 538090 995424
rect 527548 990820 527600 990826
rect 527548 990762 527600 990768
rect 526904 990752 526956 990758
rect 526904 990694 526956 990700
rect 386328 990412 386380 990418
rect 386328 990354 386380 990360
rect 397644 990412 397696 990418
rect 397644 990354 397696 990360
rect 424968 990412 425020 990418
rect 424968 990354 425020 990360
rect 483020 990412 483072 990418
rect 483020 990354 483072 990360
rect 486608 990412 486660 990418
rect 486608 990354 486660 990360
rect 521660 990412 521712 990418
rect 521660 990354 521712 990360
rect 397656 990282 397684 990354
rect 154580 990276 154632 990282
rect 154580 990218 154632 990224
rect 164148 990276 164200 990282
rect 164148 990218 164200 990224
rect 397644 990276 397696 990282
rect 397644 990218 397696 990224
rect 405740 990276 405792 990282
rect 405740 990218 405792 990224
rect 405752 990146 405780 990218
rect 424980 990146 425008 990354
rect 507768 990344 507820 990350
rect 507860 990344 507912 990350
rect 507820 990292 507860 990298
rect 507768 990286 507912 990292
rect 507780 990270 507900 990286
rect 521672 990282 521700 990354
rect 537864 990282 537892 995415
rect 539217 995407 539273 995887
rect 539692 995648 539744 995654
rect 539692 995590 539744 995596
rect 539704 995466 539732 995590
rect 539704 995438 539902 995466
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 628668 995438 628717 995466
rect 629312 995438 629361 995466
rect 628668 990758 628696 995438
rect 629312 990826 629340 995438
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 632369 995407 632425 995887
rect 633013 995407 633069 995887
rect 633808 995512 633860 995518
rect 633685 995460 633808 995466
rect 633685 995454 633860 995460
rect 633685 995438 633848 995454
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 639177 995407 639233 995887
rect 639800 995438 639849 995466
rect 629300 990820 629352 990826
rect 629300 990762 629352 990768
rect 628656 990752 628708 990758
rect 628656 990694 628708 990700
rect 596088 990684 596140 990690
rect 596088 990626 596140 990632
rect 576860 990616 576912 990622
rect 576858 990584 576860 990593
rect 596100 990593 596128 990626
rect 623688 990616 623740 990622
rect 576912 990584 576914 990593
rect 560208 990548 560260 990554
rect 576858 990519 576914 990528
rect 596086 990584 596142 990593
rect 623740 990564 623912 990570
rect 623688 990558 623912 990564
rect 623700 990554 623912 990558
rect 623700 990548 623924 990554
rect 623700 990542 623872 990548
rect 596086 990519 596142 990528
rect 560208 990490 560260 990496
rect 623872 990490 623924 990496
rect 540980 990480 541032 990486
rect 540978 990448 540980 990457
rect 560220 990457 560248 990490
rect 541032 990448 541034 990457
rect 540888 990412 540940 990418
rect 540978 990383 541034 990392
rect 560206 990448 560262 990457
rect 560206 990383 560262 990392
rect 540888 990354 540940 990360
rect 540900 990282 540928 990354
rect 521660 990276 521712 990282
rect 521660 990218 521712 990224
rect 537852 990276 537904 990282
rect 537852 990218 537904 990224
rect 540888 990276 540940 990282
rect 540888 990218 540940 990224
rect 628668 990146 628696 990694
rect 629312 990146 629340 990762
rect 639800 990554 639828 995438
rect 641017 995407 641073 995887
rect 641536 995512 641588 995518
rect 641588 995460 641689 995466
rect 641536 995454 641689 995460
rect 641548 995438 641689 995454
rect 639788 990548 639840 990554
rect 639788 990490 639840 990496
rect 639800 990214 639828 990490
rect 639788 990208 639840 990214
rect 639788 990150 639840 990156
rect 79048 990140 79100 990146
rect 79048 990082 79100 990088
rect 89996 990140 90048 990146
rect 89996 990082 90048 990088
rect 405740 990140 405792 990146
rect 405740 990082 405792 990088
rect 424968 990140 425020 990146
rect 424968 990082 425020 990088
rect 628656 990140 628708 990146
rect 628656 990082 628708 990088
rect 629300 990140 629352 990146
rect 629300 990082 629352 990088
rect 45848 879850 45968 879866
rect 45836 879844 45968 879850
rect 45888 879838 45968 879844
rect 45836 879786 45888 879792
rect 44454 835272 44510 835281
rect 44454 835207 44510 835216
rect 44468 493241 44496 835207
rect 672460 828730 672488 996367
rect 672538 828744 672594 828753
rect 672460 828702 672538 828730
rect 672538 828679 672594 828688
rect 44730 828064 44786 828073
rect 44730 827999 44786 828008
rect 44744 806002 44772 827999
rect 672644 826169 672672 996503
rect 673644 990208 673696 990214
rect 673644 990150 673696 990156
rect 673552 990140 673604 990146
rect 673552 990082 673604 990088
rect 673460 990072 673512 990078
rect 673460 990014 673512 990020
rect 673472 965326 673500 990014
rect 673460 965320 673512 965326
rect 673460 965262 673512 965268
rect 673366 908168 673422 908177
rect 673366 908103 673422 908112
rect 673184 908064 673236 908070
rect 673184 908006 673236 908012
rect 673196 888826 673224 908006
rect 673184 888820 673236 888826
rect 673184 888762 673236 888768
rect 672630 826160 672686 826169
rect 672630 826095 672686 826104
rect 673274 826160 673330 826169
rect 673274 826095 673330 826104
rect 673182 823712 673238 823721
rect 673182 823647 673238 823656
rect 44548 805996 44600 806002
rect 44548 805938 44600 805944
rect 44732 805996 44784 806002
rect 44732 805938 44784 805944
rect 44560 786570 44588 805938
rect 673196 792169 673224 823647
rect 672998 792160 673054 792169
rect 672998 792095 673054 792104
rect 673182 792160 673238 792169
rect 673182 792095 673238 792104
rect 44560 786542 44772 786570
rect 44744 778274 44772 786542
rect 673012 778394 673040 792095
rect 673000 778388 673052 778394
rect 673000 778330 673052 778336
rect 44652 778246 44772 778274
rect 673092 778252 673144 778258
rect 44652 759098 44680 778246
rect 673092 778194 673144 778200
rect 673104 772818 673132 778194
rect 672816 772812 672868 772818
rect 672816 772754 672868 772760
rect 673092 772812 673144 772818
rect 673092 772754 673144 772760
rect 44560 759070 44680 759098
rect 44560 701026 44588 759070
rect 672828 753545 672856 772754
rect 672814 753536 672870 753545
rect 672814 753471 672870 753480
rect 672998 753536 673054 753545
rect 672998 753471 673054 753480
rect 673012 739770 673040 753471
rect 673000 739764 673052 739770
rect 673000 739706 673052 739712
rect 673184 739628 673236 739634
rect 673184 739570 673236 739576
rect 673196 714762 673224 739570
rect 673104 714734 673224 714762
rect 44560 700998 44680 701026
rect 44652 695502 44680 700998
rect 673104 695570 673132 714734
rect 673092 695564 673144 695570
rect 673092 695506 673144 695512
rect 673184 695564 673236 695570
rect 673184 695506 673236 695512
rect 44640 695496 44692 695502
rect 44640 695438 44692 695444
rect 44916 695496 44968 695502
rect 44916 695438 44968 695444
rect 44928 676258 44956 695438
rect 44732 676252 44784 676258
rect 44732 676194 44784 676200
rect 44916 676252 44968 676258
rect 44916 676194 44968 676200
rect 44560 662454 44588 662485
rect 44744 662454 44772 676194
rect 673196 662522 673224 695506
rect 673184 662516 673236 662522
rect 673184 662458 673236 662464
rect 44548 662448 44600 662454
rect 44732 662448 44784 662454
rect 44600 662396 44680 662402
rect 44548 662390 44680 662396
rect 44732 662390 44784 662396
rect 44560 662374 44680 662390
rect 44652 656878 44680 662374
rect 673184 662380 673236 662386
rect 673184 662322 673236 662328
rect 44640 656872 44692 656878
rect 44640 656814 44692 656820
rect 44824 656872 44876 656878
rect 44824 656814 44876 656820
rect 44836 642818 44864 656814
rect 673196 643090 673224 662322
rect 44652 642790 44864 642818
rect 673104 643062 673224 643090
rect 44652 604586 44680 642790
rect 673104 637566 673132 643062
rect 672816 637560 672868 637566
rect 672816 637502 672868 637508
rect 673092 637560 673144 637566
rect 673092 637502 673144 637508
rect 672828 618322 672856 637502
rect 672816 618316 672868 618322
rect 672816 618258 672868 618264
rect 673000 618316 673052 618322
rect 673000 618258 673052 618264
rect 673012 618225 673040 618258
rect 672998 618216 673054 618225
rect 672998 618151 673054 618160
rect 672814 618080 672870 618089
rect 672814 618015 672870 618024
rect 44640 604580 44692 604586
rect 44640 604522 44692 604528
rect 44640 604444 44692 604450
rect 44640 604386 44692 604392
rect 44652 585154 44680 604386
rect 672828 599010 672856 618015
rect 672816 599004 672868 599010
rect 672816 598946 672868 598952
rect 673092 599004 673144 599010
rect 673092 598946 673144 598952
rect 673104 585206 673132 598946
rect 44560 585126 44680 585154
rect 673092 585200 673144 585206
rect 673092 585142 673144 585148
rect 673000 585132 673052 585138
rect 44560 560289 44588 585126
rect 673000 585074 673052 585080
rect 673012 569974 673040 585074
rect 672816 569968 672868 569974
rect 672816 569910 672868 569916
rect 673000 569968 673052 569974
rect 673000 569910 673052 569916
rect 672828 560318 672856 569910
rect 672816 560312 672868 560318
rect 44546 560280 44602 560289
rect 44546 560215 44602 560224
rect 44914 560280 44970 560289
rect 672816 560254 672868 560260
rect 673000 560312 673052 560318
rect 673000 560254 673052 560260
rect 44914 560215 44970 560224
rect 44928 541006 44956 560215
rect 673012 546582 673040 560254
rect 673000 546576 673052 546582
rect 673000 546518 673052 546524
rect 673092 546372 673144 546378
rect 673092 546314 673144 546320
rect 44732 541000 44784 541006
rect 44732 540942 44784 540948
rect 44916 541000 44968 541006
rect 44916 540942 44968 540948
rect 44744 496874 44772 540942
rect 673104 527202 673132 546314
rect 673092 527196 673144 527202
rect 673092 527138 673144 527144
rect 673184 527060 673236 527066
rect 673184 527002 673236 527008
rect 673196 521626 673224 527002
rect 673184 521620 673236 521626
rect 673184 521562 673236 521568
rect 673288 511465 673316 826095
rect 673090 511456 673146 511465
rect 673090 511391 673146 511400
rect 673274 511456 673330 511465
rect 673274 511391 673330 511400
rect 672998 509144 673054 509153
rect 672998 509079 673054 509088
rect 44548 496868 44600 496874
rect 44548 496810 44600 496816
rect 44732 496868 44784 496874
rect 44732 496810 44784 496816
rect 44454 493232 44510 493241
rect 44454 493167 44510 493176
rect 44560 488617 44588 496810
rect 44546 488608 44602 488617
rect 44546 488543 44602 488552
rect 673012 449954 673040 509079
rect 673000 449948 673052 449954
rect 673000 449890 673052 449896
rect 44362 448624 44418 448633
rect 44362 448559 44418 448568
rect 673104 427961 673132 511391
rect 673274 502344 673330 502353
rect 673274 502279 673330 502288
rect 673288 463729 673316 502279
rect 673380 483177 673408 908103
rect 673472 908070 673500 965262
rect 673564 964782 673592 990082
rect 673552 964776 673604 964782
rect 673552 964718 673604 964724
rect 673564 910790 673592 964718
rect 673656 953358 673684 990150
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 675407 965407 675887 965463
rect 675392 965320 675444 965326
rect 675392 965262 675444 965268
rect 675404 964883 675432 965262
rect 675392 964776 675444 964782
rect 675392 964718 675444 964724
rect 675404 964239 675432 964718
rect 675407 963567 675887 963623
rect 675407 963015 675887 963071
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 675407 961175 675887 961231
rect 675407 960531 675887 960587
rect 675312 959901 675418 959929
rect 673644 953352 673696 953358
rect 673644 953294 673696 953300
rect 673552 910784 673604 910790
rect 673552 910726 673604 910732
rect 673460 908064 673512 908070
rect 673460 908006 673512 908012
rect 673460 888820 673512 888826
rect 673460 888762 673512 888768
rect 673472 888729 673500 888762
rect 673458 888720 673514 888729
rect 673458 888655 673514 888664
rect 673564 875566 673592 910726
rect 673552 875560 673604 875566
rect 673552 875502 673604 875508
rect 673656 875090 673684 953294
rect 675312 951810 675340 959901
rect 675407 959243 675887 959299
rect 675407 958691 675887 958747
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 675407 956207 675887 956263
rect 675407 954367 675887 954423
rect 675404 953358 675432 953751
rect 675392 953352 675444 953358
rect 675392 953294 675444 953300
rect 675407 952527 675887 952583
rect 675404 951810 675432 951932
rect 675312 951782 675432 951810
rect 677874 918640 677930 918649
rect 677930 918598 678086 918626
rect 677874 918575 677930 918584
rect 677598 915376 677654 915385
rect 677598 915311 677654 915320
rect 677612 912801 677640 915311
rect 677796 913974 678046 914002
rect 677598 912792 677654 912801
rect 677598 912727 677654 912736
rect 677796 910790 677824 913974
rect 678018 913716 678046 913974
rect 677874 912792 677930 912801
rect 677874 912727 677930 912736
rect 677784 910784 677836 910790
rect 677784 910726 677836 910732
rect 677888 908177 677916 912727
rect 677874 908168 677930 908177
rect 677874 908103 677930 908112
rect 677782 907760 677838 907769
rect 677838 907718 678086 907746
rect 677782 907695 677838 907704
rect 675298 888720 675354 888729
rect 675298 888655 675354 888664
rect 675312 875697 675340 888655
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675220 875669 675418 875697
rect 673644 875084 673696 875090
rect 673644 875026 673696 875032
rect 673644 874948 673696 874954
rect 673644 874890 673696 874896
rect 673656 865026 673684 874890
rect 675220 869446 675248 875669
rect 675392 875560 675444 875566
rect 675392 875502 675444 875508
rect 675404 875039 675432 875502
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675887 872031
rect 675407 871331 675887 871387
rect 675404 870210 675432 870740
rect 675312 870182 675432 870210
rect 673736 869440 673788 869446
rect 673736 869382 673788 869388
rect 675208 869440 675260 869446
rect 675208 869382 675260 869388
rect 673644 865020 673696 865026
rect 673644 864962 673696 864968
rect 673748 855522 673776 869382
rect 673828 865020 673880 865026
rect 673828 864962 673880 864968
rect 673656 855494 673776 855522
rect 673656 850082 673684 855494
rect 673564 850054 673684 850082
rect 673564 836330 673592 850054
rect 673552 836324 673604 836330
rect 673552 836266 673604 836272
rect 673644 836256 673696 836262
rect 673644 836198 673696 836204
rect 673656 830822 673684 836198
rect 673552 830816 673604 830822
rect 673552 830758 673604 830764
rect 673644 830816 673696 830822
rect 673644 830758 673696 830764
rect 673564 821098 673592 830758
rect 673552 821092 673604 821098
rect 673552 821034 673604 821040
rect 673644 785324 673696 785330
rect 673644 785266 673696 785272
rect 673460 774920 673512 774926
rect 673460 774862 673512 774868
rect 673472 730182 673500 774862
rect 673552 768664 673604 768670
rect 673552 768606 673604 768612
rect 673564 741946 673592 768606
rect 673552 741940 673604 741946
rect 673552 741882 673604 741888
rect 673656 741402 673684 785266
rect 673840 774926 673868 864962
rect 675312 862730 675340 870182
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865167 675887 865223
rect 675392 865020 675444 865026
rect 675392 864962 675444 864968
rect 675404 864551 675432 864962
rect 675407 863327 675887 863383
rect 675312 862702 675418 862730
rect 676126 828744 676182 828753
rect 676126 828679 676182 828688
rect 676140 823721 676168 828679
rect 676126 823712 676182 823721
rect 676126 823647 676182 823656
rect 674104 821092 674156 821098
rect 674104 821034 674156 821040
rect 674116 797638 674144 821034
rect 674104 797632 674156 797638
rect 674104 797574 674156 797580
rect 675300 797632 675352 797638
rect 675300 797574 675352 797580
rect 675312 786497 675340 797574
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675312 786486 675418 786497
rect 674012 786480 674064 786486
rect 674012 786422 674064 786428
rect 675300 786480 675418 786486
rect 675352 786469 675418 786480
rect 675300 786422 675352 786428
rect 673828 774920 673880 774926
rect 673828 774862 673880 774868
rect 674024 768670 674052 786422
rect 675312 786386 675340 786422
rect 675404 785330 675432 785839
rect 675392 785324 675444 785330
rect 675392 785266 675444 785272
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675887 782831
rect 675407 782131 675887 782187
rect 675312 781510 675418 781538
rect 675312 773514 675340 781510
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 775967 675887 776023
rect 675404 774926 675432 775351
rect 675392 774920 675444 774926
rect 675392 774862 675444 774868
rect 675407 774127 675887 774183
rect 675312 773486 675418 773514
rect 674012 768664 674064 768670
rect 674012 768606 674064 768612
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 674196 741940 674248 741946
rect 674196 741882 674248 741888
rect 675392 741940 675444 741946
rect 675392 741882 675444 741888
rect 673644 741396 673696 741402
rect 673644 741338 673696 741344
rect 673460 730176 673512 730182
rect 673460 730118 673512 730124
rect 673472 685409 673500 730118
rect 673828 730040 673880 730046
rect 673828 729982 673880 729988
rect 673644 695972 673696 695978
rect 673644 695914 673696 695920
rect 673552 695360 673604 695366
rect 673552 695302 673604 695308
rect 673458 685400 673514 685409
rect 673458 685335 673514 685344
rect 673472 639742 673500 685335
rect 673564 651166 673592 695302
rect 673656 651778 673684 695914
rect 673840 695366 673868 729982
rect 674208 720458 674236 741882
rect 675404 741483 675432 741882
rect 675392 741396 675444 741402
rect 675392 741338 675444 741344
rect 675404 740874 675432 741338
rect 675128 740860 675432 740874
rect 675128 740846 675418 740860
rect 675128 730046 675156 740846
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675887 737831
rect 675407 737131 675887 737187
rect 675312 736494 675418 736522
rect 675116 730040 675168 730046
rect 675116 729982 675168 729988
rect 675312 729042 675340 736494
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 730967 675887 731023
rect 675404 730182 675432 730351
rect 675392 730176 675444 730182
rect 675392 730118 675444 730124
rect 675407 729127 675887 729183
rect 675312 729014 675432 729042
rect 675404 728484 675432 729014
rect 674012 720452 674064 720458
rect 674012 720394 674064 720400
rect 674196 720452 674248 720458
rect 674196 720394 674248 720400
rect 674024 710734 674052 720394
rect 674012 710728 674064 710734
rect 674012 710670 674064 710676
rect 675300 710728 675352 710734
rect 675300 710670 675352 710676
rect 675312 696497 675340 710670
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675312 696483 675418 696497
rect 675312 696469 675432 696483
rect 675404 695978 675432 696469
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675404 695366 675432 695844
rect 673828 695360 673880 695366
rect 673828 695302 673880 695308
rect 675392 695360 675444 695366
rect 675392 695302 675444 695308
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675887 692831
rect 675407 692131 675887 692187
rect 675312 691614 675432 691642
rect 675312 683525 675340 691614
rect 675404 691492 675432 691614
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 685967 675887 686023
rect 675390 685400 675446 685409
rect 675390 685335 675446 685344
rect 675407 684127 675887 684183
rect 675312 683497 675418 683525
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 673644 651772 673696 651778
rect 673644 651714 673696 651720
rect 675392 651772 675444 651778
rect 675392 651714 675444 651720
rect 673552 651160 673604 651166
rect 673552 651102 673604 651108
rect 673460 639736 673512 639742
rect 673460 639678 673512 639684
rect 673472 594930 673500 639678
rect 673564 605674 673592 651102
rect 673656 606762 673684 651714
rect 675404 651283 675432 651714
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675404 650639 675432 651102
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675887 647631
rect 675407 646931 675887 646987
rect 675404 645810 675432 646340
rect 675312 645782 675432 645810
rect 675312 638330 675340 645782
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 640767 675887 640823
rect 675404 639742 675432 640151
rect 675392 639736 675444 639742
rect 675392 639678 675444 639684
rect 675407 638927 675887 638983
rect 675312 638302 675418 638330
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 673644 606756 673696 606762
rect 673644 606698 673696 606704
rect 675392 606756 675444 606762
rect 675392 606698 675444 606704
rect 673552 605668 673604 605674
rect 673552 605610 673604 605616
rect 673564 604450 673592 605610
rect 673552 604444 673604 604450
rect 673552 604386 673604 604392
rect 673460 594924 673512 594930
rect 673460 594866 673512 594872
rect 673472 550526 673500 594866
rect 673552 565888 673604 565894
rect 673552 565830 673604 565836
rect 673564 559978 673592 565830
rect 673656 561542 673684 606698
rect 675404 606283 675432 606698
rect 675300 605668 675352 605674
rect 675352 605625 675418 605653
rect 675300 605610 675352 605616
rect 675407 604967 675887 605023
rect 673828 604444 673880 604450
rect 675407 604415 675887 604471
rect 673828 604386 673880 604392
rect 673840 585154 673868 604386
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675887 602631
rect 675407 601931 675887 601987
rect 675312 601310 675418 601338
rect 675312 593314 675340 601310
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 595767 675887 595823
rect 675404 594930 675432 595151
rect 675392 594924 675444 594930
rect 675392 594866 675444 594872
rect 675407 593927 675887 593983
rect 675312 593286 675418 593314
rect 673840 585126 673960 585154
rect 673932 565894 673960 585126
rect 673920 565888 673972 565894
rect 673920 565830 673972 565836
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 673644 561536 673696 561542
rect 673644 561478 673696 561484
rect 675392 561536 675444 561542
rect 675392 561478 675444 561484
rect 675404 561068 675432 561478
rect 675404 559978 675432 560439
rect 673552 559972 673604 559978
rect 673552 559914 673604 559920
rect 673920 559972 673972 559978
rect 673920 559914 673972 559920
rect 675392 559972 675444 559978
rect 675392 559914 675444 559920
rect 673460 550520 673512 550526
rect 673460 550462 673512 550468
rect 673932 522986 673960 559914
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675887 557431
rect 675407 556731 675887 556787
rect 675312 556101 675418 556129
rect 675312 548125 675340 556101
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 550567 675887 550623
rect 675392 550520 675444 550526
rect 675392 550462 675444 550468
rect 675404 549951 675432 550462
rect 675407 548727 675887 548783
rect 675312 548097 675418 548125
rect 673736 522980 673788 522986
rect 673736 522922 673788 522928
rect 673920 522980 673972 522986
rect 673920 522922 673972 522928
rect 673748 511850 673776 522922
rect 676128 521620 676180 521626
rect 676128 521562 676180 521568
rect 676140 514185 676168 521562
rect 676126 514176 676182 514185
rect 676126 514111 676182 514120
rect 673656 511822 673776 511850
rect 673656 502353 673684 511822
rect 676140 509153 676168 514111
rect 676126 509144 676182 509153
rect 676126 509079 676182 509088
rect 673642 502344 673698 502353
rect 673642 502279 673698 502288
rect 673366 483168 673422 483177
rect 673366 483103 673422 483112
rect 673366 483032 673422 483041
rect 673366 482967 673422 482976
rect 673380 467537 673408 482967
rect 678058 477592 678114 477601
rect 678058 477527 678114 477536
rect 678072 470778 678100 477527
rect 677888 470764 678100 470778
rect 677888 470750 678086 470764
rect 677888 469985 677916 470750
rect 677874 469976 677930 469985
rect 677874 469911 677930 469920
rect 673366 467528 673422 467537
rect 673366 467463 673422 467472
rect 677704 465990 678032 466018
rect 673274 463720 673330 463729
rect 673274 463655 673330 463664
rect 673458 463720 673514 463729
rect 677704 463690 677732 465990
rect 673458 463655 673514 463664
rect 673736 463684 673788 463690
rect 673472 463593 673500 463655
rect 673736 463626 673788 463632
rect 677692 463684 677744 463690
rect 677692 463626 677744 463632
rect 673748 463593 673776 463626
rect 673458 463584 673514 463593
rect 673458 463519 673514 463528
rect 673734 463584 673790 463593
rect 673734 463519 673790 463528
rect 673368 449948 673420 449954
rect 673368 449890 673420 449896
rect 673090 427952 673146 427961
rect 673090 427887 673146 427896
rect 673380 420889 673408 449890
rect 673748 444417 673776 463519
rect 677704 459870 678086 459898
rect 673550 444408 673606 444417
rect 673550 444343 673606 444352
rect 673734 444408 673790 444417
rect 673734 444343 673790 444352
rect 673564 430658 673592 444343
rect 677704 440230 677732 459870
rect 676220 440224 676272 440230
rect 676220 440166 676272 440172
rect 677692 440224 677744 440230
rect 677692 440166 677744 440172
rect 673564 430630 673684 430658
rect 673656 430522 673684 430630
rect 673564 430494 673684 430522
rect 673366 420880 673422 420889
rect 673366 420815 673422 420824
rect 672816 412548 672868 412554
rect 672816 412490 672868 412496
rect 672828 411210 672856 412490
rect 673564 411346 673592 430494
rect 676232 412554 676260 440166
rect 677414 427952 677470 427961
rect 677414 427887 677470 427896
rect 677428 425762 677456 427887
rect 677598 425776 677654 425785
rect 677428 425734 677598 425762
rect 677598 425711 677654 425720
rect 676220 412548 676272 412554
rect 676220 412490 676272 412496
rect 672736 411182 672856 411210
rect 673472 411318 673592 411346
rect 672736 405686 672764 411182
rect 672540 405680 672592 405686
rect 672540 405622 672592 405628
rect 672724 405680 672776 405686
rect 672724 405622 672776 405628
rect 672552 386442 672580 405622
rect 673472 401606 673500 411318
rect 673460 401600 673512 401606
rect 673460 401542 673512 401548
rect 675300 401600 675352 401606
rect 675300 401542 675352 401548
rect 672540 386436 672592 386442
rect 672540 386378 672592 386384
rect 672816 386436 672868 386442
rect 672816 386378 672868 386384
rect 672828 372586 672856 386378
rect 673552 384056 673604 384062
rect 673552 383998 673604 384004
rect 672644 372558 672856 372586
rect 672644 353394 672672 372558
rect 672632 353388 672684 353394
rect 672632 353330 672684 353336
rect 672540 353252 672592 353258
rect 672540 353194 672592 353200
rect 672552 347750 672580 353194
rect 672540 347744 672592 347750
rect 672540 347686 672592 347692
rect 672724 347744 672776 347750
rect 672724 347686 672776 347692
rect 672736 328506 672764 347686
rect 673564 338745 673592 383998
rect 675312 383253 675340 401542
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675392 384056 675444 384062
rect 675392 383998 675444 384004
rect 675404 383860 675432 383998
rect 675312 383239 675418 383253
rect 675312 383225 675432 383239
rect 675404 382770 675432 383225
rect 673644 382764 673696 382770
rect 673644 382706 673696 382712
rect 675392 382764 675444 382770
rect 675392 382706 675444 382712
rect 673550 338736 673606 338745
rect 673550 338671 673606 338680
rect 672448 328500 672500 328506
rect 672448 328442 672500 328448
rect 672724 328500 672776 328506
rect 672724 328442 672776 328448
rect 672460 314786 672488 328442
rect 672538 314800 672594 314809
rect 672460 314758 672538 314786
rect 672538 314735 672594 314744
rect 672538 314528 672594 314537
rect 672538 314463 672594 314472
rect 672552 309126 672580 314463
rect 672540 309120 672592 309126
rect 672540 309062 672592 309068
rect 672816 309120 672868 309126
rect 672816 309062 672868 309068
rect 672828 289882 672856 309062
rect 673460 304972 673512 304978
rect 673460 304914 673512 304920
rect 672632 289876 672684 289882
rect 672632 289818 672684 289824
rect 672816 289876 672868 289882
rect 672816 289818 672868 289824
rect 672644 276060 672672 289818
rect 673472 283082 673500 304914
rect 673564 293298 673592 338671
rect 673656 338570 673684 382706
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 380175 675887 380231
rect 675407 379531 675887 379587
rect 675312 378901 675418 378929
rect 673828 372360 673880 372366
rect 673828 372302 673880 372308
rect 673644 338564 673696 338570
rect 673644 338506 673696 338512
rect 673656 293554 673684 338506
rect 673840 327146 673868 372302
rect 675312 370925 675340 378901
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675404 372366 675432 372751
rect 675392 372360 675444 372366
rect 675392 372302 675444 372308
rect 675407 371527 675887 371583
rect 675312 370897 675418 370925
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675390 338736 675446 338745
rect 675390 338671 675446 338680
rect 675392 338564 675444 338570
rect 675392 338506 675444 338512
rect 675404 338028 675432 338506
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675887 335031
rect 675407 334331 675887 334387
rect 675312 333701 675418 333729
rect 673828 327140 673880 327146
rect 673828 327082 673880 327088
rect 673840 304978 673868 327082
rect 675312 325725 675340 333701
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675404 327146 675432 327556
rect 675392 327140 675444 327146
rect 675392 327082 675444 327088
rect 675407 326327 675887 326383
rect 675312 325697 675418 325725
rect 673828 304972 673880 304978
rect 673828 304914 673880 304920
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 673644 293548 673696 293554
rect 673644 293490 673696 293496
rect 675024 293548 675076 293554
rect 675024 293490 675076 293496
rect 673564 293270 673868 293298
rect 673840 293214 673868 293270
rect 673828 293208 673880 293214
rect 673828 293150 673880 293156
rect 673460 283076 673512 283082
rect 673460 283018 673512 283024
rect 672644 276032 672764 276060
rect 672736 256714 672764 276032
rect 673736 266348 673788 266354
rect 673736 266290 673788 266296
rect 672552 256686 672764 256714
rect 672552 231849 672580 256686
rect 673644 247512 673696 247518
rect 673644 247454 673696 247460
rect 672538 231840 672594 231849
rect 672538 231775 672594 231784
rect 672906 231840 672962 231849
rect 672906 231775 672962 231784
rect 672920 212566 672948 231775
rect 672724 212560 672776 212566
rect 672724 212502 672776 212508
rect 672908 212560 672960 212566
rect 672908 212502 672960 212508
rect 672736 198762 672764 212502
rect 673552 203924 673604 203930
rect 673552 203866 673604 203872
rect 673460 203380 673512 203386
rect 673460 203322 673512 203328
rect 672540 198756 672592 198762
rect 672540 198698 672592 198704
rect 672724 198756 672776 198762
rect 672724 198698 672776 198704
rect 44640 195900 44692 195906
rect 44640 195842 44692 195848
rect 44652 193225 44680 195842
rect 672552 193225 672580 198698
rect 44454 193216 44510 193225
rect 44454 193151 44510 193160
rect 44638 193216 44694 193225
rect 44638 193151 44694 193160
rect 672538 193216 672594 193225
rect 672538 193151 672594 193160
rect 672906 193216 672962 193225
rect 672906 193151 672962 193160
rect 44468 173942 44496 193151
rect 672920 173942 672948 193151
rect 44456 173936 44508 173942
rect 44456 173878 44508 173884
rect 44732 173936 44784 173942
rect 44732 173878 44784 173884
rect 672724 173936 672776 173942
rect 672724 173878 672776 173884
rect 672908 173936 672960 173942
rect 672908 173878 672960 173884
rect 44744 160206 44772 173878
rect 44732 160200 44784 160206
rect 44732 160142 44784 160148
rect 672736 160138 672764 173878
rect 672540 160132 672592 160138
rect 672540 160074 672592 160080
rect 672724 160132 672776 160138
rect 672724 160074 672776 160080
rect 44640 160064 44692 160070
rect 44640 160006 44692 160012
rect 44652 154562 44680 160006
rect 44640 154556 44692 154562
rect 44640 154498 44692 154504
rect 44732 154556 44784 154562
rect 44732 154498 44784 154504
rect 44744 140826 44772 154498
rect 44732 140820 44784 140826
rect 44732 140762 44784 140768
rect 44640 140752 44692 140758
rect 44640 140694 44692 140700
rect 672552 140706 672580 160074
rect 673472 157350 673500 203322
rect 673564 158370 673592 203866
rect 673656 203386 673684 247454
rect 673748 237726 673776 266290
rect 673840 248198 673868 293150
rect 675036 293049 675064 293490
rect 675404 293214 675432 293692
rect 675392 293208 675444 293214
rect 675392 293150 675444 293156
rect 675022 293040 675078 293049
rect 675022 292975 675078 292984
rect 675206 293040 675262 293049
rect 675206 292975 675262 292984
rect 675390 293040 675446 293049
rect 675390 292975 675446 292984
rect 674932 283076 674984 283082
rect 674932 283018 674984 283024
rect 673920 276072 673972 276078
rect 673920 276014 673972 276020
rect 673828 248192 673880 248198
rect 673828 248134 673880 248140
rect 673736 237720 673788 237726
rect 673736 237662 673788 237668
rect 673644 203380 673696 203386
rect 673644 203322 673696 203328
rect 673748 192409 673776 237662
rect 673840 203930 673868 248134
rect 673932 247518 673960 276014
rect 674944 266354 674972 283018
rect 675220 276078 675248 292975
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675887 290031
rect 675407 289331 675887 289387
rect 675312 288701 675418 288729
rect 675312 280725 675340 288701
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675392 283076 675444 283082
rect 675392 283018 675444 283024
rect 675404 282540 675432 283018
rect 675407 281327 675887 281383
rect 675312 280697 675418 280725
rect 675208 276072 675260 276078
rect 675208 276014 675260 276020
rect 674932 266348 674984 266354
rect 674932 266290 674984 266296
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675404 248198 675432 248676
rect 675392 248192 675444 248198
rect 675392 248134 675444 248140
rect 675404 247518 675432 248039
rect 673920 247512 673972 247518
rect 673920 247454 673972 247460
rect 675392 247512 675444 247518
rect 675392 247454 675444 247460
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675887 245031
rect 675407 244331 675887 244387
rect 675312 243701 675418 243729
rect 675312 235725 675340 243701
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675392 237720 675444 237726
rect 675392 237662 675444 237668
rect 675404 237524 675432 237662
rect 675407 236327 675887 236383
rect 675312 235697 675418 235725
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 673828 203924 673880 203930
rect 673828 203866 673880 203872
rect 675392 203924 675444 203930
rect 675392 203866 675444 203872
rect 675404 203483 675432 203866
rect 675392 203380 675444 203386
rect 675392 203322 675444 203328
rect 675404 202844 675432 203322
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675887 199831
rect 675407 199131 675887 199187
rect 675312 198614 675432 198642
rect 673734 192400 673790 192409
rect 673734 192335 673790 192344
rect 673748 192030 673776 192335
rect 673736 192024 673788 192030
rect 673736 191966 673788 191972
rect 674012 192024 674064 192030
rect 674012 191966 674064 191972
rect 674024 173942 674052 191966
rect 675312 190525 675340 198614
rect 675404 198492 675432 198614
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675390 192400 675446 192409
rect 675390 192335 675446 192344
rect 675407 191127 675887 191183
rect 675312 190497 675418 190525
rect 673828 173936 673880 173942
rect 673828 173878 673880 173884
rect 674012 173936 674064 173942
rect 674012 173878 674064 173884
rect 673840 160138 673868 173878
rect 675407 160295 675887 160351
rect 673644 160132 673696 160138
rect 673644 160074 673696 160080
rect 673828 160132 673880 160138
rect 673828 160074 673880 160080
rect 673552 158364 673604 158370
rect 673552 158306 673604 158312
rect 673460 157344 673512 157350
rect 673460 157286 673512 157292
rect 44652 135266 44680 140694
rect 672552 140678 672672 140706
rect 44652 135238 44772 135266
rect 44744 121582 44772 135238
rect 44732 121576 44784 121582
rect 44732 121518 44784 121524
rect 44640 121440 44692 121446
rect 44640 121382 44692 121388
rect 672644 121394 672672 140678
rect 44178 120184 44234 120193
rect 44178 120119 44234 120128
rect 42338 115968 42394 115977
rect 42338 115903 42394 115912
rect 44192 110537 44220 120119
rect 44178 110528 44234 110537
rect 44178 110463 44234 110472
rect 44652 102082 44680 121382
rect 672644 121366 672764 121394
rect 672736 115938 672764 121366
rect 672724 115932 672776 115938
rect 672724 115874 672776 115880
rect 672816 115932 672868 115938
rect 672816 115874 672868 115880
rect 45466 110528 45522 110537
rect 45466 110463 45522 110472
rect 44560 102054 44680 102082
rect 44560 96626 44588 102054
rect 44272 96620 44324 96626
rect 44272 96562 44324 96568
rect 44548 96620 44600 96626
rect 44548 96562 44600 96568
rect 44284 77314 44312 96562
rect 44272 77308 44324 77314
rect 44272 77250 44324 77256
rect 44364 77308 44416 77314
rect 44364 77250 44416 77256
rect 44270 75848 44326 75857
rect 44376 75834 44404 77250
rect 44326 75806 44404 75834
rect 44270 75783 44326 75792
rect 44284 73273 44312 75783
rect 44270 73264 44326 73273
rect 44270 73199 44326 73208
rect 44284 68241 44312 73199
rect 44270 68232 44326 68241
rect 44270 68167 44326 68176
rect 42708 64660 42760 64666
rect 42708 64602 42760 64608
rect 42248 45688 42300 45694
rect 42248 45630 42300 45636
rect 42720 45626 42748 64602
rect 45480 47938 45508 110463
rect 672828 102202 672856 115874
rect 673472 112130 673500 157286
rect 673564 112810 673592 158306
rect 673656 147898 673684 160074
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675404 158370 675432 158508
rect 675392 158364 675444 158370
rect 675392 158306 675444 158312
rect 675404 157350 675432 157828
rect 675392 157344 675444 157350
rect 675392 157286 675444 157292
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675887 154831
rect 675407 154131 675887 154187
rect 675312 153501 675418 153529
rect 673644 147892 673696 147898
rect 673644 147834 673696 147840
rect 674012 147892 674064 147898
rect 674012 147834 674064 147840
rect 674024 140706 674052 147834
rect 675312 145525 675340 153501
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675392 147892 675444 147898
rect 675392 147834 675444 147840
rect 675404 147356 675432 147834
rect 675407 146127 675887 146183
rect 675312 145497 675418 145525
rect 673932 140678 674052 140706
rect 673932 121530 673960 140678
rect 673840 121502 673960 121530
rect 673552 112804 673604 112810
rect 673552 112746 673604 112752
rect 673460 112124 673512 112130
rect 673460 112066 673512 112072
rect 672816 102196 672868 102202
rect 672816 102138 672868 102144
rect 672724 102128 672776 102134
rect 672724 102070 672776 102076
rect 672736 96642 672764 102070
rect 672736 96614 672856 96642
rect 672828 82958 672856 96614
rect 672816 82952 672868 82958
rect 672816 82894 672868 82900
rect 672816 82748 672868 82754
rect 672816 82690 672868 82696
rect 45558 68232 45614 68241
rect 45558 68167 45614 68176
rect 45468 47932 45520 47938
rect 45468 47874 45520 47880
rect 45572 47802 45600 68167
rect 179420 47932 179472 47938
rect 179420 47874 179472 47880
rect 518808 47932 518860 47938
rect 518808 47874 518860 47880
rect 45560 47796 45612 47802
rect 45560 47738 45612 47744
rect 149060 47796 149112 47802
rect 149060 47738 149112 47744
rect 86316 47728 86368 47734
rect 86316 47670 86368 47676
rect 86328 47394 86356 47670
rect 86316 47388 86368 47394
rect 86316 47330 86368 47336
rect 42708 45620 42760 45626
rect 42708 45562 42760 45568
rect 86328 40225 86356 47330
rect 149072 47122 149100 47738
rect 179432 47530 179460 47874
rect 189172 47864 189224 47870
rect 189172 47806 189224 47812
rect 179420 47524 179472 47530
rect 179420 47466 179472 47472
rect 154578 47152 154634 47161
rect 149060 47116 149112 47122
rect 154578 47087 154580 47096
rect 149060 47058 149112 47064
rect 154632 47087 154634 47096
rect 173806 47152 173862 47161
rect 173806 47087 173862 47096
rect 188528 47116 188580 47122
rect 154580 47058 154632 47064
rect 145104 45688 145156 45694
rect 145104 45630 145156 45636
rect 140964 45620 141016 45626
rect 140964 45562 141016 45568
rect 140976 44198 141004 45562
rect 145116 44266 145144 45630
rect 145104 44260 145156 44266
rect 145104 44202 145156 44208
rect 140964 44192 141016 44198
rect 140964 44134 141016 44140
rect 133098 40248 133150 40254
rect 86314 40216 86370 40225
rect 133098 40190 133150 40196
rect 140976 40202 141004 44134
rect 143816 40248 143868 40254
rect 86314 40151 86370 40160
rect 133110 39984 133138 40190
rect 140976 40174 141036 40202
rect 145116 40202 145144 44202
rect 149072 40361 149100 47058
rect 173820 47054 173848 47087
rect 188528 47058 188580 47064
rect 173808 47048 173860 47054
rect 173808 46990 173860 46996
rect 186688 46980 186740 46986
rect 186688 46922 186740 46928
rect 186700 41820 186728 46922
rect 187327 41713 187383 42193
rect 188540 41820 188568 47058
rect 189184 41834 189212 47806
rect 212538 47696 212594 47705
rect 212538 47631 212540 47640
rect 212592 47631 212594 47640
rect 231582 47696 231638 47705
rect 231582 47631 231638 47640
rect 270498 47696 270554 47705
rect 270498 47631 270500 47640
rect 212540 47602 212592 47608
rect 195980 47592 196032 47598
rect 195980 47534 196032 47540
rect 198648 47592 198700 47598
rect 198740 47592 198792 47598
rect 198700 47540 198740 47546
rect 198648 47534 198792 47540
rect 192852 47116 192904 47122
rect 192852 47058 192904 47064
rect 189264 41880 189316 41886
rect 189184 41828 189264 41834
rect 191104 41880 191156 41886
rect 189184 41822 189316 41828
rect 191038 41828 191104 41834
rect 192300 41880 192352 41886
rect 191038 41822 191156 41828
rect 192234 41828 192300 41834
rect 192234 41822 192352 41828
rect 189184 41820 189304 41822
rect 189198 41806 189304 41820
rect 191038 41806 191144 41822
rect 192234 41806 192340 41822
rect 192864 41820 192892 47058
rect 194692 46980 194744 46986
rect 194692 46922 194744 46928
rect 193522 41818 193628 41834
rect 193522 41812 193640 41818
rect 193522 41806 193588 41812
rect 193588 41754 193640 41760
rect 194043 41713 194099 42193
rect 194704 41820 194732 46922
rect 195336 44260 195388 44266
rect 195336 44202 195388 44208
rect 195348 41834 195376 44202
rect 195428 41880 195480 41886
rect 195348 41828 195428 41834
rect 195348 41822 195480 41828
rect 195348 41820 195468 41822
rect 195992 41820 196020 47534
rect 198660 47518 198780 47534
rect 231596 47410 231624 47631
rect 270552 47631 270554 47640
rect 289634 47696 289690 47705
rect 289634 47631 289690 47640
rect 270500 47602 270552 47608
rect 231768 47524 231820 47530
rect 231768 47466 231820 47472
rect 251180 47524 251232 47530
rect 251180 47466 251232 47472
rect 270408 47524 270460 47530
rect 270408 47466 270460 47472
rect 231780 47410 231808 47466
rect 199016 47388 199068 47394
rect 199016 47330 199068 47336
rect 201408 47388 201460 47394
rect 231596 47382 231808 47410
rect 251192 47394 251220 47466
rect 270420 47394 270448 47466
rect 289648 47410 289676 47631
rect 303620 47592 303672 47598
rect 303620 47534 303672 47540
rect 304540 47592 304592 47598
rect 304540 47534 304592 47540
rect 359372 47592 359424 47598
rect 359372 47534 359424 47540
rect 361488 47592 361540 47598
rect 361488 47534 361540 47540
rect 289728 47456 289780 47462
rect 289648 47404 289728 47410
rect 289648 47398 289780 47404
rect 251180 47388 251232 47394
rect 201408 47330 201460 47336
rect 251180 47330 251232 47336
rect 270408 47388 270460 47394
rect 289648 47382 289768 47398
rect 303632 47394 303660 47534
rect 303620 47388 303672 47394
rect 270408 47330 270460 47336
rect 303620 47330 303672 47336
rect 195362 41806 195468 41820
rect 196452 41818 198504 41834
rect 199028 41820 199056 47330
rect 199660 47320 199712 47326
rect 199660 47262 199712 47268
rect 199568 41880 199620 41886
rect 199672 41834 199700 47262
rect 200856 47184 200908 47190
rect 200856 47126 200908 47132
rect 200868 41834 200896 47126
rect 201420 47122 201448 47330
rect 285588 47320 285640 47326
rect 285588 47262 285640 47268
rect 217968 47252 218020 47258
rect 217968 47194 218020 47200
rect 240140 47252 240192 47258
rect 240140 47194 240192 47200
rect 201408 47116 201460 47122
rect 201408 47058 201460 47064
rect 217980 47054 218008 47194
rect 201592 47048 201644 47054
rect 201592 46990 201644 46996
rect 217968 47048 218020 47054
rect 217968 46990 218020 46996
rect 201604 41834 201632 46990
rect 199620 41828 199700 41834
rect 199568 41822 199700 41828
rect 199580 41820 199700 41822
rect 200132 41820 200896 41834
rect 196440 41812 198516 41818
rect 196492 41806 198464 41812
rect 196440 41754 196492 41760
rect 199580 41806 199686 41820
rect 200132 41818 200882 41820
rect 200120 41812 200882 41818
rect 198464 41754 198516 41760
rect 200172 41806 200882 41812
rect 201526 41806 201632 41834
rect 200120 41754 200172 41760
rect 149058 40352 149114 40361
rect 149058 40287 149114 40296
rect 143816 40190 143868 40196
rect 141008 40118 141036 40174
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143072 40112 143124 40118
rect 143072 40054 143124 40060
rect 143356 40112 143408 40118
rect 143356 40054 143408 40060
rect 141008 39984 141036 40054
rect 143084 39984 143112 40054
rect 143368 39916 143396 40054
rect 143828 39916 143856 40190
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 145091 39706 145143 40000
rect 240152 39953 240180 47194
rect 242900 47184 242952 47190
rect 242900 47126 242952 47132
rect 242912 45558 242940 47126
rect 285600 47122 285628 47262
rect 299480 47184 299532 47190
rect 299480 47126 299532 47132
rect 247408 47116 247460 47122
rect 247408 47058 247460 47064
rect 285588 47116 285640 47122
rect 285588 47058 285640 47064
rect 242900 45552 242952 45558
rect 242900 45494 242952 45500
rect 240138 39944 240194 39953
rect 240138 39879 240194 39888
rect 242912 39817 242940 45494
rect 241242 39808 241298 39817
rect 241242 39743 241298 39752
rect 242898 39808 242954 39817
rect 242898 39743 242954 39752
rect 241256 39372 241284 39743
rect 247420 39581 247448 47058
rect 297732 45552 297784 45558
rect 297732 45494 297784 45500
rect 254032 44192 254084 44198
rect 254032 44134 254084 44140
rect 253940 41608 253992 41614
rect 253940 41550 253992 41556
rect 253952 39953 253980 41550
rect 253938 39944 253994 39953
rect 253938 39879 253994 39888
rect 254044 39710 254072 44134
rect 296904 41948 296956 41954
rect 296904 41890 296956 41896
rect 296916 41834 296944 41890
rect 297744 41834 297772 45494
rect 299492 42022 299520 47126
rect 303896 47116 303948 47122
rect 303896 47058 303948 47064
rect 299480 42016 299532 42022
rect 299480 41958 299532 41964
rect 302240 42016 302292 42022
rect 302240 41958 302292 41964
rect 297916 41880 297968 41886
rect 295311 41818 295472 41834
rect 295311 41812 295484 41818
rect 295311 41806 295432 41812
rect 296916 41806 297151 41834
rect 297744 41828 297916 41834
rect 297744 41822 297968 41828
rect 299492 41834 299520 41958
rect 300676 41880 300728 41886
rect 297744 41806 297956 41822
rect 299492 41806 299635 41834
rect 302252 41834 302280 41958
rect 300728 41828 302280 41834
rect 300676 41822 302280 41828
rect 300688 41806 302280 41822
rect 295432 41754 295484 41760
rect 302643 41713 302699 42193
rect 303908 41834 303936 47058
rect 304552 41834 304580 47534
rect 307576 47320 307628 47326
rect 307576 47262 307628 47268
rect 305736 47184 305788 47190
rect 305736 47126 305788 47132
rect 305000 42016 305052 42022
rect 305000 41958 305052 41964
rect 305012 41834 305040 41958
rect 305748 41834 305776 47126
rect 303172 41818 303315 41834
rect 303160 41812 303315 41818
rect 303212 41806 303315 41812
rect 303908 41806 303959 41834
rect 304552 41806 304603 41834
rect 305012 41818 305316 41834
rect 305012 41812 305328 41818
rect 305012 41806 305276 41812
rect 303160 41754 303212 41760
rect 305748 41806 305799 41834
rect 306443 41818 306604 41834
rect 306443 41812 306616 41818
rect 306443 41806 306564 41812
rect 305276 41754 305328 41760
rect 306564 41754 306616 41760
rect 306967 41713 307023 42193
rect 307588 41834 307616 47262
rect 309416 47252 309468 47258
rect 309416 47194 309468 47200
rect 352564 47252 352616 47258
rect 352564 47194 352616 47200
rect 308220 47116 308272 47122
rect 308220 47058 308272 47064
rect 308232 41834 308260 47058
rect 309428 41834 309456 47194
rect 351920 47184 351972 47190
rect 351920 47126 351972 47132
rect 307588 41806 307639 41834
rect 308232 41806 308283 41834
rect 308692 41818 309479 41834
rect 308680 41812 309479 41818
rect 308732 41806 309479 41812
rect 308680 41754 308732 41760
rect 310095 41713 310151 42193
rect 351932 41834 351960 47126
rect 352576 41970 352604 47194
rect 358728 47116 358780 47122
rect 358728 47058 358780 47064
rect 352576 41954 352696 41970
rect 352576 41948 352708 41954
rect 352576 41942 352656 41948
rect 352012 41880 352064 41886
rect 350106 41818 350212 41834
rect 351932 41828 352012 41834
rect 351932 41822 352064 41828
rect 351932 41820 352052 41822
rect 352576 41820 352604 41942
rect 352656 41890 352708 41896
rect 355508 41948 355560 41954
rect 355508 41890 355560 41896
rect 356980 41948 357032 41954
rect 356980 41890 357032 41896
rect 354312 41880 354364 41886
rect 355520 41834 355548 41890
rect 356992 41834 357020 41890
rect 354364 41828 354430 41834
rect 354312 41822 354430 41828
rect 350106 41812 350224 41818
rect 350106 41806 350172 41812
rect 351946 41806 352052 41820
rect 354324 41806 354430 41822
rect 355520 41806 357020 41834
rect 350172 41754 350224 41760
rect 357443 41713 357499 42193
rect 358004 41818 358110 41834
rect 358740 41820 358768 47058
rect 359384 41820 359412 47534
rect 361500 47394 361528 47534
rect 416780 47524 416832 47530
rect 416780 47466 416832 47472
rect 364156 47456 364208 47462
rect 364156 47398 364208 47404
rect 361488 47388 361540 47394
rect 361488 47330 361540 47336
rect 364168 47326 364196 47398
rect 414204 47388 414256 47394
rect 414204 47330 414256 47336
rect 362408 47320 362460 47326
rect 362408 47262 362460 47268
rect 364156 47320 364208 47326
rect 364156 47262 364208 47268
rect 406752 47320 406804 47326
rect 406752 47262 406804 47268
rect 360568 47184 360620 47190
rect 360568 47126 360620 47132
rect 359832 41948 359884 41954
rect 359832 41890 359884 41896
rect 359844 41834 359872 41890
rect 360476 41880 360528 41886
rect 357992 41812 358110 41818
rect 358044 41806 358110 41812
rect 359844 41806 359950 41834
rect 360580 41834 360608 47126
rect 361120 41948 361172 41954
rect 361120 41890 361172 41896
rect 360528 41828 360608 41834
rect 360476 41822 360608 41828
rect 360488 41820 360608 41822
rect 361132 41834 361160 41890
rect 360488 41806 360594 41820
rect 361132 41806 361238 41834
rect 357992 41754 358044 41760
rect 361767 41713 361823 42193
rect 362420 41820 362448 47262
rect 364248 47252 364300 47258
rect 364248 47194 364300 47200
rect 363052 47116 363104 47122
rect 363052 47058 363104 47064
rect 363064 41820 363092 47058
rect 364260 41834 364288 47194
rect 406764 47190 406792 47262
rect 407396 47252 407448 47258
rect 407396 47194 407448 47200
rect 406752 47184 406804 47190
rect 406752 47126 406804 47132
rect 363524 41820 364288 41834
rect 363524 41818 364274 41820
rect 363512 41812 364274 41818
rect 363564 41806 364274 41812
rect 363512 41754 363564 41760
rect 364895 41713 364951 42193
rect 404938 41818 405044 41834
rect 404938 41812 405056 41818
rect 404938 41806 405004 41812
rect 405004 41754 405056 41760
rect 405527 41713 405583 42193
rect 406764 41820 406792 47126
rect 407408 41970 407436 47194
rect 413560 47116 413612 47122
rect 413560 47058 413612 47064
rect 411536 42016 411588 42022
rect 407408 41954 407528 41970
rect 411588 41964 411760 41970
rect 411536 41958 411760 41964
rect 407408 41948 407540 41954
rect 407408 41942 407488 41948
rect 407408 41820 407436 41942
rect 407488 41890 407540 41896
rect 410248 41948 410300 41954
rect 410248 41890 410300 41896
rect 411168 41948 411220 41954
rect 411548 41942 411760 41958
rect 411168 41890 411220 41896
rect 409328 41880 409380 41886
rect 409262 41828 409328 41834
rect 409262 41822 409380 41828
rect 410260 41834 410288 41890
rect 411180 41834 411208 41890
rect 409262 41806 409368 41822
rect 410260 41806 410458 41834
rect 411102 41806 411208 41834
rect 411732 41820 411760 41942
rect 412243 41834 412299 42193
rect 412364 41880 412416 41886
rect 412243 41828 412364 41834
rect 412243 41822 412416 41828
rect 412243 41806 412404 41822
rect 412744 41818 412942 41834
rect 413572 41820 413600 47058
rect 414216 41820 414244 47330
rect 416792 47258 416820 47466
rect 417976 47388 418028 47394
rect 417976 47330 418028 47336
rect 418068 47388 418120 47394
rect 418068 47330 418120 47336
rect 471980 47388 472032 47394
rect 471980 47330 472032 47336
rect 416780 47252 416832 47258
rect 416780 47194 416832 47200
rect 417240 47252 417292 47258
rect 417240 47194 417292 47200
rect 414572 42016 414624 42022
rect 414572 41958 414624 41964
rect 415860 42016 415912 42022
rect 415860 41958 415912 41964
rect 414584 41834 414612 41958
rect 415492 41880 415544 41886
rect 412732 41812 412942 41818
rect 412243 41713 412299 41806
rect 412784 41806 412942 41812
rect 414584 41806 414782 41834
rect 415426 41828 415492 41834
rect 415426 41822 415544 41828
rect 415872 41834 415900 41958
rect 415426 41806 415532 41822
rect 415872 41806 416070 41834
rect 412732 41754 412784 41760
rect 416567 41713 416623 42193
rect 417252 41820 417280 47194
rect 417988 47122 418016 47330
rect 418080 47258 418108 47330
rect 461492 47320 461544 47326
rect 461492 47262 461544 47268
rect 418068 47252 418120 47258
rect 418068 47194 418120 47200
rect 419080 47252 419132 47258
rect 419080 47194 419132 47200
rect 417884 47116 417936 47122
rect 417884 47058 417936 47064
rect 417976 47116 418028 47122
rect 417976 47058 418028 47064
rect 417896 41820 417924 47058
rect 418252 42016 418304 42022
rect 418252 41958 418304 41964
rect 418264 41834 418292 41958
rect 419092 41834 419120 47194
rect 418264 41820 419120 41834
rect 419540 41880 419592 41886
rect 419695 41834 419751 42193
rect 459836 41880 459888 41886
rect 419592 41828 419751 41834
rect 419540 41822 419751 41828
rect 418264 41806 419106 41820
rect 419552 41806 419751 41822
rect 459711 41828 459836 41834
rect 459711 41822 459888 41828
rect 459711 41806 459876 41822
rect 419695 41713 419751 41806
rect 460327 41713 460383 42193
rect 461504 41834 461532 47262
rect 462136 47252 462188 47258
rect 462136 47194 462188 47200
rect 462148 41834 462176 47194
rect 468300 47184 468352 47190
rect 468300 47126 468352 47132
rect 466368 42016 466420 42022
rect 466368 41958 466420 41964
rect 462320 41948 462372 41954
rect 462320 41890 462372 41896
rect 465080 41948 465132 41954
rect 465080 41890 465132 41896
rect 466000 41948 466052 41954
rect 466000 41890 466052 41896
rect 462332 41834 462360 41890
rect 465092 41834 465120 41890
rect 466012 41834 466040 41890
rect 461504 41806 461551 41834
rect 462148 41806 462360 41834
rect 464035 41818 464200 41834
rect 464035 41812 464212 41818
rect 464035 41806 464160 41812
rect 465092 41806 465231 41834
rect 465875 41806 466040 41834
rect 466380 41834 466408 41958
rect 467043 41834 467099 42193
rect 467564 41880 467616 41886
rect 466380 41806 466519 41834
rect 467043 41818 467236 41834
rect 468312 41834 468340 47126
rect 468944 47116 468996 47122
rect 468944 47058 468996 47064
rect 468484 41880 468536 41886
rect 467616 41828 467715 41834
rect 467564 41822 467715 41828
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 464160 41754 464212 41760
rect 467043 41713 467099 41806
rect 467576 41806 467715 41822
rect 468312 41828 468484 41834
rect 468312 41822 468536 41828
rect 468956 41834 468984 47058
rect 469404 42016 469456 42022
rect 469404 41958 469456 41964
rect 470692 42016 470744 42022
rect 470692 41958 470744 41964
rect 469416 41834 469444 41958
rect 470704 41834 470732 41958
rect 468312 41806 468524 41822
rect 468956 41806 469003 41834
rect 469416 41806 469555 41834
rect 470060 41818 470199 41834
rect 470048 41812 470199 41818
rect 467196 41754 467248 41760
rect 470100 41806 470199 41812
rect 470704 41806 470843 41834
rect 470048 41754 470100 41760
rect 471367 41713 471423 42193
rect 471992 41834 472020 47330
rect 518820 47326 518848 47874
rect 527456 47864 527508 47870
rect 527456 47806 527508 47812
rect 526812 47388 526864 47394
rect 526812 47330 526864 47336
rect 516324 47320 516376 47326
rect 516324 47262 516376 47268
rect 518808 47320 518860 47326
rect 518808 47262 518860 47268
rect 473820 47252 473872 47258
rect 473820 47194 473872 47200
rect 473084 42016 473136 42022
rect 473084 41958 473136 41964
rect 472532 41880 472584 41886
rect 471992 41806 472039 41834
rect 473096 41834 473124 41958
rect 473832 41834 473860 47194
rect 514484 46980 514536 46986
rect 514484 46922 514536 46928
rect 474372 41948 474424 41954
rect 474372 41890 474424 41896
rect 474384 41834 474412 41890
rect 474495 41834 474551 42193
rect 472584 41828 472683 41834
rect 472532 41822 472683 41828
rect 472544 41806 472683 41822
rect 473096 41806 473879 41834
rect 474384 41806 474551 41834
rect 514496 41820 514524 46922
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 516336 41820 516364 47262
rect 516968 47252 517020 47258
rect 516968 47194 517020 47200
rect 516980 41834 517008 47194
rect 523776 47116 523828 47122
rect 523776 47058 523828 47064
rect 522488 46980 522540 46986
rect 522488 46922 522540 46928
rect 518900 41880 518952 41886
rect 516980 41820 517100 41834
rect 516994 41818 517100 41820
rect 518834 41828 518900 41834
rect 518834 41822 518952 41828
rect 516994 41812 517112 41818
rect 516994 41806 517060 41812
rect 518834 41806 518940 41822
rect 520030 41818 520136 41834
rect 520030 41812 520148 41818
rect 520030 41806 520096 41812
rect 517060 41754 517112 41760
rect 520096 41754 520148 41760
rect 520647 41713 520703 42193
rect 521318 41818 521424 41834
rect 521318 41812 521436 41818
rect 521318 41806 521384 41812
rect 521384 41754 521436 41760
rect 521843 41713 521899 42193
rect 522500 41820 522528 46922
rect 523224 41948 523276 41954
rect 523224 41890 523276 41896
rect 523236 41834 523264 41890
rect 523158 41806 523264 41834
rect 523788 41820 523816 47058
rect 526824 46986 526852 47330
rect 527468 47190 527496 47806
rect 672828 47802 672856 82690
rect 528652 47796 528704 47802
rect 528652 47738 528704 47744
rect 672816 47796 672868 47802
rect 672816 47738 672868 47744
rect 527456 47184 527508 47190
rect 527456 47126 527508 47132
rect 526812 46980 526864 46986
rect 526812 46922 526864 46928
rect 524880 41880 524932 41886
rect 524354 41818 524460 41834
rect 524971 41834 525027 42193
rect 524932 41828 525027 41834
rect 524880 41822 525027 41828
rect 524354 41812 524472 41818
rect 524354 41806 524420 41812
rect 524892 41806 525027 41822
rect 525642 41818 525748 41834
rect 525642 41812 525760 41818
rect 525642 41806 525708 41812
rect 524420 41754 524472 41760
rect 524971 41713 525027 41806
rect 525708 41754 525760 41760
rect 526167 41713 526223 42193
rect 526824 41820 526852 46922
rect 527468 41970 527496 47126
rect 527376 41954 527496 41970
rect 527364 41948 527496 41954
rect 527416 41942 527496 41948
rect 527364 41890 527416 41896
rect 527468 41820 527496 41942
rect 528664 41834 528692 47738
rect 569132 47116 569184 47122
rect 569132 47058 569184 47064
rect 527928 41820 528692 41834
rect 527928 41818 528678 41820
rect 527916 41812 528678 41818
rect 527968 41806 528678 41812
rect 527916 41754 527968 41760
rect 529295 41713 529351 42193
rect 252100 39704 252152 39710
rect 252100 39646 252152 39652
rect 254032 39704 254084 39710
rect 254032 39646 254084 39652
rect 247342 39553 247448 39581
rect 252112 39372 252140 39646
rect 569144 39644 569172 47058
rect 634820 46980 634872 46986
rect 634820 46922 634872 46928
rect 579160 45552 579212 45558
rect 579160 45494 579212 45500
rect 569224 44192 569276 44198
rect 569224 44134 569276 44140
rect 569236 40225 569264 44134
rect 579172 40225 579200 45494
rect 622950 40488 623006 40497
rect 622950 40423 623006 40432
rect 569222 40216 569278 40225
rect 569222 40151 569278 40160
rect 579158 40216 579214 40225
rect 579158 40151 579214 40160
rect 579172 39644 579200 40151
rect 622964 39681 622992 40423
rect 634832 40225 634860 46922
rect 673472 45558 673500 112066
rect 673564 47870 673592 112746
rect 673840 102202 673868 121502
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675404 112810 675432 113283
rect 675392 112804 675444 112810
rect 675392 112746 675444 112752
rect 675404 112130 675432 112639
rect 675392 112124 675444 112130
rect 675392 112066 675444 112072
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 109575 675887 109631
rect 675407 108931 675887 108987
rect 675312 108310 675418 108338
rect 673644 102196 673696 102202
rect 673644 102138 673696 102144
rect 673828 102196 673880 102202
rect 673828 102138 673880 102144
rect 673656 102066 673684 102138
rect 673644 102060 673696 102066
rect 673644 102002 673696 102008
rect 673656 47938 673684 102002
rect 675312 100314 675340 108310
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675404 102066 675432 102151
rect 675392 102060 675444 102066
rect 675392 102002 675444 102008
rect 675407 100927 675887 100983
rect 675312 100286 675418 100314
rect 673644 47932 673696 47938
rect 673644 47874 673696 47880
rect 673552 47864 673604 47870
rect 673552 47806 673604 47812
rect 673460 45552 673512 45558
rect 673460 45494 673512 45500
rect 632978 40216 633034 40225
rect 632978 40151 633034 40160
rect 634818 40216 634874 40225
rect 634818 40151 634874 40160
rect 622950 39672 623006 39681
rect 632992 39644 633020 40151
rect 622950 39607 623006 39616
<< via2 >>
rect 333518 997600 333574 997656
rect 45926 996512 45982 996568
rect 45466 990120 45522 990176
rect 39670 908112 39726 908168
rect 40406 907976 40462 908032
rect 40406 888936 40462 888992
rect 40130 879960 40186 880016
rect 41418 875064 41474 875120
rect 39854 837528 39910 837584
rect 39854 832632 39910 832688
rect 39670 827464 39726 827520
rect 39762 492904 39818 492960
rect 39946 455368 40002 455424
rect 39670 451832 39726 451888
rect 39670 440952 39726 441008
rect 42246 400152 42302 400208
rect 42614 400152 42670 400208
rect 39762 120128 39818 120184
rect 41418 115912 41474 115968
rect 39394 84224 39450 84280
rect 44362 917224 44418 917280
rect 160098 990664 160154 990720
rect 173806 990664 173862 990720
rect 193218 990548 193274 990584
rect 193218 990528 193220 990548
rect 193220 990528 193272 990548
rect 193272 990528 193274 990548
rect 212446 990548 212502 990584
rect 212446 990528 212448 990548
rect 212448 990528 212500 990548
rect 212500 990528 212502 990548
rect 672630 996512 672686 996568
rect 585690 996376 585746 996432
rect 672446 996376 672502 996432
rect 537850 995424 537906 995480
rect 538034 995424 538090 995480
rect 576858 990564 576860 990584
rect 576860 990564 576912 990584
rect 576912 990564 576914 990584
rect 576858 990528 576914 990564
rect 596086 990528 596142 990584
rect 540978 990428 540980 990448
rect 540980 990428 541032 990448
rect 541032 990428 541034 990448
rect 540978 990392 541034 990428
rect 560206 990392 560262 990448
rect 44454 835216 44510 835272
rect 672538 828688 672594 828744
rect 44730 828008 44786 828064
rect 673366 908112 673422 908168
rect 672630 826104 672686 826160
rect 673274 826104 673330 826160
rect 673182 823656 673238 823712
rect 672998 792104 673054 792160
rect 673182 792104 673238 792160
rect 672814 753480 672870 753536
rect 672998 753480 673054 753536
rect 672998 618160 673054 618216
rect 672814 618024 672870 618080
rect 44546 560224 44602 560280
rect 44914 560224 44970 560280
rect 673090 511400 673146 511456
rect 673274 511400 673330 511456
rect 672998 509088 673054 509144
rect 44454 493176 44510 493232
rect 44546 488552 44602 488608
rect 44362 448568 44418 448624
rect 673274 502288 673330 502344
rect 673458 888664 673514 888720
rect 677874 918584 677930 918640
rect 677598 915320 677654 915376
rect 677598 912736 677654 912792
rect 677874 912736 677930 912792
rect 677874 908112 677930 908168
rect 677782 907704 677838 907760
rect 675298 888664 675354 888720
rect 676126 828688 676182 828744
rect 676126 823656 676182 823712
rect 673458 685344 673514 685400
rect 675390 685344 675446 685400
rect 676126 514120 676182 514176
rect 676126 509088 676182 509144
rect 673642 502288 673698 502344
rect 673366 483112 673422 483168
rect 673366 482976 673422 483032
rect 678058 477536 678114 477592
rect 677874 469920 677930 469976
rect 673366 467472 673422 467528
rect 673274 463664 673330 463720
rect 673458 463664 673514 463720
rect 673458 463528 673514 463584
rect 673734 463528 673790 463584
rect 673090 427896 673146 427952
rect 673550 444352 673606 444408
rect 673734 444352 673790 444408
rect 673366 420824 673422 420880
rect 677414 427896 677470 427952
rect 677598 425720 677654 425776
rect 673550 338680 673606 338736
rect 672538 314744 672594 314800
rect 672538 314472 672594 314528
rect 675390 338680 675446 338736
rect 672538 231784 672594 231840
rect 672906 231784 672962 231840
rect 44454 193160 44510 193216
rect 44638 193160 44694 193216
rect 672538 193160 672594 193216
rect 672906 193160 672962 193216
rect 675022 292984 675078 293040
rect 675206 292984 675262 293040
rect 675390 292984 675446 293040
rect 673734 192344 673790 192400
rect 675390 192344 675446 192400
rect 44178 120128 44234 120184
rect 42338 115912 42394 115968
rect 44178 110472 44234 110528
rect 45466 110472 45522 110528
rect 44270 75792 44326 75848
rect 44270 73208 44326 73264
rect 44270 68176 44326 68232
rect 45558 68176 45614 68232
rect 154578 47116 154634 47152
rect 154578 47096 154580 47116
rect 154580 47096 154632 47116
rect 154632 47096 154634 47116
rect 173806 47096 173862 47152
rect 86314 40160 86370 40216
rect 212538 47660 212594 47696
rect 212538 47640 212540 47660
rect 212540 47640 212592 47660
rect 212592 47640 212594 47660
rect 231582 47640 231638 47696
rect 270498 47660 270554 47696
rect 270498 47640 270500 47660
rect 270500 47640 270552 47660
rect 270552 47640 270554 47660
rect 289634 47640 289690 47696
rect 149058 40296 149114 40352
rect 240138 39888 240194 39944
rect 241242 39752 241298 39808
rect 242898 39752 242954 39808
rect 253938 39888 253994 39944
rect 622950 40432 623006 40488
rect 569222 40160 569278 40216
rect 579158 40160 579214 40216
rect 632978 40160 633034 40216
rect 634818 40160 634874 40216
rect 622950 39616 623006 39672
<< metal3 >>
rect 333513 997658 333579 997661
rect 333500 997656 333579 997658
rect 333500 997600 333518 997656
rect 333574 997600 333579 997656
rect 333500 997598 333579 997600
rect 333513 997595 333579 997598
rect 45921 996570 45987 996573
rect 341014 996570 341074 997628
rect 580796 997598 581746 997658
rect 581686 997522 581746 997598
rect 585734 997522 585794 997628
rect 581686 997462 585794 997522
rect 585734 997114 585794 997462
rect 585734 997054 585978 997114
rect 45921 996568 341074 996570
rect 45921 996512 45926 996568
rect 45982 996512 341074 996568
rect 45921 996510 341074 996512
rect 585918 996570 585978 997054
rect 672625 996570 672691 996573
rect 585918 996568 672691 996570
rect 585918 996512 672630 996568
rect 672686 996512 672691 996568
rect 585918 996510 672691 996512
rect 45921 996507 45987 996510
rect 672625 996507 672691 996510
rect 585685 996434 585751 996437
rect 672441 996434 672507 996437
rect 585685 996432 672507 996434
rect 585685 996376 585690 996432
rect 585746 996376 672446 996432
rect 672502 996376 672507 996432
rect 585685 996374 672507 996376
rect 585685 996371 585751 996374
rect 672441 996371 672507 996374
rect 537845 995482 537911 995485
rect 538029 995482 538095 995485
rect 537845 995480 538095 995482
rect 537845 995424 537850 995480
rect 537906 995424 538034 995480
rect 538090 995424 538095 995480
rect 537845 995422 538095 995424
rect 537845 995419 537911 995422
rect 538029 995419 538095 995422
rect 160093 990722 160159 990725
rect 173801 990722 173867 990725
rect 160093 990720 173867 990722
rect 160093 990664 160098 990720
rect 160154 990664 173806 990720
rect 173862 990664 173867 990720
rect 160093 990662 173867 990664
rect 160093 990659 160159 990662
rect 173801 990659 173867 990662
rect 193213 990586 193279 990589
rect 212441 990586 212507 990589
rect 193213 990584 212507 990586
rect 193213 990528 193218 990584
rect 193274 990528 212446 990584
rect 212502 990528 212507 990584
rect 193213 990526 212507 990528
rect 193213 990523 193279 990526
rect 212441 990523 212507 990526
rect 576853 990586 576919 990589
rect 596081 990586 596147 990589
rect 576853 990584 596147 990586
rect 576853 990528 576858 990584
rect 576914 990528 596086 990584
rect 596142 990528 596147 990584
rect 576853 990526 596147 990528
rect 576853 990523 576919 990526
rect 596081 990523 596147 990526
rect 540973 990450 541039 990453
rect 560201 990450 560267 990453
rect 540973 990448 560267 990450
rect 540973 990392 540978 990448
rect 541034 990392 560206 990448
rect 560262 990392 560267 990448
rect 540973 990390 560267 990392
rect 540973 990387 541039 990390
rect 560201 990387 560267 990390
rect 45461 990178 45527 990181
rect 676254 990178 676260 990180
rect 45461 990176 676260 990178
rect 45461 990120 45466 990176
rect 45522 990120 676260 990176
rect 45461 990118 676260 990120
rect 45461 990115 45527 990118
rect 676254 990116 676260 990118
rect 676324 990116 676330 990180
rect 39468 922254 39866 922314
rect 39806 921770 39866 922254
rect 39438 921710 39866 921770
rect 39438 919730 39498 921710
rect 39438 919700 39866 919730
rect 39468 919670 39866 919700
rect 39806 919322 39866 919670
rect 39438 919262 39866 919322
rect 39438 917282 39498 919262
rect 677542 918580 677548 918644
rect 677612 918642 677618 918644
rect 677869 918642 677935 918645
rect 677612 918640 677935 918642
rect 677612 918584 677874 918640
rect 677930 918584 677935 918640
rect 677612 918582 677935 918584
rect 677612 918580 677618 918582
rect 677869 918579 677935 918582
rect 44357 917282 44423 917285
rect 39438 917280 44423 917282
rect 39438 917252 44362 917280
rect 39468 917224 44362 917252
rect 44418 917224 44423 917280
rect 39468 917222 44423 917224
rect 44357 917219 44423 917222
rect 677593 915378 677659 915381
rect 677593 915376 678132 915378
rect 677593 915320 677598 915376
rect 677654 915320 678132 915376
rect 677593 915318 678132 915320
rect 677593 915315 677659 915318
rect 677593 912794 677659 912797
rect 677869 912794 677935 912797
rect 677593 912792 678132 912794
rect 677593 912736 677598 912792
rect 677654 912736 677874 912792
rect 677930 912736 678132 912792
rect 677593 912734 678132 912736
rect 677593 912731 677659 912734
rect 677869 912731 677935 912734
rect 39665 908170 39731 908173
rect 40534 908170 40540 908172
rect 39665 908168 40540 908170
rect 39665 908112 39670 908168
rect 39726 908112 40540 908168
rect 39665 908110 40540 908112
rect 39665 908107 39731 908110
rect 40534 908108 40540 908110
rect 40604 908108 40610 908172
rect 673361 908170 673427 908173
rect 677869 908170 677935 908173
rect 673361 908168 678162 908170
rect 673361 908112 673366 908168
rect 673422 908112 677874 908168
rect 677930 908112 678162 908168
rect 673361 908110 678162 908112
rect 673361 908107 673427 908110
rect 677869 908107 677935 908110
rect 40401 908034 40467 908037
rect 40534 908034 40540 908036
rect 40401 908032 40540 908034
rect 40401 907976 40406 908032
rect 40462 907976 40540 908032
rect 40401 907974 40540 907976
rect 40401 907971 40467 907974
rect 40534 907972 40540 907974
rect 40604 907972 40610 908036
rect 676254 907700 676260 907764
rect 676324 907762 676330 907764
rect 677777 907762 677843 907765
rect 676324 907760 677843 907762
rect 676324 907704 677782 907760
rect 677838 907704 677843 907760
rect 678102 907732 678162 908110
rect 676324 907702 677843 907704
rect 676324 907700 676330 907702
rect 677777 907699 677843 907702
rect 40401 888994 40467 888997
rect 40358 888992 40467 888994
rect 40358 888936 40406 888992
rect 40462 888936 40467 888992
rect 40358 888931 40467 888936
rect 40358 888860 40418 888931
rect 40350 888796 40356 888860
rect 40420 888796 40426 888860
rect 673453 888722 673519 888725
rect 675293 888722 675359 888725
rect 673453 888720 675359 888722
rect 673453 888664 673458 888720
rect 673514 888664 675298 888720
rect 675354 888664 675359 888720
rect 673453 888662 675359 888664
rect 673453 888659 673519 888662
rect 675293 888659 675359 888662
rect 40125 880018 40191 880021
rect 39652 880016 40191 880018
rect 39652 879960 40130 880016
rect 40186 879960 40191 880016
rect 39652 879958 40191 879960
rect 40125 879955 40191 879958
rect 41413 875122 41479 875125
rect 39652 875120 41479 875122
rect 39652 875064 41418 875120
rect 41474 875064 41479 875120
rect 39652 875062 41479 875064
rect 41413 875059 41479 875062
rect 39982 855810 39988 855812
rect 39806 855750 39988 855810
rect 39806 855540 39866 855750
rect 39982 855748 39988 855750
rect 40052 855748 40058 855812
rect 39798 855476 39804 855540
rect 39868 855476 39874 855540
rect 39849 837588 39915 837589
rect 39798 837586 39804 837588
rect 39758 837526 39804 837586
rect 39868 837584 39915 837588
rect 39910 837528 39915 837584
rect 39798 837524 39804 837526
rect 39868 837524 39915 837528
rect 39849 837523 39915 837524
rect 44449 835274 44515 835277
rect 39652 835272 44515 835274
rect 39652 835216 44454 835272
rect 44510 835216 44515 835272
rect 39652 835214 44515 835216
rect 44449 835211 44515 835214
rect 39849 832690 39915 832693
rect 39982 832690 39988 832692
rect 39849 832688 39988 832690
rect 39849 832632 39854 832688
rect 39910 832632 39988 832688
rect 39849 832630 39988 832632
rect 39849 832627 39915 832630
rect 39982 832628 39988 832630
rect 40052 832628 40058 832692
rect 672533 828746 672599 828749
rect 676121 828746 676187 828749
rect 672533 828744 677794 828746
rect 672533 828688 672538 828744
rect 672594 828688 676126 828744
rect 676182 828688 677794 828744
rect 672533 828686 677794 828688
rect 672533 828683 672599 828686
rect 676121 828683 676187 828686
rect 677734 828580 677794 828686
rect 44725 828066 44791 828069
rect 39806 828064 44791 828066
rect 39806 828008 44730 828064
rect 44786 828008 44791 828064
rect 39806 828006 44791 828008
rect 39806 827794 39866 828006
rect 44725 828003 44791 828006
rect 39652 827734 39866 827794
rect 39665 827522 39731 827525
rect 39806 827522 39866 827734
rect 39665 827520 39866 827522
rect 39665 827464 39670 827520
rect 39726 827464 39866 827520
rect 39665 827462 39866 827464
rect 39665 827459 39731 827462
rect 672625 826162 672691 826165
rect 673269 826162 673335 826165
rect 672625 826160 677764 826162
rect 672625 826104 672630 826160
rect 672686 826104 673274 826160
rect 673330 826104 677764 826160
rect 672625 826102 677764 826104
rect 672625 826099 672691 826102
rect 673269 826099 673335 826102
rect 673177 823714 673243 823717
rect 676121 823714 676187 823717
rect 673177 823712 677764 823714
rect 673177 823656 673182 823712
rect 673238 823656 676126 823712
rect 676182 823656 677764 823712
rect 673177 823654 677764 823656
rect 673177 823651 673243 823654
rect 676121 823651 676187 823654
rect 40350 797676 40356 797740
rect 40420 797676 40426 797740
rect 40358 797604 40418 797676
rect 40350 797540 40356 797604
rect 40420 797540 40426 797604
rect 40350 792100 40356 792164
rect 40420 792162 40426 792164
rect 40534 792162 40540 792164
rect 40420 792102 40540 792162
rect 40420 792100 40426 792102
rect 40534 792100 40540 792102
rect 40604 792100 40610 792164
rect 672993 792162 673059 792165
rect 673177 792162 673243 792165
rect 672993 792160 673243 792162
rect 672993 792104 672998 792160
rect 673054 792104 673182 792160
rect 673238 792104 673243 792160
rect 672993 792102 673243 792104
rect 672993 792099 673059 792102
rect 673177 792099 673243 792102
rect 40534 778562 40540 778564
rect 40358 778502 40540 778562
rect 40358 778292 40418 778502
rect 40534 778500 40540 778502
rect 40604 778500 40610 778564
rect 40350 778228 40356 778292
rect 40420 778228 40426 778292
rect 40350 763132 40356 763196
rect 40420 763194 40426 763196
rect 40718 763194 40724 763196
rect 40420 763134 40724 763194
rect 40420 763132 40426 763134
rect 40718 763132 40724 763134
rect 40788 763132 40794 763196
rect 40350 753476 40356 753540
rect 40420 753538 40426 753540
rect 40718 753538 40724 753540
rect 40420 753478 40724 753538
rect 40420 753476 40426 753478
rect 40718 753476 40724 753478
rect 40788 753476 40794 753540
rect 672809 753538 672875 753541
rect 672993 753538 673059 753541
rect 672809 753536 673059 753538
rect 672809 753480 672814 753536
rect 672870 753480 672998 753536
rect 673054 753480 673059 753536
rect 672809 753478 673059 753480
rect 672809 753475 672875 753478
rect 672993 753475 673059 753478
rect 40350 750620 40356 750684
rect 40420 750682 40426 750684
rect 40420 750622 40602 750682
rect 40420 750620 40426 750622
rect 40350 750348 40356 750412
rect 40420 750410 40426 750412
rect 40542 750410 40602 750622
rect 40420 750350 40602 750410
rect 40420 750348 40426 750350
rect 40166 731308 40172 731372
rect 40236 731308 40242 731372
rect 40174 731234 40234 731308
rect 40718 731234 40724 731236
rect 40174 731174 40724 731234
rect 40718 731172 40724 731174
rect 40788 731172 40794 731236
rect 40350 712268 40356 712332
rect 40420 712330 40426 712332
rect 40718 712330 40724 712332
rect 40420 712270 40724 712330
rect 40420 712268 40426 712270
rect 40718 712268 40724 712270
rect 40788 712268 40794 712332
rect 40350 702068 40356 702132
rect 40420 702130 40426 702132
rect 40902 702130 40908 702132
rect 40420 702070 40908 702130
rect 40420 702068 40426 702070
rect 40902 702068 40908 702070
rect 40972 702068 40978 702132
rect 40534 695268 40540 695332
rect 40604 695330 40610 695332
rect 40902 695330 40908 695332
rect 40604 695270 40908 695330
rect 40604 695268 40610 695270
rect 40902 695268 40908 695270
rect 40972 695268 40978 695332
rect 673453 685402 673519 685405
rect 675385 685402 675451 685405
rect 673453 685400 675451 685402
rect 673453 685344 673458 685400
rect 673514 685344 675390 685400
rect 675446 685344 675451 685400
rect 673453 685342 675451 685344
rect 673453 685339 673519 685342
rect 675385 685339 675451 685342
rect 40166 673372 40172 673436
rect 40236 673434 40242 673436
rect 40534 673434 40540 673436
rect 40236 673374 40540 673434
rect 40236 673372 40242 673374
rect 40534 673372 40540 673374
rect 40604 673372 40610 673436
rect 40534 654394 40540 654396
rect 40174 654334 40540 654394
rect 40174 654260 40234 654334
rect 40534 654332 40540 654334
rect 40604 654332 40610 654396
rect 40166 654196 40172 654260
rect 40236 654196 40242 654260
rect 40350 634748 40356 634812
rect 40420 634810 40426 634812
rect 40902 634810 40908 634812
rect 40420 634750 40908 634810
rect 40420 634748 40426 634750
rect 40902 634748 40908 634750
rect 40972 634748 40978 634812
rect 672993 618218 673059 618221
rect 672993 618216 673194 618218
rect 672993 618160 672998 618216
rect 673054 618160 673194 618216
rect 672993 618158 673194 618160
rect 672993 618155 673059 618158
rect 672809 618082 672875 618085
rect 673134 618082 673194 618158
rect 672809 618080 673194 618082
rect 672809 618024 672814 618080
rect 672870 618024 673194 618080
rect 672809 618022 673194 618024
rect 672809 618019 672875 618022
rect 40534 598980 40540 599044
rect 40604 599042 40610 599044
rect 40902 599042 40908 599044
rect 40604 598982 40908 599042
rect 40604 598980 40610 598982
rect 40902 598980 40908 598982
rect 40972 598980 40978 599044
rect 40166 565932 40172 565996
rect 40236 565932 40242 565996
rect 40174 565724 40234 565932
rect 40166 565660 40172 565724
rect 40236 565660 40242 565724
rect 44541 560282 44607 560285
rect 44909 560282 44975 560285
rect 44541 560280 44975 560282
rect 44541 560224 44546 560280
rect 44602 560224 44914 560280
rect 44970 560224 44975 560280
rect 44541 560222 44975 560224
rect 44541 560219 44607 560222
rect 44909 560219 44975 560222
rect 40166 550564 40172 550628
rect 40236 550626 40242 550628
rect 40534 550626 40540 550628
rect 40236 550566 40540 550626
rect 40236 550564 40242 550566
rect 40534 550564 40540 550566
rect 40604 550564 40610 550628
rect 40534 540908 40540 540972
rect 40604 540970 40610 540972
rect 40902 540970 40908 540972
rect 40604 540910 40908 540970
rect 40604 540908 40610 540910
rect 40902 540908 40908 540910
rect 40972 540908 40978 540972
rect 40902 521930 40908 521932
rect 40174 521870 40908 521930
rect 40174 521796 40234 521870
rect 40902 521868 40908 521870
rect 40972 521868 40978 521932
rect 40166 521732 40172 521796
rect 40236 521732 40242 521796
rect 676121 514178 676187 514181
rect 676121 514176 677794 514178
rect 676121 514120 676126 514176
rect 676182 514120 677794 514176
rect 676121 514118 677794 514120
rect 676121 514115 676187 514118
rect 677734 514012 677794 514118
rect 673085 511458 673151 511461
rect 673269 511458 673335 511461
rect 673085 511456 677764 511458
rect 673085 511400 673090 511456
rect 673146 511400 673274 511456
rect 673330 511400 677764 511456
rect 673085 511398 677764 511400
rect 673085 511395 673151 511398
rect 673269 511395 673335 511398
rect 672993 509146 673059 509149
rect 676121 509146 676187 509149
rect 672993 509144 677764 509146
rect 672993 509088 672998 509144
rect 673054 509088 676126 509144
rect 676182 509088 677764 509144
rect 672993 509086 677764 509088
rect 672993 509083 673059 509086
rect 676121 509083 676187 509086
rect 40166 508058 40172 508060
rect 39990 507998 40172 508058
rect 39990 507788 40050 507998
rect 40166 507996 40172 507998
rect 40236 507996 40242 508060
rect 39982 507724 39988 507788
rect 40052 507724 40058 507788
rect 673269 502346 673335 502349
rect 673637 502346 673703 502349
rect 673269 502344 673703 502346
rect 673269 502288 673274 502344
rect 673330 502288 673642 502344
rect 673698 502288 673703 502344
rect 673269 502286 673703 502288
rect 673269 502283 673335 502286
rect 673637 502283 673703 502286
rect 44449 493234 44515 493237
rect 39652 493232 44515 493234
rect 39652 493176 44454 493232
rect 44510 493176 44515 493232
rect 39652 493174 44515 493176
rect 39806 492965 39866 493174
rect 44449 493171 44515 493174
rect 39757 492960 39866 492965
rect 39757 492904 39762 492960
rect 39818 492904 39866 492960
rect 39757 492902 39866 492904
rect 39757 492899 39823 492902
rect 44541 488610 44607 488613
rect 39806 488608 44607 488610
rect 39806 488552 44546 488608
rect 44602 488552 44607 488608
rect 39806 488550 44607 488552
rect 39806 488338 39866 488550
rect 44541 488547 44607 488550
rect 39652 488278 39866 488338
rect 673361 483170 673427 483173
rect 673318 483168 673427 483170
rect 673318 483112 673366 483168
rect 673422 483112 673427 483168
rect 673318 483107 673427 483112
rect 673318 483037 673378 483107
rect 673318 483032 673427 483037
rect 673318 482976 673366 483032
rect 673422 482976 673427 483032
rect 673318 482974 673427 482976
rect 673361 482971 673427 482974
rect 677542 477532 677548 477596
rect 677612 477594 677618 477596
rect 678053 477594 678119 477597
rect 677612 477592 678119 477594
rect 677612 477536 678058 477592
rect 678114 477536 678119 477592
rect 677612 477534 678119 477536
rect 677612 477532 677618 477534
rect 678053 477531 678119 477534
rect 677869 469978 677935 469981
rect 677869 469976 678132 469978
rect 677869 469920 677874 469976
rect 677930 469920 678132 469976
rect 677869 469918 678132 469920
rect 677869 469915 677935 469918
rect 673361 467530 673427 467533
rect 673361 467528 678132 467530
rect 673361 467472 673366 467528
rect 673422 467500 678132 467528
rect 673422 467472 678162 467500
rect 673361 467470 678162 467472
rect 673361 467467 673427 467470
rect 678102 465052 678162 467470
rect 673269 463722 673335 463725
rect 673453 463722 673519 463725
rect 673269 463720 673519 463722
rect 673269 463664 673274 463720
rect 673330 463664 673458 463720
rect 673514 463664 673519 463720
rect 673269 463662 673519 463664
rect 673269 463659 673335 463662
rect 673453 463659 673519 463662
rect 673453 463586 673519 463589
rect 673729 463586 673795 463589
rect 673453 463584 673795 463586
rect 673453 463528 673458 463584
rect 673514 463528 673734 463584
rect 673790 463528 673795 463584
rect 673453 463526 673795 463528
rect 673453 463523 673519 463526
rect 673729 463523 673795 463526
rect 39941 455426 40007 455429
rect 40166 455426 40172 455428
rect 39941 455424 40172 455426
rect 39941 455368 39946 455424
rect 40002 455368 40172 455424
rect 39941 455366 40172 455368
rect 39941 455363 40007 455366
rect 40166 455364 40172 455366
rect 40236 455364 40242 455428
rect 39665 451890 39731 451893
rect 40166 451890 40172 451892
rect 39665 451888 40172 451890
rect 39665 451832 39670 451888
rect 39726 451832 40172 451888
rect 39665 451830 40172 451832
rect 39665 451827 39731 451830
rect 40166 451828 40172 451830
rect 40236 451828 40242 451892
rect 44357 448626 44423 448629
rect 39468 448624 44423 448626
rect 39468 448596 44362 448624
rect 39438 448568 44362 448596
rect 44418 448568 44423 448624
rect 39438 448566 44423 448568
rect 39438 446012 39498 448566
rect 44357 448563 44423 448566
rect 673545 444410 673611 444413
rect 673729 444410 673795 444413
rect 673545 444408 673795 444410
rect 673545 444352 673550 444408
rect 673606 444352 673734 444408
rect 673790 444352 673795 444408
rect 673545 444350 673795 444352
rect 673545 444347 673611 444350
rect 673729 444347 673795 444350
rect 39665 441010 39731 441013
rect 39468 441008 39731 441010
rect 39468 440952 39670 441008
rect 39726 440952 39731 441008
rect 39468 440950 39731 440952
rect 39665 440947 39731 440950
rect 673085 427954 673151 427957
rect 677409 427954 677475 427957
rect 673085 427952 677475 427954
rect 673085 427896 673090 427952
rect 673146 427896 677414 427952
rect 677470 427896 677475 427952
rect 673085 427894 677475 427896
rect 673085 427891 673151 427894
rect 677409 427891 677475 427894
rect 677593 425778 677659 425781
rect 677593 425776 677764 425778
rect 677593 425720 677598 425776
rect 677654 425720 677764 425776
rect 677593 425718 677764 425720
rect 677593 425715 677659 425718
rect 673361 420882 673427 420885
rect 673361 420880 677764 420882
rect 673361 420824 673366 420880
rect 673422 420824 677764 420880
rect 673361 420822 677764 420824
rect 673361 420819 673427 420822
rect 42241 400210 42307 400213
rect 42609 400210 42675 400213
rect 42241 400208 42675 400210
rect 42241 400152 42246 400208
rect 42302 400152 42614 400208
rect 42670 400152 42675 400208
rect 42241 400150 42675 400152
rect 42241 400147 42307 400150
rect 42609 400147 42675 400150
rect 673545 338738 673611 338741
rect 675385 338738 675451 338741
rect 673545 338736 675451 338738
rect 673545 338680 673550 338736
rect 673606 338680 675390 338736
rect 675446 338680 675451 338736
rect 673545 338678 675451 338680
rect 673545 338675 673611 338678
rect 675385 338675 675451 338678
rect 672533 314802 672599 314805
rect 672533 314800 672642 314802
rect 672533 314744 672538 314800
rect 672594 314744 672642 314800
rect 672533 314739 672642 314744
rect 672582 314533 672642 314739
rect 672533 314528 672642 314533
rect 672533 314472 672538 314528
rect 672594 314472 672642 314528
rect 672533 314470 672642 314472
rect 672533 314467 672599 314470
rect 675017 293042 675083 293045
rect 675201 293042 675267 293045
rect 675385 293042 675451 293045
rect 675017 293040 675451 293042
rect 675017 292984 675022 293040
rect 675078 292984 675206 293040
rect 675262 292984 675390 293040
rect 675446 292984 675451 293040
rect 675017 292982 675451 292984
rect 675017 292979 675083 292982
rect 675201 292979 675267 292982
rect 675385 292979 675451 292982
rect 672533 231842 672599 231845
rect 672901 231842 672967 231845
rect 672533 231840 672967 231842
rect 672533 231784 672538 231840
rect 672594 231784 672906 231840
rect 672962 231784 672967 231840
rect 672533 231782 672967 231784
rect 672533 231779 672599 231782
rect 672901 231779 672967 231782
rect 44449 193218 44515 193221
rect 44633 193218 44699 193221
rect 44449 193216 44699 193218
rect 44449 193160 44454 193216
rect 44510 193160 44638 193216
rect 44694 193160 44699 193216
rect 44449 193158 44699 193160
rect 44449 193155 44515 193158
rect 44633 193155 44699 193158
rect 672533 193218 672599 193221
rect 672901 193218 672967 193221
rect 672533 193216 672967 193218
rect 672533 193160 672538 193216
rect 672594 193160 672906 193216
rect 672962 193160 672967 193216
rect 672533 193158 672967 193160
rect 672533 193155 672599 193158
rect 672901 193155 672967 193158
rect 673729 192402 673795 192405
rect 675385 192402 675451 192405
rect 673729 192400 675451 192402
rect 673729 192344 673734 192400
rect 673790 192344 675390 192400
rect 675446 192344 675451 192400
rect 673729 192342 675451 192344
rect 673729 192339 673795 192342
rect 675385 192339 675451 192342
rect 39757 120186 39823 120189
rect 44173 120186 44239 120189
rect 39757 120184 44239 120186
rect 39757 120128 39762 120184
rect 39818 120128 44178 120184
rect 44234 120128 44239 120184
rect 39757 120126 44239 120128
rect 39757 120123 39823 120126
rect 44173 120123 44239 120126
rect 41413 115970 41479 115973
rect 42333 115970 42399 115973
rect 39806 115968 42399 115970
rect 39806 115912 41418 115968
rect 41474 115912 42338 115968
rect 42394 115912 42399 115968
rect 39806 115910 42399 115912
rect 39806 115562 39866 115910
rect 41413 115907 41479 115910
rect 42333 115907 42399 115910
rect 39622 115502 39866 115562
rect 39622 115396 39682 115502
rect 44173 110530 44239 110533
rect 45461 110530 45527 110533
rect 39652 110528 45527 110530
rect 39652 110472 44178 110528
rect 44234 110472 45466 110528
rect 45522 110472 45527 110528
rect 39652 110470 45527 110472
rect 44173 110467 44239 110470
rect 45461 110467 45527 110470
rect 39389 84282 39455 84285
rect 40166 84282 40172 84284
rect 39389 84280 40172 84282
rect 39389 84224 39394 84280
rect 39450 84224 40172 84280
rect 39389 84222 40172 84224
rect 39389 84219 39455 84222
rect 40166 84220 40172 84222
rect 40236 84220 40242 84284
rect 44265 75850 44331 75853
rect 39438 75848 44331 75850
rect 39438 75792 44270 75848
rect 44326 75792 44331 75848
rect 39438 75790 44331 75792
rect 39438 75684 39498 75790
rect 44265 75787 44331 75790
rect 44265 73266 44331 73269
rect 39468 73264 44331 73266
rect 39468 73208 44270 73264
rect 44326 73208 44331 73264
rect 39468 73206 44331 73208
rect 44265 73203 44331 73206
rect 44265 68234 44331 68237
rect 45553 68234 45619 68237
rect 39468 68232 45619 68234
rect 39468 68176 44270 68232
rect 44326 68176 45558 68232
rect 45614 68176 45619 68232
rect 39468 68174 45619 68176
rect 44265 68171 44331 68174
rect 45553 68171 45619 68174
rect 212533 47698 212599 47701
rect 231577 47698 231643 47701
rect 212533 47696 231643 47698
rect 212533 47640 212538 47696
rect 212594 47640 231582 47696
rect 231638 47640 231643 47696
rect 212533 47638 231643 47640
rect 212533 47635 212599 47638
rect 231577 47635 231643 47638
rect 270493 47698 270559 47701
rect 289629 47698 289695 47701
rect 270493 47696 289695 47698
rect 270493 47640 270498 47696
rect 270554 47640 289634 47696
rect 289690 47640 289695 47696
rect 270493 47638 289695 47640
rect 270493 47635 270559 47638
rect 289629 47635 289695 47638
rect 154573 47154 154639 47157
rect 173801 47154 173867 47157
rect 154573 47152 173867 47154
rect 154573 47096 154578 47152
rect 154634 47096 173806 47152
rect 173862 47096 173867 47152
rect 154573 47094 173867 47096
rect 154573 47091 154639 47094
rect 173801 47091 173867 47094
rect 622945 40490 623011 40493
rect 84334 40488 623011 40490
rect 84334 40432 622950 40488
rect 623006 40432 623011 40488
rect 84334 40430 623011 40432
rect 84334 40218 84394 40430
rect 622945 40427 623011 40430
rect 149053 40354 149119 40357
rect 145838 40352 149119 40354
rect 145838 40296 149058 40352
rect 149114 40296 149119 40352
rect 145838 40294 149119 40296
rect 84150 40158 84394 40218
rect 86309 40218 86375 40221
rect 86309 40216 86602 40218
rect 86309 40160 86314 40216
rect 86370 40160 86602 40216
rect 86309 40158 86602 40160
rect 84150 39644 84210 40158
rect 86309 40155 86375 40158
rect 86542 39810 86602 40158
rect 86542 39750 88994 39810
rect 86542 39644 86602 39750
rect 88934 39644 88994 39750
rect 141667 38031 141813 39999
rect 145838 39967 145898 40294
rect 149053 40291 149119 40294
rect 569217 40218 569283 40221
rect 579153 40218 579219 40221
rect 569174 40216 579219 40218
rect 569174 40160 569222 40216
rect 569278 40160 579158 40216
rect 579214 40160 579219 40216
rect 569174 40158 579219 40160
rect 569174 40155 569283 40158
rect 579153 40155 579219 40158
rect 632973 40218 633039 40221
rect 634813 40218 634879 40221
rect 632973 40216 634879 40218
rect 632973 40160 632978 40216
rect 633034 40160 634818 40216
rect 634874 40160 634879 40216
rect 632973 40158 634879 40160
rect 632973 40155 633039 40158
rect 634813 40155 634879 40158
rect 240133 39946 240199 39949
rect 253933 39946 253999 39949
rect 240133 39944 246498 39946
rect 240133 39888 240138 39944
rect 240194 39888 246498 39944
rect 240133 39886 246498 39888
rect 240133 39883 240199 39886
rect 241237 39810 241303 39813
rect 242893 39810 242959 39813
rect 241156 39808 242959 39810
rect 241156 39752 241242 39808
rect 241298 39752 242898 39808
rect 242954 39752 242959 39808
rect 241156 39750 242959 39752
rect 241237 39747 241346 39750
rect 242893 39747 242959 39750
rect 241286 39372 241346 39747
rect 246438 39538 246498 39886
rect 248830 39944 253999 39946
rect 248830 39888 253938 39944
rect 253994 39888 253999 39944
rect 248830 39886 253999 39888
rect 248830 39538 248890 39886
rect 253933 39883 253999 39886
rect 569174 39644 569234 40155
rect 622945 39674 623011 39677
rect 622945 39672 623116 39674
rect 622945 39616 622950 39672
rect 623006 39616 623116 39672
rect 622945 39614 623116 39616
rect 622945 39611 623011 39614
rect 246438 39478 248890 39538
rect 246438 39372 246498 39478
rect 248830 39372 248890 39478
<< via3 >>
rect 676260 990116 676324 990180
rect 677548 918580 677612 918644
rect 40540 908108 40604 908172
rect 40540 907972 40604 908036
rect 676260 907700 676324 907764
rect 40356 888796 40420 888860
rect 39988 855748 40052 855812
rect 39804 855476 39868 855540
rect 39804 837584 39868 837588
rect 39804 837528 39854 837584
rect 39854 837528 39868 837584
rect 39804 837524 39868 837528
rect 39988 832628 40052 832692
rect 40356 797676 40420 797740
rect 40356 797540 40420 797604
rect 40356 792100 40420 792164
rect 40540 792100 40604 792164
rect 40540 778500 40604 778564
rect 40356 778228 40420 778292
rect 40356 763132 40420 763196
rect 40724 763132 40788 763196
rect 40356 753476 40420 753540
rect 40724 753476 40788 753540
rect 40356 750620 40420 750684
rect 40356 750348 40420 750412
rect 40172 731308 40236 731372
rect 40724 731172 40788 731236
rect 40356 712268 40420 712332
rect 40724 712268 40788 712332
rect 40356 702068 40420 702132
rect 40908 702068 40972 702132
rect 40540 695268 40604 695332
rect 40908 695268 40972 695332
rect 40172 673372 40236 673436
rect 40540 673372 40604 673436
rect 40540 654332 40604 654396
rect 40172 654196 40236 654260
rect 40356 634748 40420 634812
rect 40908 634748 40972 634812
rect 40540 598980 40604 599044
rect 40908 598980 40972 599044
rect 40172 565932 40236 565996
rect 40172 565660 40236 565724
rect 40172 550564 40236 550628
rect 40540 550564 40604 550628
rect 40540 540908 40604 540972
rect 40908 540908 40972 540972
rect 40908 521868 40972 521932
rect 40172 521732 40236 521796
rect 40172 507996 40236 508060
rect 39988 507724 40052 507788
rect 677548 477532 677612 477596
rect 40172 455364 40236 455428
rect 40172 451828 40236 451892
rect 40172 84220 40236 84284
<< metal4 >>
rect 676259 990180 676325 990181
rect 676259 990116 676260 990180
rect 676324 990116 676325 990180
rect 676259 990115 676325 990116
rect 40539 908172 40605 908173
rect 40539 908108 40540 908172
rect 40604 908108 40605 908172
rect 40539 908107 40605 908108
rect 40542 908037 40602 908107
rect 40539 908036 40605 908037
rect 40539 907972 40540 908036
rect 40604 907972 40605 908036
rect 40539 907971 40605 907972
rect 676262 907765 676322 990115
rect 677547 918644 677613 918645
rect 677547 918580 677548 918644
rect 677612 918580 677613 918644
rect 677547 918579 677613 918580
rect 676259 907764 676325 907765
rect 676259 907700 676260 907764
rect 676324 907700 676325 907764
rect 676259 907699 676325 907700
rect 40355 888860 40421 888861
rect 40355 888796 40356 888860
rect 40420 888796 40421 888860
rect 40355 888795 40421 888796
rect 40358 874850 40418 888795
rect 39990 874790 40418 874850
rect 39990 855813 40050 874790
rect 39987 855812 40053 855813
rect 39987 855748 39988 855812
rect 40052 855748 40053 855812
rect 39987 855747 40053 855748
rect 39803 855540 39869 855541
rect 39803 855476 39804 855540
rect 39868 855476 39869 855540
rect 39803 855475 39869 855476
rect 39806 837589 39866 855475
rect 39803 837588 39869 837589
rect 39803 837524 39804 837588
rect 39868 837524 39869 837588
rect 39803 837523 39869 837524
rect 39987 832692 40053 832693
rect 39987 832628 39988 832692
rect 40052 832628 40053 832692
rect 39987 832627 40053 832628
rect 39990 817050 40050 832627
rect 39990 816990 40418 817050
rect 40358 797741 40418 816990
rect 40355 797740 40421 797741
rect 40355 797676 40356 797740
rect 40420 797676 40421 797740
rect 40355 797675 40421 797676
rect 40355 797604 40421 797605
rect 40355 797540 40356 797604
rect 40420 797540 40421 797604
rect 40355 797539 40421 797540
rect 40358 792165 40418 797539
rect 40355 792164 40421 792165
rect 40355 792100 40356 792164
rect 40420 792100 40421 792164
rect 40355 792099 40421 792100
rect 40539 792164 40605 792165
rect 40539 792100 40540 792164
rect 40604 792100 40605 792164
rect 40539 792099 40605 792100
rect 40542 778565 40602 792099
rect 40539 778564 40605 778565
rect 40539 778500 40540 778564
rect 40604 778500 40605 778564
rect 40539 778499 40605 778500
rect 40355 778292 40421 778293
rect 40355 778228 40356 778292
rect 40420 778228 40421 778292
rect 40355 778227 40421 778228
rect 40358 763197 40418 778227
rect 40355 763196 40421 763197
rect 40355 763132 40356 763196
rect 40420 763132 40421 763196
rect 40355 763131 40421 763132
rect 40723 763196 40789 763197
rect 40723 763132 40724 763196
rect 40788 763132 40789 763196
rect 40723 763131 40789 763132
rect 40726 753541 40786 763131
rect 40355 753540 40421 753541
rect 40355 753476 40356 753540
rect 40420 753476 40421 753540
rect 40355 753475 40421 753476
rect 40723 753540 40789 753541
rect 40723 753476 40724 753540
rect 40788 753476 40789 753540
rect 40723 753475 40789 753476
rect 40358 750685 40418 753475
rect 40355 750684 40421 750685
rect 40355 750620 40356 750684
rect 40420 750620 40421 750684
rect 40355 750619 40421 750620
rect 40355 750412 40421 750413
rect 40355 750410 40356 750412
rect 40174 750350 40356 750410
rect 40174 731373 40234 750350
rect 40355 750348 40356 750350
rect 40420 750348 40421 750412
rect 40355 750347 40421 750348
rect 40171 731372 40237 731373
rect 40171 731308 40172 731372
rect 40236 731308 40237 731372
rect 40171 731307 40237 731308
rect 40723 731236 40789 731237
rect 40723 731172 40724 731236
rect 40788 731172 40789 731236
rect 40723 731171 40789 731172
rect 40726 712333 40786 731171
rect 40355 712332 40421 712333
rect 40355 712330 40356 712332
rect 40174 712270 40356 712330
rect 40174 702130 40234 712270
rect 40355 712268 40356 712270
rect 40420 712268 40421 712332
rect 40355 712267 40421 712268
rect 40723 712332 40789 712333
rect 40723 712268 40724 712332
rect 40788 712268 40789 712332
rect 40723 712267 40789 712268
rect 40355 702132 40421 702133
rect 40355 702130 40356 702132
rect 40174 702070 40356 702130
rect 40355 702068 40356 702070
rect 40420 702068 40421 702132
rect 40355 702067 40421 702068
rect 40907 702132 40973 702133
rect 40907 702068 40908 702132
rect 40972 702068 40973 702132
rect 40907 702067 40973 702068
rect 40910 695333 40970 702067
rect 40539 695332 40605 695333
rect 40539 695268 40540 695332
rect 40604 695268 40605 695332
rect 40539 695267 40605 695268
rect 40907 695332 40973 695333
rect 40907 695268 40908 695332
rect 40972 695268 40973 695332
rect 40907 695267 40973 695268
rect 40542 676290 40602 695267
rect 40174 676230 40602 676290
rect 40174 673437 40234 676230
rect 40171 673436 40237 673437
rect 40171 673372 40172 673436
rect 40236 673372 40237 673436
rect 40171 673371 40237 673372
rect 40539 673436 40605 673437
rect 40539 673372 40540 673436
rect 40604 673372 40605 673436
rect 40539 673371 40605 673372
rect 40542 654397 40602 673371
rect 40539 654396 40605 654397
rect 40539 654332 40540 654396
rect 40604 654332 40605 654396
rect 40539 654331 40605 654332
rect 40171 654260 40237 654261
rect 40171 654196 40172 654260
rect 40236 654196 40237 654260
rect 40171 654195 40237 654196
rect 40174 642970 40234 654195
rect 39990 642910 40234 642970
rect 39990 637530 40050 642910
rect 39990 637470 40418 637530
rect 40358 634813 40418 637470
rect 40355 634812 40421 634813
rect 40355 634748 40356 634812
rect 40420 634748 40421 634812
rect 40355 634747 40421 634748
rect 40907 634812 40973 634813
rect 40907 634748 40908 634812
rect 40972 634748 40973 634812
rect 40907 634747 40973 634748
rect 40910 599045 40970 634747
rect 40539 599044 40605 599045
rect 40539 598980 40540 599044
rect 40604 598980 40605 599044
rect 40539 598979 40605 598980
rect 40907 599044 40973 599045
rect 40907 598980 40908 599044
rect 40972 598980 40973 599044
rect 40907 598979 40973 598980
rect 40542 585170 40602 598979
rect 40174 585110 40602 585170
rect 40174 565997 40234 585110
rect 40171 565996 40237 565997
rect 40171 565932 40172 565996
rect 40236 565932 40237 565996
rect 40171 565931 40237 565932
rect 40171 565724 40237 565725
rect 40171 565660 40172 565724
rect 40236 565660 40237 565724
rect 40171 565659 40237 565660
rect 40174 550629 40234 565659
rect 40171 550628 40237 550629
rect 40171 550564 40172 550628
rect 40236 550564 40237 550628
rect 40171 550563 40237 550564
rect 40539 550628 40605 550629
rect 40539 550564 40540 550628
rect 40604 550564 40605 550628
rect 40539 550563 40605 550564
rect 40542 540973 40602 550563
rect 40539 540972 40605 540973
rect 40539 540908 40540 540972
rect 40604 540908 40605 540972
rect 40539 540907 40605 540908
rect 40907 540972 40973 540973
rect 40907 540908 40908 540972
rect 40972 540908 40973 540972
rect 40907 540907 40973 540908
rect 40910 521933 40970 540907
rect 40907 521932 40973 521933
rect 40907 521868 40908 521932
rect 40972 521868 40973 521932
rect 40907 521867 40973 521868
rect 40171 521796 40237 521797
rect 40171 521732 40172 521796
rect 40236 521732 40237 521796
rect 40171 521731 40237 521732
rect 40174 508061 40234 521731
rect 40171 508060 40237 508061
rect 40171 507996 40172 508060
rect 40236 507996 40237 508060
rect 40171 507995 40237 507996
rect 39987 507788 40053 507789
rect 39987 507724 39988 507788
rect 40052 507724 40053 507788
rect 39987 507723 40053 507724
rect 39990 488610 40050 507723
rect 39990 488550 40234 488610
rect 40174 455429 40234 488550
rect 677550 477597 677610 918579
rect 677547 477596 677613 477597
rect 677547 477532 677548 477596
rect 677612 477532 677613 477596
rect 677547 477531 677613 477532
rect 40171 455428 40237 455429
rect 40171 455364 40172 455428
rect 40236 455364 40237 455428
rect 40171 455363 40237 455364
rect 40171 451892 40237 451893
rect 40171 451828 40172 451892
rect 40236 451828 40237 451892
rect 40171 451827 40237 451828
rect 40174 84285 40234 451827
rect 40171 84284 40237 84285
rect 40171 84220 40172 84284
rect 40236 84220 40237 84284
rect 40171 84219 40237 84220
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334620 1018402 347160 1030924
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 576820 1018402 589360 1030924
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6086 913863 19572 925191
rect 698028 909409 711514 920737
rect 698512 863640 711002 876160
rect 6675 828820 19197 841360
rect 698402 819640 710924 832180
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 6675 484220 19197 496760
rect 698028 461609 711514 472937
rect 6086 442663 19572 453991
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6675 111420 19197 123960
rect 698512 101240 711002 113760
rect 6086 69863 19572 81191
rect 80040 6675 92580 19197
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243009 6086 254337 19572
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 624040 6675 636580 19197
use sky130_ef_io__corner_pad  user1_corner
timestamp 1606789654
transform 1 0 677600 0 1 996800
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_173
timestamp 1606789654
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1606789654
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_175
timestamp 1606789654
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_176
timestamp 1606789654
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_816
timestamp 1606789654
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_817
timestamp 1606789654
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_818
timestamp 1606789654
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_811
timestamp 1606789654
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_812
timestamp 1606789654
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_813
timestamp 1606789654
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_814
timestamp 1606789654
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_815
timestamp 1606789654
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1606789654
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_165
timestamp 1606789654
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_166
timestamp 1606789654
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_167
timestamp 1606789654
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_168
timestamp 1606789654
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_169
timestamp 1606789654
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1606789654
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_171
timestamp 1606789654
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_172
timestamp 1606789654
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[15\]
timestamp 1606789654
transform 1 0 626000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_160
timestamp 1606789654
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_161
timestamp 1606789654
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_162
timestamp 1606789654
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_156
timestamp 1606789654
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1606789654
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1606789654
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_159
timestamp 1606789654
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_152
timestamp 1606789654
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_153
timestamp 1606789654
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_154
timestamp 1606789654
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_155
timestamp 1606789654
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1606789654
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1606789654
transform 1 0 575600 0 1 998007
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1606789654
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1606789654
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_146
timestamp 1606789654
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_147
timestamp 1606789654
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_148
timestamp 1606789654
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_149
timestamp 1606789654
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_141
timestamp 1606789654
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_142
timestamp 1606789654
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_143
timestamp 1606789654
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1606789654
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_139
timestamp 1606789654
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_140
timestamp 1606789654
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[16\]
timestamp 1606789654
transform 1 0 524200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_134
timestamp 1606789654
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_135
timestamp 1606789654
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_136
timestamp 1606789654
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_130
timestamp 1606789654
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1606789654
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1606789654
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_133
timestamp 1606789654
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_127
timestamp 1606789654
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_128
timestamp 1606789654
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_129
timestamp 1606789654
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1606789654
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_126
timestamp 1606789654
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[17\]
timestamp 1606789654
transform 1 0 472800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1606789654
transform 1 0 465200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_119
timestamp 1606789654
transform 1 0 469200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_120
timestamp 1606789654
transform 1 0 471200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_121
timestamp 1606789654
transform 1 0 472200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_122
timestamp 1606789654
transform 1 0 472400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_123
timestamp 1606789654
transform 1 0 472600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_117
timestamp 1606789654
transform 1 0 461200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_116
timestamp 1606789654
transform 1 0 457200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1606789654
transform 1 0 453200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1606789654
transform 1 0 449200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1606789654
transform 1 0 445200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1606789654
transform 1 0 441200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_107
timestamp 1606789654
transform 1 0 434800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_108
timestamp 1606789654
transform 1 0 435000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0
timestamp 1606789654
transform 1 0 435200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_0
timestamp 1606789654
transform 1 0 436200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1606789654
transform 1 0 437200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_105
timestamp 1606789654
transform 1 0 431800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_106
timestamp 1606789654
transform 1 0 433800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1606789654
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1606789654
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1606789654
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1606789654
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_97
timestamp 1606789654
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1606789654
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1606789654
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1606789654
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[0\]
timestamp 1606789654
transform 1 0 383800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_92
timestamp 1606789654
transform 1 0 380400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_93
timestamp 1606789654
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_94
timestamp 1606789654
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1606789654
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_84
timestamp 1606789654
transform 1 0 348400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_85
timestamp 1606789654
transform 1 0 352400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1606789654
transform 1 0 356400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1606789654
transform 1 0 360400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1606789654
transform 1 0 364400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1606789654
transform 1 0 368400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1606789654
transform 1 0 372400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1606789654
transform 1 0 376400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[0\]
timestamp 1606789654
transform 1 0 333400 0 1 998007
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1606789654
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1606789654
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1606789654
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1606789654
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1606789654
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1606789654
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1606789654
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1606789654
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1606789654
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1606789654
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1606789654
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1606789654
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[1\]
timestamp 1606789654
transform 1 0 282000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1606789654
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1606789654
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1606789654
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1606789654
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1606789654
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1606789654
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1606789654
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1606789654
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1606789654
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1606789654
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1606789654
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1606789654
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1606789654
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[2\]
timestamp 1606789654
transform 1 0 230400 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1606789654
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1606789654
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1606789654
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1606789654
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1606789654
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1606789654
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1606789654
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1606789654
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1606789654
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1606789654
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1606789654
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1606789654
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[3\]
timestamp 1606789654
transform 1 0 179000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1606789654
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1606789654
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1606789654
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1606789654
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1606789654
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1606789654
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1606789654
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1606789654
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1606789654
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1606789654
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1606789654
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1606789654
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[4\]
timestamp 1606789654
transform 1 0 127600 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1606789654
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1606789654
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1606789654
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1606789654
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1606789654
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1606789654
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1606789654
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1606789654
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1606789654
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1606789654
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1606789654
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1606789654
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[5\]
timestamp 1606789654
transform 1 0 76200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_14
timestamp 1606789654
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15
timestamp 1606789654
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1606789654
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1606789654
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1606789654
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1606789654
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13
timestamp 1606789654
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1606789654
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1606789654
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1606789654
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1606789654
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1606789654
transform 0 -1 40800 1 0 997600
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_5
timestamp 1606789654
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_608
timestamp 1606789654
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_609
timestamp 1606789654
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_610
timestamp 1606789654
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_611
timestamp 1606789654
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_603
timestamp 1606789654
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_604
timestamp 1606789654
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1606789654
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1606789654
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1606789654
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[14\]
timestamp 1606789654
transform 0 1 675407 -1 0 967600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1606789654
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1606789654
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1606789654
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1606789654
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1606789654
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_808
timestamp 1606789654
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_810
timestamp 1606789654
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_602
timestamp 1606789654
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[6\]
timestamp 1606789654
transform 0 -1 42193 1 0 954200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1606789654
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_598
timestamp 1606789654
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_599
timestamp 1606789654
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_600
timestamp 1606789654
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_593
timestamp 1606789654
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_594
timestamp 1606789654
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1606789654
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1606789654
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_801
timestamp 1606789654
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_802
timestamp 1606789654
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user1_vccd_lvclamp_pad
timestamp 1606789654
transform 0 1 678007 -1 0 922600
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1606789654
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_798
timestamp 1606789654
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_799
timestamp 1606789654
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_793
timestamp 1606789654
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1606789654
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1606789654
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1606789654
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_592
timestamp 1606789654
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  user2_vccd_lvclamp_pad
timestamp 1606789654
transform 0 -1 39593 1 0 912000
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1606789654
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_588
timestamp 1606789654
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_589
timestamp 1606789654
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_590
timestamp 1606789654
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_583
timestamp 1606789654
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_584
timestamp 1606789654
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1606789654
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1606789654
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[13\]
timestamp 1606789654
transform 0 1 675407 -1 0 878400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1606789654
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1606789654
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1606789654
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1606789654
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_789
timestamp 1606789654
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_791
timestamp 1606789654
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_792
timestamp 1606789654
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_582
timestamp 1606789654
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1606789654
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1606789654
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_578
timestamp 1606789654
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_579
timestamp 1606789654
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_580
timestamp 1606789654
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_573
timestamp 1606789654
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_574
timestamp 1606789654
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1606789654
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1606789654
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1606789654
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1606789654
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1606789654
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1606789654
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_779
timestamp 1606789654
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_780
timestamp 1606789654
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_782
timestamp 1606789654
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_783
timestamp 1606789654
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1606789654
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_572
timestamp 1606789654
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user2_vssa_hvclamp_pad
timestamp 1606789654
transform 0 -1 39593 1 0 827600
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1606789654
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_568
timestamp 1606789654
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_569
timestamp 1606789654
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_570
timestamp 1606789654
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_563
timestamp 1606789654
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_564
timestamp 1606789654
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1606789654
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1606789654
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[12\]
timestamp 1606789654
transform 0 1 675407 -1 0 789200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1606789654
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1606789654
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1606789654
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_770
timestamp 1606789654
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_772
timestamp 1606789654
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_773
timestamp 1606789654
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_774
timestamp 1606789654
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1606789654
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_562
timestamp 1606789654
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[7\]
timestamp 1606789654
transform 0 -1 42193 1 0 784400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1606789654
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_558
timestamp 1606789654
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_559
timestamp 1606789654
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_560
timestamp 1606789654
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_553
timestamp 1606789654
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_554
timestamp 1606789654
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1606789654
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1606789654
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[11\]
timestamp 1606789654
transform 0 1 675407 -1 0 744200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1606789654
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1606789654
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_761
timestamp 1606789654
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_763
timestamp 1606789654
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_764
timestamp 1606789654
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1606789654
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1606789654
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_552
timestamp 1606789654
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[8\]
timestamp 1606789654
transform 0 -1 42193 1 0 741200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1606789654
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_548
timestamp 1606789654
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_549
timestamp 1606789654
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_550
timestamp 1606789654
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_543
timestamp 1606789654
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_544
timestamp 1606789654
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1606789654
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1606789654
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[10\]
timestamp 1606789654
transform 0 1 675407 -1 0 699200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1606789654
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_751
timestamp 1606789654
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_752
timestamp 1606789654
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_754
timestamp 1606789654
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_755
timestamp 1606789654
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1606789654
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1606789654
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1606789654
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[9\]
timestamp 1606789654
transform 0 -1 42193 1 0 698000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_534
timestamp 1606789654
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1606789654
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1606789654
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1606789654
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_538
timestamp 1606789654
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_539
timestamp 1606789654
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_540
timestamp 1606789654
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_542
timestamp 1606789654
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[9\]
timestamp 1606789654
transform 0 1 675407 -1 0 654000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1606789654
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_742
timestamp 1606789654
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_744
timestamp 1606789654
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_745
timestamp 1606789654
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_746
timestamp 1606789654
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1606789654
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1606789654
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1606789654
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_532
timestamp 1606789654
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_533
timestamp 1606789654
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[10\]
timestamp 1606789654
transform 0 -1 42193 1 0 654800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_528
timestamp 1606789654
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_529
timestamp 1606789654
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_530
timestamp 1606789654
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_524
timestamp 1606789654
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1606789654
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1606789654
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1606789654
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[8\]
timestamp 1606789654
transform 0 1 675407 -1 0 609000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_732
timestamp 1606789654
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_733
timestamp 1606789654
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_735
timestamp 1606789654
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_736
timestamp 1606789654
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1606789654
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1606789654
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1606789654
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1606789654
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_522
timestamp 1606789654
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_523
timestamp 1606789654
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[11\]
timestamp 1606789654
transform 0 -1 42193 1 0 611600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_518
timestamp 1606789654
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_519
timestamp 1606789654
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_520
timestamp 1606789654
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_514
timestamp 1606789654
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1606789654
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1606789654
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1606789654
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_725
timestamp 1606789654
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_726
timestamp 1606789654
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_727
timestamp 1606789654
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1606789654
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1606789654
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1606789654
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1606789654
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_512
timestamp 1606789654
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_513
timestamp 1606789654
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[12\]
timestamp 1606789654
transform 0 -1 42193 1 0 568400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_508
timestamp 1606789654
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_509
timestamp 1606789654
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_510
timestamp 1606789654
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_504
timestamp 1606789654
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1606789654
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1606789654
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1606789654
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[7\]
timestamp 1606789654
transform 0 1 675407 -1 0 563800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_716
timestamp 1606789654
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_717
timestamp 1606789654
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1606789654
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1606789654
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1606789654
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1606789654
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1606789654
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_723
timestamp 1606789654
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[13\]
timestamp 1606789654
transform 0 -1 42193 1 0 525200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1606789654
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1606789654
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1606789654
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_498
timestamp 1606789654
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_499
timestamp 1606789654
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_500
timestamp 1606789654
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_502
timestamp 1606789654
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_503
timestamp 1606789654
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1606789654
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_707
timestamp 1606789654
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_708
timestamp 1606789654
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1606789654
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1606789654
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1606789654
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1606789654
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1606789654
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_714
timestamp 1606789654
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_492
timestamp 1606789654
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_493
timestamp 1606789654
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_494
timestamp 1606789654
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  user2_vdda_hvclamp_pad
timestamp 1606789654
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_488
timestamp 1606789654
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_489
timestamp 1606789654
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_490
timestamp 1606789654
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1606789654
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1606789654
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1606789654
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user1_vssd_lvclmap_pad
timestamp 1606789654
transform 0 1 678007 -1 0 474800
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1606789654
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_704
timestamp 1606789654
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_705
timestamp 1606789654
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_699
timestamp 1606789654
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1606789654
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1606789654
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1606789654
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_697
timestamp 1606789654
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_698
timestamp 1606789654
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_482
timestamp 1606789654
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_483
timestamp 1606789654
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_484
timestamp 1606789654
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  user2_vssd_lvclmap_pad
timestamp 1606789654
transform 0 -1 39593 1 0 440800
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_478
timestamp 1606789654
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_479
timestamp 1606789654
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_480
timestamp 1606789654
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1606789654
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1606789654
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1606789654
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1606789654
transform 0 1 678007 -1 0 430600
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_688
timestamp 1606789654
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_689
timestamp 1606789654
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1606789654
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1606789654
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1606789654
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1606789654
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1606789654
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_695
timestamp 1606789654
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_472
timestamp 1606789654
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_473
timestamp 1606789654
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_474
timestamp 1606789654
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[14\]
timestamp 1606789654
transform 0 -1 42193 1 0 397600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_5um  FILLER_469
timestamp 1606789654
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_470
timestamp 1606789654
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1606789654
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1606789654
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1606789654
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_468
timestamp 1606789654
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[6\]
timestamp 1606789654
transform 0 1 675407 -1 0 386600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_686
timestamp 1606789654
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1606789654
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1606789654
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1606789654
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_685
timestamp 1606789654
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_678
timestamp 1606789654
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_679
timestamp 1606789654
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_680
timestamp 1606789654
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1606789654
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_462
timestamp 1606789654
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_463
timestamp 1606789654
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_464
timestamp 1606789654
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[15\]
timestamp 1606789654
transform 0 -1 42193 1 0 354400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_460
timestamp 1606789654
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1606789654
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1606789654
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1606789654
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_458
timestamp 1606789654
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_459
timestamp 1606789654
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[5\]
timestamp 1606789654
transform 0 1 675407 -1 0 341400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_669
timestamp 1606789654
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_670
timestamp 1606789654
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1606789654
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1606789654
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1606789654
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1606789654
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1606789654
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_676
timestamp 1606789654
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_453
timestamp 1606789654
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_454
timestamp 1606789654
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_452
timestamp 1606789654
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[16\]
timestamp 1606789654
transform 0 -1 42193 1 0 311200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1606789654
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1606789654
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1606789654
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_448
timestamp 1606789654
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_449
timestamp 1606789654
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_450
timestamp 1606789654
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[4\]
timestamp 1606789654
transform 0 1 675407 -1 0 296400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_661
timestamp 1606789654
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1606789654
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1606789654
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1606789654
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1606789654
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1606789654
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_667
timestamp 1606789654
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[17\]
timestamp 1606789654
transform 0 -1 42193 1 0 268000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1606789654
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1606789654
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_438
timestamp 1606789654
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_439
timestamp 1606789654
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_440
timestamp 1606789654
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_442
timestamp 1606789654
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_443
timestamp 1606789654
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_444
timestamp 1606789654
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[3\]
timestamp 1606789654
transform 0 1 675407 -1 0 251400
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_652
timestamp 1606789654
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1606789654
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1606789654
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1606789654
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1606789654
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_657
timestamp 1606789654
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_658
timestamp 1606789654
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_660
timestamp 1606789654
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_433
timestamp 1606789654
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_434
timestamp 1606789654
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1606789654
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_432
timestamp 1606789654
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[18\]
timestamp 1606789654
transform 0 -1 42193 1 0 224800
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1606789654
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1606789654
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_428
timestamp 1606789654
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_429
timestamp 1606789654
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_430
timestamp 1606789654
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[2\]
timestamp 1606789654
transform 0 1 675407 -1 0 206200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1606789654
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1606789654
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1606789654
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1606789654
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1606789654
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_648
timestamp 1606789654
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_650
timestamp 1606789654
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_651
timestamp 1606789654
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_423
timestamp 1606789654
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_424
timestamp 1606789654
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1606789654
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_422
timestamp 1606789654
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area2_io_pad\[19\]
timestamp 1606789654
transform 0 -1 42193 1 0 181600
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1606789654
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1606789654
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_418
timestamp 1606789654
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_419
timestamp 1606789654
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_420
timestamp 1606789654
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[1\]
timestamp 1606789654
transform 0 1 675407 -1 0 161200
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1606789654
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1606789654
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1606789654
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1606789654
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_638
timestamp 1606789654
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_639
timestamp 1606789654
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_641
timestamp 1606789654
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_642
timestamp 1606789654
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1606789654
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_414
timestamp 1606789654
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_413
timestamp 1606789654
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_408
timestamp 1606789654
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_409
timestamp 1606789654
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1606789654
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_2
timestamp 1606789654
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_412
timestamp 1606789654
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_407
timestamp 1606789654
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1606789654
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1606789654
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_404
timestamp 1606789654
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_403
timestamp 1606789654
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_402
timestamp 1606789654
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  mprj_pads.area1_io_pad\[0\]
timestamp 1606789654
transform 0 1 675407 -1 0 116000
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1606789654
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1606789654
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1606789654
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_629
timestamp 1606789654
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_631
timestamp 1606789654
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_632
timestamp 1606789654
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_633
timestamp 1606789654
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_401
timestamp 1606789654
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__vddio_hvc_pad  mgmt_vddio_hvclamp_pad\[0\]
timestamp 1606789654
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1606789654
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_397
timestamp 1606789654
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_398
timestamp 1606789654
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_399
timestamp 1606789654
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_392
timestamp 1606789654
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_393
timestamp 1606789654
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1606789654
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1606789654
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1606789654
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1606789654
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_623
timestamp 1606789654
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_622
timestamp 1606789654
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_619
timestamp 1606789654
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1
timestamp 1606789654
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vccd_slice_5um  disconnect_vccd_1
timestamp 1606789654
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1606789654
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1606789654
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1606789654
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1606789654
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_614
timestamp 1606789654
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_613
timestamp 1606789654
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_391
timestamp 1606789654
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__vccd_lvc_pad  mgmt_vccd_lvclamp_pad
timestamp 1606789654
transform 0 -1 39593 1 0 68000
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1606789654
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_387
timestamp 1606789654
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_388
timestamp 1606789654
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_389
timestamp 1606789654
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_382
timestamp 1606789654
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_383
timestamp 1606789654
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1606789654
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1606789654
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[1\]
timestamp 1606789654
transform 0 1 676800 -1 0 40000
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_5um  FILLER_377
timestamp 1606789654
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_378
timestamp 1606789654
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_379
timestamp 1606789654
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_380
timestamp 1606789654
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_612
timestamp 1606789654
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_376
timestamp 1606789654
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1606789654
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1606789654
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1606789654
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1606789654
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1606789654
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1606789654
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_368
timestamp 1606789654
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1606789654
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_365
timestamp 1606789654
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_366
timestamp 1606789654
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_367
timestamp 1606789654
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_364
timestamp 1606789654
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vdda_hvc_pad  mgmt_vdda_hvclamp_pad
timestamp 1606789654
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_360
timestamp 1606789654
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1606789654
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_362
timestamp 1606789654
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1606789654
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1606789654
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_358
timestamp 1606789654
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_359
timestamp 1606789654
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_350
timestamp 1606789654
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_351
timestamp 1606789654
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1606789654
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1606789654
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1606789654
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1606789654
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_347
timestamp 1606789654
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_348
timestamp 1606789654
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_349
timestamp 1606789654
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__vssio_hvc_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1606789654
transform -1 0 584000 0 -1 39593
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_342
timestamp 1606789654
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_343
timestamp 1606789654
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1606789654
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_345
timestamp 1606789654
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1606789654
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1606789654
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1606789654
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_341
timestamp 1606789654
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1606789654
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1606789654
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_330
timestamp 1606789654
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_331
timestamp 1606789654
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_332
timestamp 1606789654
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_333
timestamp 1606789654
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_334
timestamp 1606789654
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1606789654
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  gpio_pad
timestamp 1606789654
transform -1 0 530200 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_324
timestamp 1606789654
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_325
timestamp 1606789654
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_326
timestamp 1606789654
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1606789654
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_328
timestamp 1606789654
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1606789654
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1606789654
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1606789654
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1606789654
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1606789654
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_315
timestamp 1606789654
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_316
timestamp 1606789654
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_317
timestamp 1606789654
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1606789654
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_314
timestamp 1606789654
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_313
timestamp 1606789654
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io1_pad
timestamp 1606789654
transform -1 0 475400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_10um  FILLER_308
timestamp 1606789654
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_309
timestamp 1606789654
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1606789654
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_311
timestamp 1606789654
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1606789654
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1606789654
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1606789654
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_307
timestamp 1606789654
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_297
timestamp 1606789654
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_298
timestamp 1606789654
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_299
timestamp 1606789654
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_300
timestamp 1606789654
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1606789654
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1606789654
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1606789654
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_296
timestamp 1606789654
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_io0_pad
timestamp 1606789654
transform -1 0 420600 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_290
timestamp 1606789654
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_291
timestamp 1606789654
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_292
timestamp 1606789654
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1606789654
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_294
timestamp 1606789654
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1606789654
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1606789654
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1606789654
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1606789654
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_281
timestamp 1606789654
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_282
timestamp 1606789654
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_283
timestamp 1606789654
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1606789654
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1606789654
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_279
timestamp 1606789654
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_280
timestamp 1606789654
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_clk_pad
timestamp 1606789654
transform -1 0 365800 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1606789654
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_273
timestamp 1606789654
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_274
timestamp 1606789654
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_275
timestamp 1606789654
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1606789654
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_277
timestamp 1606789654
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1606789654
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1606789654
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1606789654
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1606789654
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_264
timestamp 1606789654
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_265
timestamp 1606789654
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_266
timestamp 1606789654
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1606789654
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_263
timestamp 1606789654
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_262
timestamp 1606789654
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  flash_csb_pad
timestamp 1606789654
transform -1 0 311000 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_20um  FILLER_256
timestamp 1606789654
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_257
timestamp 1606789654
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_258
timestamp 1606789654
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1606789654
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_260
timestamp 1606789654
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1606789654
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1606789654
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1606789654
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1606789654
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_245
timestamp 1606789654
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_246
timestamp 1606789654
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_247
timestamp 1606789654
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_248
timestamp 1606789654
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_249
timestamp 1606789654
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1606789654
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1606789654
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssd_lvc_pad  mgmt_vssd_lvclmap_pad
timestamp 1606789654
transform -1 0 256200 0 -1 39593
box 0 -46 15000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_243
timestamp 1606789654
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1606789654
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_239
timestamp 1606789654
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_240
timestamp 1606789654
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_241
timestamp 1606789654
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1606789654
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1606789654
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1606789654
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1606789654
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1606789654
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_228
timestamp 1606789654
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_229
timestamp 1606789654
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_230
timestamp 1606789654
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_231
timestamp 1606789654
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_232
timestamp 1606789654
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1606789654
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__gpiov2_pad_wrapped  clock_pad
timestamp 1606789654
transform -1 0 202400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1606789654
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_226
timestamp 1606789654
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1606789654
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1606789654
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_222
timestamp 1606789654
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_223
timestamp 1606789654
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_224
timestamp 1606789654
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1606789654
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1606789654
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1606789654
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_211
timestamp 1606789654
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_212
timestamp 1606789654
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_213
timestamp 1606789654
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_214
timestamp 1606789654
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_215
timestamp 1606789654
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1606789654
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_fd_io__top_xres4v2  resetb_pad
timestamp 1606789654
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__com_bus_slice_10um  FILLER_206
timestamp 1606789654
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_207
timestamp 1606789654
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1606789654
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_209
timestamp 1606789654
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_205
timestamp 1606789654
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1606789654
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1606789654
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1606789654
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1606789654
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1606789654
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_197
timestamp 1606789654
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_198
timestamp 1606789654
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1606789654
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_195
timestamp 1606789654
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_196
timestamp 1606789654
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_194
timestamp 1606789654
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__vssa_hvc_pad  mgmt_vssa_hvclamp_pad
timestamp 1606789654
transform -1 0 93800 0 -1 39593
box 0 -434 15000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_189
timestamp 1606789654
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_190
timestamp 1606789654
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1606789654
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_192
timestamp 1606789654
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1606789654
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1606789654
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1606789654
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_188
timestamp 1606789654
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_178
timestamp 1606789654
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_179
timestamp 1606789654
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_180
timestamp 1606789654
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_181
timestamp 1606789654
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1
timestamp 1606789654
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1606789654
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3
timestamp 1606789654
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__corner_pad  mgmt_corner\[0\]
timestamp 1606789654
transform -1 0 40000 0 -1 40800
box -271 -204 40000 40800
use sky130_ef_io__com_bus_slice_20um  FILLER_177
timestamp 1606789654
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_381
timestamp 1606789654
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 4 clock
port 1 nsew
rlabel metal2 s 187327 41713 187383 42193 4 clock_core
port 2 nsew
rlabel metal2 s 194043 41713 194099 42193 4 por
port 3 nsew
rlabel metal5 s 351040 6598 363560 19088 4 flash_clk
port 4 nsew
rlabel metal2 s 361767 41713 361823 42193 4 flash_clk_core
port 5 nsew
rlabel metal2 s 357443 41713 357499 42193 4 flash_clk_ieb_core
port 6 nsew
rlabel metal2 s 364895 41713 364951 42193 4 flash_clk_oeb_core
port 7 nsew
rlabel metal5 s 296240 6598 308760 19088 4 flash_csb
port 8 nsew
rlabel metal2 s 306967 41713 307023 42193 4 flash_csb_core
port 9 nsew
rlabel metal2 s 302643 41713 302699 42193 4 flash_csb_ieb_core
port 10 nsew
rlabel metal2 s 310095 41713 310151 42193 4 flash_csb_oeb_core
port 11 nsew
rlabel metal5 s 405840 6598 418360 19088 4 flash_io0
port 12 nsew
rlabel metal2 s 405527 41713 405583 42193 4 flash_io0_di_core
port 13 nsew
rlabel metal2 s 416567 41713 416623 42193 4 flash_io0_do_core
port 14 nsew
rlabel metal2 s 412243 41713 412299 42193 4 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 419695 41713 419751 42193 4 flash_io0_oeb_core
port 16 nsew
rlabel metal5 s 460640 6598 473160 19088 4 flash_io1
port 17 nsew
rlabel metal2 s 460327 41713 460383 42193 4 flash_io1_di_core
port 18 nsew
rlabel metal2 s 471367 41713 471423 42193 4 flash_io1_do_core
port 19 nsew
rlabel metal2 s 467043 41713 467099 42193 4 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 474495 41713 474551 42193 4 flash_io1_oeb_core
port 21 nsew
rlabel metal5 s 515440 6598 527960 19088 4 gpio
port 22 nsew
rlabel metal2 s 515127 41713 515183 42193 4 gpio_in_core
port 23 nsew
rlabel metal2 s 521843 41713 521899 42193 4 gpio_inenb_core
port 24 nsew
rlabel metal2 s 520647 41713 520703 42193 4 gpio_mode0_core
port 25 nsew
rlabel metal2 s 524971 41713 525027 42193 4 gpio_mode1_core
port 26 nsew
rlabel metal2 s 526167 41713 526223 42193 4 gpio_out_core
port 27 nsew
rlabel metal2 s 529295 41713 529351 42193 4 gpio_outenb_core
port 28 nsew
rlabel metal5 s 6086 69863 19572 81191 4 vccd
port 29 nsew
rlabel metal5 s 624040 6675 636580 19197 4 vdda
port 30 nsew
rlabel metal5 s 6675 111420 19197 123960 4 vddio
port 31 nsew
rlabel metal5 s 80040 6675 92580 19197 4 vssa
port 32 nsew
rlabel metal5 s 243009 6086 254337 19572 4 vssd
port 33 nsew
rlabel metal5 s 334620 1018402 347160 1030924 4 vssio
port 34 nsew
rlabel metal5 s 698512 101240 711002 113760 4 mprj_io[0]
port 35 nsew
rlabel metal2 s 675407 105803 675887 105859 4 mprj_io_analog_en[0]
port 36 nsew
rlabel metal2 s 675407 107091 675887 107147 4 mprj_io_analog_pol[0]
port 37 nsew
rlabel metal2 s 675407 110127 675887 110183 4 mprj_io_analog_sel[0]
port 38 nsew
rlabel metal2 s 675407 106447 675887 106503 4 mprj_io_dm[0]
port 39 nsew
rlabel metal2 s 675407 104607 675887 104663 4 mprj_io_dm[1]
port 40 nsew
rlabel metal2 s 675407 110771 675887 110827 4 mprj_io_dm[2]
port 41 nsew
rlabel metal2 s 675407 108931 675887 108987 4 mprj_io_enh[0]
port 42 nsew
rlabel metal2 s 675407 109575 675887 109631 4 mprj_io_hldh_n[0]
port 43 nsew
rlabel metal2 s 675407 111415 675887 111471 4 mprj_io_holdover[0]
port 44 nsew
rlabel metal2 s 675407 114451 675887 114507 4 mprj_io_ib_mode_sel[0]
port 45 nsew
rlabel metal2 s 675407 107643 675887 107699 4 mprj_io_inp_dis[0]
port 46 nsew
rlabel metal2 s 675407 115095 675887 115151 4 mprj_io_oeb[0]
port 47 nsew
rlabel metal2 s 675407 111967 675887 112023 4 mprj_io_out[0]
port 48 nsew
rlabel metal2 s 675407 102767 675887 102823 4 mprj_io_slow_sel[0]
port 49 nsew
rlabel metal2 s 675407 113807 675887 113863 4 mprj_io_vtrip_sel[0]
port 50 nsew
rlabel metal2 s 675407 100927 675887 100983 4 mprj_io_in[0]
port 51 nsew
rlabel metal5 s 698512 684440 711002 696960 4 mprj_io[10]
port 52 nsew
rlabel metal2 s 675407 689003 675887 689059 4 mprj_io_analog_en[10]
port 53 nsew
rlabel metal2 s 675407 690291 675887 690347 4 mprj_io_analog_pol[10]
port 54 nsew
rlabel metal2 s 675407 693327 675887 693383 4 mprj_io_analog_sel[10]
port 55 nsew
rlabel metal2 s 675407 689647 675887 689703 4 mprj_io_dm[30]
port 56 nsew
rlabel metal2 s 675407 687807 675887 687863 4 mprj_io_dm[31]
port 57 nsew
rlabel metal2 s 675407 693971 675887 694027 4 mprj_io_dm[32]
port 58 nsew
rlabel metal2 s 675407 692131 675887 692187 4 mprj_io_enh[10]
port 59 nsew
rlabel metal2 s 675407 692775 675887 692831 4 mprj_io_hldh_n[10]
port 60 nsew
rlabel metal2 s 675407 694615 675887 694671 4 mprj_io_holdover[10]
port 61 nsew
rlabel metal2 s 675407 697651 675887 697707 4 mprj_io_ib_mode_sel[10]
port 62 nsew
rlabel metal2 s 675407 690843 675887 690899 4 mprj_io_inp_dis[10]
port 63 nsew
rlabel metal2 s 675407 698295 675887 698351 4 mprj_io_oeb[10]
port 64 nsew
rlabel metal2 s 675407 695167 675887 695223 4 mprj_io_out[10]
port 65 nsew
rlabel metal2 s 675407 685967 675887 686023 4 mprj_io_slow_sel[10]
port 66 nsew
rlabel metal2 s 675407 697007 675887 697063 4 mprj_io_vtrip_sel[10]
port 67 nsew
rlabel metal2 s 675407 684127 675887 684183 4 mprj_io_in[10]
port 68 nsew
rlabel metal5 s 698512 729440 711002 741960 4 mprj_io[11]
port 69 nsew
rlabel metal2 s 675407 734003 675887 734059 4 mprj_io_analog_en[11]
port 70 nsew
rlabel metal2 s 675407 735291 675887 735347 4 mprj_io_analog_pol[11]
port 71 nsew
rlabel metal2 s 675407 738327 675887 738383 4 mprj_io_analog_sel[11]
port 72 nsew
rlabel metal2 s 675407 734647 675887 734703 4 mprj_io_dm[33]
port 73 nsew
rlabel metal2 s 675407 732807 675887 732863 4 mprj_io_dm[34]
port 74 nsew
rlabel metal2 s 675407 738971 675887 739027 4 mprj_io_dm[35]
port 75 nsew
rlabel metal2 s 675407 737131 675887 737187 4 mprj_io_enh[11]
port 76 nsew
rlabel metal2 s 675407 737775 675887 737831 4 mprj_io_hldh_n[11]
port 77 nsew
rlabel metal2 s 675407 739615 675887 739671 4 mprj_io_holdover[11]
port 78 nsew
rlabel metal2 s 675407 742651 675887 742707 4 mprj_io_ib_mode_sel[11]
port 79 nsew
rlabel metal2 s 675407 735843 675887 735899 4 mprj_io_inp_dis[11]
port 80 nsew
rlabel metal2 s 675407 743295 675887 743351 4 mprj_io_oeb[11]
port 81 nsew
rlabel metal2 s 675407 740167 675887 740223 4 mprj_io_out[11]
port 82 nsew
rlabel metal2 s 675407 730967 675887 731023 4 mprj_io_slow_sel[11]
port 83 nsew
rlabel metal2 s 675407 742007 675887 742063 4 mprj_io_vtrip_sel[11]
port 84 nsew
rlabel metal2 s 675407 729127 675887 729183 4 mprj_io_in[11]
port 85 nsew
rlabel metal5 s 698512 774440 711002 786960 4 mprj_io[12]
port 86 nsew
rlabel metal2 s 675407 779003 675887 779059 4 mprj_io_analog_en[12]
port 87 nsew
rlabel metal2 s 675407 780291 675887 780347 4 mprj_io_analog_pol[12]
port 88 nsew
rlabel metal2 s 675407 783327 675887 783383 4 mprj_io_analog_sel[12]
port 89 nsew
rlabel metal2 s 675407 779647 675887 779703 4 mprj_io_dm[36]
port 90 nsew
rlabel metal2 s 675407 777807 675887 777863 4 mprj_io_dm[37]
port 91 nsew
rlabel metal2 s 675407 783971 675887 784027 4 mprj_io_dm[38]
port 92 nsew
rlabel metal2 s 675407 782131 675887 782187 4 mprj_io_enh[12]
port 93 nsew
rlabel metal2 s 675407 782775 675887 782831 4 mprj_io_hldh_n[12]
port 94 nsew
rlabel metal2 s 675407 784615 675887 784671 4 mprj_io_holdover[12]
port 95 nsew
rlabel metal2 s 675407 787651 675887 787707 4 mprj_io_ib_mode_sel[12]
port 96 nsew
rlabel metal2 s 675407 780843 675887 780899 4 mprj_io_inp_dis[12]
port 97 nsew
rlabel metal2 s 675407 788295 675887 788351 4 mprj_io_oeb[12]
port 98 nsew
rlabel metal2 s 675407 785167 675887 785223 4 mprj_io_out[12]
port 99 nsew
rlabel metal2 s 675407 775967 675887 776023 4 mprj_io_slow_sel[12]
port 100 nsew
rlabel metal2 s 675407 787007 675887 787063 4 mprj_io_vtrip_sel[12]
port 101 nsew
rlabel metal2 s 675407 774127 675887 774183 4 mprj_io_in[12]
port 102 nsew
rlabel metal5 s 698512 863640 711002 876160 4 mprj_io[13]
port 103 nsew
rlabel metal2 s 675407 868203 675887 868259 4 mprj_io_analog_en[13]
port 104 nsew
rlabel metal2 s 675407 869491 675887 869547 4 mprj_io_analog_pol[13]
port 105 nsew
rlabel metal2 s 675407 872527 675887 872583 4 mprj_io_analog_sel[13]
port 106 nsew
rlabel metal2 s 675407 868847 675887 868903 4 mprj_io_dm[39]
port 107 nsew
rlabel metal2 s 675407 867007 675887 867063 4 mprj_io_dm[40]
port 108 nsew
rlabel metal2 s 675407 873171 675887 873227 4 mprj_io_dm[41]
port 109 nsew
rlabel metal2 s 675407 871331 675887 871387 4 mprj_io_enh[13]
port 110 nsew
rlabel metal2 s 675407 871975 675887 872031 4 mprj_io_hldh_n[13]
port 111 nsew
rlabel metal2 s 675407 873815 675887 873871 4 mprj_io_holdover[13]
port 112 nsew
rlabel metal2 s 675407 876851 675887 876907 4 mprj_io_ib_mode_sel[13]
port 113 nsew
rlabel metal2 s 675407 870043 675887 870099 4 mprj_io_inp_dis[13]
port 114 nsew
rlabel metal2 s 675407 877495 675887 877551 4 mprj_io_oeb[13]
port 115 nsew
rlabel metal2 s 675407 874367 675887 874423 4 mprj_io_out[13]
port 116 nsew
rlabel metal2 s 675407 865167 675887 865223 4 mprj_io_slow_sel[13]
port 117 nsew
rlabel metal2 s 675407 876207 675887 876263 4 mprj_io_vtrip_sel[13]
port 118 nsew
rlabel metal2 s 675407 863327 675887 863383 4 mprj_io_in[13]
port 119 nsew
rlabel metal5 s 698512 952840 711002 965360 4 mprj_io[14]
port 120 nsew
rlabel metal2 s 675407 957403 675887 957459 4 mprj_io_analog_en[14]
port 121 nsew
rlabel metal2 s 675407 958691 675887 958747 4 mprj_io_analog_pol[14]
port 122 nsew
rlabel metal2 s 675407 961727 675887 961783 4 mprj_io_analog_sel[14]
port 123 nsew
rlabel metal2 s 675407 958047 675887 958103 4 mprj_io_dm[42]
port 124 nsew
rlabel metal2 s 675407 956207 675887 956263 4 mprj_io_dm[43]
port 125 nsew
rlabel metal2 s 675407 962371 675887 962427 4 mprj_io_dm[44]
port 126 nsew
rlabel metal2 s 675407 960531 675887 960587 4 mprj_io_enh[14]
port 127 nsew
rlabel metal2 s 675407 961175 675887 961231 4 mprj_io_hldh_n[14]
port 128 nsew
rlabel metal2 s 675407 963015 675887 963071 4 mprj_io_holdover[14]
port 129 nsew
rlabel metal2 s 675407 966051 675887 966107 4 mprj_io_ib_mode_sel[14]
port 130 nsew
rlabel metal2 s 675407 959243 675887 959299 4 mprj_io_inp_dis[14]
port 131 nsew
rlabel metal2 s 675407 966695 675887 966751 4 mprj_io_oeb[14]
port 132 nsew
rlabel metal2 s 675407 963567 675887 963623 4 mprj_io_out[14]
port 133 nsew
rlabel metal2 s 675407 954367 675887 954423 4 mprj_io_slow_sel[14]
port 134 nsew
rlabel metal2 s 675407 965407 675887 965463 4 mprj_io_vtrip_sel[14]
port 135 nsew
rlabel metal2 s 675407 952527 675887 952583 4 mprj_io_in[14]
port 136 nsew
rlabel metal5 s 628240 1018512 640760 1031002 4 mprj_io[15]
port 137 nsew
rlabel metal2 s 636141 995407 636197 995887 4 mprj_io_analog_en[15]
port 138 nsew
rlabel metal2 s 634853 995407 634909 995887 4 mprj_io_analog_pol[15]
port 139 nsew
rlabel metal2 s 631817 995407 631873 995887 4 mprj_io_analog_sel[15]
port 140 nsew
rlabel metal2 s 635497 995407 635553 995887 4 mprj_io_dm[45]
port 141 nsew
rlabel metal2 s 637337 995407 637393 995887 4 mprj_io_dm[46]
port 142 nsew
rlabel metal2 s 631173 995407 631229 995887 4 mprj_io_dm[47]
port 143 nsew
rlabel metal2 s 633013 995407 633069 995887 4 mprj_io_enh[15]
port 144 nsew
rlabel metal2 s 632369 995407 632425 995887 4 mprj_io_hldh_n[15]
port 145 nsew
rlabel metal2 s 630529 995407 630585 995887 4 mprj_io_holdover[15]
port 146 nsew
rlabel metal2 s 627493 995407 627549 995887 4 mprj_io_ib_mode_sel[15]
port 147 nsew
rlabel metal2 s 634301 995407 634357 995887 4 mprj_io_inp_dis[15]
port 148 nsew
rlabel metal2 s 626849 995407 626905 995887 4 mprj_io_oeb[15]
port 149 nsew
rlabel metal2 s 629977 995407 630033 995887 4 mprj_io_out[15]
port 150 nsew
rlabel metal2 s 639177 995407 639233 995887 4 mprj_io_slow_sel[15]
port 151 nsew
rlabel metal2 s 628137 995407 628193 995887 4 mprj_io_vtrip_sel[15]
port 152 nsew
rlabel metal2 s 641017 995407 641073 995887 4 mprj_io_in[15]
port 153 nsew
rlabel metal5 s 526440 1018512 538960 1031002 4 mprj_io[16]
port 154 nsew
rlabel metal2 s 534341 995407 534397 995887 4 mprj_io_analog_en[16]
port 155 nsew
rlabel metal2 s 533053 995407 533109 995887 4 mprj_io_analog_pol[16]
port 156 nsew
rlabel metal2 s 530017 995407 530073 995887 4 mprj_io_analog_sel[16]
port 157 nsew
rlabel metal2 s 533697 995407 533753 995887 4 mprj_io_dm[48]
port 158 nsew
rlabel metal2 s 535537 995407 535593 995887 4 mprj_io_dm[49]
port 159 nsew
rlabel metal2 s 529373 995407 529429 995887 4 mprj_io_dm[50]
port 160 nsew
rlabel metal2 s 531213 995407 531269 995887 4 mprj_io_enh[16]
port 161 nsew
rlabel metal2 s 530569 995407 530625 995887 4 mprj_io_hldh_n[16]
port 162 nsew
rlabel metal2 s 528729 995407 528785 995887 4 mprj_io_holdover[16]
port 163 nsew
rlabel metal2 s 525693 995407 525749 995887 4 mprj_io_ib_mode_sel[16]
port 164 nsew
rlabel metal2 s 532501 995407 532557 995887 4 mprj_io_inp_dis[16]
port 165 nsew
rlabel metal2 s 525049 995407 525105 995887 4 mprj_io_oeb[16]
port 166 nsew
rlabel metal2 s 528177 995407 528233 995887 4 mprj_io_out[16]
port 167 nsew
rlabel metal2 s 537377 995407 537433 995887 4 mprj_io_slow_sel[16]
port 168 nsew
rlabel metal2 s 526337 995407 526393 995887 4 mprj_io_vtrip_sel[16]
port 169 nsew
rlabel metal2 s 539217 995407 539273 995887 4 mprj_io_in[16]
port 170 nsew
rlabel metal5 s 475040 1018512 487560 1031002 4 mprj_io[17]
port 171 nsew
rlabel metal2 s 482941 995407 482997 995887 4 mprj_io_analog_en[17]
port 172 nsew
rlabel metal2 s 481653 995407 481709 995887 4 mprj_io_analog_pol[17]
port 173 nsew
rlabel metal2 s 478617 995407 478673 995887 4 mprj_io_analog_sel[17]
port 174 nsew
rlabel metal2 s 482297 995407 482353 995887 4 mprj_io_dm[51]
port 175 nsew
rlabel metal2 s 484137 995407 484193 995887 4 mprj_io_dm[52]
port 176 nsew
rlabel metal2 s 477973 995407 478029 995887 4 mprj_io_dm[53]
port 177 nsew
rlabel metal2 s 479813 995407 479869 995887 4 mprj_io_enh[17]
port 178 nsew
rlabel metal2 s 479169 995407 479225 995887 4 mprj_io_hldh_n[17]
port 179 nsew
rlabel metal2 s 477329 995407 477385 995887 4 mprj_io_holdover[17]
port 180 nsew
rlabel metal2 s 474293 995407 474349 995887 4 mprj_io_ib_mode_sel[17]
port 181 nsew
rlabel metal2 s 481101 995407 481157 995887 4 mprj_io_inp_dis[17]
port 182 nsew
rlabel metal2 s 473649 995407 473705 995887 4 mprj_io_oeb[17]
port 183 nsew
rlabel metal2 s 476777 995407 476833 995887 4 mprj_io_out[17]
port 184 nsew
rlabel metal2 s 485977 995407 486033 995887 4 mprj_io_slow_sel[17]
port 185 nsew
rlabel metal2 s 474937 995407 474993 995887 4 mprj_io_vtrip_sel[17]
port 186 nsew
rlabel metal2 s 487817 995407 487873 995887 4 mprj_io_in[17]
port 187 nsew
rlabel metal5 s 698512 146440 711002 158960 4 mprj_io[1]
port 188 nsew
rlabel metal2 s 675407 151003 675887 151059 4 mprj_io_analog_en[1]
port 189 nsew
rlabel metal2 s 675407 152291 675887 152347 4 mprj_io_analog_pol[1]
port 190 nsew
rlabel metal2 s 675407 155327 675887 155383 4 mprj_io_analog_sel[1]
port 191 nsew
rlabel metal2 s 675407 151647 675887 151703 4 mprj_io_dm[3]
port 192 nsew
rlabel metal2 s 675407 149807 675887 149863 4 mprj_io_dm[4]
port 193 nsew
rlabel metal2 s 675407 155971 675887 156027 4 mprj_io_dm[5]
port 194 nsew
rlabel metal2 s 675407 154131 675887 154187 4 mprj_io_enh[1]
port 195 nsew
rlabel metal2 s 675407 154775 675887 154831 4 mprj_io_hldh_n[1]
port 196 nsew
rlabel metal2 s 675407 156615 675887 156671 4 mprj_io_holdover[1]
port 197 nsew
rlabel metal2 s 675407 159651 675887 159707 4 mprj_io_ib_mode_sel[1]
port 198 nsew
rlabel metal2 s 675407 152843 675887 152899 4 mprj_io_inp_dis[1]
port 199 nsew
rlabel metal2 s 675407 160295 675887 160351 4 mprj_io_oeb[1]
port 200 nsew
rlabel metal2 s 675407 157167 675887 157223 4 mprj_io_out[1]
port 201 nsew
rlabel metal2 s 675407 147967 675887 148023 4 mprj_io_slow_sel[1]
port 202 nsew
rlabel metal2 s 675407 159007 675887 159063 4 mprj_io_vtrip_sel[1]
port 203 nsew
rlabel metal2 s 675407 146127 675887 146183 4 mprj_io_in[1]
port 204 nsew
rlabel metal5 s 698512 191440 711002 203960 4 mprj_io[2]
port 205 nsew
rlabel metal2 s 675407 196003 675887 196059 4 mprj_io_analog_en[2]
port 206 nsew
rlabel metal2 s 675407 197291 675887 197347 4 mprj_io_analog_pol[2]
port 207 nsew
rlabel metal2 s 675407 200327 675887 200383 4 mprj_io_analog_sel[2]
port 208 nsew
rlabel metal2 s 675407 196647 675887 196703 4 mprj_io_dm[6]
port 209 nsew
rlabel metal2 s 675407 194807 675887 194863 4 mprj_io_dm[7]
port 210 nsew
rlabel metal2 s 675407 200971 675887 201027 4 mprj_io_dm[8]
port 211 nsew
rlabel metal2 s 675407 199131 675887 199187 4 mprj_io_enh[2]
port 212 nsew
rlabel metal2 s 675407 199775 675887 199831 4 mprj_io_hldh_n[2]
port 213 nsew
rlabel metal2 s 675407 201615 675887 201671 4 mprj_io_holdover[2]
port 214 nsew
rlabel metal2 s 675407 204651 675887 204707 4 mprj_io_ib_mode_sel[2]
port 215 nsew
rlabel metal2 s 675407 197843 675887 197899 4 mprj_io_inp_dis[2]
port 216 nsew
rlabel metal2 s 675407 205295 675887 205351 4 mprj_io_oeb[2]
port 217 nsew
rlabel metal2 s 675407 202167 675887 202223 4 mprj_io_out[2]
port 218 nsew
rlabel metal2 s 675407 192967 675887 193023 4 mprj_io_slow_sel[2]
port 219 nsew
rlabel metal2 s 675407 204007 675887 204063 4 mprj_io_vtrip_sel[2]
port 220 nsew
rlabel metal2 s 675407 191127 675887 191183 4 mprj_io_in[2]
port 221 nsew
rlabel metal5 s 698512 236640 711002 249160 4 mprj_io[3]
port 222 nsew
rlabel metal2 s 675407 241203 675887 241259 4 mprj_io_analog_en[3]
port 223 nsew
rlabel metal2 s 675407 242491 675887 242547 4 mprj_io_analog_pol[3]
port 224 nsew
rlabel metal2 s 675407 245527 675887 245583 4 mprj_io_analog_sel[3]
port 225 nsew
rlabel metal2 s 675407 240007 675887 240063 4 mprj_io_dm[10]
port 226 nsew
rlabel metal2 s 675407 246171 675887 246227 4 mprj_io_dm[11]
port 227 nsew
rlabel metal2 s 675407 241847 675887 241903 4 mprj_io_dm[9]
port 228 nsew
rlabel metal2 s 675407 244331 675887 244387 4 mprj_io_enh[3]
port 229 nsew
rlabel metal2 s 675407 244975 675887 245031 4 mprj_io_hldh_n[3]
port 230 nsew
rlabel metal2 s 675407 246815 675887 246871 4 mprj_io_holdover[3]
port 231 nsew
rlabel metal2 s 675407 249851 675887 249907 4 mprj_io_ib_mode_sel[3]
port 232 nsew
rlabel metal2 s 675407 243043 675887 243099 4 mprj_io_inp_dis[3]
port 233 nsew
rlabel metal2 s 675407 250495 675887 250551 4 mprj_io_oeb[3]
port 234 nsew
rlabel metal2 s 675407 247367 675887 247423 4 mprj_io_out[3]
port 235 nsew
rlabel metal2 s 675407 238167 675887 238223 4 mprj_io_slow_sel[3]
port 236 nsew
rlabel metal2 s 675407 249207 675887 249263 4 mprj_io_vtrip_sel[3]
port 237 nsew
rlabel metal2 s 675407 236327 675887 236383 4 mprj_io_in[3]
port 238 nsew
rlabel metal5 s 698512 281640 711002 294160 4 mprj_io[4]
port 239 nsew
rlabel metal2 s 675407 286203 675887 286259 4 mprj_io_analog_en[4]
port 240 nsew
rlabel metal2 s 675407 287491 675887 287547 4 mprj_io_analog_pol[4]
port 241 nsew
rlabel metal2 s 675407 290527 675887 290583 4 mprj_io_analog_sel[4]
port 242 nsew
rlabel metal2 s 675407 286847 675887 286903 4 mprj_io_dm[12]
port 243 nsew
rlabel metal2 s 675407 285007 675887 285063 4 mprj_io_dm[13]
port 244 nsew
rlabel metal2 s 675407 291171 675887 291227 4 mprj_io_dm[14]
port 245 nsew
rlabel metal2 s 675407 289331 675887 289387 4 mprj_io_enh[4]
port 246 nsew
rlabel metal2 s 675407 289975 675887 290031 4 mprj_io_hldh_n[4]
port 247 nsew
rlabel metal2 s 675407 291815 675887 291871 4 mprj_io_holdover[4]
port 248 nsew
rlabel metal2 s 675407 294851 675887 294907 4 mprj_io_ib_mode_sel[4]
port 249 nsew
rlabel metal2 s 675407 288043 675887 288099 4 mprj_io_inp_dis[4]
port 250 nsew
rlabel metal2 s 675407 295495 675887 295551 4 mprj_io_oeb[4]
port 251 nsew
rlabel metal2 s 675407 292367 675887 292423 4 mprj_io_out[4]
port 252 nsew
rlabel metal2 s 675407 283167 675887 283223 4 mprj_io_slow_sel[4]
port 253 nsew
rlabel metal2 s 675407 294207 675887 294263 4 mprj_io_vtrip_sel[4]
port 254 nsew
rlabel metal2 s 675407 281327 675887 281383 4 mprj_io_in[4]
port 255 nsew
rlabel metal5 s 698512 326640 711002 339160 4 mprj_io[5]
port 256 nsew
rlabel metal2 s 675407 331203 675887 331259 4 mprj_io_analog_en[5]
port 257 nsew
rlabel metal2 s 675407 332491 675887 332547 4 mprj_io_analog_pol[5]
port 258 nsew
rlabel metal2 s 675407 335527 675887 335583 4 mprj_io_analog_sel[5]
port 259 nsew
rlabel metal2 s 675407 331847 675887 331903 4 mprj_io_dm[15]
port 260 nsew
rlabel metal2 s 675407 330007 675887 330063 4 mprj_io_dm[16]
port 261 nsew
rlabel metal2 s 675407 336171 675887 336227 4 mprj_io_dm[17]
port 262 nsew
rlabel metal2 s 675407 334331 675887 334387 4 mprj_io_enh[5]
port 263 nsew
rlabel metal2 s 675407 334975 675887 335031 4 mprj_io_hldh_n[5]
port 264 nsew
rlabel metal2 s 675407 336815 675887 336871 4 mprj_io_holdover[5]
port 265 nsew
rlabel metal2 s 675407 339851 675887 339907 4 mprj_io_ib_mode_sel[5]
port 266 nsew
rlabel metal2 s 675407 333043 675887 333099 4 mprj_io_inp_dis[5]
port 267 nsew
rlabel metal2 s 675407 340495 675887 340551 4 mprj_io_oeb[5]
port 268 nsew
rlabel metal2 s 675407 337367 675887 337423 4 mprj_io_out[5]
port 269 nsew
rlabel metal2 s 675407 328167 675887 328223 4 mprj_io_slow_sel[5]
port 270 nsew
rlabel metal2 s 675407 339207 675887 339263 4 mprj_io_vtrip_sel[5]
port 271 nsew
rlabel metal2 s 675407 326327 675887 326383 4 mprj_io_in[5]
port 272 nsew
rlabel metal5 s 698512 371840 711002 384360 4 mprj_io[6]
port 273 nsew
rlabel metal2 s 675407 376403 675887 376459 4 mprj_io_analog_en[6]
port 274 nsew
rlabel metal2 s 675407 377691 675887 377747 4 mprj_io_analog_pol[6]
port 275 nsew
rlabel metal2 s 675407 380727 675887 380783 4 mprj_io_analog_sel[6]
port 276 nsew
rlabel metal2 s 675407 377047 675887 377103 4 mprj_io_dm[18]
port 277 nsew
rlabel metal2 s 675407 375207 675887 375263 4 mprj_io_dm[19]
port 278 nsew
rlabel metal2 s 675407 381371 675887 381427 4 mprj_io_dm[20]
port 279 nsew
rlabel metal2 s 675407 379531 675887 379587 4 mprj_io_enh[6]
port 280 nsew
rlabel metal2 s 675407 380175 675887 380231 4 mprj_io_hldh_n[6]
port 281 nsew
rlabel metal2 s 675407 382015 675887 382071 4 mprj_io_holdover[6]
port 282 nsew
rlabel metal2 s 675407 385051 675887 385107 4 mprj_io_ib_mode_sel[6]
port 283 nsew
rlabel metal2 s 675407 378243 675887 378299 4 mprj_io_inp_dis[6]
port 284 nsew
rlabel metal2 s 675407 385695 675887 385751 4 mprj_io_oeb[6]
port 285 nsew
rlabel metal2 s 675407 382567 675887 382623 4 mprj_io_out[6]
port 286 nsew
rlabel metal2 s 675407 373367 675887 373423 4 mprj_io_slow_sel[6]
port 287 nsew
rlabel metal2 s 675407 384407 675887 384463 4 mprj_io_vtrip_sel[6]
port 288 nsew
rlabel metal2 s 675407 371527 675887 371583 4 mprj_io_in[6]
port 289 nsew
rlabel metal5 s 698512 549040 711002 561560 4 mprj_io[7]
port 290 nsew
rlabel metal2 s 675407 553603 675887 553659 4 mprj_io_analog_en[7]
port 291 nsew
rlabel metal2 s 675407 554891 675887 554947 4 mprj_io_analog_pol[7]
port 292 nsew
rlabel metal2 s 675407 557927 675887 557983 4 mprj_io_analog_sel[7]
port 293 nsew
rlabel metal2 s 675407 554247 675887 554303 4 mprj_io_dm[21]
port 294 nsew
rlabel metal2 s 675407 552407 675887 552463 4 mprj_io_dm[22]
port 295 nsew
rlabel metal2 s 675407 558571 675887 558627 4 mprj_io_dm[23]
port 296 nsew
rlabel metal2 s 675407 556731 675887 556787 4 mprj_io_enh[7]
port 297 nsew
rlabel metal2 s 675407 557375 675887 557431 4 mprj_io_hldh_n[7]
port 298 nsew
rlabel metal2 s 675407 559215 675887 559271 4 mprj_io_holdover[7]
port 299 nsew
rlabel metal2 s 675407 562251 675887 562307 4 mprj_io_ib_mode_sel[7]
port 300 nsew
rlabel metal2 s 675407 555443 675887 555499 4 mprj_io_inp_dis[7]
port 301 nsew
rlabel metal2 s 675407 562895 675887 562951 4 mprj_io_oeb[7]
port 302 nsew
rlabel metal2 s 675407 559767 675887 559823 4 mprj_io_out[7]
port 303 nsew
rlabel metal2 s 675407 550567 675887 550623 4 mprj_io_slow_sel[7]
port 304 nsew
rlabel metal2 s 675407 561607 675887 561663 4 mprj_io_vtrip_sel[7]
port 305 nsew
rlabel metal2 s 675407 548727 675887 548783 4 mprj_io_in[7]
port 306 nsew
rlabel metal5 s 698512 594240 711002 606760 4 mprj_io[8]
port 307 nsew
rlabel metal2 s 675407 598803 675887 598859 4 mprj_io_analog_en[8]
port 308 nsew
rlabel metal2 s 675407 600091 675887 600147 4 mprj_io_analog_pol[8]
port 309 nsew
rlabel metal2 s 675407 603127 675887 603183 4 mprj_io_analog_sel[8]
port 310 nsew
rlabel metal2 s 675407 599447 675887 599503 4 mprj_io_dm[24]
port 311 nsew
rlabel metal2 s 675407 597607 675887 597663 4 mprj_io_dm[25]
port 312 nsew
rlabel metal2 s 675407 603771 675887 603827 4 mprj_io_dm[26]
port 313 nsew
rlabel metal2 s 675407 601931 675887 601987 4 mprj_io_enh[8]
port 314 nsew
rlabel metal2 s 675407 602575 675887 602631 4 mprj_io_hldh_n[8]
port 315 nsew
rlabel metal2 s 675407 604415 675887 604471 4 mprj_io_holdover[8]
port 316 nsew
rlabel metal2 s 675407 607451 675887 607507 4 mprj_io_ib_mode_sel[8]
port 317 nsew
rlabel metal2 s 675407 600643 675887 600699 4 mprj_io_inp_dis[8]
port 318 nsew
rlabel metal2 s 675407 608095 675887 608151 4 mprj_io_oeb[8]
port 319 nsew
rlabel metal2 s 675407 604967 675887 605023 4 mprj_io_out[8]
port 320 nsew
rlabel metal2 s 675407 595767 675887 595823 4 mprj_io_slow_sel[8]
port 321 nsew
rlabel metal2 s 675407 606807 675887 606863 4 mprj_io_vtrip_sel[8]
port 322 nsew
rlabel metal2 s 675407 593927 675887 593983 4 mprj_io_in[8]
port 323 nsew
rlabel metal5 s 698512 639240 711002 651760 4 mprj_io[9]
port 324 nsew
rlabel metal2 s 675407 643803 675887 643859 4 mprj_io_analog_en[9]
port 325 nsew
rlabel metal2 s 675407 645091 675887 645147 4 mprj_io_analog_pol[9]
port 326 nsew
rlabel metal2 s 675407 648127 675887 648183 4 mprj_io_analog_sel[9]
port 327 nsew
rlabel metal2 s 675407 644447 675887 644503 4 mprj_io_dm[27]
port 328 nsew
rlabel metal2 s 675407 642607 675887 642663 4 mprj_io_dm[28]
port 329 nsew
rlabel metal2 s 675407 648771 675887 648827 4 mprj_io_dm[29]
port 330 nsew
rlabel metal2 s 675407 646931 675887 646987 4 mprj_io_enh[9]
port 331 nsew
rlabel metal2 s 675407 647575 675887 647631 4 mprj_io_hldh_n[9]
port 332 nsew
rlabel metal2 s 675407 649415 675887 649471 4 mprj_io_holdover[9]
port 333 nsew
rlabel metal2 s 675407 652451 675887 652507 4 mprj_io_ib_mode_sel[9]
port 334 nsew
rlabel metal2 s 675407 645643 675887 645699 4 mprj_io_inp_dis[9]
port 335 nsew
rlabel metal2 s 675407 653095 675887 653151 4 mprj_io_oeb[9]
port 336 nsew
rlabel metal2 s 675407 649967 675887 650023 4 mprj_io_out[9]
port 337 nsew
rlabel metal2 s 675407 640767 675887 640823 4 mprj_io_slow_sel[9]
port 338 nsew
rlabel metal2 s 675407 651807 675887 651863 4 mprj_io_vtrip_sel[9]
port 339 nsew
rlabel metal2 s 675407 638927 675887 638983 4 mprj_io_in[9]
port 340 nsew
rlabel metal5 s 386040 1018512 398560 1031002 4 mprj_io[18]
port 341 nsew
rlabel metal2 s 393941 995407 393997 995887 4 mprj_io_analog_en[18]
port 342 nsew
rlabel metal2 s 392653 995407 392709 995887 4 mprj_io_analog_pol[18]
port 343 nsew
rlabel metal2 s 389617 995407 389673 995887 4 mprj_io_analog_sel[18]
port 344 nsew
rlabel metal2 s 393297 995407 393353 995887 4 mprj_io_dm[54]
port 345 nsew
rlabel metal2 s 395137 995407 395193 995887 4 mprj_io_dm[55]
port 346 nsew
rlabel metal2 s 388973 995407 389029 995887 4 mprj_io_dm[56]
port 347 nsew
rlabel metal2 s 390813 995407 390869 995887 4 mprj_io_enh[18]
port 348 nsew
rlabel metal2 s 390169 995407 390225 995887 4 mprj_io_hldh_n[18]
port 349 nsew
rlabel metal2 s 388329 995407 388385 995887 4 mprj_io_holdover[18]
port 350 nsew
rlabel metal2 s 385293 995407 385349 995887 4 mprj_io_ib_mode_sel[18]
port 351 nsew
rlabel metal2 s 392101 995407 392157 995887 4 mprj_io_inp_dis[18]
port 352 nsew
rlabel metal2 s 384649 995407 384705 995887 4 mprj_io_oeb[18]
port 353 nsew
rlabel metal2 s 387777 995407 387833 995887 4 mprj_io_out[18]
port 354 nsew
rlabel metal2 s 396977 995407 397033 995887 4 mprj_io_slow_sel[18]
port 355 nsew
rlabel metal2 s 385937 995407 385993 995887 4 mprj_io_vtrip_sel[18]
port 356 nsew
rlabel metal2 s 398817 995407 398873 995887 4 mprj_io_in[18]
port 357 nsew
rlabel metal5 s 6598 657040 19088 669560 4 mprj_io[28]
port 358 nsew
rlabel metal2 s 41713 664941 42193 664997 4 mprj_io_analog_en[28]
port 359 nsew
rlabel metal2 s 41713 663653 42193 663709 4 mprj_io_analog_pol[28]
port 360 nsew
rlabel metal2 s 41713 660617 42193 660673 4 mprj_io_analog_sel[28]
port 361 nsew
rlabel metal2 s 41713 664297 42193 664353 4 mprj_io_dm[84]
port 362 nsew
rlabel metal2 s 41713 666137 42193 666193 4 mprj_io_dm[85]
port 363 nsew
rlabel metal2 s 41713 659973 42193 660029 4 mprj_io_dm[86]
port 364 nsew
rlabel metal2 s 41713 661813 42193 661869 4 mprj_io_enh[28]
port 365 nsew
rlabel metal2 s 41713 661169 42193 661225 4 mprj_io_hldh_n[28]
port 366 nsew
rlabel metal2 s 41713 659329 42193 659385 4 mprj_io_holdover[28]
port 367 nsew
rlabel metal2 s 41713 656293 42193 656349 4 mprj_io_ib_mode_sel[28]
port 368 nsew
rlabel metal2 s 41713 663101 42193 663157 4 mprj_io_inp_dis[28]
port 369 nsew
rlabel metal2 s 41713 655649 42193 655705 4 mprj_io_oeb[28]
port 370 nsew
rlabel metal2 s 41713 658777 42193 658833 4 mprj_io_out[28]
port 371 nsew
rlabel metal2 s 41713 667977 42193 668033 4 mprj_io_slow_sel[28]
port 372 nsew
rlabel metal2 s 41713 656937 42193 656993 4 mprj_io_vtrip_sel[28]
port 373 nsew
rlabel metal2 s 41713 669817 42193 669873 4 mprj_io_in[28]
port 374 nsew
rlabel metal5 s 6598 613840 19088 626360 4 mprj_io[29]
port 375 nsew
rlabel metal2 s 41713 621741 42193 621797 4 mprj_io_analog_en[29]
port 376 nsew
rlabel metal2 s 41713 620453 42193 620509 4 mprj_io_analog_pol[29]
port 377 nsew
rlabel metal2 s 41713 617417 42193 617473 4 mprj_io_analog_sel[29]
port 378 nsew
rlabel metal2 s 41713 621097 42193 621153 4 mprj_io_dm[87]
port 379 nsew
rlabel metal2 s 41713 622937 42193 622993 4 mprj_io_dm[88]
port 380 nsew
rlabel metal2 s 41713 616773 42193 616829 4 mprj_io_dm[89]
port 381 nsew
rlabel metal2 s 41713 618613 42193 618669 4 mprj_io_enh[29]
port 382 nsew
rlabel metal2 s 41713 617969 42193 618025 4 mprj_io_hldh_n[29]
port 383 nsew
rlabel metal2 s 41713 616129 42193 616185 4 mprj_io_holdover[29]
port 384 nsew
rlabel metal2 s 41713 613093 42193 613149 4 mprj_io_ib_mode_sel[29]
port 385 nsew
rlabel metal2 s 41713 619901 42193 619957 4 mprj_io_inp_dis[29]
port 386 nsew
rlabel metal2 s 41713 612449 42193 612505 4 mprj_io_oeb[29]
port 387 nsew
rlabel metal2 s 41713 615577 42193 615633 4 mprj_io_out[29]
port 388 nsew
rlabel metal2 s 41713 624777 42193 624833 4 mprj_io_slow_sel[29]
port 389 nsew
rlabel metal2 s 41713 613737 42193 613793 4 mprj_io_vtrip_sel[29]
port 390 nsew
rlabel metal2 s 41713 626617 42193 626673 4 mprj_io_in[29]
port 391 nsew
rlabel metal5 s 6598 570640 19088 583160 4 mprj_io[30]
port 392 nsew
rlabel metal2 s 41713 578541 42193 578597 4 mprj_io_analog_en[30]
port 393 nsew
rlabel metal2 s 41713 577253 42193 577309 4 mprj_io_analog_pol[30]
port 394 nsew
rlabel metal2 s 41713 574217 42193 574273 4 mprj_io_analog_sel[30]
port 395 nsew
rlabel metal2 s 41713 577897 42193 577953 4 mprj_io_dm[90]
port 396 nsew
rlabel metal2 s 41713 579737 42193 579793 4 mprj_io_dm[91]
port 397 nsew
rlabel metal2 s 41713 573573 42193 573629 4 mprj_io_dm[92]
port 398 nsew
rlabel metal2 s 41713 575413 42193 575469 4 mprj_io_enh[30]
port 399 nsew
rlabel metal2 s 41713 574769 42193 574825 4 mprj_io_hldh_n[30]
port 400 nsew
rlabel metal2 s 41713 572929 42193 572985 4 mprj_io_holdover[30]
port 401 nsew
rlabel metal2 s 41713 569893 42193 569949 4 mprj_io_ib_mode_sel[30]
port 402 nsew
rlabel metal2 s 41713 576701 42193 576757 4 mprj_io_inp_dis[30]
port 403 nsew
rlabel metal2 s 41713 569249 42193 569305 4 mprj_io_oeb[30]
port 404 nsew
rlabel metal2 s 41713 572377 42193 572433 4 mprj_io_out[30]
port 405 nsew
rlabel metal2 s 41713 581577 42193 581633 4 mprj_io_slow_sel[30]
port 406 nsew
rlabel metal2 s 41713 570537 42193 570593 4 mprj_io_vtrip_sel[30]
port 407 nsew
rlabel metal2 s 41713 583417 42193 583473 4 mprj_io_in[30]
port 408 nsew
rlabel metal5 s 6598 527440 19088 539960 4 mprj_io[31]
port 409 nsew
rlabel metal2 s 41713 535341 42193 535397 4 mprj_io_analog_en[31]
port 410 nsew
rlabel metal2 s 41713 534053 42193 534109 4 mprj_io_analog_pol[31]
port 411 nsew
rlabel metal2 s 41713 531017 42193 531073 4 mprj_io_analog_sel[31]
port 412 nsew
rlabel metal2 s 41713 534697 42193 534753 4 mprj_io_dm[93]
port 413 nsew
rlabel metal2 s 41713 536537 42193 536593 4 mprj_io_dm[94]
port 414 nsew
rlabel metal2 s 41713 530373 42193 530429 4 mprj_io_dm[95]
port 415 nsew
rlabel metal2 s 41713 532213 42193 532269 4 mprj_io_enh[31]
port 416 nsew
rlabel metal2 s 41713 531569 42193 531625 4 mprj_io_hldh_n[31]
port 417 nsew
rlabel metal2 s 41713 529729 42193 529785 4 mprj_io_holdover[31]
port 418 nsew
rlabel metal2 s 41713 526693 42193 526749 4 mprj_io_ib_mode_sel[31]
port 419 nsew
rlabel metal2 s 41713 533501 42193 533557 4 mprj_io_inp_dis[31]
port 420 nsew
rlabel metal2 s 41713 526049 42193 526105 4 mprj_io_oeb[31]
port 421 nsew
rlabel metal2 s 41713 529177 42193 529233 4 mprj_io_out[31]
port 422 nsew
rlabel metal2 s 41713 538377 42193 538433 4 mprj_io_slow_sel[31]
port 423 nsew
rlabel metal2 s 41713 527337 42193 527393 4 mprj_io_vtrip_sel[31]
port 424 nsew
rlabel metal2 s 41713 540217 42193 540273 4 mprj_io_in[31]
port 425 nsew
rlabel metal5 s 6598 399840 19088 412360 4 mprj_io[32]
port 426 nsew
rlabel metal2 s 41713 407741 42193 407797 4 mprj_io_analog_en[32]
port 427 nsew
rlabel metal2 s 41713 406453 42193 406509 4 mprj_io_analog_pol[32]
port 428 nsew
rlabel metal2 s 41713 403417 42193 403473 4 mprj_io_analog_sel[32]
port 429 nsew
rlabel metal2 s 41713 407097 42193 407153 4 mprj_io_dm[96]
port 430 nsew
rlabel metal2 s 41713 408937 42193 408993 4 mprj_io_dm[97]
port 431 nsew
rlabel metal2 s 41713 402773 42193 402829 4 mprj_io_dm[98]
port 432 nsew
rlabel metal2 s 41713 404613 42193 404669 4 mprj_io_enh[32]
port 433 nsew
rlabel metal2 s 41713 403969 42193 404025 4 mprj_io_hldh_n[32]
port 434 nsew
rlabel metal2 s 41713 402129 42193 402185 4 mprj_io_holdover[32]
port 435 nsew
rlabel metal2 s 41713 399093 42193 399149 4 mprj_io_ib_mode_sel[32]
port 436 nsew
rlabel metal2 s 41713 405901 42193 405957 4 mprj_io_inp_dis[32]
port 437 nsew
rlabel metal2 s 41713 398449 42193 398505 4 mprj_io_oeb[32]
port 438 nsew
rlabel metal2 s 41713 401577 42193 401633 4 mprj_io_out[32]
port 439 nsew
rlabel metal2 s 41713 410777 42193 410833 4 mprj_io_slow_sel[32]
port 440 nsew
rlabel metal2 s 41713 399737 42193 399793 4 mprj_io_vtrip_sel[32]
port 441 nsew
rlabel metal2 s 41713 412617 42193 412673 4 mprj_io_in[32]
port 442 nsew
rlabel metal5 s 6598 356640 19088 369160 4 mprj_io[33]
port 443 nsew
rlabel metal2 s 41713 364541 42193 364597 4 mprj_io_analog_en[33]
port 444 nsew
rlabel metal2 s 41713 363253 42193 363309 4 mprj_io_analog_pol[33]
port 445 nsew
rlabel metal2 s 41713 360217 42193 360273 4 mprj_io_analog_sel[33]
port 446 nsew
rlabel metal2 s 41713 365737 42193 365793 4 mprj_io_dm[100]
port 447 nsew
rlabel metal2 s 41713 359573 42193 359629 4 mprj_io_dm[101]
port 448 nsew
rlabel metal2 s 41713 363897 42193 363953 4 mprj_io_dm[99]
port 449 nsew
rlabel metal2 s 41713 361413 42193 361469 4 mprj_io_enh[33]
port 450 nsew
rlabel metal2 s 41713 360769 42193 360825 4 mprj_io_hldh_n[33]
port 451 nsew
rlabel metal2 s 41713 358929 42193 358985 4 mprj_io_holdover[33]
port 452 nsew
rlabel metal2 s 41713 355893 42193 355949 4 mprj_io_ib_mode_sel[33]
port 453 nsew
rlabel metal2 s 41713 362701 42193 362757 4 mprj_io_inp_dis[33]
port 454 nsew
rlabel metal2 s 41713 355249 42193 355305 4 mprj_io_oeb[33]
port 455 nsew
rlabel metal2 s 41713 358377 42193 358433 4 mprj_io_out[33]
port 456 nsew
rlabel metal2 s 41713 367577 42193 367633 4 mprj_io_slow_sel[33]
port 457 nsew
rlabel metal2 s 41713 356537 42193 356593 4 mprj_io_vtrip_sel[33]
port 458 nsew
rlabel metal2 s 41713 369417 42193 369473 4 mprj_io_in[33]
port 459 nsew
rlabel metal5 s 6598 313440 19088 325960 4 mprj_io[34]
port 460 nsew
rlabel metal2 s 41713 321341 42193 321397 4 mprj_io_analog_en[34]
port 461 nsew
rlabel metal2 s 41713 320053 42193 320109 4 mprj_io_analog_pol[34]
port 462 nsew
rlabel metal2 s 41713 317017 42193 317073 4 mprj_io_analog_sel[34]
port 463 nsew
rlabel metal2 s 41713 320697 42193 320753 4 mprj_io_dm[102]
port 464 nsew
rlabel metal2 s 41713 322537 42193 322593 4 mprj_io_dm[103]
port 465 nsew
rlabel metal2 s 41713 316373 42193 316429 4 mprj_io_dm[104]
port 466 nsew
rlabel metal2 s 41713 318213 42193 318269 4 mprj_io_enh[34]
port 467 nsew
rlabel metal2 s 41713 317569 42193 317625 4 mprj_io_hldh_n[34]
port 468 nsew
rlabel metal2 s 41713 315729 42193 315785 4 mprj_io_holdover[34]
port 469 nsew
rlabel metal2 s 41713 312693 42193 312749 4 mprj_io_ib_mode_sel[34]
port 470 nsew
rlabel metal2 s 41713 319501 42193 319557 4 mprj_io_inp_dis[34]
port 471 nsew
rlabel metal2 s 41713 312049 42193 312105 4 mprj_io_oeb[34]
port 472 nsew
rlabel metal2 s 41713 315177 42193 315233 4 mprj_io_out[34]
port 473 nsew
rlabel metal2 s 41713 324377 42193 324433 4 mprj_io_slow_sel[34]
port 474 nsew
rlabel metal2 s 41713 313337 42193 313393 4 mprj_io_vtrip_sel[34]
port 475 nsew
rlabel metal2 s 41713 326217 42193 326273 4 mprj_io_in[34]
port 476 nsew
rlabel metal5 s 6598 270240 19088 282760 4 mprj_io[35]
port 477 nsew
rlabel metal2 s 41713 278141 42193 278197 4 mprj_io_analog_en[35]
port 478 nsew
rlabel metal2 s 41713 276853 42193 276909 4 mprj_io_analog_pol[35]
port 479 nsew
rlabel metal2 s 41713 273817 42193 273873 4 mprj_io_analog_sel[35]
port 480 nsew
rlabel metal2 s 41713 277497 42193 277553 4 mprj_io_dm[105]
port 481 nsew
rlabel metal2 s 41713 279337 42193 279393 4 mprj_io_dm[106]
port 482 nsew
rlabel metal2 s 41713 273173 42193 273229 4 mprj_io_dm[107]
port 483 nsew
rlabel metal2 s 41713 275013 42193 275069 4 mprj_io_enh[35]
port 484 nsew
rlabel metal2 s 41713 274369 42193 274425 4 mprj_io_hldh_n[35]
port 485 nsew
rlabel metal2 s 41713 272529 42193 272585 4 mprj_io_holdover[35]
port 486 nsew
rlabel metal2 s 41713 269493 42193 269549 4 mprj_io_ib_mode_sel[35]
port 487 nsew
rlabel metal2 s 41713 276301 42193 276357 4 mprj_io_inp_dis[35]
port 488 nsew
rlabel metal2 s 41713 268849 42193 268905 4 mprj_io_oeb[35]
port 489 nsew
rlabel metal2 s 41713 271977 42193 272033 4 mprj_io_out[35]
port 490 nsew
rlabel metal2 s 41713 281177 42193 281233 4 mprj_io_slow_sel[35]
port 491 nsew
rlabel metal2 s 41713 270137 42193 270193 4 mprj_io_vtrip_sel[35]
port 492 nsew
rlabel metal2 s 41713 283017 42193 283073 4 mprj_io_in[35]
port 493 nsew
rlabel metal5 s 6598 227040 19088 239560 4 mprj_io[36]
port 494 nsew
rlabel metal2 s 41713 234941 42193 234997 4 mprj_io_analog_en[36]
port 495 nsew
rlabel metal2 s 41713 233653 42193 233709 4 mprj_io_analog_pol[36]
port 496 nsew
rlabel metal2 s 41713 230617 42193 230673 4 mprj_io_analog_sel[36]
port 497 nsew
rlabel metal2 s 41713 234297 42193 234353 4 mprj_io_dm[108]
port 498 nsew
rlabel metal2 s 41713 236137 42193 236193 4 mprj_io_dm[109]
port 499 nsew
rlabel metal2 s 41713 229973 42193 230029 4 mprj_io_dm[110]
port 500 nsew
rlabel metal2 s 41713 231813 42193 231869 4 mprj_io_enh[36]
port 501 nsew
rlabel metal2 s 41713 231169 42193 231225 4 mprj_io_hldh_n[36]
port 502 nsew
rlabel metal2 s 41713 229329 42193 229385 4 mprj_io_holdover[36]
port 503 nsew
rlabel metal2 s 41713 226293 42193 226349 4 mprj_io_ib_mode_sel[36]
port 504 nsew
rlabel metal2 s 41713 233101 42193 233157 4 mprj_io_inp_dis[36]
port 505 nsew
rlabel metal2 s 41713 225649 42193 225705 4 mprj_io_oeb[36]
port 506 nsew
rlabel metal2 s 41713 228777 42193 228833 4 mprj_io_out[36]
port 507 nsew
rlabel metal2 s 41713 237977 42193 238033 4 mprj_io_slow_sel[36]
port 508 nsew
rlabel metal2 s 41713 226937 42193 226993 4 mprj_io_vtrip_sel[36]
port 509 nsew
rlabel metal2 s 41713 239817 42193 239873 4 mprj_io_in[36]
port 510 nsew
rlabel metal5 s 6598 183840 19088 196360 4 mprj_io[37]
port 511 nsew
rlabel metal2 s 41713 191741 42193 191797 4 mprj_io_analog_en[37]
port 512 nsew
rlabel metal2 s 41713 190453 42193 190509 4 mprj_io_analog_pol[37]
port 513 nsew
rlabel metal2 s 41713 187417 42193 187473 4 mprj_io_analog_sel[37]
port 514 nsew
rlabel metal2 s 41713 191097 42193 191153 4 mprj_io_dm[111]
port 515 nsew
rlabel metal2 s 41713 192937 42193 192993 4 mprj_io_dm[112]
port 516 nsew
rlabel metal2 s 41713 186773 42193 186829 4 mprj_io_dm[113]
port 517 nsew
rlabel metal2 s 41713 188613 42193 188669 4 mprj_io_enh[37]
port 518 nsew
rlabel metal2 s 41713 187969 42193 188025 4 mprj_io_hldh_n[37]
port 519 nsew
rlabel metal2 s 41713 186129 42193 186185 4 mprj_io_holdover[37]
port 520 nsew
rlabel metal2 s 41713 183093 42193 183149 4 mprj_io_ib_mode_sel[37]
port 521 nsew
rlabel metal2 s 41713 189901 42193 189957 4 mprj_io_inp_dis[37]
port 522 nsew
rlabel metal2 s 41713 182449 42193 182505 4 mprj_io_oeb[37]
port 523 nsew
rlabel metal2 s 41713 185577 42193 185633 4 mprj_io_out[37]
port 524 nsew
rlabel metal2 s 41713 194777 42193 194833 4 mprj_io_slow_sel[37]
port 525 nsew
rlabel metal2 s 41713 183737 42193 183793 4 mprj_io_vtrip_sel[37]
port 526 nsew
rlabel metal2 s 41713 196617 42193 196673 4 mprj_io_in[37]
port 527 nsew
rlabel metal5 s 284240 1018512 296760 1031002 4 mprj_io[19]
port 528 nsew
rlabel metal2 s 292141 995407 292197 995887 4 mprj_io_analog_en[19]
port 529 nsew
rlabel metal2 s 290853 995407 290909 995887 4 mprj_io_analog_pol[19]
port 530 nsew
rlabel metal2 s 287817 995407 287873 995887 4 mprj_io_analog_sel[19]
port 531 nsew
rlabel metal2 s 291497 995407 291553 995887 4 mprj_io_dm[57]
port 532 nsew
rlabel metal2 s 293337 995407 293393 995887 4 mprj_io_dm[58]
port 533 nsew
rlabel metal2 s 287173 995407 287229 995887 4 mprj_io_dm[59]
port 534 nsew
rlabel metal2 s 289013 995407 289069 995887 4 mprj_io_enh[19]
port 535 nsew
rlabel metal2 s 288369 995407 288425 995887 4 mprj_io_hldh_n[19]
port 536 nsew
rlabel metal2 s 286529 995407 286585 995887 4 mprj_io_holdover[19]
port 537 nsew
rlabel metal2 s 283493 995407 283549 995887 4 mprj_io_ib_mode_sel[19]
port 538 nsew
rlabel metal2 s 290301 995407 290357 995887 4 mprj_io_inp_dis[19]
port 539 nsew
rlabel metal2 s 282849 995407 282905 995887 4 mprj_io_oeb[19]
port 540 nsew
rlabel metal2 s 285977 995407 286033 995887 4 mprj_io_out[19]
port 541 nsew
rlabel metal2 s 295177 995407 295233 995887 4 mprj_io_slow_sel[19]
port 542 nsew
rlabel metal2 s 284137 995407 284193 995887 4 mprj_io_vtrip_sel[19]
port 543 nsew
rlabel metal2 s 297017 995407 297073 995887 4 mprj_io_in[19]
port 544 nsew
rlabel metal5 s 232640 1018512 245160 1031002 4 mprj_io[20]
port 545 nsew
rlabel metal2 s 240541 995407 240597 995887 4 mprj_io_analog_en[20]
port 546 nsew
rlabel metal2 s 239253 995407 239309 995887 4 mprj_io_analog_pol[20]
port 547 nsew
rlabel metal2 s 236217 995407 236273 995887 4 mprj_io_analog_sel[20]
port 548 nsew
rlabel metal2 s 239897 995407 239953 995887 4 mprj_io_dm[60]
port 549 nsew
rlabel metal2 s 241737 995407 241793 995887 4 mprj_io_dm[61]
port 550 nsew
rlabel metal2 s 235573 995407 235629 995887 4 mprj_io_dm[62]
port 551 nsew
rlabel metal2 s 237413 995407 237469 995887 4 mprj_io_enh[20]
port 552 nsew
rlabel metal2 s 236769 995407 236825 995887 4 mprj_io_hldh_n[20]
port 553 nsew
rlabel metal2 s 234929 995407 234985 995887 4 mprj_io_holdover[20]
port 554 nsew
rlabel metal2 s 231893 995407 231949 995887 4 mprj_io_ib_mode_sel[20]
port 555 nsew
rlabel metal2 s 238701 995407 238757 995887 4 mprj_io_inp_dis[20]
port 556 nsew
rlabel metal2 s 231249 995407 231305 995887 4 mprj_io_oeb[20]
port 557 nsew
rlabel metal2 s 234377 995407 234433 995887 4 mprj_io_out[20]
port 558 nsew
rlabel metal2 s 243577 995407 243633 995887 4 mprj_io_slow_sel[20]
port 559 nsew
rlabel metal2 s 232537 995407 232593 995887 4 mprj_io_vtrip_sel[20]
port 560 nsew
rlabel metal2 s 245417 995407 245473 995887 4 mprj_io_in[20]
port 561 nsew
rlabel metal5 s 181240 1018512 193760 1031002 4 mprj_io[21]
port 562 nsew
rlabel metal2 s 189141 995407 189197 995887 4 mprj_io_analog_en[21]
port 563 nsew
rlabel metal2 s 187853 995407 187909 995887 4 mprj_io_analog_pol[21]
port 564 nsew
rlabel metal2 s 184817 995407 184873 995887 4 mprj_io_analog_sel[21]
port 565 nsew
rlabel metal2 s 188497 995407 188553 995887 4 mprj_io_dm[63]
port 566 nsew
rlabel metal2 s 190337 995407 190393 995887 4 mprj_io_dm[64]
port 567 nsew
rlabel metal2 s 184173 995407 184229 995887 4 mprj_io_dm[65]
port 568 nsew
rlabel metal2 s 186013 995407 186069 995887 4 mprj_io_enh[21]
port 569 nsew
rlabel metal2 s 185369 995407 185425 995887 4 mprj_io_hldh_n[21]
port 570 nsew
rlabel metal2 s 183529 995407 183585 995887 4 mprj_io_holdover[21]
port 571 nsew
rlabel metal2 s 180493 995407 180549 995887 4 mprj_io_ib_mode_sel[21]
port 572 nsew
rlabel metal2 s 187301 995407 187357 995887 4 mprj_io_inp_dis[21]
port 573 nsew
rlabel metal2 s 179849 995407 179905 995887 4 mprj_io_oeb[21]
port 574 nsew
rlabel metal2 s 182977 995407 183033 995887 4 mprj_io_out[21]
port 575 nsew
rlabel metal2 s 192177 995407 192233 995887 4 mprj_io_slow_sel[21]
port 576 nsew
rlabel metal2 s 181137 995407 181193 995887 4 mprj_io_vtrip_sel[21]
port 577 nsew
rlabel metal2 s 194017 995407 194073 995887 4 mprj_io_in[21]
port 578 nsew
rlabel metal5 s 129840 1018512 142360 1031002 4 mprj_io[22]
port 579 nsew
rlabel metal2 s 137741 995407 137797 995887 4 mprj_io_analog_en[22]
port 580 nsew
rlabel metal2 s 136453 995407 136509 995887 4 mprj_io_analog_pol[22]
port 581 nsew
rlabel metal2 s 133417 995407 133473 995887 4 mprj_io_analog_sel[22]
port 582 nsew
rlabel metal2 s 137097 995407 137153 995887 4 mprj_io_dm[66]
port 583 nsew
rlabel metal2 s 138937 995407 138993 995887 4 mprj_io_dm[67]
port 584 nsew
rlabel metal2 s 132773 995407 132829 995887 4 mprj_io_dm[68]
port 585 nsew
rlabel metal2 s 134613 995407 134669 995887 4 mprj_io_enh[22]
port 586 nsew
rlabel metal2 s 133969 995407 134025 995887 4 mprj_io_hldh_n[22]
port 587 nsew
rlabel metal2 s 132129 995407 132185 995887 4 mprj_io_holdover[22]
port 588 nsew
rlabel metal2 s 129093 995407 129149 995887 4 mprj_io_ib_mode_sel[22]
port 589 nsew
rlabel metal2 s 135901 995407 135957 995887 4 mprj_io_inp_dis[22]
port 590 nsew
rlabel metal2 s 128449 995407 128505 995887 4 mprj_io_oeb[22]
port 591 nsew
rlabel metal2 s 131577 995407 131633 995887 4 mprj_io_out[22]
port 592 nsew
rlabel metal2 s 140777 995407 140833 995887 4 mprj_io_slow_sel[22]
port 593 nsew
rlabel metal2 s 129737 995407 129793 995887 4 mprj_io_vtrip_sel[22]
port 594 nsew
rlabel metal2 s 142617 995407 142673 995887 4 mprj_io_in[22]
port 595 nsew
rlabel metal5 s 78440 1018512 90960 1031002 4 mprj_io[23]
port 596 nsew
rlabel metal2 s 86341 995407 86397 995887 4 mprj_io_analog_en[23]
port 597 nsew
rlabel metal2 s 85053 995407 85109 995887 4 mprj_io_analog_pol[23]
port 598 nsew
rlabel metal2 s 82017 995407 82073 995887 4 mprj_io_analog_sel[23]
port 599 nsew
rlabel metal2 s 85697 995407 85753 995887 4 mprj_io_dm[69]
port 600 nsew
rlabel metal2 s 87537 995407 87593 995887 4 mprj_io_dm[70]
port 601 nsew
rlabel metal2 s 81373 995407 81429 995887 4 mprj_io_dm[71]
port 602 nsew
rlabel metal2 s 83213 995407 83269 995887 4 mprj_io_enh[23]
port 603 nsew
rlabel metal2 s 82569 995407 82625 995887 4 mprj_io_hldh_n[23]
port 604 nsew
rlabel metal2 s 80729 995407 80785 995887 4 mprj_io_holdover[23]
port 605 nsew
rlabel metal2 s 77693 995407 77749 995887 4 mprj_io_ib_mode_sel[23]
port 606 nsew
rlabel metal2 s 84501 995407 84557 995887 4 mprj_io_inp_dis[23]
port 607 nsew
rlabel metal2 s 77049 995407 77105 995887 4 mprj_io_oeb[23]
port 608 nsew
rlabel metal2 s 80177 995407 80233 995887 4 mprj_io_out[23]
port 609 nsew
rlabel metal2 s 89377 995407 89433 995887 4 mprj_io_slow_sel[23]
port 610 nsew
rlabel metal2 s 78337 995407 78393 995887 4 mprj_io_vtrip_sel[23]
port 611 nsew
rlabel metal2 s 91217 995407 91273 995887 4 mprj_io_in[23]
port 612 nsew
rlabel metal5 s 6598 956440 19088 968960 4 mprj_io[24]
port 613 nsew
rlabel metal2 s 41713 964341 42193 964397 4 mprj_io_analog_en[24]
port 614 nsew
rlabel metal2 s 41713 963053 42193 963109 4 mprj_io_analog_pol[24]
port 615 nsew
rlabel metal2 s 41713 960017 42193 960073 4 mprj_io_analog_sel[24]
port 616 nsew
rlabel metal2 s 41713 963697 42193 963753 4 mprj_io_dm[72]
port 617 nsew
rlabel metal2 s 41713 965537 42193 965593 4 mprj_io_dm[73]
port 618 nsew
rlabel metal2 s 41713 959373 42193 959429 4 mprj_io_dm[74]
port 619 nsew
rlabel metal2 s 41713 961213 42193 961269 4 mprj_io_enh[24]
port 620 nsew
rlabel metal2 s 41713 960569 42193 960625 4 mprj_io_hldh_n[24]
port 621 nsew
rlabel metal2 s 41713 958729 42193 958785 4 mprj_io_holdover[24]
port 622 nsew
rlabel metal2 s 41713 955693 42193 955749 4 mprj_io_ib_mode_sel[24]
port 623 nsew
rlabel metal2 s 41713 962501 42193 962557 4 mprj_io_inp_dis[24]
port 624 nsew
rlabel metal2 s 41713 955049 42193 955105 4 mprj_io_oeb[24]
port 625 nsew
rlabel metal2 s 41713 958177 42193 958233 4 mprj_io_out[24]
port 626 nsew
rlabel metal2 s 41713 967377 42193 967433 4 mprj_io_slow_sel[24]
port 627 nsew
rlabel metal2 s 41713 956337 42193 956393 4 mprj_io_vtrip_sel[24]
port 628 nsew
rlabel metal2 s 41713 969217 42193 969273 4 mprj_io_in[24]
port 629 nsew
rlabel metal5 s 6598 786640 19088 799160 4 mprj_io[25]
port 630 nsew
rlabel metal2 s 41713 794541 42193 794597 4 mprj_io_analog_en[25]
port 631 nsew
rlabel metal2 s 41713 793253 42193 793309 4 mprj_io_analog_pol[25]
port 632 nsew
rlabel metal2 s 41713 790217 42193 790273 4 mprj_io_analog_sel[25]
port 633 nsew
rlabel metal2 s 41713 793897 42193 793953 4 mprj_io_dm[75]
port 634 nsew
rlabel metal2 s 41713 795737 42193 795793 4 mprj_io_dm[76]
port 635 nsew
rlabel metal2 s 41713 789573 42193 789629 4 mprj_io_dm[77]
port 636 nsew
rlabel metal2 s 41713 791413 42193 791469 4 mprj_io_enh[25]
port 637 nsew
rlabel metal2 s 41713 790769 42193 790825 4 mprj_io_hldh_n[25]
port 638 nsew
rlabel metal2 s 41713 788929 42193 788985 4 mprj_io_holdover[25]
port 639 nsew
rlabel metal2 s 41713 785893 42193 785949 4 mprj_io_ib_mode_sel[25]
port 640 nsew
rlabel metal2 s 41713 792701 42193 792757 4 mprj_io_inp_dis[25]
port 641 nsew
rlabel metal2 s 41713 785249 42193 785305 4 mprj_io_oeb[25]
port 642 nsew
rlabel metal2 s 41713 788377 42193 788433 4 mprj_io_out[25]
port 643 nsew
rlabel metal2 s 41713 797577 42193 797633 4 mprj_io_slow_sel[25]
port 644 nsew
rlabel metal2 s 41713 786537 42193 786593 4 mprj_io_vtrip_sel[25]
port 645 nsew
rlabel metal2 s 41713 799417 42193 799473 4 mprj_io_in[25]
port 646 nsew
rlabel metal5 s 6598 743440 19088 755960 4 mprj_io[26]
port 647 nsew
rlabel metal2 s 41713 751341 42193 751397 4 mprj_io_analog_en[26]
port 648 nsew
rlabel metal2 s 41713 750053 42193 750109 4 mprj_io_analog_pol[26]
port 649 nsew
rlabel metal2 s 41713 747017 42193 747073 4 mprj_io_analog_sel[26]
port 650 nsew
rlabel metal2 s 41713 750697 42193 750753 4 mprj_io_dm[78]
port 651 nsew
rlabel metal2 s 41713 752537 42193 752593 4 mprj_io_dm[79]
port 652 nsew
rlabel metal2 s 41713 746373 42193 746429 4 mprj_io_dm[80]
port 653 nsew
rlabel metal2 s 41713 748213 42193 748269 4 mprj_io_enh[26]
port 654 nsew
rlabel metal2 s 41713 747569 42193 747625 4 mprj_io_hldh_n[26]
port 655 nsew
rlabel metal2 s 41713 745729 42193 745785 4 mprj_io_holdover[26]
port 656 nsew
rlabel metal2 s 41713 742693 42193 742749 4 mprj_io_ib_mode_sel[26]
port 657 nsew
rlabel metal2 s 41713 749501 42193 749557 4 mprj_io_inp_dis[26]
port 658 nsew
rlabel metal2 s 41713 742049 42193 742105 4 mprj_io_oeb[26]
port 659 nsew
rlabel metal2 s 41713 745177 42193 745233 4 mprj_io_out[26]
port 660 nsew
rlabel metal2 s 41713 754377 42193 754433 4 mprj_io_slow_sel[26]
port 661 nsew
rlabel metal2 s 41713 743337 42193 743393 4 mprj_io_vtrip_sel[26]
port 662 nsew
rlabel metal2 s 41713 756217 42193 756273 4 mprj_io_in[26]
port 663 nsew
rlabel metal5 s 6598 700240 19088 712760 4 mprj_io[27]
port 664 nsew
rlabel metal2 s 41713 708141 42193 708197 4 mprj_io_analog_en[27]
port 665 nsew
rlabel metal2 s 41713 706853 42193 706909 4 mprj_io_analog_pol[27]
port 666 nsew
rlabel metal2 s 41713 703817 42193 703873 4 mprj_io_analog_sel[27]
port 667 nsew
rlabel metal2 s 41713 707497 42193 707553 4 mprj_io_dm[81]
port 668 nsew
rlabel metal2 s 41713 709337 42193 709393 4 mprj_io_dm[82]
port 669 nsew
rlabel metal2 s 41713 703173 42193 703229 4 mprj_io_dm[83]
port 670 nsew
rlabel metal2 s 41713 705013 42193 705069 4 mprj_io_enh[27]
port 671 nsew
rlabel metal2 s 41713 704369 42193 704425 4 mprj_io_hldh_n[27]
port 672 nsew
rlabel metal2 s 41713 702529 42193 702585 4 mprj_io_holdover[27]
port 673 nsew
rlabel metal2 s 41713 699493 42193 699549 4 mprj_io_ib_mode_sel[27]
port 674 nsew
rlabel metal2 s 41713 706301 42193 706357 4 mprj_io_inp_dis[27]
port 675 nsew
rlabel metal2 s 41713 698849 42193 698905 4 mprj_io_oeb[27]
port 676 nsew
rlabel metal2 s 41713 701977 42193 702033 4 mprj_io_out[27]
port 677 nsew
rlabel metal2 s 41713 711177 42193 711233 4 mprj_io_slow_sel[27]
port 678 nsew
rlabel metal2 s 41713 700137 42193 700193 4 mprj_io_vtrip_sel[27]
port 679 nsew
rlabel metal2 s 41713 713017 42193 713073 4 mprj_io_in[27]
port 680 nsew
rlabel metal2 s 145091 39706 145143 40000 4 porb_h
port 681 nsew
rlabel metal5 s 136713 7143 144149 18309 4 resetb
port 682 nsew
rlabel metal3 s 141667 38031 141813 39999 4 resetb_core_h
port 683 nsew
rlabel metal5 s 698028 909409 711514 920737 4 vccd1
port 684 nsew
rlabel metal5 s 698402 819640 710924 832180 4 vdda1
port 685 nsew
rlabel metal5 s 576820 1018402 589360 1030924 4 vssa1
port 686 nsew
rlabel metal5 s 698028 461609 711514 472937 4 vssd1
port 687 nsew
rlabel metal5 s 6086 913863 19572 925191 4 vccd2
port 688 nsew
rlabel metal5 s 6675 484220 19197 496760 4 vdda2
port 689 nsew
rlabel metal5 s 6675 828820 19197 841360 4 vssa2
port 690 nsew
rlabel metal5 s 6086 442663 19572 453991 4 vssd2
port 691 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
string GDS_FILE chip_io.gds
string GDS_END 35112252
string GDS_START 34578978
<< end >>
