// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module storage(mgmt_clk, mgmt_ena_ro, VPWR, VGND, mgmt_addr, mgmt_addr_ro, mgmt_ena, mgmt_rdata, mgmt_rdata_ro, mgmt_wdata, mgmt_wen, mgmt_wen_mask);
  input VGND;
  input VPWR;
  wire _NC1;
  wire _NC10;
  wire _NC11;
  wire _NC12;
  wire _NC13;
  wire _NC14;
  wire _NC15;
  wire _NC16;
  wire _NC17;
  wire _NC18;
  wire _NC19;
  wire _NC2;
  wire _NC20;
  wire _NC21;
  wire _NC22;
  wire _NC23;
  wire _NC24;
  wire _NC25;
  wire _NC26;
  wire _NC27;
  wire _NC28;
  wire _NC29;
  wire _NC3;
  wire _NC30;
  wire _NC31;
  wire _NC32;
  wire _NC33;
  wire _NC34;
  wire _NC35;
  wire _NC36;
  wire _NC37;
  wire _NC38;
  wire _NC39;
  wire _NC4;
  wire _NC40;
  wire _NC5;
  wire _NC6;
  wire _NC7;
  wire _NC8;
  wire _NC9;
  input [7:0] mgmt_addr;
  input [7:0] mgmt_addr_ro;
  input mgmt_clk;
  input [1:0] mgmt_ena;
  input mgmt_ena_ro;
  output [63:0] mgmt_rdata;
  output [31:0] mgmt_rdata_ro;
  input [31:0] mgmt_wdata;
  input [1:0] mgmt_wen;
  input [7:0] mgmt_wen_mask;
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[0]  (
    .DIODE(mgmt_addr[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[1]  (
    .DIODE(mgmt_addr[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[2]  (
    .DIODE(mgmt_addr[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[3]  (
    .DIODE(mgmt_addr[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[4]  (
    .DIODE(mgmt_addr[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[5]  (
    .DIODE(mgmt_addr[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[6]  (
    .DIODE(mgmt_addr[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr0[7]  (
    .DIODE(mgmt_addr[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[0]  (
    .DIODE(mgmt_addr_ro[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[1]  (
    .DIODE(mgmt_addr_ro[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[2]  (
    .DIODE(mgmt_addr_ro[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[3]  (
    .DIODE(mgmt_addr_ro[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[4]  (
    .DIODE(mgmt_addr_ro[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[5]  (
    .DIODE(mgmt_addr_ro[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[6]  (
    .DIODE(mgmt_addr_ro[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_addr1[7]  (
    .DIODE(mgmt_addr_ro[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_0_clk0 (
    .DIODE(mgmt_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_0_clk1 (
    .DIODE(mgmt_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_0_csb0 (
    .DIODE(mgmt_ena[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_0_csb1 (
    .DIODE(mgmt_ena_ro),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[0]  (
    .DIODE(mgmt_wdata[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[10]  (
    .DIODE(mgmt_wdata[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[11]  (
    .DIODE(mgmt_wdata[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[12]  (
    .DIODE(mgmt_wdata[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[13]  (
    .DIODE(mgmt_wdata[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[14]  (
    .DIODE(mgmt_wdata[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[15]  (
    .DIODE(mgmt_wdata[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[16]  (
    .DIODE(mgmt_wdata[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[17]  (
    .DIODE(mgmt_wdata[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[18]  (
    .DIODE(mgmt_wdata[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[19]  (
    .DIODE(mgmt_wdata[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[1]  (
    .DIODE(mgmt_wdata[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[20]  (
    .DIODE(mgmt_wdata[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[21]  (
    .DIODE(mgmt_wdata[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[22]  (
    .DIODE(mgmt_wdata[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[23]  (
    .DIODE(mgmt_wdata[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[24]  (
    .DIODE(mgmt_wdata[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[25]  (
    .DIODE(mgmt_wdata[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[26]  (
    .DIODE(mgmt_wdata[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[27]  (
    .DIODE(mgmt_wdata[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[28]  (
    .DIODE(mgmt_wdata[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[29]  (
    .DIODE(mgmt_wdata[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[2]  (
    .DIODE(mgmt_wdata[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[30]  (
    .DIODE(mgmt_wdata[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[31]  (
    .DIODE(mgmt_wdata[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[3]  (
    .DIODE(mgmt_wdata[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[4]  (
    .DIODE(mgmt_wdata[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[5]  (
    .DIODE(mgmt_wdata[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[6]  (
    .DIODE(mgmt_wdata[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[7]  (
    .DIODE(mgmt_wdata[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[8]  (
    .DIODE(mgmt_wdata[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_din0[9]  (
    .DIODE(mgmt_wdata[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_0_web0 (
    .DIODE(mgmt_wen[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_wmask0[0]  (
    .DIODE(mgmt_wen_mask[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_wmask0[1]  (
    .DIODE(mgmt_wen_mask[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_wmask0[2]  (
    .DIODE(mgmt_wen_mask[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_0_wmask0[3]  (
    .DIODE(mgmt_wen_mask[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[0]  (
    .DIODE(mgmt_addr[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[1]  (
    .DIODE(mgmt_addr[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[2]  (
    .DIODE(mgmt_addr[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[3]  (
    .DIODE(mgmt_addr[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[4]  (
    .DIODE(mgmt_addr[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[5]  (
    .DIODE(mgmt_addr[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[6]  (
    .DIODE(mgmt_addr[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_addr0[7]  (
    .DIODE(mgmt_addr[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_1_clk0 (
    .DIODE(mgmt_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_1_csb0 (
    .DIODE(mgmt_ena[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[0]  (
    .DIODE(mgmt_wdata[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[10]  (
    .DIODE(mgmt_wdata[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[11]  (
    .DIODE(mgmt_wdata[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[12]  (
    .DIODE(mgmt_wdata[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[13]  (
    .DIODE(mgmt_wdata[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[14]  (
    .DIODE(mgmt_wdata[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[15]  (
    .DIODE(mgmt_wdata[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[16]  (
    .DIODE(mgmt_wdata[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[17]  (
    .DIODE(mgmt_wdata[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[18]  (
    .DIODE(mgmt_wdata[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[19]  (
    .DIODE(mgmt_wdata[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[1]  (
    .DIODE(mgmt_wdata[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[20]  (
    .DIODE(mgmt_wdata[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[21]  (
    .DIODE(mgmt_wdata[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[22]  (
    .DIODE(mgmt_wdata[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[23]  (
    .DIODE(mgmt_wdata[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[24]  (
    .DIODE(mgmt_wdata[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[25]  (
    .DIODE(mgmt_wdata[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[26]  (
    .DIODE(mgmt_wdata[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[27]  (
    .DIODE(mgmt_wdata[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[28]  (
    .DIODE(mgmt_wdata[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[29]  (
    .DIODE(mgmt_wdata[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[2]  (
    .DIODE(mgmt_wdata[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[30]  (
    .DIODE(mgmt_wdata[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[31]  (
    .DIODE(mgmt_wdata[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[3]  (
    .DIODE(mgmt_wdata[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[4]  (
    .DIODE(mgmt_wdata[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[5]  (
    .DIODE(mgmt_wdata[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[6]  (
    .DIODE(mgmt_wdata[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[7]  (
    .DIODE(mgmt_wdata[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[8]  (
    .DIODE(mgmt_wdata[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_din0[9]  (
    .DIODE(mgmt_wdata[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 ANTENNA_SRAM_1_web0 (
    .DIODE(mgmt_wen[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_wmask0[0]  (
    .DIODE(mgmt_wen_mask[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_wmask0[1]  (
    .DIODE(mgmt_wen_mask[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_wmask0[2]  (
    .DIODE(mgmt_wen_mask[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__diode_2 \ANTENNA_SRAM_1_wmask0[3]  (
    .DIODE(mgmt_wen_mask[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_19 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_916 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_928 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_100_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_100_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_100_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_100_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_100_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_100_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_101_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_101_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_101_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_102_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_102_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_102_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_102_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_102_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_102_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_103_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_103_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_103_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_104_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_104_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_104_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_104_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_104_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_104_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_105_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_105_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_105_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_106_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_106_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_106_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_106_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_106_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_106_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_107_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_107_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_107_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_108_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_108_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_108_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_108_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_108_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_108_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_109_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_109_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_109_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_10_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_10_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_10_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_110_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_110_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_110_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_110_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_110_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_110_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_111_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_111_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_111_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_112_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_112_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_112_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_112_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_112_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_112_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_113_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_113_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_113_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_114_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_114_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_114_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_114_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_114_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_114_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_115_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_115_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_115_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_116_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_116_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_116_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_116_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_116_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_116_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_117_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_117_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_117_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_118_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_118_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_118_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_118_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_118_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_118_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_119_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_119_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_119_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_11_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_11_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_120_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_120_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_120_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_120_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_120_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_120_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_121_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_121_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_121_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_122_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_122_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_122_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_122_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_122_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_122_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_123_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_123_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_123_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_124_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_124_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_124_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_124_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_124_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_124_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_125_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_125_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_125_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_126_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_126_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_126_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_126_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_126_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_126_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_127_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_127_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_127_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_128_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_128_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_128_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_128_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_128_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_128_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_129_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_129_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_129_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_12_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_130_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_130_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_130_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_130_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_130_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_130_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_131_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_131_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_131_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_132_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_132_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_132_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_132_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_132_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_132_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_133_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_133_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_133_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_134_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_134_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_134_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_134_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_134_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_134_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_135_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_135_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_135_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_136_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_136_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_136_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_136_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_136_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_136_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_137_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_137_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_137_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_138_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_138_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_138_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_138_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_138_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_138_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_139_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_139_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_139_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_140_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_140_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_140_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_140_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_140_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_140_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_141_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_141_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_141_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_142_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_142_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_142_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_142_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_142_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_142_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_143_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_143_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_143_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_143_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_143_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_144_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_144_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_144_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_144_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_144_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_144_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_145_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_145_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_145_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_146_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_146_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_146_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_146_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_146_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_146_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_147_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_147_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_147_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_147_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_147_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_148_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_148_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_148_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_148_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_148_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_148_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_149_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_149_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_149_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_149_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_149_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_14_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_150_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_150_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_150_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_150_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_150_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_150_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_151_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_151_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_151_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_152_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_152_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_152_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_152_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_152_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_152_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_153_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_153_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_153_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_154_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_154_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_154_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_154_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_154_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_154_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_155_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_155_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_155_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_156_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_156_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_156_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_156_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_156_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_156_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_157_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_157_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_157_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_157_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_157_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_158_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_158_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_158_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_158_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_158_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_158_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_159_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_159_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_159_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_159_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_159_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_160_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_160_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_160_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_160_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_160_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_160_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_161_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_161_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_161_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_162_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_162_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_162_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_162_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_162_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_162_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_163_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_163_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_163_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_164_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_164_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_164_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_164_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_164_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_164_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_165_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_165_936 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_165_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_166_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_166_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_166_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_166_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_166_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_166_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_167_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_167_936 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_167_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_168_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_168_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_168_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_168_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_168_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_168_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_169_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_169_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_169_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_16_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_16_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_170_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_170_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_170_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_170_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_170_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_170_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_171_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_171_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_171_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_171_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_171_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_172_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_172_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_172_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_172_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_172_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_172_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_172_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_172_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_173_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_173_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_173_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_173_31 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_173_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_173_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_173_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_916 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_173_928 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_173_940 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_173_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_11 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_19 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_174_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_174_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_174_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_916 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_174_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_174_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_19 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_31 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_175_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_916 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_175_928 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_175_940 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_175_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_176_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_176_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_176_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_176_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_176_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_176_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_176_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_176_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_177_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_177_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_177_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_177_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_177_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_178_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_178_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_178_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_178_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_178_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_178_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_179_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_179_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_179_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_17_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_180_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_180_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_180_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_180_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_180_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_180_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_181_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_181_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_181_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_182_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_182_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_182_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_182_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_182_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_182_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_183_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_183_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_183_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_184_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_184_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_184_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_184_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_184_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_184_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_185_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_185_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_185_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_186_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_186_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_186_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_186_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_186_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_186_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_187_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_187_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_187_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_188_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_188_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_188_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_188_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_188_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_188_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_189_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_189_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_189_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_18_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_18_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_190_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_190_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_190_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_190_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_190_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_190_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_191_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_191_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_191_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_192_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_192_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_192_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_192_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_192_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_192_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_193_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_193_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_193_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_194_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_194_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_194_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_194_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_194_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_194_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_195_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_195_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_195_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_196_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_196_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_196_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_196_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_196_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_196_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_197_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_197_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_197_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_198_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_198_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_198_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_198_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_198_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_198_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_199_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_199_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_199_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_11 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_19 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_31 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_7 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_916 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_936 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_200_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_200_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_200_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_200_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_200_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_200_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_201_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_201_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_201_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_202_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_202_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_202_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_202_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_202_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_202_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_203_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_203_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_203_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_204_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_204_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_204_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_204_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_204_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_204_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_205_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_205_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_205_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_206_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_206_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_206_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_206_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_206_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_206_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_207_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_207_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_207_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_207_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_207_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_208_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_208_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_208_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_208_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_208_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_208_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_209_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_209_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_209_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_20_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_20_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_20_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_20_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_20_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_210_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_210_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_210_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_210_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_210_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_210_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_211_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_211_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_211_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_212_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_212_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_212_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_212_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_212_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_212_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_212_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_212_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_212_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_212_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_213_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_213_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_213_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_213_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_213_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_213_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_213_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_213_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_214_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_214_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_214_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_214_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_214_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_214_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_214_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_214_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_214_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_214_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_215_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_215_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_215_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_215_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_215_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_215_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_215_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_215_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_216_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_216_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_216_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_216_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_216_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_216_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_216_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_216_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_216_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_216_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_217_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_217_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_217_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_217_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_217_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_217_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_217_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_217_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_218_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_218_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_218_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_218_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_218_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_218_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_218_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_218_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_218_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_218_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_219_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_219_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_219_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_219_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_219_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_219_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_219_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_219_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_21_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_21_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_21_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_220_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_220_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_220_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_220_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_220_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_220_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_220_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_220_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_220_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_220_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_221_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_221_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_221_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_221_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_221_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_221_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_221_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_221_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_222_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_222_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_222_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_222_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_222_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_222_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_222_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_222_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_222_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_222_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_223_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_223_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_223_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_223_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_223_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_223_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_223_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_223_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_224_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_224_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_224_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_224_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_224_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_224_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_224_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_224_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_224_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_224_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_225_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_225_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_225_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_225_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_225_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_225_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_225_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_225_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_226_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_226_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_226_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_226_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_226_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_226_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_226_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_226_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_226_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_226_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_227_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_227_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_227_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_227_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_227_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_227_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_227_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_227_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_228_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_228_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_228_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_228_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_228_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_228_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_228_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_228_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_228_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_228_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_229_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_229_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_229_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_229_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_229_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_229_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_229_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_229_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_22_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_22_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_22_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_22_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_22_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_230_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_230_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_230_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_230_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_230_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_230_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_230_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_230_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_230_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_230_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_231_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_231_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_231_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_231_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_231_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_231_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_231_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_231_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_232_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_232_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_232_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_232_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_232_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_232_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_232_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_232_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_232_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_232_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_233_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_233_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_233_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_233_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_233_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_233_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_233_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_233_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_234_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_234_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_234_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_234_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_234_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_234_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_234_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_234_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_234_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_234_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_235_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_235_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_235_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_235_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_235_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_235_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_235_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_235_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_236_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_236_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_236_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_236_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_236_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_236_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_236_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_236_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_236_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_236_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_237_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_237_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_237_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_237_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_237_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_237_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_237_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_237_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_238_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_238_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_238_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_238_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_238_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_238_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_238_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_238_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_238_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_238_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_239_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_239_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_239_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_239_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_239_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_239_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_239_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_239_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_23_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_23_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_23_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_240_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_240_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_240_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_240_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_240_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_240_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_240_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_240_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_240_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_240_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_241_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_241_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_241_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_241_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_241_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_241_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_241_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_241_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_242_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_242_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_242_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_242_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_242_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_242_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_242_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_242_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_242_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_242_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_243_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_243_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_243_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_243_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_243_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_243_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_243_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_243_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_244_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_244_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_244_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_244_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_244_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_244_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_244_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_244_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_244_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_244_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_245_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_245_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_245_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_245_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_245_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_245_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_245_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_245_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_246_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_246_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_246_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_246_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_246_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_246_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_246_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_246_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_246_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_246_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_247_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_247_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_247_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_247_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_247_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_247_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_247_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_247_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_248_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_248_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_248_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_248_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_248_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_248_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_248_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_248_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_248_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_248_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_249_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_249_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_249_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_249_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_249_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_249_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_249_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_249_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_24_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_24_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_24_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_24_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_24_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_250_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_250_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_250_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_250_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_250_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_250_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_250_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_250_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_250_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_250_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_251_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_251_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_251_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_251_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_251_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_251_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_251_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_251_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_252_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_252_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_252_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_252_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_252_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_252_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_252_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_252_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_252_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_252_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_253_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_253_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_253_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_253_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_253_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_253_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_253_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_253_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_254_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_254_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_254_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_254_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_254_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_254_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_254_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_254_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_254_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_254_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_255_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_255_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_255_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_255_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_255_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_255_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_255_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_255_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_256_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_256_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_256_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_256_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_256_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_256_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_256_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_256_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_256_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_256_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_257_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_257_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_257_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_257_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_257_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_257_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_257_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_257_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_258_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_258_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_258_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_258_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_258_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_258_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_258_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_258_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_258_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_258_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_259_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_259_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_259_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_259_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_259_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_259_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_259_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_259_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_25_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_25_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_25_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_260_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_260_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_260_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_260_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_260_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_260_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_260_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_260_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_260_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_260_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_261_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_261_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_261_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_261_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_261_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_261_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_261_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_261_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_262_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_262_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_262_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_262_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_262_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_262_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_262_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_262_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_262_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_262_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_263_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_263_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_263_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_263_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_263_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_263_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_263_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_263_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_264_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_264_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_264_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_264_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_264_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_264_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_264_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_264_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_264_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_264_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_265_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_265_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_265_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_265_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_265_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_265_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_265_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_265_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_266_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_266_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_266_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_266_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_266_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_266_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_266_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_266_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_266_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_266_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_267_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_267_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_267_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_267_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_267_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_267_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_267_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_267_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_268_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_268_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_268_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_268_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_268_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_268_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_268_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_268_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_268_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_268_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_269_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_269_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_269_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_269_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_269_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_269_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_269_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_269_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_26_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_26_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_26_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_26_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_26_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_270_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_270_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_270_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_270_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_270_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_270_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_270_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_270_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_270_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_270_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_271_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_271_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_271_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_271_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_271_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_271_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_271_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_271_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_272_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_272_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_272_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_272_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_272_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_272_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_272_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_272_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_272_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_272_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_273_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_273_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_273_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_273_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_273_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_273_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_273_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_273_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_274_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_274_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_274_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_274_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_274_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_274_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_274_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_274_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_274_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_274_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_275_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_275_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_275_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_275_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_275_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_275_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_275_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_275_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_276_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_276_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_276_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_276_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_276_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_276_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_276_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_276_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_276_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_276_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_277_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_277_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_277_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_277_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_277_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_277_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_277_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_277_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_278_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_278_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_278_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_278_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_278_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_278_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_278_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_278_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_278_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_278_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_279_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_279_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_279_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_279_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_279_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_279_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_279_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_279_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_27_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_27_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_27_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_280_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_280_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_280_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_280_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_280_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_280_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_280_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_280_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_280_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_280_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_281_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_281_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_281_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_281_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_281_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_281_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_281_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_281_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_282_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_282_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_282_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_282_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_282_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_282_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_282_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_282_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_282_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_282_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_283_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_283_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_283_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_283_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_283_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_283_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_283_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_283_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_284_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_284_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_284_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_284_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_284_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_284_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_284_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_284_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_284_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_284_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_285_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_285_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_285_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_285_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_285_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_285_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_285_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_285_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_286_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_286_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_286_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_286_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_286_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_286_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_286_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_286_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_286_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_286_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_287_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_287_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_287_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_287_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_287_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_287_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_287_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_287_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_288_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_288_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_288_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_288_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_288_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_288_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_288_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_288_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_288_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_288_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_289_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_289_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_289_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_289_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_289_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_289_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_289_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_289_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_28_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_28_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_28_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_28_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_28_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_28_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_290_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_290_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_290_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_290_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_290_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_290_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_290_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_290_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_290_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_290_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_291_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_291_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_291_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_291_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_291_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_291_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_291_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_291_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_292_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_292_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_292_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_292_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_292_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_292_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_292_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_292_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_292_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_292_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_293_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_293_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_293_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_293_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_293_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_293_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_293_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_293_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_294_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_294_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_294_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_294_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_294_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_294_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_294_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_294_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_294_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_294_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_295_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_295_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_295_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_295_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_295_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_295_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_295_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_295_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_296_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_296_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_296_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_296_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_296_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_296_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_296_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_296_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_296_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_296_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_297_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_297_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_297_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_297_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_297_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_297_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_297_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_297_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_298_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_298_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_298_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_298_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_298_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_298_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_298_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_298_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_298_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_298_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_299_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_299_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_299_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_299_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_299_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_299_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_299_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_299_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_29_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_29_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_29_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_11 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_19 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_916 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_300_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_300_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_300_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_300_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_300_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_300_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_300_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_300_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_300_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_300_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_301_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_301_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_301_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_301_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_301_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_301_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_301_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_301_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_302_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_302_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_302_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_302_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_302_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_302_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_302_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_302_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_302_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_302_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_303_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_303_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_303_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_303_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_303_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_303_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_303_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_303_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_304_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_304_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_304_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_304_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_304_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_304_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_304_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_304_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_304_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_304_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_305_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_305_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_305_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_305_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_305_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_305_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_305_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_305_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_306_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_306_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_306_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_306_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_306_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_306_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_306_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_306_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_306_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_306_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_307_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_307_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_307_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_307_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_307_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_307_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_307_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_307_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_308_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_308_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_308_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_308_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_308_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_308_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_308_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_308_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_308_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_308_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_309_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_309_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_309_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_309_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_309_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_309_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_309_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_309_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_30_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_30_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_30_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_30_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_30_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_30_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_310_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_310_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_310_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_310_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_310_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_310_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_310_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_310_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_310_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_310_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_311_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_311_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_311_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_311_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_311_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_311_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_311_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_311_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_312_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_312_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_312_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_312_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_312_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_312_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_312_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_312_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_312_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_312_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_313_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_313_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_313_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_313_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_313_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_313_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_313_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_313_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_314_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_314_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_314_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_314_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_314_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_314_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_314_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_314_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_314_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_314_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_315_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_315_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_315_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_315_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_315_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_315_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_315_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_315_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_316_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_316_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_316_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_316_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_316_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_316_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_316_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_316_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_316_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_316_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_317_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_317_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_317_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_317_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_317_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_317_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_317_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_317_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_318_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_318_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_318_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_318_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_318_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_318_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_318_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_318_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_318_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_318_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_319_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_319_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_319_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_319_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_319_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_319_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_319_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_319_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_319_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_31_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_31_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_31_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_320_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_320_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_320_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_320_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_320_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_320_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_320_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_320_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_320_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_320_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_321_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_321_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_321_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_321_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_321_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_321_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_321_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_321_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_321_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_322_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_322_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_322_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_322_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_322_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_322_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_322_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_322_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_322_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_322_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_323_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_323_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_323_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_323_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_323_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_323_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_323_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_323_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_324_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_324_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_324_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_324_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_324_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_324_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_324_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_324_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_324_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_324_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_325_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_325_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_325_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_325_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_325_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_325_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_325_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_325_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_325_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_326_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_326_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_326_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_326_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_326_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_326_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_326_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_326_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_326_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_326_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_327_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_327_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_327_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_327_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_327_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_327_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_327_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_327_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_327_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_328_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_328_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_328_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_328_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_328_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_328_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_328_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_328_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_328_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_328_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_329_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_329_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_329_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_329_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_329_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_329_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_329_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_329_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_32_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_32_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_32_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_32_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_32_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_32_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_330_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_330_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_330_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_330_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_330_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_330_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_330_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_330_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_330_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_330_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_331_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_331_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_331_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_331_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_331_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_331_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_331_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_331_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_332_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_332_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_332_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_332_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_332_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_332_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_332_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_332_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_332_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_332_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_333_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_333_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_333_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_333_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_333_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_333_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_333_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_333_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_334_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_334_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_334_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_334_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_334_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_334_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_334_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_334_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_334_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_334_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_335_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_335_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_335_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_335_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_335_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_335_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_335_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_335_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_336_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_336_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_336_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_336_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_336_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_336_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_336_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_336_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_336_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_336_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_337_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_337_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_337_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_337_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_337_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_337_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_337_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_337_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_338_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_338_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_338_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_338_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_338_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_338_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_338_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_338_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_338_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_338_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_339_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_339_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_339_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_339_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_339_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_339_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_339_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_339_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_33_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_33_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_33_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_340_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_340_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_340_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_340_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_340_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_340_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_340_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_340_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_340_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_340_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_34_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_34_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_34_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_34_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_34_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_34_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_35_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_35_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_35_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_36_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_36_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_36_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_36_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_36_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_36_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_37_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_37_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_37_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_37_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_37_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_38_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_38_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_38_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_38_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_38_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_38_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_39_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_39_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_39_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_31 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_936 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_40_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_40_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_40_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_40_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_40_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_40_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_41_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_41_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_41_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_42_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_42_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_42_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_42_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_42_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_42_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_43_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_43_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_43_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_44_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_44_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_44_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_44_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_44_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_44_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_45_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_45_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_45_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_46_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_46_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_46_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_46_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_46_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_46_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_47_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_47_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_47_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_48_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_48_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_48_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_48_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_48_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_48_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_49_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_49_936 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_49_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_4_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_50_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_50_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_50_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_50_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_50_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_50_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_51_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_51_936 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 FILLER_51_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_52_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_52_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_52_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_52_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_52_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_52_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_53_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_53_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_53_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_54_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_54_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_54_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_54_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_54_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_54_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_55_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_55_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_55_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_56_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_56_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_56_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_56_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_56_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_56_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_57_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_57_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_57_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_58_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_58_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_58_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_58_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_58_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_58_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_59_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_59_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_59_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_5_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_5_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_60_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_60_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_60_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_60_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_60_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_60_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_61_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_61_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_61_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_62_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_62_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_62_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_62_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_62_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_62_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_63_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_63_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_63_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_64_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_64_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_64_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_64_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_64_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_64_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_65_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_65_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_65_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_66_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_66_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_66_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_66_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_66_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_66_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_67_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_67_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_67_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_68_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_68_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_68_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_68_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_68_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_68_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_69_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_69_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_69_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_70_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_70_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_70_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_70_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_70_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_70_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_71_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_71_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_71_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_72_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_72_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_72_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_72_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_72_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_72_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_73_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_73_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_73_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_74_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_74_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_74_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_74_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_74_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_74_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_75_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_75_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_75_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_76_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_76_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_76_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_76_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_76_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_76_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_77_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_77_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_77_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_78_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_78_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_78_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_78_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_78_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_78_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_79_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_79_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_79_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_7_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_7_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_80_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_80_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_80_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_80_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_80_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_80_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_81_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_81_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_81_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_82_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_82_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_82_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_82_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_82_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_82_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_83_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_83_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_83_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_84_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_84_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_84_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_84_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_84_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_84_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_85_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_85_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_85_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_86_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_86_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_86_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_86_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_86_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_86_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_87_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_87_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_87_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_88_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_88_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_88_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_88_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_88_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_88_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_89_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_89_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_89_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_8_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_90_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_90_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_90_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_90_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_90_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_90_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_91_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_91_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_91_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_92_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_92_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_92_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_92_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_92_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_92_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_93_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_93_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_93_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_94_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_94_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_94_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_94_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_94_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_94_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_95_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_95_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_95_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_96_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_96_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_96_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_96_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_96_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_96_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_97_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_97_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_97_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_98_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_98_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_98_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_4 FILLER_98_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_98_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_2 FILLER_98_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_99_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_99_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_99_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_12 FILLER_9_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_6 FILLER_9_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_10 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_100 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1000 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1001 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1002 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1003 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1004 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1005 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1006 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1007 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1008 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1009 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_101 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1010 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1011 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1012 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1013 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1014 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1015 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1016 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1017 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1018 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1019 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_102 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1020 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1021 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1022 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1023 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1024 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1025 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1026 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1027 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1028 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1029 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_103 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1030 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1031 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1032 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1033 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1034 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1035 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1036 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1037 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1038 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1039 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_104 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1040 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1041 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1042 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1043 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1044 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1045 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1046 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1047 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1048 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1049 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_105 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1050 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1051 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1052 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1053 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1054 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1055 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1056 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1057 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1058 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1059 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_106 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1060 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1061 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1062 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1063 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1064 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1065 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1066 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1067 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1068 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1069 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_107 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1070 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1071 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1072 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1073 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1074 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1075 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1076 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1077 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1078 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1079 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_108 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1080 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1081 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1082 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1083 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1084 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1085 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1086 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1087 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1088 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1089 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_109 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1090 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1091 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1092 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1093 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1094 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1095 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1096 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1097 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1098 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1099 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_11 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_110 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1100 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1101 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1102 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1103 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1104 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1105 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1106 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1107 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1108 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1109 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_111 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1110 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1111 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1112 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1113 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1114 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1115 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1116 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1117 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1118 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1119 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_112 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1120 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1121 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1122 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1123 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1124 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1125 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1126 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1127 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1128 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1129 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_113 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1130 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1131 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1132 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1133 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1134 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1135 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1136 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1137 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1138 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1139 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_114 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1140 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1141 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1142 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1143 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1144 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1145 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1146 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1147 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1148 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1149 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_115 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1150 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1151 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1152 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1153 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1154 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1155 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1156 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1157 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1158 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1159 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_116 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1160 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1161 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1162 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1163 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1164 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1165 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1166 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1167 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1168 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1169 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_117 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1170 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1171 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1172 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1173 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1174 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1175 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1176 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1177 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1178 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1179 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_118 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1180 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1181 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1182 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1183 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1184 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1185 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1186 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1187 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1188 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1189 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_119 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1190 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1191 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1192 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1193 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1194 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1195 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1196 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1197 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1198 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1199 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_12 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_120 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1200 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1201 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1202 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1203 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1204 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1205 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1206 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1207 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1208 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1209 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_121 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1210 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1211 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1212 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1213 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1214 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1215 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1216 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1217 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1218 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1219 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_122 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1220 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1221 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1222 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1223 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1224 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1225 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1226 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1227 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1228 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1229 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_123 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1230 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1231 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1232 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1233 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1234 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1235 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1236 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1237 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1238 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1239 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_124 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1240 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1241 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1242 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1243 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1244 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1245 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1246 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1247 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1248 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1249 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_125 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1250 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1251 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1252 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1253 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1254 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1255 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1256 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1257 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1258 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1259 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_126 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1260 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1261 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1262 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1263 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1264 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1265 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1266 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1267 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1268 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1269 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_127 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1270 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1271 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1272 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1273 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1274 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1275 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1276 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1277 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1278 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1279 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_128 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1280 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1281 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1282 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1283 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1284 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1285 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1286 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1287 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1288 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1289 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_129 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1290 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1291 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1292 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1293 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1294 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1295 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1296 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1297 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1298 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1299 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_13 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_130 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1300 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1301 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1302 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1303 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1304 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1305 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1306 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1307 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1308 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1309 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_131 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1310 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1311 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1312 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1313 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1314 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1315 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1316 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1317 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1318 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1319 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_132 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1320 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1321 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1322 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1323 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1324 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1325 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1326 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1327 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1328 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1329 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_133 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1330 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1331 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1332 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1333 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1334 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1335 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1336 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1337 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1338 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1339 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_134 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1340 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1341 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1342 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1343 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1344 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1345 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1346 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1347 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1348 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1349 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_135 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1350 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1351 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1352 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1353 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1354 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1355 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1356 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1357 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1358 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1359 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_136 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1360 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1361 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1362 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_1363 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_137 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_138 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_139 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_14 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_140 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_141 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_142 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_143 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_144 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_145 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_146 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_147 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_148 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_149 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_15 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_150 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_151 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_152 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_153 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_154 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_155 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_156 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_157 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_158 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_159 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_16 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_160 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_161 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_162 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_163 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_164 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_165 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_166 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_167 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_168 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_169 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_17 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_170 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 (
    .VGND(VGND),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_171 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_172 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_173 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_174 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_175 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_176 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_177 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_178 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_179 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_18 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_180 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_181 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_182 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_183 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_184 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_185 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_186 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_187 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_188 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_189 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_19 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_190 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_191 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_192 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_193 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_194 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_195 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_196 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_197 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_198 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_199 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_20 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_200 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_201 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_202 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_203 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_204 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_205 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_206 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_207 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_208 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_209 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_21 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_210 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_211 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_212 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_213 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_214 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_215 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_216 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_217 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_218 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_219 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_22 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_220 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_221 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_222 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_223 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_224 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_225 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_226 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_227 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_228 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_229 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_23 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_230 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_231 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_232 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_233 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_234 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_235 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_236 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_237 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_238 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_239 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_24 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_240 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_241 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_242 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_243 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_244 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_245 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_246 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_247 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_248 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_249 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_25 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_250 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_251 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_252 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_253 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_254 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_255 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_256 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_257 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_258 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_259 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_26 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_260 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_261 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_262 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_263 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_264 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_265 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_266 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_267 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_268 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_269 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_27 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_270 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_271 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_272 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_273 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_274 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_275 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_276 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_277 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_278 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_279 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_28 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_280 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_281 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_282 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_283 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_284 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_285 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_286 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_287 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_288 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_289 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_29 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_290 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_291 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_292 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_293 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_294 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_295 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_296 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_297 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_298 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_299 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_30 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_300 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_301 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_302 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_303 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_304 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_305 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_306 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_307 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_308 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_309 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_31 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_310 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_311 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_312 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_313 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_314 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_315 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_316 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_317 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_318 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_319 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_32 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_320 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_321 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_322 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_323 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_324 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_325 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_326 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_327 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_328 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_329 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_33 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_330 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_331 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_332 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_333 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_334 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_335 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_336 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_337 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_338 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_339 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_34 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_340 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_341 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_342 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_343 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_344 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_345 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_346 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_347 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_348 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_349 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_35 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_350 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_351 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_352 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_353 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_354 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_355 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_356 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_357 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_358 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_359 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_36 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_360 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_361 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_362 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_363 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_364 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_365 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_366 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_367 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_368 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_369 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_37 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_370 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_371 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_372 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_373 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_374 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_375 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_376 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_377 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_378 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_379 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_38 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_380 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_381 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_382 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_383 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_384 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_385 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_386 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_387 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_388 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_389 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_39 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_390 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_391 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_392 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_393 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_394 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_395 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_396 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_397 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_398 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_399 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_40 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_400 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_401 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_402 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_403 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_404 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_405 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_406 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_407 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_408 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_409 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_41 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_410 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_411 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_412 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_413 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_414 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_415 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_416 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_417 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_418 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_419 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_42 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_420 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_421 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_422 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_423 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_424 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_425 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_426 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_427 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_428 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_429 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_43 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_430 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_431 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_432 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_433 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_434 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_435 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_436 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_437 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_438 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_439 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_44 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_440 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_441 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_442 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_443 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_444 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_445 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_446 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_447 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_448 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_449 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_45 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_450 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_451 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_452 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_453 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_454 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_455 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_456 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_457 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_458 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_459 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_46 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_460 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_461 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_462 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_463 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_464 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_465 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_466 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_467 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_468 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_469 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_47 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_470 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_471 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_472 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_473 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_474 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_475 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_476 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_477 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_478 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_479 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_48 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_480 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_481 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_482 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_483 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_484 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_485 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_486 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_487 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_488 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_489 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_49 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_490 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_491 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_492 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_493 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_494 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_495 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_496 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_497 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_498 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_499 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_50 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_500 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_501 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_502 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_503 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_504 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_505 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_506 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_507 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_508 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_509 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_51 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_510 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_511 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_512 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_513 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_514 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_515 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_516 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_517 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_518 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_519 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_52 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_520 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_521 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_522 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_523 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_524 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_525 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_526 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_527 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_528 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_529 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_53 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_530 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_531 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_532 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_533 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_534 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_535 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_536 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_537 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_538 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_539 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_54 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_540 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_541 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_542 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_543 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_544 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_545 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_546 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_547 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_548 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_549 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_55 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_550 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_551 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_552 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_553 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_554 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_555 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_556 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_557 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_558 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_559 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_56 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_560 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_561 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_562 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_563 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_564 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_565 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_566 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_567 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_568 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_569 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_57 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_570 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_571 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_572 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_573 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_574 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_575 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_576 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_577 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_578 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_579 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_58 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_580 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_581 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_582 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_583 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_584 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_585 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_586 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_587 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_588 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_589 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_59 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_590 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_591 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_592 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_593 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_594 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_595 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_596 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_597 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_598 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_599 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_60 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_600 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_601 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_602 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_603 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_604 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_605 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_606 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_607 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_608 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_609 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_61 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_610 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_611 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_612 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_613 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_614 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_615 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_616 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_617 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_618 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_619 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_62 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_620 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_621 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_622 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_623 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_624 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_625 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_626 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_627 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_628 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_629 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_63 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_630 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_631 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_632 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_633 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_634 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_635 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_636 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_637 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_638 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_639 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_64 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_640 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_641 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_642 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_643 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_644 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_645 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_646 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_647 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_648 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_649 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_65 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_650 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_651 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_652 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_653 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_654 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_655 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_656 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_657 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_658 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_659 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_66 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_660 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_661 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_662 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_663 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_664 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_665 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_666 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_667 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_668 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_669 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_67 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_670 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_671 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_672 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_673 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_674 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_675 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_676 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_677 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_678 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_679 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_68 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_680 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_681 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_682 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_683 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_684 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_685 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_686 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_687 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_688 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_689 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_69 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_690 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_691 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_692 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_693 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_694 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_695 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_696 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_697 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_698 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_699 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_70 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_700 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_701 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_702 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_703 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_704 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_705 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_706 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_707 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_708 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_709 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_71 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_710 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_711 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_712 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_713 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_714 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_715 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_716 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_717 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_718 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_719 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_72 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_720 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_721 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_722 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_723 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_724 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_725 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_726 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_727 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_728 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_729 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_73 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_730 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_731 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_732 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_733 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_734 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_735 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_736 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_737 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_738 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_739 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_74 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_740 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_741 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_742 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_743 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_744 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_745 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_746 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_747 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_748 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_749 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_75 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_750 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_751 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_752 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_753 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_754 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_755 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_756 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_757 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_758 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_759 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_76 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_760 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_761 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_762 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_763 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_764 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_765 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_766 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_767 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_768 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_769 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_77 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_770 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_771 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_772 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_773 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_774 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_775 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_776 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_777 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_778 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_779 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_78 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_780 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_781 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_782 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_783 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_784 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_785 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_786 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_787 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_788 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_789 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_79 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_790 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_791 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_792 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_793 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_794 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_795 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_796 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_797 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_798 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_799 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_8 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_80 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_800 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_801 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_802 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_803 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_804 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_805 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_806 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_807 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_808 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_809 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_81 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_810 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_811 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_812 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_813 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_814 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_815 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_816 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_817 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_818 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_819 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_82 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_820 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_821 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_822 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_823 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_824 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_825 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_826 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_827 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_828 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_829 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_83 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_830 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_831 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_832 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_833 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_834 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_835 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_836 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_837 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_838 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_839 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_84 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_840 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_841 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_842 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_843 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_844 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_845 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_846 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_847 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_848 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_849 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_85 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_850 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_851 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_852 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_853 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_854 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_855 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_856 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_857 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_858 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_859 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_86 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_860 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_861 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_862 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_863 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_864 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_865 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_866 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_867 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_868 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_869 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_87 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_870 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_871 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_872 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_873 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_874 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_875 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_876 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_877 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_878 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_879 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_88 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_880 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_881 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_882 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_883 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_884 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_885 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_886 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_887 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_888 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_889 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_89 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_890 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_891 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_892 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_893 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_894 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_895 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_896 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_897 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_898 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_899 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_9 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_90 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_900 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_901 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_902 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_903 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_904 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_905 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_906 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_907 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_908 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_909 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_91 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_910 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_911 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_912 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_913 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_914 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_915 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_916 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_917 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_918 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_919 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_92 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_920 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_921 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_922 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_923 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_924 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_925 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_926 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_927 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_928 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_929 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_93 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_930 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_931 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_932 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_933 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_934 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_935 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_936 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_937 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_938 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_939 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_94 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_940 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_941 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_942 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_943 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_944 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_945 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_946 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_947 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_948 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_949 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_95 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_950 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_951 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_952 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_953 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_954 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_955 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_956 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_957 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_958 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_959 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_96 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_960 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_961 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_962 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_963 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_964 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_965 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_966 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_967 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_968 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_969 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_97 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_970 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_971 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_972 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_973 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_974 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_975 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_976 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_977 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_978 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_979 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_98 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_980 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_981 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_982 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_983 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_984 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_985 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_986 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_987 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_988 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_989 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_99 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_990 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_991 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_992 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_993 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_994 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_995 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_996 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_997 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_998 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sky130_fd_sc_hd__decap_3 PHY_999 (
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR)
  );
  sram_1rw1r_32_256_8_sky130 SRAM_0 (
    .addr0(mgmt_addr),
    .addr1(mgmt_addr_ro),
    .clk0(mgmt_clk),
    .clk1(mgmt_clk),
    .csb0(mgmt_ena[0]),
    .csb1(mgmt_ena_ro),
    .din0(mgmt_wdata),
    .dout0(mgmt_rdata[31:0]),
    .dout1(mgmt_rdata_ro),
    .gnd(VGND),
    .vdd(VPWR),
    .web0(mgmt_wen[0]),
    .wmask0(mgmt_wen_mask[3:0])
  );
  sram_1rw1r_32_256_8_sky130 SRAM_1 (
    .addr0(mgmt_addr),
    .addr1({ _NC1, _NC2, _NC3, _NC4, _NC5, _NC6, _NC7, _NC8 }),
    .clk0(mgmt_clk),
    .csb0(mgmt_ena[1]),
    .din0(mgmt_wdata),
    .dout0(mgmt_rdata[63:32]),
    .dout1({ _NC9, _NC10, _NC11, _NC12, _NC13, _NC14, _NC15, _NC16, _NC17, _NC18, _NC19, _NC20, _NC21, _NC22, _NC23, _NC24, _NC25, _NC26, _NC27, _NC28, _NC29, _NC30, _NC31, _NC32, _NC33, _NC34, _NC35, _NC36, _NC37, _NC38, _NC39, _NC40 }),
    .gnd(VGND),
    .vdd(VPWR),
    .web0(mgmt_wen[1]),
    .wmask0(mgmt_wen_mask[7:4])
  );
endmodule
