VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 598.760 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.860 596.000 2.140 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.640 596.000 159.920 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.280 596.000 175.560 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.920 596.000 191.200 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.020 596.000 207.300 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.660 596.000 222.940 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.300 596.000 238.580 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.400 596.000 254.680 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.040 596.000 270.320 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.680 596.000 285.960 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.780 596.000 302.060 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.500 596.000 17.780 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.420 596.000 317.700 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.060 596.000 333.340 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.700 596.000 348.980 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.800 596.000 365.080 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.440 596.000 380.720 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.080 596.000 396.360 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.180 596.000 412.460 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.820 596.000 428.100 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.460 596.000 443.740 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.560 596.000 459.840 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.140 596.000 33.420 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.200 596.000 475.480 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.840 596.000 491.120 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.940 596.000 507.220 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.580 596.000 522.860 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.220 596.000 538.500 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.320 596.000 554.600 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.960 596.000 570.240 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.600 596.000 585.880 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.780 596.000 49.060 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.880 596.000 65.160 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.520 596.000 80.800 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.160 596.000 96.440 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.260 596.000 112.540 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.900 596.000 128.180 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.540 596.000 143.820 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.920 596.000 7.200 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.700 596.000 164.980 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.340 596.000 180.620 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.440 596.000 196.720 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.080 596.000 212.360 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.720 596.000 228.000 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.820 596.000 244.100 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.460 596.000 259.740 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.100 596.000 275.380 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.200 596.000 291.480 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.840 596.000 307.120 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.560 596.000 22.840 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.480 596.000 322.760 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.580 596.000 338.860 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.220 596.000 354.500 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.860 596.000 370.140 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.960 596.000 386.240 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.600 596.000 401.880 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.240 596.000 417.520 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.880 596.000 433.160 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.980 596.000 449.260 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.620 596.000 464.900 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.660 596.000 38.940 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.260 596.000 480.540 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.360 596.000 496.640 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.000 596.000 512.280 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.640 596.000 527.920 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.740 596.000 544.020 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.380 596.000 559.660 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.020 596.000 575.300 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.120 596.000 591.400 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.300 596.000 54.580 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.940 596.000 70.220 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.040 596.000 86.320 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.680 596.000 101.960 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.320 596.000 117.600 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.960 596.000 133.240 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.060 596.000 149.340 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.980 596.000 12.260 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.220 596.000 170.500 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.860 596.000 186.140 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.500 596.000 201.780 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.140 596.000 217.420 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.240 596.000 233.520 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.880 596.000 249.160 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.520 596.000 264.800 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.620 596.000 280.900 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.260 596.000 296.540 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.900 596.000 312.180 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.080 596.000 28.360 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.000 596.000 328.280 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.640 596.000 343.920 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.280 596.000 359.560 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.380 596.000 375.660 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.020 596.000 391.300 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.660 596.000 406.940 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.760 596.000 423.040 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.400 596.000 438.680 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.040 596.000 454.320 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.140 596.000 470.420 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.720 596.000 44.000 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.780 596.000 486.060 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.420 596.000 501.700 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.060 596.000 517.340 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.160 596.000 533.440 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.800 596.000 549.080 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.440 596.000 564.720 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.540 596.000 580.820 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.180 596.000 596.460 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.360 596.000 59.640 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.460 596.000 75.740 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.100 596.000 91.380 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.740 596.000 107.020 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.840 596.000 123.120 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.480 596.000 138.760 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.120 596.000 154.400 600.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.740 0.000 130.020 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.820 0.000 497.100 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.500 0.000 500.780 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.180 0.000 504.460 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.860 0.000 508.140 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.540 0.000 511.820 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.220 0.000 515.500 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.900 0.000 519.180 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.580 0.000 522.860 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.260 0.000 526.540 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.940 0.000 530.220 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.080 0.000 166.360 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.620 0.000 533.900 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.300 0.000 537.580 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.980 0.000 541.260 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.660 0.000 544.940 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.340 0.000 548.620 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.020 0.000 552.300 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.700 0.000 555.980 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.380 0.000 559.660 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.060 0.000 563.340 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.740 0.000 567.020 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.760 0.000 170.040 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.420 0.000 570.700 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.100 0.000 574.380 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.780 0.000 578.060 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.460 0.000 581.740 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.140 0.000 585.420 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.820 0.000 589.100 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.500 0.000 592.780 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.180 0.000 596.460 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.440 0.000 173.720 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.120 0.000 177.400 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.800 0.000 181.080 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.480 0.000 184.760 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.160 0.000 188.440 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.840 0.000 192.120 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.520 0.000 195.800 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.200 0.000 199.480 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.420 0.000 133.700 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.880 0.000 203.160 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.560 0.000 206.840 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.240 0.000 210.520 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.920 0.000 214.200 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.600 0.000 217.880 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.280 0.000 221.560 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.960 0.000 225.240 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.640 0.000 228.920 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.320 0.000 232.600 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.000 0.000 236.280 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.100 0.000 137.380 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.680 0.000 239.960 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.360 0.000 243.640 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.040 0.000 247.320 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.720 0.000 251.000 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.400 0.000 254.680 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.080 0.000 258.360 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.760 0.000 262.040 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.440 0.000 265.720 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.120 0.000 269.400 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.800 0.000 273.080 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.780 0.000 141.060 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.480 0.000 276.760 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.160 0.000 280.440 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.840 0.000 284.120 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.520 0.000 287.800 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.200 0.000 291.480 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.880 0.000 295.160 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.560 0.000 298.840 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.240 0.000 302.520 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.920 0.000 306.200 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.600 0.000 309.880 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.460 0.000 144.740 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.280 0.000 313.560 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.960 0.000 317.240 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.640 0.000 320.920 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.320 0.000 324.600 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.000 0.000 328.280 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.680 0.000 331.960 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.360 0.000 335.640 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.040 0.000 339.320 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.720 0.000 343.000 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.400 0.000 346.680 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.140 0.000 148.420 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.080 0.000 350.360 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.760 0.000 354.040 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.440 0.000 357.720 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.120 0.000 361.400 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.800 0.000 365.080 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.480 0.000 368.760 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.160 0.000 372.440 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.380 0.000 375.660 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.060 0.000 379.340 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.740 0.000 383.020 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.360 0.000 151.640 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.420 0.000 386.700 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.100 0.000 390.380 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.780 0.000 394.060 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.460 0.000 397.740 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.140 0.000 401.420 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.820 0.000 405.100 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.500 0.000 408.780 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.180 0.000 412.460 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.860 0.000 416.140 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.540 0.000 419.820 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.040 0.000 155.320 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.220 0.000 423.500 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.900 0.000 427.180 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.580 0.000 430.860 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.260 0.000 434.540 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.940 0.000 438.220 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.620 0.000 441.900 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.300 0.000 445.580 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.980 0.000 449.260 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.660 0.000 452.940 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.340 0.000 456.620 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.720 0.000 159.000 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.020 0.000 460.300 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.700 0.000 463.980 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.380 0.000 467.660 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.060 0.000 471.340 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.740 0.000 475.020 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.420 0.000 478.700 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.100 0.000 482.380 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.780 0.000 486.060 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.460 0.000 489.740 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.140 0.000 493.420 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.400 0.000 162.680 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.660 0.000 130.940 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.200 0.000 498.480 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.880 0.000 502.160 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.560 0.000 505.840 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.240 0.000 509.520 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.920 0.000 513.200 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.600 0.000 516.880 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.280 0.000 520.560 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.960 0.000 524.240 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.180 0.000 527.460 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.860 0.000 531.140 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.460 0.000 167.740 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.540 0.000 534.820 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.220 0.000 538.500 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.900 0.000 542.180 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.580 0.000 545.860 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.260 0.000 549.540 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.940 0.000 553.220 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.620 0.000 556.900 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.300 0.000 560.580 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.980 0.000 564.260 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.660 0.000 567.940 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.140 0.000 171.420 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.340 0.000 571.620 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.020 0.000 575.300 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.700 0.000 578.980 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.380 0.000 582.660 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.060 0.000 586.340 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.740 0.000 590.020 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.420 0.000 593.700 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.100 0.000 597.380 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.820 0.000 175.100 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.500 0.000 178.780 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.180 0.000 182.460 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.860 0.000 186.140 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.540 0.000 189.820 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.220 0.000 193.500 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.900 0.000 197.180 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.580 0.000 200.860 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.340 0.000 134.620 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.260 0.000 204.540 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.940 0.000 208.220 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.620 0.000 211.900 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.300 0.000 215.580 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.980 0.000 219.260 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.660 0.000 222.940 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.340 0.000 226.620 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.020 0.000 230.300 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.700 0.000 233.980 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.380 0.000 237.660 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.020 0.000 138.300 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.060 0.000 241.340 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.740 0.000 245.020 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.420 0.000 248.700 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.100 0.000 252.380 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.780 0.000 256.060 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.460 0.000 259.740 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.140 0.000 263.420 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.820 0.000 267.100 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.500 0.000 270.780 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.180 0.000 274.460 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.700 0.000 141.980 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.860 0.000 278.140 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.540 0.000 281.820 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.220 0.000 285.500 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.900 0.000 289.180 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.580 0.000 292.860 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.260 0.000 296.540 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.940 0.000 300.220 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.160 0.000 303.440 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.840 0.000 307.120 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.520 0.000 310.800 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.380 0.000 145.660 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.200 0.000 314.480 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.880 0.000 318.160 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.560 0.000 321.840 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.240 0.000 325.520 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.920 0.000 329.200 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.600 0.000 332.880 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.280 0.000 336.560 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.960 0.000 340.240 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.640 0.000 343.920 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.320 0.000 347.600 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.060 0.000 149.340 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.000 0.000 351.280 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.680 0.000 354.960 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.360 0.000 358.640 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.040 0.000 362.320 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.720 0.000 366.000 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.400 0.000 369.680 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.080 0.000 373.360 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.760 0.000 377.040 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.440 0.000 380.720 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.120 0.000 384.400 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.740 0.000 153.020 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.800 0.000 388.080 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.480 0.000 391.760 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.160 0.000 395.440 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.840 0.000 399.120 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.520 0.000 402.800 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.200 0.000 406.480 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.880 0.000 410.160 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.560 0.000 413.840 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.240 0.000 417.520 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.920 0.000 421.200 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.420 0.000 156.700 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.600 0.000 424.880 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.280 0.000 428.560 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.960 0.000 432.240 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.640 0.000 435.920 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.320 0.000 439.600 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.000 0.000 443.280 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.680 0.000 446.960 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.360 0.000 450.640 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.040 0.000 454.320 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.720 0.000 458.000 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.100 0.000 160.380 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.400 0.000 461.680 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.080 0.000 465.360 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.760 0.000 469.040 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.440 0.000 472.720 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.120 0.000 476.400 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.800 0.000 480.080 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.480 0.000 483.760 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.160 0.000 487.440 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.840 0.000 491.120 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.520 0.000 494.800 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.780 0.000 164.060 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.040 0.000 132.320 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.120 0.000 499.400 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.800 0.000 503.080 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.480 0.000 506.760 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.160 0.000 510.440 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.840 0.000 514.120 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.520 0.000 517.800 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.200 0.000 521.480 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.880 0.000 525.160 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.560 0.000 528.840 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.240 0.000 532.520 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.840 0.000 169.120 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.920 0.000 536.200 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.600 0.000 539.880 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.280 0.000 543.560 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.960 0.000 547.240 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.640 0.000 550.920 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.320 0.000 554.600 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.000 0.000 558.280 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.680 0.000 561.960 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.360 0.000 565.640 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.040 0.000 569.320 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.520 0.000 172.800 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.720 0.000 573.000 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.400 0.000 576.680 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.080 0.000 580.360 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.760 0.000 584.040 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.440 0.000 587.720 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.120 0.000 591.400 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.800 0.000 595.080 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.480 0.000 598.760 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.200 0.000 176.480 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.880 0.000 180.160 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.560 0.000 183.840 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.240 0.000 187.520 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.920 0.000 191.200 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.600 0.000 194.880 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.280 0.000 198.560 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.960 0.000 202.240 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.720 0.000 136.000 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.640 0.000 205.920 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.320 0.000 209.600 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.000 0.000 213.280 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.680 0.000 216.960 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.360 0.000 220.640 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.040 0.000 224.320 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.260 0.000 227.540 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.940 0.000 231.220 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.620 0.000 234.900 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.300 0.000 238.580 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.400 0.000 139.680 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.980 0.000 242.260 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.660 0.000 245.940 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.340 0.000 249.620 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.020 0.000 253.300 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.700 0.000 256.980 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.380 0.000 260.660 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.060 0.000 264.340 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.740 0.000 268.020 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.420 0.000 271.700 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.100 0.000 275.380 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.080 0.000 143.360 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.780 0.000 279.060 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.460 0.000 282.740 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.140 0.000 286.420 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.820 0.000 290.100 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.500 0.000 293.780 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.180 0.000 297.460 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.860 0.000 301.140 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.540 0.000 304.820 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.220 0.000 308.500 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.900 0.000 312.180 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.760 0.000 147.040 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.580 0.000 315.860 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.260 0.000 319.540 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.940 0.000 323.220 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.620 0.000 326.900 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.300 0.000 330.580 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.980 0.000 334.260 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.660 0.000 337.940 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.340 0.000 341.620 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.020 0.000 345.300 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.700 0.000 348.980 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.440 0.000 150.720 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.380 0.000 352.660 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.060 0.000 356.340 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.740 0.000 360.020 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.420 0.000 363.700 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.100 0.000 367.380 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.780 0.000 371.060 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.460 0.000 374.740 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.140 0.000 378.420 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.820 0.000 382.100 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.500 0.000 385.780 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.120 0.000 154.400 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.180 0.000 389.460 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.860 0.000 393.140 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.540 0.000 396.820 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.220 0.000 400.500 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.900 0.000 404.180 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.580 0.000 407.860 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.260 0.000 411.540 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.940 0.000 415.220 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.620 0.000 418.900 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.300 0.000 422.580 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.800 0.000 158.080 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.980 0.000 426.260 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.660 0.000 429.940 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.340 0.000 433.620 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.020 0.000 437.300 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.700 0.000 440.980 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.380 0.000 444.660 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.060 0.000 448.340 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.280 0.000 451.560 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.960 0.000 455.240 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.640 0.000 458.920 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.480 0.000 161.760 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.320 0.000 462.600 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.000 0.000 466.280 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.680 0.000 469.960 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.360 0.000 473.640 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.040 0.000 477.320 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.720 0.000 481.000 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.400 0.000 484.680 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.080 0.000 488.360 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.760 0.000 492.040 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.440 0.000 495.720 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.160 0.000 165.440 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.940 0.000 1.220 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.320 0.000 2.600 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.920 0.000 7.200 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.780 0.000 49.060 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.460 0.000 52.740 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.140 0.000 56.420 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.820 0.000 60.100 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.500 0.000 63.780 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.180 0.000 67.460 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.860 0.000 71.140 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.540 0.000 74.820 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.220 0.000 78.500 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.900 0.000 82.180 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.980 0.000 12.260 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.580 0.000 85.860 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.260 0.000 89.540 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.940 0.000 93.220 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.620 0.000 96.900 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.300 0.000 100.580 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.980 0.000 104.260 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.660 0.000 107.940 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.340 0.000 111.620 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.020 0.000 115.300 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.700 0.000 118.980 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.040 0.000 17.320 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.380 0.000 122.660 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.060 0.000 126.340 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.640 0.000 21.920 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.700 0.000 26.980 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.380 0.000 30.660 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.060 0.000 34.340 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.740 0.000 38.020 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.420 0.000 41.700 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.100 0.000 45.380 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.240 0.000 3.520 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.300 0.000 8.580 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.160 0.000 50.440 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.840 0.000 54.120 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.520 0.000 57.800 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.200 0.000 61.480 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.880 0.000 65.160 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.560 0.000 68.840 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.240 0.000 72.520 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.460 0.000 75.740 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.140 0.000 79.420 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.820 0.000 83.100 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.360 0.000 13.640 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.500 0.000 86.780 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.180 0.000 90.460 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.860 0.000 94.140 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.540 0.000 97.820 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.220 0.000 101.500 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.900 0.000 105.180 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.580 0.000 108.860 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.260 0.000 112.540 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.940 0.000 116.220 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.620 0.000 119.900 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.960 0.000 18.240 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.300 0.000 123.580 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.980 0.000 127.260 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.020 0.000 23.300 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.080 0.000 28.360 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.760 0.000 32.040 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.440 0.000 35.720 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.120 0.000 39.400 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.800 0.000 43.080 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.480 0.000 46.760 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.680 0.000 9.960 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.080 0.000 51.360 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.760 0.000 55.040 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.440 0.000 58.720 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.120 0.000 62.400 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.800 0.000 66.080 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.480 0.000 69.760 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.160 0.000 73.440 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.840 0.000 77.120 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.520 0.000 80.800 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.200 0.000 84.480 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.280 0.000 14.560 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.880 0.000 88.160 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.560 0.000 91.840 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.240 0.000 95.520 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.920 0.000 99.200 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.600 0.000 102.880 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.280 0.000 106.560 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.960 0.000 110.240 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.640 0.000 113.920 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.320 0.000 117.600 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.000 0.000 121.280 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.340 0.000 19.620 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.680 0.000 124.960 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.360 0.000 128.640 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.400 0.000 24.680 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.000 0.000 29.280 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.680 0.000 32.960 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.360 0.000 36.640 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.040 0.000 40.320 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.400 0.000 47.680 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.600 0.000 10.880 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.660 0.000 15.940 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.720 0.000 21.000 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.320 0.000 25.600 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.620 0.000 4.900 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.000 0.000 6.280 4.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.310 10.640 482.910 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 327.710 10.640 329.310 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.110 10.640 175.710 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.510 10.640 22.110 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.110 10.640 559.710 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 404.510 10.640 406.110 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 250.910 10.640 252.510 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.310 10.640 98.910 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 484.610 10.880 486.210 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.010 10.880 332.610 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.410 10.880 179.010 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.810 10.880 25.410 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.410 10.880 563.010 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 407.810 10.880 409.410 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.210 10.880 255.810 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 100.610 10.880 102.210 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 487.910 10.880 489.510 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.310 10.880 335.910 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 180.710 10.880 182.310 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.110 10.880 28.710 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 564.710 10.880 566.310 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.110 10.880 412.710 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 257.510 10.880 259.110 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 103.910 10.880 105.510 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.210 10.880 492.810 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 337.610 10.880 339.210 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.010 10.880 185.610 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.410 10.880 32.010 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.010 10.880 569.610 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.410 10.880 416.010 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 260.810 10.880 262.410 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.210 10.880 108.810 587.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 4.990 6.885 593.790 587.605 ;
      LAYER met1 ;
        RECT 0.000 5.480 597.400 595.640 ;
      LAYER met2 ;
        RECT 0.030 595.720 1.580 596.000 ;
        RECT 2.420 595.720 6.640 596.000 ;
        RECT 7.480 595.720 11.700 596.000 ;
        RECT 12.540 595.720 17.220 596.000 ;
        RECT 18.060 595.720 22.280 596.000 ;
        RECT 23.120 595.720 27.800 596.000 ;
        RECT 28.640 595.720 32.860 596.000 ;
        RECT 33.700 595.720 38.380 596.000 ;
        RECT 39.220 595.720 43.440 596.000 ;
        RECT 44.280 595.720 48.500 596.000 ;
        RECT 49.340 595.720 54.020 596.000 ;
        RECT 54.860 595.720 59.080 596.000 ;
        RECT 59.920 595.720 64.600 596.000 ;
        RECT 65.440 595.720 69.660 596.000 ;
        RECT 70.500 595.720 75.180 596.000 ;
        RECT 76.020 595.720 80.240 596.000 ;
        RECT 81.080 595.720 85.760 596.000 ;
        RECT 86.600 595.720 90.820 596.000 ;
        RECT 91.660 595.720 95.880 596.000 ;
        RECT 96.720 595.720 101.400 596.000 ;
        RECT 102.240 595.720 106.460 596.000 ;
        RECT 107.300 595.720 111.980 596.000 ;
        RECT 112.820 595.720 117.040 596.000 ;
        RECT 117.880 595.720 122.560 596.000 ;
        RECT 123.400 595.720 127.620 596.000 ;
        RECT 128.460 595.720 132.680 596.000 ;
        RECT 133.520 595.720 138.200 596.000 ;
        RECT 139.040 595.720 143.260 596.000 ;
        RECT 144.100 595.720 148.780 596.000 ;
        RECT 149.620 595.720 153.840 596.000 ;
        RECT 154.680 595.720 159.360 596.000 ;
        RECT 160.200 595.720 164.420 596.000 ;
        RECT 165.260 595.720 169.940 596.000 ;
        RECT 170.780 595.720 175.000 596.000 ;
        RECT 175.840 595.720 180.060 596.000 ;
        RECT 180.900 595.720 185.580 596.000 ;
        RECT 186.420 595.720 190.640 596.000 ;
        RECT 191.480 595.720 196.160 596.000 ;
        RECT 197.000 595.720 201.220 596.000 ;
        RECT 202.060 595.720 206.740 596.000 ;
        RECT 207.580 595.720 211.800 596.000 ;
        RECT 212.640 595.720 216.860 596.000 ;
        RECT 217.700 595.720 222.380 596.000 ;
        RECT 223.220 595.720 227.440 596.000 ;
        RECT 228.280 595.720 232.960 596.000 ;
        RECT 233.800 595.720 238.020 596.000 ;
        RECT 238.860 595.720 243.540 596.000 ;
        RECT 244.380 595.720 248.600 596.000 ;
        RECT 249.440 595.720 254.120 596.000 ;
        RECT 254.960 595.720 259.180 596.000 ;
        RECT 260.020 595.720 264.240 596.000 ;
        RECT 265.080 595.720 269.760 596.000 ;
        RECT 270.600 595.720 274.820 596.000 ;
        RECT 275.660 595.720 280.340 596.000 ;
        RECT 281.180 595.720 285.400 596.000 ;
        RECT 286.240 595.720 290.920 596.000 ;
        RECT 291.760 595.720 295.980 596.000 ;
        RECT 296.820 595.720 301.500 596.000 ;
        RECT 302.340 595.720 306.560 596.000 ;
        RECT 307.400 595.720 311.620 596.000 ;
        RECT 312.460 595.720 317.140 596.000 ;
        RECT 317.980 595.720 322.200 596.000 ;
        RECT 323.040 595.720 327.720 596.000 ;
        RECT 328.560 595.720 332.780 596.000 ;
        RECT 333.620 595.720 338.300 596.000 ;
        RECT 339.140 595.720 343.360 596.000 ;
        RECT 344.200 595.720 348.420 596.000 ;
        RECT 349.260 595.720 353.940 596.000 ;
        RECT 354.780 595.720 359.000 596.000 ;
        RECT 359.840 595.720 364.520 596.000 ;
        RECT 365.360 595.720 369.580 596.000 ;
        RECT 370.420 595.720 375.100 596.000 ;
        RECT 375.940 595.720 380.160 596.000 ;
        RECT 381.000 595.720 385.680 596.000 ;
        RECT 386.520 595.720 390.740 596.000 ;
        RECT 391.580 595.720 395.800 596.000 ;
        RECT 396.640 595.720 401.320 596.000 ;
        RECT 402.160 595.720 406.380 596.000 ;
        RECT 407.220 595.720 411.900 596.000 ;
        RECT 412.740 595.720 416.960 596.000 ;
        RECT 417.800 595.720 422.480 596.000 ;
        RECT 423.320 595.720 427.540 596.000 ;
        RECT 428.380 595.720 432.600 596.000 ;
        RECT 433.440 595.720 438.120 596.000 ;
        RECT 438.960 595.720 443.180 596.000 ;
        RECT 444.020 595.720 448.700 596.000 ;
        RECT 449.540 595.720 453.760 596.000 ;
        RECT 454.600 595.720 459.280 596.000 ;
        RECT 460.120 595.720 464.340 596.000 ;
        RECT 465.180 595.720 469.860 596.000 ;
        RECT 470.700 595.720 474.920 596.000 ;
        RECT 475.760 595.720 479.980 596.000 ;
        RECT 480.820 595.720 485.500 596.000 ;
        RECT 486.340 595.720 490.560 596.000 ;
        RECT 491.400 595.720 496.080 596.000 ;
        RECT 496.920 595.720 501.140 596.000 ;
        RECT 501.980 595.720 506.660 596.000 ;
        RECT 507.500 595.720 511.720 596.000 ;
        RECT 512.560 595.720 516.780 596.000 ;
        RECT 517.620 595.720 522.300 596.000 ;
        RECT 523.140 595.720 527.360 596.000 ;
        RECT 528.200 595.720 532.880 596.000 ;
        RECT 533.720 595.720 537.940 596.000 ;
        RECT 538.780 595.720 543.460 596.000 ;
        RECT 544.300 595.720 548.520 596.000 ;
        RECT 549.360 595.720 554.040 596.000 ;
        RECT 554.880 595.720 559.100 596.000 ;
        RECT 559.940 595.720 564.160 596.000 ;
        RECT 565.000 595.720 569.680 596.000 ;
        RECT 570.520 595.720 574.740 596.000 ;
        RECT 575.580 595.720 580.260 596.000 ;
        RECT 581.100 595.720 585.320 596.000 ;
        RECT 586.160 595.720 590.840 596.000 ;
        RECT 591.680 595.720 595.900 596.000 ;
        RECT 596.740 595.720 597.370 596.000 ;
        RECT 0.030 4.280 597.370 595.720 ;
        RECT 0.580 4.000 0.660 4.280 ;
        RECT 1.500 4.000 2.040 4.280 ;
        RECT 2.880 4.000 2.960 4.280 ;
        RECT 3.800 4.000 4.340 4.280 ;
        RECT 5.180 4.000 5.720 4.280 ;
        RECT 6.560 4.000 6.640 4.280 ;
        RECT 7.480 4.000 8.020 4.280 ;
        RECT 8.860 4.000 9.400 4.280 ;
        RECT 10.240 4.000 10.320 4.280 ;
        RECT 11.160 4.000 11.700 4.280 ;
        RECT 12.540 4.000 13.080 4.280 ;
        RECT 13.920 4.000 14.000 4.280 ;
        RECT 14.840 4.000 15.380 4.280 ;
        RECT 16.220 4.000 16.760 4.280 ;
        RECT 17.600 4.000 17.680 4.280 ;
        RECT 18.520 4.000 19.060 4.280 ;
        RECT 19.900 4.000 20.440 4.280 ;
        RECT 21.280 4.000 21.360 4.280 ;
        RECT 22.200 4.000 22.740 4.280 ;
        RECT 23.580 4.000 24.120 4.280 ;
        RECT 24.960 4.000 25.040 4.280 ;
        RECT 25.880 4.000 26.420 4.280 ;
        RECT 27.260 4.000 27.800 4.280 ;
        RECT 28.640 4.000 28.720 4.280 ;
        RECT 29.560 4.000 30.100 4.280 ;
        RECT 30.940 4.000 31.480 4.280 ;
        RECT 32.320 4.000 32.400 4.280 ;
        RECT 33.240 4.000 33.780 4.280 ;
        RECT 34.620 4.000 35.160 4.280 ;
        RECT 36.000 4.000 36.080 4.280 ;
        RECT 36.920 4.000 37.460 4.280 ;
        RECT 38.300 4.000 38.840 4.280 ;
        RECT 39.680 4.000 39.760 4.280 ;
        RECT 40.600 4.000 41.140 4.280 ;
        RECT 41.980 4.000 42.520 4.280 ;
        RECT 43.360 4.000 43.440 4.280 ;
        RECT 44.280 4.000 44.820 4.280 ;
        RECT 45.660 4.000 46.200 4.280 ;
        RECT 47.040 4.000 47.120 4.280 ;
        RECT 47.960 4.000 48.500 4.280 ;
        RECT 49.340 4.000 49.880 4.280 ;
        RECT 50.720 4.000 50.800 4.280 ;
        RECT 51.640 4.000 52.180 4.280 ;
        RECT 53.020 4.000 53.560 4.280 ;
        RECT 54.400 4.000 54.480 4.280 ;
        RECT 55.320 4.000 55.860 4.280 ;
        RECT 56.700 4.000 57.240 4.280 ;
        RECT 58.080 4.000 58.160 4.280 ;
        RECT 59.000 4.000 59.540 4.280 ;
        RECT 60.380 4.000 60.920 4.280 ;
        RECT 61.760 4.000 61.840 4.280 ;
        RECT 62.680 4.000 63.220 4.280 ;
        RECT 64.060 4.000 64.600 4.280 ;
        RECT 65.440 4.000 65.520 4.280 ;
        RECT 66.360 4.000 66.900 4.280 ;
        RECT 67.740 4.000 68.280 4.280 ;
        RECT 69.120 4.000 69.200 4.280 ;
        RECT 70.040 4.000 70.580 4.280 ;
        RECT 71.420 4.000 71.960 4.280 ;
        RECT 72.800 4.000 72.880 4.280 ;
        RECT 73.720 4.000 74.260 4.280 ;
        RECT 75.100 4.000 75.180 4.280 ;
        RECT 76.020 4.000 76.560 4.280 ;
        RECT 77.400 4.000 77.940 4.280 ;
        RECT 78.780 4.000 78.860 4.280 ;
        RECT 79.700 4.000 80.240 4.280 ;
        RECT 81.080 4.000 81.620 4.280 ;
        RECT 82.460 4.000 82.540 4.280 ;
        RECT 83.380 4.000 83.920 4.280 ;
        RECT 84.760 4.000 85.300 4.280 ;
        RECT 86.140 4.000 86.220 4.280 ;
        RECT 87.060 4.000 87.600 4.280 ;
        RECT 88.440 4.000 88.980 4.280 ;
        RECT 89.820 4.000 89.900 4.280 ;
        RECT 90.740 4.000 91.280 4.280 ;
        RECT 92.120 4.000 92.660 4.280 ;
        RECT 93.500 4.000 93.580 4.280 ;
        RECT 94.420 4.000 94.960 4.280 ;
        RECT 95.800 4.000 96.340 4.280 ;
        RECT 97.180 4.000 97.260 4.280 ;
        RECT 98.100 4.000 98.640 4.280 ;
        RECT 99.480 4.000 100.020 4.280 ;
        RECT 100.860 4.000 100.940 4.280 ;
        RECT 101.780 4.000 102.320 4.280 ;
        RECT 103.160 4.000 103.700 4.280 ;
        RECT 104.540 4.000 104.620 4.280 ;
        RECT 105.460 4.000 106.000 4.280 ;
        RECT 106.840 4.000 107.380 4.280 ;
        RECT 108.220 4.000 108.300 4.280 ;
        RECT 109.140 4.000 109.680 4.280 ;
        RECT 110.520 4.000 111.060 4.280 ;
        RECT 111.900 4.000 111.980 4.280 ;
        RECT 112.820 4.000 113.360 4.280 ;
        RECT 114.200 4.000 114.740 4.280 ;
        RECT 115.580 4.000 115.660 4.280 ;
        RECT 116.500 4.000 117.040 4.280 ;
        RECT 117.880 4.000 118.420 4.280 ;
        RECT 119.260 4.000 119.340 4.280 ;
        RECT 120.180 4.000 120.720 4.280 ;
        RECT 121.560 4.000 122.100 4.280 ;
        RECT 122.940 4.000 123.020 4.280 ;
        RECT 123.860 4.000 124.400 4.280 ;
        RECT 125.240 4.000 125.780 4.280 ;
        RECT 126.620 4.000 126.700 4.280 ;
        RECT 127.540 4.000 128.080 4.280 ;
        RECT 128.920 4.000 129.460 4.280 ;
        RECT 130.300 4.000 130.380 4.280 ;
        RECT 131.220 4.000 131.760 4.280 ;
        RECT 132.600 4.000 133.140 4.280 ;
        RECT 133.980 4.000 134.060 4.280 ;
        RECT 134.900 4.000 135.440 4.280 ;
        RECT 136.280 4.000 136.820 4.280 ;
        RECT 137.660 4.000 137.740 4.280 ;
        RECT 138.580 4.000 139.120 4.280 ;
        RECT 139.960 4.000 140.500 4.280 ;
        RECT 141.340 4.000 141.420 4.280 ;
        RECT 142.260 4.000 142.800 4.280 ;
        RECT 143.640 4.000 144.180 4.280 ;
        RECT 145.020 4.000 145.100 4.280 ;
        RECT 145.940 4.000 146.480 4.280 ;
        RECT 147.320 4.000 147.860 4.280 ;
        RECT 148.700 4.000 148.780 4.280 ;
        RECT 149.620 4.000 150.160 4.280 ;
        RECT 151.000 4.000 151.080 4.280 ;
        RECT 151.920 4.000 152.460 4.280 ;
        RECT 153.300 4.000 153.840 4.280 ;
        RECT 154.680 4.000 154.760 4.280 ;
        RECT 155.600 4.000 156.140 4.280 ;
        RECT 156.980 4.000 157.520 4.280 ;
        RECT 158.360 4.000 158.440 4.280 ;
        RECT 159.280 4.000 159.820 4.280 ;
        RECT 160.660 4.000 161.200 4.280 ;
        RECT 162.040 4.000 162.120 4.280 ;
        RECT 162.960 4.000 163.500 4.280 ;
        RECT 164.340 4.000 164.880 4.280 ;
        RECT 165.720 4.000 165.800 4.280 ;
        RECT 166.640 4.000 167.180 4.280 ;
        RECT 168.020 4.000 168.560 4.280 ;
        RECT 169.400 4.000 169.480 4.280 ;
        RECT 170.320 4.000 170.860 4.280 ;
        RECT 171.700 4.000 172.240 4.280 ;
        RECT 173.080 4.000 173.160 4.280 ;
        RECT 174.000 4.000 174.540 4.280 ;
        RECT 175.380 4.000 175.920 4.280 ;
        RECT 176.760 4.000 176.840 4.280 ;
        RECT 177.680 4.000 178.220 4.280 ;
        RECT 179.060 4.000 179.600 4.280 ;
        RECT 180.440 4.000 180.520 4.280 ;
        RECT 181.360 4.000 181.900 4.280 ;
        RECT 182.740 4.000 183.280 4.280 ;
        RECT 184.120 4.000 184.200 4.280 ;
        RECT 185.040 4.000 185.580 4.280 ;
        RECT 186.420 4.000 186.960 4.280 ;
        RECT 187.800 4.000 187.880 4.280 ;
        RECT 188.720 4.000 189.260 4.280 ;
        RECT 190.100 4.000 190.640 4.280 ;
        RECT 191.480 4.000 191.560 4.280 ;
        RECT 192.400 4.000 192.940 4.280 ;
        RECT 193.780 4.000 194.320 4.280 ;
        RECT 195.160 4.000 195.240 4.280 ;
        RECT 196.080 4.000 196.620 4.280 ;
        RECT 197.460 4.000 198.000 4.280 ;
        RECT 198.840 4.000 198.920 4.280 ;
        RECT 199.760 4.000 200.300 4.280 ;
        RECT 201.140 4.000 201.680 4.280 ;
        RECT 202.520 4.000 202.600 4.280 ;
        RECT 203.440 4.000 203.980 4.280 ;
        RECT 204.820 4.000 205.360 4.280 ;
        RECT 206.200 4.000 206.280 4.280 ;
        RECT 207.120 4.000 207.660 4.280 ;
        RECT 208.500 4.000 209.040 4.280 ;
        RECT 209.880 4.000 209.960 4.280 ;
        RECT 210.800 4.000 211.340 4.280 ;
        RECT 212.180 4.000 212.720 4.280 ;
        RECT 213.560 4.000 213.640 4.280 ;
        RECT 214.480 4.000 215.020 4.280 ;
        RECT 215.860 4.000 216.400 4.280 ;
        RECT 217.240 4.000 217.320 4.280 ;
        RECT 218.160 4.000 218.700 4.280 ;
        RECT 219.540 4.000 220.080 4.280 ;
        RECT 220.920 4.000 221.000 4.280 ;
        RECT 221.840 4.000 222.380 4.280 ;
        RECT 223.220 4.000 223.760 4.280 ;
        RECT 224.600 4.000 224.680 4.280 ;
        RECT 225.520 4.000 226.060 4.280 ;
        RECT 226.900 4.000 226.980 4.280 ;
        RECT 227.820 4.000 228.360 4.280 ;
        RECT 229.200 4.000 229.740 4.280 ;
        RECT 230.580 4.000 230.660 4.280 ;
        RECT 231.500 4.000 232.040 4.280 ;
        RECT 232.880 4.000 233.420 4.280 ;
        RECT 234.260 4.000 234.340 4.280 ;
        RECT 235.180 4.000 235.720 4.280 ;
        RECT 236.560 4.000 237.100 4.280 ;
        RECT 237.940 4.000 238.020 4.280 ;
        RECT 238.860 4.000 239.400 4.280 ;
        RECT 240.240 4.000 240.780 4.280 ;
        RECT 241.620 4.000 241.700 4.280 ;
        RECT 242.540 4.000 243.080 4.280 ;
        RECT 243.920 4.000 244.460 4.280 ;
        RECT 245.300 4.000 245.380 4.280 ;
        RECT 246.220 4.000 246.760 4.280 ;
        RECT 247.600 4.000 248.140 4.280 ;
        RECT 248.980 4.000 249.060 4.280 ;
        RECT 249.900 4.000 250.440 4.280 ;
        RECT 251.280 4.000 251.820 4.280 ;
        RECT 252.660 4.000 252.740 4.280 ;
        RECT 253.580 4.000 254.120 4.280 ;
        RECT 254.960 4.000 255.500 4.280 ;
        RECT 256.340 4.000 256.420 4.280 ;
        RECT 257.260 4.000 257.800 4.280 ;
        RECT 258.640 4.000 259.180 4.280 ;
        RECT 260.020 4.000 260.100 4.280 ;
        RECT 260.940 4.000 261.480 4.280 ;
        RECT 262.320 4.000 262.860 4.280 ;
        RECT 263.700 4.000 263.780 4.280 ;
        RECT 264.620 4.000 265.160 4.280 ;
        RECT 266.000 4.000 266.540 4.280 ;
        RECT 267.380 4.000 267.460 4.280 ;
        RECT 268.300 4.000 268.840 4.280 ;
        RECT 269.680 4.000 270.220 4.280 ;
        RECT 271.060 4.000 271.140 4.280 ;
        RECT 271.980 4.000 272.520 4.280 ;
        RECT 273.360 4.000 273.900 4.280 ;
        RECT 274.740 4.000 274.820 4.280 ;
        RECT 275.660 4.000 276.200 4.280 ;
        RECT 277.040 4.000 277.580 4.280 ;
        RECT 278.420 4.000 278.500 4.280 ;
        RECT 279.340 4.000 279.880 4.280 ;
        RECT 280.720 4.000 281.260 4.280 ;
        RECT 282.100 4.000 282.180 4.280 ;
        RECT 283.020 4.000 283.560 4.280 ;
        RECT 284.400 4.000 284.940 4.280 ;
        RECT 285.780 4.000 285.860 4.280 ;
        RECT 286.700 4.000 287.240 4.280 ;
        RECT 288.080 4.000 288.620 4.280 ;
        RECT 289.460 4.000 289.540 4.280 ;
        RECT 290.380 4.000 290.920 4.280 ;
        RECT 291.760 4.000 292.300 4.280 ;
        RECT 293.140 4.000 293.220 4.280 ;
        RECT 294.060 4.000 294.600 4.280 ;
        RECT 295.440 4.000 295.980 4.280 ;
        RECT 296.820 4.000 296.900 4.280 ;
        RECT 297.740 4.000 298.280 4.280 ;
        RECT 299.120 4.000 299.660 4.280 ;
        RECT 300.500 4.000 300.580 4.280 ;
        RECT 301.420 4.000 301.960 4.280 ;
        RECT 302.800 4.000 302.880 4.280 ;
        RECT 303.720 4.000 304.260 4.280 ;
        RECT 305.100 4.000 305.640 4.280 ;
        RECT 306.480 4.000 306.560 4.280 ;
        RECT 307.400 4.000 307.940 4.280 ;
        RECT 308.780 4.000 309.320 4.280 ;
        RECT 310.160 4.000 310.240 4.280 ;
        RECT 311.080 4.000 311.620 4.280 ;
        RECT 312.460 4.000 313.000 4.280 ;
        RECT 313.840 4.000 313.920 4.280 ;
        RECT 314.760 4.000 315.300 4.280 ;
        RECT 316.140 4.000 316.680 4.280 ;
        RECT 317.520 4.000 317.600 4.280 ;
        RECT 318.440 4.000 318.980 4.280 ;
        RECT 319.820 4.000 320.360 4.280 ;
        RECT 321.200 4.000 321.280 4.280 ;
        RECT 322.120 4.000 322.660 4.280 ;
        RECT 323.500 4.000 324.040 4.280 ;
        RECT 324.880 4.000 324.960 4.280 ;
        RECT 325.800 4.000 326.340 4.280 ;
        RECT 327.180 4.000 327.720 4.280 ;
        RECT 328.560 4.000 328.640 4.280 ;
        RECT 329.480 4.000 330.020 4.280 ;
        RECT 330.860 4.000 331.400 4.280 ;
        RECT 332.240 4.000 332.320 4.280 ;
        RECT 333.160 4.000 333.700 4.280 ;
        RECT 334.540 4.000 335.080 4.280 ;
        RECT 335.920 4.000 336.000 4.280 ;
        RECT 336.840 4.000 337.380 4.280 ;
        RECT 338.220 4.000 338.760 4.280 ;
        RECT 339.600 4.000 339.680 4.280 ;
        RECT 340.520 4.000 341.060 4.280 ;
        RECT 341.900 4.000 342.440 4.280 ;
        RECT 343.280 4.000 343.360 4.280 ;
        RECT 344.200 4.000 344.740 4.280 ;
        RECT 345.580 4.000 346.120 4.280 ;
        RECT 346.960 4.000 347.040 4.280 ;
        RECT 347.880 4.000 348.420 4.280 ;
        RECT 349.260 4.000 349.800 4.280 ;
        RECT 350.640 4.000 350.720 4.280 ;
        RECT 351.560 4.000 352.100 4.280 ;
        RECT 352.940 4.000 353.480 4.280 ;
        RECT 354.320 4.000 354.400 4.280 ;
        RECT 355.240 4.000 355.780 4.280 ;
        RECT 356.620 4.000 357.160 4.280 ;
        RECT 358.000 4.000 358.080 4.280 ;
        RECT 358.920 4.000 359.460 4.280 ;
        RECT 360.300 4.000 360.840 4.280 ;
        RECT 361.680 4.000 361.760 4.280 ;
        RECT 362.600 4.000 363.140 4.280 ;
        RECT 363.980 4.000 364.520 4.280 ;
        RECT 365.360 4.000 365.440 4.280 ;
        RECT 366.280 4.000 366.820 4.280 ;
        RECT 367.660 4.000 368.200 4.280 ;
        RECT 369.040 4.000 369.120 4.280 ;
        RECT 369.960 4.000 370.500 4.280 ;
        RECT 371.340 4.000 371.880 4.280 ;
        RECT 372.720 4.000 372.800 4.280 ;
        RECT 373.640 4.000 374.180 4.280 ;
        RECT 375.020 4.000 375.100 4.280 ;
        RECT 375.940 4.000 376.480 4.280 ;
        RECT 377.320 4.000 377.860 4.280 ;
        RECT 378.700 4.000 378.780 4.280 ;
        RECT 379.620 4.000 380.160 4.280 ;
        RECT 381.000 4.000 381.540 4.280 ;
        RECT 382.380 4.000 382.460 4.280 ;
        RECT 383.300 4.000 383.840 4.280 ;
        RECT 384.680 4.000 385.220 4.280 ;
        RECT 386.060 4.000 386.140 4.280 ;
        RECT 386.980 4.000 387.520 4.280 ;
        RECT 388.360 4.000 388.900 4.280 ;
        RECT 389.740 4.000 389.820 4.280 ;
        RECT 390.660 4.000 391.200 4.280 ;
        RECT 392.040 4.000 392.580 4.280 ;
        RECT 393.420 4.000 393.500 4.280 ;
        RECT 394.340 4.000 394.880 4.280 ;
        RECT 395.720 4.000 396.260 4.280 ;
        RECT 397.100 4.000 397.180 4.280 ;
        RECT 398.020 4.000 398.560 4.280 ;
        RECT 399.400 4.000 399.940 4.280 ;
        RECT 400.780 4.000 400.860 4.280 ;
        RECT 401.700 4.000 402.240 4.280 ;
        RECT 403.080 4.000 403.620 4.280 ;
        RECT 404.460 4.000 404.540 4.280 ;
        RECT 405.380 4.000 405.920 4.280 ;
        RECT 406.760 4.000 407.300 4.280 ;
        RECT 408.140 4.000 408.220 4.280 ;
        RECT 409.060 4.000 409.600 4.280 ;
        RECT 410.440 4.000 410.980 4.280 ;
        RECT 411.820 4.000 411.900 4.280 ;
        RECT 412.740 4.000 413.280 4.280 ;
        RECT 414.120 4.000 414.660 4.280 ;
        RECT 415.500 4.000 415.580 4.280 ;
        RECT 416.420 4.000 416.960 4.280 ;
        RECT 417.800 4.000 418.340 4.280 ;
        RECT 419.180 4.000 419.260 4.280 ;
        RECT 420.100 4.000 420.640 4.280 ;
        RECT 421.480 4.000 422.020 4.280 ;
        RECT 422.860 4.000 422.940 4.280 ;
        RECT 423.780 4.000 424.320 4.280 ;
        RECT 425.160 4.000 425.700 4.280 ;
        RECT 426.540 4.000 426.620 4.280 ;
        RECT 427.460 4.000 428.000 4.280 ;
        RECT 428.840 4.000 429.380 4.280 ;
        RECT 430.220 4.000 430.300 4.280 ;
        RECT 431.140 4.000 431.680 4.280 ;
        RECT 432.520 4.000 433.060 4.280 ;
        RECT 433.900 4.000 433.980 4.280 ;
        RECT 434.820 4.000 435.360 4.280 ;
        RECT 436.200 4.000 436.740 4.280 ;
        RECT 437.580 4.000 437.660 4.280 ;
        RECT 438.500 4.000 439.040 4.280 ;
        RECT 439.880 4.000 440.420 4.280 ;
        RECT 441.260 4.000 441.340 4.280 ;
        RECT 442.180 4.000 442.720 4.280 ;
        RECT 443.560 4.000 444.100 4.280 ;
        RECT 444.940 4.000 445.020 4.280 ;
        RECT 445.860 4.000 446.400 4.280 ;
        RECT 447.240 4.000 447.780 4.280 ;
        RECT 448.620 4.000 448.700 4.280 ;
        RECT 449.540 4.000 450.080 4.280 ;
        RECT 450.920 4.000 451.000 4.280 ;
        RECT 451.840 4.000 452.380 4.280 ;
        RECT 453.220 4.000 453.760 4.280 ;
        RECT 454.600 4.000 454.680 4.280 ;
        RECT 455.520 4.000 456.060 4.280 ;
        RECT 456.900 4.000 457.440 4.280 ;
        RECT 458.280 4.000 458.360 4.280 ;
        RECT 459.200 4.000 459.740 4.280 ;
        RECT 460.580 4.000 461.120 4.280 ;
        RECT 461.960 4.000 462.040 4.280 ;
        RECT 462.880 4.000 463.420 4.280 ;
        RECT 464.260 4.000 464.800 4.280 ;
        RECT 465.640 4.000 465.720 4.280 ;
        RECT 466.560 4.000 467.100 4.280 ;
        RECT 467.940 4.000 468.480 4.280 ;
        RECT 469.320 4.000 469.400 4.280 ;
        RECT 470.240 4.000 470.780 4.280 ;
        RECT 471.620 4.000 472.160 4.280 ;
        RECT 473.000 4.000 473.080 4.280 ;
        RECT 473.920 4.000 474.460 4.280 ;
        RECT 475.300 4.000 475.840 4.280 ;
        RECT 476.680 4.000 476.760 4.280 ;
        RECT 477.600 4.000 478.140 4.280 ;
        RECT 478.980 4.000 479.520 4.280 ;
        RECT 480.360 4.000 480.440 4.280 ;
        RECT 481.280 4.000 481.820 4.280 ;
        RECT 482.660 4.000 483.200 4.280 ;
        RECT 484.040 4.000 484.120 4.280 ;
        RECT 484.960 4.000 485.500 4.280 ;
        RECT 486.340 4.000 486.880 4.280 ;
        RECT 487.720 4.000 487.800 4.280 ;
        RECT 488.640 4.000 489.180 4.280 ;
        RECT 490.020 4.000 490.560 4.280 ;
        RECT 491.400 4.000 491.480 4.280 ;
        RECT 492.320 4.000 492.860 4.280 ;
        RECT 493.700 4.000 494.240 4.280 ;
        RECT 495.080 4.000 495.160 4.280 ;
        RECT 496.000 4.000 496.540 4.280 ;
        RECT 497.380 4.000 497.920 4.280 ;
        RECT 498.760 4.000 498.840 4.280 ;
        RECT 499.680 4.000 500.220 4.280 ;
        RECT 501.060 4.000 501.600 4.280 ;
        RECT 502.440 4.000 502.520 4.280 ;
        RECT 503.360 4.000 503.900 4.280 ;
        RECT 504.740 4.000 505.280 4.280 ;
        RECT 506.120 4.000 506.200 4.280 ;
        RECT 507.040 4.000 507.580 4.280 ;
        RECT 508.420 4.000 508.960 4.280 ;
        RECT 509.800 4.000 509.880 4.280 ;
        RECT 510.720 4.000 511.260 4.280 ;
        RECT 512.100 4.000 512.640 4.280 ;
        RECT 513.480 4.000 513.560 4.280 ;
        RECT 514.400 4.000 514.940 4.280 ;
        RECT 515.780 4.000 516.320 4.280 ;
        RECT 517.160 4.000 517.240 4.280 ;
        RECT 518.080 4.000 518.620 4.280 ;
        RECT 519.460 4.000 520.000 4.280 ;
        RECT 520.840 4.000 520.920 4.280 ;
        RECT 521.760 4.000 522.300 4.280 ;
        RECT 523.140 4.000 523.680 4.280 ;
        RECT 524.520 4.000 524.600 4.280 ;
        RECT 525.440 4.000 525.980 4.280 ;
        RECT 526.820 4.000 526.900 4.280 ;
        RECT 527.740 4.000 528.280 4.280 ;
        RECT 529.120 4.000 529.660 4.280 ;
        RECT 530.500 4.000 530.580 4.280 ;
        RECT 531.420 4.000 531.960 4.280 ;
        RECT 532.800 4.000 533.340 4.280 ;
        RECT 534.180 4.000 534.260 4.280 ;
        RECT 535.100 4.000 535.640 4.280 ;
        RECT 536.480 4.000 537.020 4.280 ;
        RECT 537.860 4.000 537.940 4.280 ;
        RECT 538.780 4.000 539.320 4.280 ;
        RECT 540.160 4.000 540.700 4.280 ;
        RECT 541.540 4.000 541.620 4.280 ;
        RECT 542.460 4.000 543.000 4.280 ;
        RECT 543.840 4.000 544.380 4.280 ;
        RECT 545.220 4.000 545.300 4.280 ;
        RECT 546.140 4.000 546.680 4.280 ;
        RECT 547.520 4.000 548.060 4.280 ;
        RECT 548.900 4.000 548.980 4.280 ;
        RECT 549.820 4.000 550.360 4.280 ;
        RECT 551.200 4.000 551.740 4.280 ;
        RECT 552.580 4.000 552.660 4.280 ;
        RECT 553.500 4.000 554.040 4.280 ;
        RECT 554.880 4.000 555.420 4.280 ;
        RECT 556.260 4.000 556.340 4.280 ;
        RECT 557.180 4.000 557.720 4.280 ;
        RECT 558.560 4.000 559.100 4.280 ;
        RECT 559.940 4.000 560.020 4.280 ;
        RECT 560.860 4.000 561.400 4.280 ;
        RECT 562.240 4.000 562.780 4.280 ;
        RECT 563.620 4.000 563.700 4.280 ;
        RECT 564.540 4.000 565.080 4.280 ;
        RECT 565.920 4.000 566.460 4.280 ;
        RECT 567.300 4.000 567.380 4.280 ;
        RECT 568.220 4.000 568.760 4.280 ;
        RECT 569.600 4.000 570.140 4.280 ;
        RECT 570.980 4.000 571.060 4.280 ;
        RECT 571.900 4.000 572.440 4.280 ;
        RECT 573.280 4.000 573.820 4.280 ;
        RECT 574.660 4.000 574.740 4.280 ;
        RECT 575.580 4.000 576.120 4.280 ;
        RECT 576.960 4.000 577.500 4.280 ;
        RECT 578.340 4.000 578.420 4.280 ;
        RECT 579.260 4.000 579.800 4.280 ;
        RECT 580.640 4.000 581.180 4.280 ;
        RECT 582.020 4.000 582.100 4.280 ;
        RECT 582.940 4.000 583.480 4.280 ;
        RECT 584.320 4.000 584.860 4.280 ;
        RECT 585.700 4.000 585.780 4.280 ;
        RECT 586.620 4.000 587.160 4.280 ;
        RECT 588.000 4.000 588.540 4.280 ;
        RECT 589.380 4.000 589.460 4.280 ;
        RECT 590.300 4.000 590.840 4.280 ;
        RECT 591.680 4.000 592.220 4.280 ;
        RECT 593.060 4.000 593.140 4.280 ;
        RECT 593.980 4.000 594.520 4.280 ;
        RECT 595.360 4.000 595.900 4.280 ;
        RECT 596.740 4.000 596.820 4.280 ;
      LAYER met3 ;
        RECT 0.915 4.255 559.710 587.685 ;
      LAYER met4 ;
        RECT 95.445 11.055 96.910 76.665 ;
        RECT 99.310 11.055 100.210 76.665 ;
        RECT 102.610 11.055 103.510 76.665 ;
        RECT 105.910 11.055 106.810 76.665 ;
        RECT 109.210 11.055 173.710 76.665 ;
        RECT 176.110 11.055 177.010 76.665 ;
        RECT 179.410 11.055 180.310 76.665 ;
        RECT 182.710 11.055 183.610 76.665 ;
        RECT 186.010 11.055 208.015 76.665 ;
  END
END user_proj_example
END LIBRARY

