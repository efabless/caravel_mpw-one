VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_control_block
  CLASS BLOCK ;
  FOREIGN gpio_control_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 70.000 ;
  PIN mgmt_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 5.480 170.000 6.080 ;
    END
  END mgmt_gpio_in
  PIN mgmt_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 8.200 170.000 8.800 ;
    END
  END mgmt_gpio_oeb
  PIN mgmt_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 10.920 170.000 11.520 ;
    END
  END mgmt_gpio_out
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 2.760 170.000 3.360 ;
    END
  END one
  PIN pad_gpio_ana_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 13.640 170.000 14.240 ;
    END
  END pad_gpio_ana_en
  PIN pad_gpio_ana_pol
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 16.360 170.000 16.960 ;
    END
  END pad_gpio_ana_pol
  PIN pad_gpio_ana_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 19.080 170.000 19.680 ;
    END
  END pad_gpio_ana_sel
  PIN pad_gpio_dm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 21.800 170.000 22.400 ;
    END
  END pad_gpio_dm[0]
  PIN pad_gpio_dm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 24.520 170.000 25.120 ;
    END
  END pad_gpio_dm[1]
  PIN pad_gpio_dm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 27.240 170.000 27.840 ;
    END
  END pad_gpio_dm[2]
  PIN pad_gpio_holdover
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 29.960 170.000 30.560 ;
    END
  END pad_gpio_holdover
  PIN pad_gpio_ib_mode_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 32.680 170.000 33.280 ;
    END
  END pad_gpio_ib_mode_sel
  PIN pad_gpio_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 35.400 170.000 36.000 ;
    END
  END pad_gpio_in
  PIN pad_gpio_inenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 38.120 170.000 38.720 ;
    END
  END pad_gpio_inenb
  PIN pad_gpio_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 40.840 170.000 41.440 ;
    END
  END pad_gpio_out
  PIN pad_gpio_outenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 43.560 170.000 44.160 ;
    END
  END pad_gpio_outenb
  PIN pad_gpio_slow_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 46.280 170.000 46.880 ;
    END
  END pad_gpio_slow_sel
  PIN pad_gpio_vtrip_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 49.000 170.000 49.600 ;
    END
  END pad_gpio_vtrip_sel
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 51.720 170.000 52.320 ;
    END
  END resetn
  PIN serial_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 54.440 170.000 55.040 ;
    END
  END serial_clock
  PIN serial_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 57.160 170.000 57.760 ;
    END
  END serial_data_in
  PIN serial_data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 59.880 170.000 60.480 ;
    END
  END serial_data_out
  PIN user_gpio_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 62.600 170.000 63.200 ;
    END
  END user_gpio_in
  PIN user_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 65.320 170.000 65.920 ;
    END
  END user_gpio_oeb
  PIN user_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 68.040 170.000 68.640 ;
    END
  END user_gpio_out
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 0.720 170.000 1.320 ;
    END
  END zero
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.300 4.780 26.900 63.220 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.300 4.780 11.900 63.220 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 36.620 8.080 38.220 59.920 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.800 8.080 3.400 59.920 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 1.800 58.320 38.220 59.920 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -1.500 50.580 41.520 52.180 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -1.500 34.580 41.520 36.180 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -1.500 18.580 41.520 20.180 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 1.800 8.080 38.220 9.680 ;
    END
  END vccd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.920 4.780 41.520 63.220 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 17.800 4.780 19.400 63.220 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -1.500 4.780 0.100 63.220 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -1.500 61.620 41.520 63.220 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -1.500 42.580 41.520 44.180 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -1.500 26.580 41.520 28.180 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -1.500 4.780 41.520 6.380 ;
    END
  END vssd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.800 -1.820 31.400 69.820 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.800 -1.820 16.400 69.820 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 43.220 1.480 44.820 66.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -4.800 1.480 -3.200 66.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -4.800 64.920 44.820 66.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -8.100 39.080 48.120 40.680 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -8.100 23.080 48.120 24.680 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -4.800 1.480 44.820 3.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.520 -1.820 48.120 69.820 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 22.300 -1.820 23.900 69.820 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -8.100 -1.820 -6.500 69.820 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -8.100 68.220 48.120 69.820 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -8.100 47.080 48.120 48.680 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -8.100 31.080 48.120 32.680 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -8.100 -1.820 48.120 -0.220 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 0.460 10.795 35.420 57.205 ;
      LAYER met1 ;
        RECT 0.000 5.820 132.410 62.860 ;
      LAYER met2 ;
        RECT 0.000 0.835 132.390 68.525 ;
      LAYER met3 ;
        RECT 0.000 10.715 26.900 57.360 ;
  END
END gpio_control_block
END LIBRARY

