*** This is a chip_io smoke test with transient supply ramps

* Most models come from here:
.lib ../../../../../../../pdks/sky130A-xyce/libs.tech/xyce/sky130.lib.spice tt
*.inc ../../../../../../../pdks/sky130A-xyce/libs.tech/xyce/all.spice

* Include chip_io .subckt extracted using Calibre:
.include ./chip_io-extracted.spice

* This device is also missing from the libraries:
.include ./sky130_fd_io__condiode.spice
.include ./sky130_fd_pr__model__parasitic__diode_ps2nw.spice 
.include ./sky130_fd_pr__model__parasitic__diode_pw2dn.spice
.include ./sky130_fd_pr__model__parasitic__diode_ps2dn.spice
.include ./sky130_fd_pr__diode_pd2nw_05v5.spice
.include ./sky130_fd_pr__diode_pw2nd_11v0.spice

***************************************

*********************
Xchip_io  mprj_io_oeb[24] mprj_io_ib_mode_sel[24] mprj_io_vtrip_sel[24] mprj_io_out[24] mprj_io_holdover[24] mprj_io_dm[74] mprj_io_analog_sel[24] mprj_io_hldh_n[24] mprj_io_enh[24] mprj_io_inp_dis[24] mprj_io_analog_pol[24] mprj_io_dm[72] mprj_io_analog_en[24] mprj_io_dm[73] mprj_analog_io[17] mprj_io_slow_sel[24] mprj_io_in[24] porb_h mprj_io_oeb[23] mprj_io_ib_mode_sel[23]
+ mprj_io_vtrip_sel[23] mprj_io_out[23] mprj_io_holdover[23] mprj_io_dm[71] mprj_io_analog_sel[23] mprj_io_hldh_n[23] mprj_io_enh[23] mprj_io_inp_dis[23] mprj_io_analog_pol[23] mprj_io_dm[69] mprj_io_analog_en[23] mprj_io_dm[70] mprj_analog_io[16] mprj_io_slow_sel[23] mprj_io_in[23] mprj_io_oeb[22] mprj_io_ib_mode_sel[22] mprj_io_vtrip_sel[22] mprj_io_out[22] mprj_io_holdover[22]
+ mprj_io_dm[68] mprj_io_analog_sel[22] mprj_io_hldh_n[22] mprj_io_enh[22] mprj_io_inp_dis[22] mprj_io_analog_pol[22] mprj_io_dm[66] mprj_io_analog_en[22] mprj_io_dm[67] mprj_analog_io[15] mprj_io_slow_sel[22] mprj_io_in[22] mprj_io_oeb[21] mprj_io_ib_mode_sel[21] mprj_io_vtrip_sel[21] mprj_io_out[21] mprj_io_holdover[21] mprj_io_dm[65] mprj_io_analog_sel[21] mprj_io_hldh_n[21]
+ mprj_io_enh[21] mprj_io_inp_dis[21] mprj_io_analog_pol[21] mprj_io_dm[63] mprj_io_analog_en[21] mprj_io_dm[64] mprj_analog_io[14] mprj_io_slow_sel[21] mprj_io_in[21] mprj_io_oeb[20] mprj_io_ib_mode_sel[20] mprj_io_vtrip_sel[20] mprj_io_out[20] mprj_io_holdover[20] mprj_io_dm[62] mprj_io_analog_sel[20] mprj_io_hldh_n[20] mprj_io_enh[20] mprj_io_inp_dis[20] mprj_io_analog_pol[20]
+ mprj_io_dm[60] mprj_io_analog_en[20] mprj_io_dm[61] mprj_analog_io[13] mprj_io_slow_sel[20] mprj_io_in[20] mprj_io_oeb[19] mprj_io_ib_mode_sel[19] mprj_io_vtrip_sel[19] mprj_io_out[19] mprj_io_holdover[19] mprj_io_dm[59] mprj_io_analog_sel[19] mprj_io_hldh_n[19] mprj_io_enh[19] mprj_io_inp_dis[19] mprj_io_analog_pol[19] mprj_io_dm[57] mprj_io_analog_en[19] mprj_io_dm[58]
+ mprj_analog_io[12] mprj_io_slow_sel[19] mprj_io_in[19] mprj_io_oeb[18] mprj_io_ib_mode_sel[18] mprj_io_vtrip_sel[18] mprj_io_out[18] mprj_io_holdover[18] mprj_io_dm[56] mprj_io_analog_sel[18] mprj_io_hldh_n[18] mprj_io_enh[18] mprj_io_inp_dis[18] mprj_io_analog_pol[18] mprj_io_dm[54] mprj_io_analog_en[18] mprj_io_dm[55] mprj_analog_io[11] mprj_io_slow_sel[18] mprj_io_in[18]
+ mprj_io_oeb[17] mprj_io_ib_mode_sel[17] mprj_io_vtrip_sel[17] mprj_io_out[17] mprj_io_holdover[17] mprj_io_dm[53] mprj_io_analog_sel[17] mprj_io_hldh_n[17] mprj_io_enh[17] mprj_io_inp_dis[17] mprj_io_analog_pol[17] mprj_io_dm[51] mprj_io_analog_en[17] mprj_io_dm[52] mprj_analog_io[10] mprj_io_slow_sel[17] mprj_io_in[17] mprj_io_oeb[16] mprj_io_ib_mode_sel[16] mprj_io_vtrip_sel[16]
+ mprj_io_out[16] mprj_io_holdover[16] mprj_io_dm[50] mprj_io_analog_sel[16] mprj_io_hldh_n[16] mprj_io_enh[16] mprj_io_inp_dis[16] mprj_io_analog_pol[16] mprj_io_dm[48] mprj_io_analog_en[16] mprj_io_dm[49] mprj_analog_io[9] mprj_io_slow_sel[16] mprj_io_in[16] mprj_io_oeb[15] mprj_io_ib_mode_sel[15] mprj_io_vtrip_sel[15] mprj_io_out[15] mprj_io_holdover[15] mprj_io_dm[47]
+ mprj_io_analog_sel[15] mprj_io_hldh_n[15] mprj_io_enh[15] mprj_io_inp_dis[15] mprj_io_analog_pol[15] mprj_io_dm[45] mprj_io_analog_en[15] mprj_io_dm[46] mprj_analog_io[8] mprj_io_slow_sel[15] mprj_io_in[15] mprj_io_in[14] mprj_io_slow_sel[14] mprj_analog_io[7] mprj_io_dm[43] mprj_io_analog_en[14] mprj_io_dm[42] mprj_io_analog_pol[14] mprj_io_inp_dis[14] mprj_io_enh[14]
+ mprj_io_hldh_n[14] mprj_io_analog_sel[14] mprj_io_dm[44] mprj_io_holdover[14] mprj_io_out[14] mprj_io_vtrip_sel[14] mprj_io_ib_mode_sel[14] mprj_io_oeb[14] mprj_io_in[13] mprj_io_slow_sel[13] mprj_analog_io[6] mprj_io_dm[40] mprj_io_analog_en[13] mprj_io_dm[39] mprj_io_analog_pol[13] mprj_io_inp_dis[13] mprj_io_enh[13] mprj_io_hldh_n[13] mprj_io_analog_sel[13] mprj_io_dm[41]
+ mprj_io_holdover[13] mprj_io_out[13] mprj_io_vtrip_sel[13] mprj_io_ib_mode_sel[13] mprj_io_oeb[13] mprj_io_oeb[31] mprj_io_ib_mode_sel[31] mprj_io_vtrip_sel[31] mprj_io_out[31] mprj_io_holdover[31] mprj_io_dm[95] mprj_io_analog_sel[31] mprj_io_hldh_n[31] mprj_io_enh[31] mprj_io_inp_dis[31] mprj_io_analog_pol[31] mprj_io_dm[93] mprj_io_analog_en[31] mprj_io_dm[94] mprj_analog_io[24]
+ mprj_io_slow_sel[31] mprj_io_in[31] mprj_io_oeb[30] mprj_io_ib_mode_sel[30] mprj_io_vtrip_sel[30] mprj_io_out[30] mprj_io_holdover[30] mprj_io_dm[92] mprj_io_analog_sel[30] mprj_io_hldh_n[30] mprj_io_enh[30] mprj_io_inp_dis[30] mprj_io_analog_pol[30] mprj_io_dm[90] mprj_io_analog_en[30] mprj_io_dm[91] mprj_analog_io[23] mprj_io_slow_sel[30] mprj_io_in[30] mprj_io_oeb[29]
+ mprj_io_ib_mode_sel[29] mprj_io_vtrip_sel[29] mprj_io_out[29] mprj_io_holdover[29] mprj_io_dm[89] mprj_io_analog_sel[29] mprj_io_hldh_n[29] mprj_io_enh[29] mprj_io_inp_dis[29] mprj_io_analog_pol[29] mprj_io_dm[87] mprj_io_analog_en[29] mprj_io_dm[88] mprj_analog_io[22] mprj_io_slow_sel[29] mprj_io_in[29] mprj_io_oeb[28] mprj_io_ib_mode_sel[28] mprj_io_vtrip_sel[28] mprj_io_out[28]
+ mprj_io_holdover[28] mprj_io_dm[86] mprj_io_analog_sel[28] mprj_io_hldh_n[28] mprj_io_enh[28] mprj_io_inp_dis[28] mprj_io_analog_pol[28] mprj_io_dm[84] mprj_io_analog_en[28] mprj_io_dm[85] mprj_analog_io[21] mprj_io_slow_sel[28] mprj_io_in[28] mprj_io_oeb[27] mprj_io_ib_mode_sel[27] mprj_io_vtrip_sel[27] mprj_io_out[27] mprj_io_holdover[27] mprj_io_dm[83] mprj_io_analog_sel[27]
+ mprj_io_hldh_n[27] mprj_io_enh[27] mprj_io_inp_dis[27] mprj_io_analog_pol[27] mprj_io_dm[81] mprj_io_analog_en[27] mprj_io_dm[82] mprj_analog_io[20] mprj_io_slow_sel[27] mprj_io_in[27] mprj_io_oeb[26] mprj_io_ib_mode_sel[26] mprj_io_vtrip_sel[26] mprj_io_out[26] mprj_io_holdover[26] mprj_io_dm[80] mprj_io_analog_sel[26] mprj_io_hldh_n[26] mprj_io_enh[26] mprj_io_inp_dis[26]
+ mprj_io_analog_pol[26] mprj_io_dm[78] mprj_io_analog_en[26] mprj_io_dm[79] mprj_analog_io[19] mprj_io_slow_sel[26] mprj_io_in[26] mprj_io_oeb[25] mprj_io_ib_mode_sel[25] mprj_io_vtrip_sel[25] mprj_io_out[25] mprj_io_holdover[25] mprj_io_dm[77] mprj_io_analog_sel[25] mprj_io_hldh_n[25] mprj_io_enh[25] mprj_io_inp_dis[25] mprj_io_analog_pol[25] mprj_io_dm[75] mprj_io_analog_en[25]
+ mprj_io_dm[76] mprj_analog_io[18] mprj_io_slow_sel[25] mprj_io_in[25] mprj_io_in[7] mprj_io_slow_sel[7] mprj_analog_io[0] mprj_io_dm[22] mprj_io_analog_en[7] mprj_io_dm[21] mprj_io_analog_pol[7] mprj_io_inp_dis[7] mprj_io_enh[7] mprj_io_hldh_n[7] mprj_io_analog_sel[7] mprj_io_dm[23] mprj_io_holdover[7] mprj_io_out[7] mprj_io_vtrip_sel[7] mprj_io_ib_mode_sel[7]
+ mprj_io_oeb[7] mprj_io_in[8] mprj_io_slow_sel[8] mprj_analog_io[1] mprj_io_dm[25] mprj_io_analog_en[8] mprj_io_dm[24] mprj_io_analog_pol[8] mprj_io_inp_dis[8] mprj_io_enh[8] mprj_io_hldh_n[8] mprj_io_analog_sel[8] mprj_io_dm[26] mprj_io_holdover[8] mprj_io_out[8] mprj_io_vtrip_sel[8] mprj_io_ib_mode_sel[8] mprj_io_oeb[8] mprj_io_in[9] mprj_io_slow_sel[9]
+ mprj_analog_io[2] mprj_io_dm[28] mprj_io_analog_en[9] mprj_io_dm[27] mprj_io_analog_pol[9] mprj_io_inp_dis[9] mprj_io_enh[9] mprj_io_hldh_n[9] mprj_io_analog_sel[9] mprj_io_dm[29] mprj_io_holdover[9] mprj_io_out[9] mprj_io_vtrip_sel[9] mprj_io_ib_mode_sel[9] mprj_io_oeb[9] mprj_io_in[10] mprj_io_slow_sel[10] mprj_analog_io[3] mprj_io_dm[31] mprj_io_analog_en[10]
+ mprj_io_dm[30] mprj_io_analog_pol[10] mprj_io_inp_dis[10] mprj_io_enh[10] mprj_io_hldh_n[10] mprj_io_analog_sel[10] mprj_io_dm[32] mprj_io_holdover[10] mprj_io_out[10] mprj_io_vtrip_sel[10] mprj_io_ib_mode_sel[10] mprj_io_oeb[10] mprj_io_in[11] mprj_io_slow_sel[11] mprj_analog_io[4] mprj_io_dm[34] mprj_io_analog_en[11] mprj_io_dm[33] mprj_io_analog_pol[11] mprj_io_inp_dis[11]
+ mprj_io_enh[11] mprj_io_hldh_n[11] mprj_io_analog_sel[11] mprj_io_dm[35] mprj_io_holdover[11] mprj_io_out[11] mprj_io_vtrip_sel[11] mprj_io_ib_mode_sel[11] mprj_io_oeb[11] mprj_io_in[12] mprj_io_slow_sel[12] mprj_analog_io[5] mprj_io_dm[37] mprj_io_analog_en[12] mprj_io_dm[36] mprj_io_analog_pol[12] mprj_io_inp_dis[12] mprj_io_enh[12] mprj_io_hldh_n[12] mprj_io_analog_sel[12]
+ mprj_io_dm[38] mprj_io_holdover[12] mprj_io_out[12] mprj_io_vtrip_sel[12] mprj_io_ib_mode_sel[12] mprj_io_oeb[12] mprj_io_oeb[37] mprj_io_ib_mode_sel[37] mprj_io_vtrip_sel[37] mprj_io_out[37] mprj_io_holdover[37] mprj_io_dm[113] mprj_io_analog_sel[37] mprj_io_hldh_n[37] mprj_io_enh[37] mprj_io_inp_dis[37] mprj_io_analog_pol[37] mprj_io_dm[111] mprj_io_analog_en[37] mprj_io_dm[112]
+ mprj_io_slow_sel[37] mprj_io_in[37] mprj_io_oeb[36] mprj_io_ib_mode_sel[36] mprj_io_vtrip_sel[36] mprj_io_out[36] mprj_io_holdover[36] mprj_io_dm[110] mprj_io_analog_sel[36] mprj_io_hldh_n[36] mprj_io_enh[36] mprj_io_inp_dis[36] mprj_io_analog_pol[36] mprj_io_dm[108] mprj_io_analog_en[36] mprj_io_dm[109] mprj_io_slow_sel[36] mprj_io_in[36] mprj_io_oeb[35] mprj_io_ib_mode_sel[35]
+ mprj_io_vtrip_sel[35] mprj_io_out[35] mprj_io_holdover[35] mprj_io_dm[107] mprj_io_analog_sel[35] mprj_io_hldh_n[35] mprj_io_enh[35] mprj_io_inp_dis[35] mprj_io_analog_pol[35] mprj_io_dm[105] mprj_io_analog_en[35] mprj_io_dm[106] mprj_analog_io[28] mprj_io_slow_sel[35] mprj_io_in[35] mprj_io_oeb[34] mprj_io_ib_mode_sel[34] mprj_io_vtrip_sel[34] mprj_io_out[34] mprj_io_holdover[34]
+ mprj_io_dm[104] mprj_io_analog_sel[34] mprj_io_hldh_n[34] mprj_io_enh[34] mprj_io_inp_dis[34] mprj_io_analog_pol[34] mprj_io_dm[102] mprj_io_analog_en[34] mprj_io_dm[103] mprj_analog_io[27] mprj_io_slow_sel[34] mprj_io_in[34] mprj_io_oeb[33] mprj_io_ib_mode_sel[33] mprj_io_vtrip_sel[33] mprj_io_out[33] mprj_io_holdover[33] mprj_io_dm[101] mprj_io_analog_sel[33] mprj_io_hldh_n[33]
+ mprj_io_enh[33] mprj_io_inp_dis[33] mprj_io_analog_pol[33] mprj_io_dm[99] mprj_io_analog_en[33] mprj_io_dm[100] mprj_analog_io[26] mprj_io_slow_sel[33] mprj_io_in[33] mprj_io_oeb[32] mprj_io_ib_mode_sel[32] mprj_io_vtrip_sel[32] mprj_io_out[32] mprj_io_holdover[32] mprj_io_dm[98] mprj_io_analog_sel[32] mprj_io_hldh_n[32] mprj_io_enh[32] mprj_io_inp_dis[32] mprj_io_analog_pol[32]
+ mprj_io_dm[96] mprj_io_analog_en[32] mprj_io_dm[97] mprj_analog_io[25] mprj_io_slow_sel[32] mprj_io_in[32] mprj_io_in[0] mprj_io_slow_sel[0] mprj_io_dm[1] mprj_io_analog_en[0] mprj_io_dm[0] mprj_io_analog_pol[0] mprj_io_inp_dis[0] mprj_io_enh[0] mprj_io_hldh_n[0] mprj_io_analog_sel[0] mprj_io_dm[2] mprj_io_holdover[0] mprj_io_out[0] mprj_io_vtrip_sel[0]
+ mprj_io_ib_mode_sel[0] mprj_io_oeb[0] mprj_io_in[1] mprj_io_slow_sel[1] mprj_io_dm[4] mprj_io_analog_en[1] mprj_io_dm[3] mprj_io_analog_pol[1] mprj_io_inp_dis[1] mprj_io_enh[1] mprj_io_hldh_n[1] mprj_io_analog_sel[1] mprj_io_dm[5] mprj_io_holdover[1] mprj_io_out[1] mprj_io_vtrip_sel[1] mprj_io_ib_mode_sel[1] mprj_io_oeb[1] mprj_io_in[2] mprj_io_slow_sel[2]
+ mprj_io_dm[7] mprj_io_analog_en[2] mprj_io_dm[6] mprj_io_analog_pol[2] mprj_io_inp_dis[2] mprj_io_enh[2] mprj_io_hldh_n[2] mprj_io_analog_sel[2] mprj_io_dm[8] mprj_io_holdover[2] mprj_io_out[2] mprj_io_vtrip_sel[2] mprj_io_ib_mode_sel[2] mprj_io_oeb[2] mprj_io_in[3] mprj_io_slow_sel[3] mprj_io_dm[10] mprj_io_analog_en[3] mprj_io_dm[9] mprj_io_analog_pol[3]
+ mprj_io_inp_dis[3] mprj_io_enh[3] mprj_io_hldh_n[3] mprj_io_analog_sel[3] mprj_io_dm[11] mprj_io_holdover[3] mprj_io_out[3] mprj_io_vtrip_sel[3] mprj_io_ib_mode_sel[3] mprj_io_oeb[3] mprj_io_in[4] mprj_io_slow_sel[4] mprj_io_dm[13] mprj_io_analog_en[4] mprj_io_dm[12] mprj_io_analog_pol[4] mprj_io_inp_dis[4] mprj_io_enh[4] mprj_io_hldh_n[4] mprj_io_analog_sel[4]
+ mprj_io_dm[14] mprj_io_holdover[4] mprj_io_out[4] mprj_io_vtrip_sel[4] mprj_io_ib_mode_sel[4] mprj_io_oeb[4] mprj_io_in[5] mprj_io_slow_sel[5] mprj_io_dm[16] mprj_io_analog_en[5] mprj_io_dm[15] mprj_io_analog_pol[5] mprj_io_inp_dis[5] mprj_io_enh[5] mprj_io_hldh_n[5] mprj_io_analog_sel[5] mprj_io_dm[17] mprj_io_holdover[5] mprj_io_out[5] mprj_io_vtrip_sel[5]
+ mprj_io_ib_mode_sel[5] mprj_io_oeb[5] mprj_io_in[6] mprj_io_slow_sel[6] mprj_io_dm[19] mprj_io_analog_en[6] mprj_io_dm[18] mprj_io_analog_pol[6] mprj_io_inp_dis[6] mprj_io_enh[6] mprj_io_hldh_n[6] mprj_io_analog_sel[6] mprj_io_dm[20] mprj_io_holdover[6] mprj_io_out[6] mprj_io_vtrip_sel[6] mprj_io_ib_mode_sel[6] mprj_io_oeb[6] clock_core por
+ flash_csb_ieb_core flash_csb_core flash_csb_oeb_core flash_clk_ieb_core flash_clk_core flash_clk_oeb_core flash_io0_di_core flash_io0_ieb_core flash_io0_do_core flash_io0_oeb_core flash_io1_di_core flash_io1_ieb_core flash_io1_do_core flash_io1_oeb_core gpio_in_core gpio_mode0_core gpio_inenb_core gpio_mode1_core gpio_out_core gpio_outenb_core
+ resetb_core_h mprj_io[24] vccd2_pad mprj_io[23] mprj_io[22] mprj_io[21] mprj_io[20] mprj_io[19] vssio_pad mprj_io[18] mprj_io[17] mprj_io[16] vssa1_pad mprj_io[15] vccd1_pad mprj_io[14] mprj_io[13] mprj_io[31] mprj_io[30] mprj_io[29]
+ mprj_io[28] mprj_io[27] mprj_io[26] mprj_io[25] vssa2_pad vdda1_pad mprj_io[7] mprj_io[8] mprj_io[9] mprj_io[10] mprj_io[11] mprj_io[12] vssd2_pad vdda2_pad vssd1_pad mprj_io[37] mprj_io[36] mprj_io[35] mprj_io[34] mprj_io[33]
+ mprj_io[32] vddio_pad mprj_io[0] mprj_io[1] mprj_io[2] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] vssa_pad clock flash_csb flash_clk flash_io0 flash_io1 gpio vdda_pad resetb vssd_pad vccd_pad
**
+ chip_io

***  

v1		vddio_pad	vdd3v3
v2		vddio_pad2	vdd3v3
v3		vssio_pad	vss3v3
v4		vssio_pad2	vss3v3
v5		vdda_pad	vdd3v3
v6		vssa_pad	vss3v3
v7		vccd_pad	vdd1v8	
v8		vssd_pad	vss1v8
v9		vdda1_pad	vdd3v3
v10		vdda1_pad2	vdd3v3
v11		vdda2_pad	vdd3v3
v12		vssa1_pad	vss3v3
v13		vssa1_pad2	vss3v3
v14		vssa2_pad	vss3v3
v15		vccd1_pad	vdd1v8
v16		vccd2_pad	vdd1v8
v17		vssd1_pad	vss1v8
v18		vssd2_pad	vss1v8

		
vvdd3v3		vdd3v3 	      	pwl	0 	2u  3.3  1m 3.3
vvss3p3		vss3v3 	      	dc	0
vvdd1v8		vdd1v8 	      	pwl 	0 	3u  1.8  1m 1.8
vvss1v8		vss1v8 	      	dc	0


.PRINT TRAN FORMAT=RAW 
+ vdd3v3    
+ vss3v3
+ vdd1v8
+ vss1v8

.TRAN 10n 2u

.END
