magic
tech sky130A
magscale 1 2
timestamp 1611263049
<< locali >>
rect 10333 8619 10367 9061
<< viali >>
rect 3525 11305 3559 11339
rect 3341 11237 3375 11271
rect 3985 11169 4019 11203
rect 4445 11169 4479 11203
rect 4721 11169 4755 11203
rect 4813 11169 4847 11203
rect 6101 11169 6135 11203
rect 1225 11101 1259 11135
rect 4997 11101 5031 11135
rect 6469 11101 6503 11135
rect 3709 11033 3743 11067
rect 4169 11033 4203 11067
rect 4537 11033 4571 11067
rect 1869 10625 1903 10659
rect 1593 10557 1627 10591
rect 3893 10557 3927 10591
rect 4353 10557 4387 10591
rect 6469 10557 6503 10591
rect 3617 10489 3651 10523
rect 4629 10489 4663 10523
rect 6377 10489 6411 10523
rect 4077 10421 4111 10455
rect 6653 10421 6687 10455
rect 1225 10081 1259 10115
rect 3709 10081 3743 10115
rect 5549 10081 5583 10115
rect 5733 10081 5767 10115
rect 6193 10081 6227 10115
rect 1501 10013 1535 10047
rect 3249 10013 3283 10047
rect 3341 10013 3375 10047
rect 5089 10013 5123 10047
rect 5825 9877 5859 9911
rect 6377 9877 6411 9911
rect 6745 9877 6779 9911
rect 6285 9673 6319 9707
rect 2053 9605 2087 9639
rect 3525 9537 3559 9571
rect 5917 9537 5951 9571
rect 1869 9469 1903 9503
rect 2697 9469 2731 9503
rect 2973 9469 3007 9503
rect 3065 9469 3099 9503
rect 3709 9469 3743 9503
rect 3893 9469 3927 9503
rect 6009 9469 6043 9503
rect 6101 9469 6135 9503
rect 2237 9401 2271 9435
rect 4169 9401 4203 9435
rect 1409 9129 1443 9163
rect 1777 9129 1811 9163
rect 2789 9129 2823 9163
rect 3157 9061 3191 9095
rect 4997 9061 5031 9095
rect 10333 9061 10367 9095
rect 1593 8993 1627 9027
rect 1685 8993 1719 9027
rect 1961 8993 1995 9027
rect 2329 8993 2363 9027
rect 5457 8993 5491 9027
rect 5733 8993 5767 9027
rect 5917 8993 5951 9027
rect 6377 8993 6411 9027
rect 2881 8925 2915 8959
rect 4905 8925 4939 8959
rect 6285 8925 6319 8959
rect 2145 8789 2179 8823
rect 2513 8789 2547 8823
rect 6653 8789 6687 8823
rect 3525 8585 3559 8619
rect 5917 8585 5951 8619
rect 6285 8585 6319 8619
rect 6745 8585 6779 8619
rect 10333 8585 10367 8619
rect 5181 8517 5215 8551
rect 1225 8449 1259 8483
rect 1501 8449 1535 8483
rect 6561 8449 6595 8483
rect 3341 8381 3375 8415
rect 3893 8381 3927 8415
rect 5733 8381 5767 8415
rect 6101 8381 6135 8415
rect 3249 8313 3283 8347
rect 6009 8041 6043 8075
rect 1501 7973 1535 8007
rect 1225 7905 1259 7939
rect 3341 7905 3375 7939
rect 4261 7905 4295 7939
rect 6101 7905 6135 7939
rect 3249 7837 3283 7871
rect 3893 7837 3927 7871
rect 3525 7701 3559 7735
rect 6285 7701 6319 7735
rect 6745 7701 6779 7735
rect 3617 7497 3651 7531
rect 6653 7497 6687 7531
rect 1593 7361 1627 7395
rect 1317 7293 1351 7327
rect 3433 7293 3467 7327
rect 3985 7293 4019 7327
rect 4353 7293 4387 7327
rect 6469 7293 6503 7327
rect 3341 7225 3375 7259
rect 4629 7225 4663 7259
rect 6377 7225 6411 7259
rect 4169 7157 4203 7191
rect 2421 6953 2455 6987
rect 3249 6885 3283 6919
rect 5917 6885 5951 6919
rect 1869 6817 1903 6851
rect 2237 6817 2271 6851
rect 5089 6817 5123 6851
rect 5457 6817 5491 6851
rect 5549 6817 5583 6851
rect 6745 6817 6779 6851
rect 2973 6749 3007 6783
rect 4997 6749 5031 6783
rect 5825 6749 5859 6783
rect 6101 6749 6135 6783
rect 2053 6613 2087 6647
rect 5273 6613 5307 6647
rect 1501 6273 1535 6307
rect 4537 6273 4571 6307
rect 1225 6205 1259 6239
rect 3433 6205 3467 6239
rect 4261 6205 4295 6239
rect 6377 6205 6411 6239
rect 3249 6137 3283 6171
rect 6285 6137 6319 6171
rect 3617 6069 3651 6103
rect 6561 6069 6595 6103
rect 5181 5865 5215 5899
rect 6745 5865 6779 5899
rect 4629 5797 4663 5831
rect 5917 5797 5951 5831
rect 1753 5729 1787 5763
rect 1894 5729 1928 5763
rect 2237 5729 2271 5763
rect 4997 5729 5031 5763
rect 5365 5729 5399 5763
rect 2605 5661 2639 5695
rect 2881 5661 2915 5695
rect 5825 5661 5859 5695
rect 6469 5661 6503 5695
rect 1593 5593 1627 5627
rect 2053 5525 2087 5559
rect 2421 5525 2455 5559
rect 4813 5525 4847 5559
rect 5549 5525 5583 5559
rect 1225 5185 1259 5219
rect 1501 5185 1535 5219
rect 3249 5185 3283 5219
rect 3341 5117 3375 5151
rect 3985 5117 4019 5151
rect 4353 5117 4387 5151
rect 4629 5117 4663 5151
rect 4997 5117 5031 5151
rect 3525 4981 3559 5015
rect 4169 4981 4203 5015
rect 4445 4981 4479 5015
rect 6745 4981 6779 5015
rect 3709 4709 3743 4743
rect 1317 4641 1351 4675
rect 3433 4641 3467 4675
rect 6009 4641 6043 4675
rect 6469 4641 6503 4675
rect 6745 4641 6779 4675
rect 1593 4573 1627 4607
rect 3341 4573 3375 4607
rect 5457 4573 5491 4607
rect 5825 4505 5859 4539
rect 5641 4437 5675 4471
rect 6469 4233 6503 4267
rect 1225 4097 1259 4131
rect 1501 4097 1535 4131
rect 3249 4097 3283 4131
rect 3893 4097 3927 4131
rect 4169 4097 4203 4131
rect 3341 4029 3375 4063
rect 5917 4029 5951 4063
rect 6101 4029 6135 4063
rect 6193 4029 6227 4063
rect 6285 4029 6319 4063
rect 3525 3893 3559 3927
rect 2145 3689 2179 3723
rect 4353 3621 4387 3655
rect 4721 3621 4755 3655
rect 6469 3621 6503 3655
rect 1961 3553 1995 3587
rect 2329 3553 2363 3587
rect 2605 3485 2639 3519
rect 4445 3485 4479 3519
rect 6745 3349 6779 3383
rect 6561 3145 6595 3179
rect 1961 3009 1995 3043
rect 3709 3009 3743 3043
rect 1685 2941 1719 2975
rect 3893 2941 3927 2975
rect 4445 2941 4479 2975
rect 4813 2941 4847 2975
rect 4077 2805 4111 2839
rect 6745 2805 6779 2839
rect 5457 2601 5491 2635
rect 5825 2601 5859 2635
rect 1961 2533 1995 2567
rect 6009 2533 6043 2567
rect 1685 2465 1719 2499
rect 3709 2465 3743 2499
rect 3893 2465 3927 2499
rect 5273 2465 5307 2499
rect 5641 2465 5675 2499
rect 6193 2465 6227 2499
rect 4997 2397 5031 2431
rect 4077 2329 4111 2363
rect 5181 2261 5215 2295
rect 6285 2261 6319 2295
<< metal1 >>
rect 6454 12452 6460 12504
rect 6512 12492 6518 12504
rect 16574 12492 16580 12504
rect 6512 12464 16580 12492
rect 6512 12452 6518 12464
rect 16574 12452 16580 12464
rect 16632 12452 16638 12504
rect 920 11450 7084 11472
rect 920 11398 3598 11450
rect 3650 11398 3662 11450
rect 3714 11398 3726 11450
rect 3778 11398 3790 11450
rect 3842 11398 7084 11450
rect 920 11376 7084 11398
rect 3513 11339 3571 11345
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 4522 11336 4528 11348
rect 3559 11308 4528 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 6822 11336 6828 11348
rect 4764 11308 6828 11336
rect 4764 11296 4770 11308
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 3326 11268 3332 11280
rect 3239 11240 3332 11268
rect 3326 11228 3332 11240
rect 3384 11268 3390 11280
rect 16574 11268 16580 11280
rect 3384 11240 16580 11268
rect 3384 11228 3390 11240
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 3970 11200 3976 11212
rect 3931 11172 3976 11200
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4522 11200 4528 11212
rect 4479 11172 4528 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 4706 11200 4712 11212
rect 4667 11172 4712 11200
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 4847 11172 6101 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 6089 11169 6101 11172
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 1213 11135 1271 11141
rect 1213 11101 1225 11135
rect 1259 11132 1271 11135
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 1259 11104 4997 11132
rect 1259 11101 1271 11104
rect 1213 11095 1271 11101
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 6454 11132 6460 11144
rect 6415 11104 6460 11132
rect 4985 11095 5043 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 3697 11067 3755 11073
rect 3697 11033 3709 11067
rect 3743 11064 3755 11067
rect 4154 11064 4160 11076
rect 3743 11036 4016 11064
rect 4115 11036 4160 11064
rect 3743 11033 3755 11036
rect 3697 11027 3755 11033
rect 3988 10996 4016 11036
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 4525 11067 4583 11073
rect 4525 11033 4537 11067
rect 4571 11064 4583 11067
rect 5442 11064 5448 11076
rect 4571 11036 5448 11064
rect 4571 11033 4583 11036
rect 4525 11027 4583 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 4706 10996 4712 11008
rect 3988 10968 4712 10996
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 920 10906 7084 10928
rect 920 10854 2098 10906
rect 2150 10854 2162 10906
rect 2214 10854 2226 10906
rect 2278 10854 2290 10906
rect 2342 10854 5098 10906
rect 5150 10854 5162 10906
rect 5214 10854 5226 10906
rect 5278 10854 5290 10906
rect 5342 10854 7084 10906
rect 920 10832 7084 10854
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 3326 10656 3332 10668
rect 1903 10628 3332 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 1210 10548 1216 10600
rect 1268 10588 1274 10600
rect 1581 10591 1639 10597
rect 1581 10588 1593 10591
rect 1268 10560 1593 10588
rect 1268 10548 1274 10560
rect 1581 10557 1593 10560
rect 1627 10557 1639 10591
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 1581 10551 1639 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4338 10588 4344 10600
rect 4299 10560 4344 10588
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 6086 10548 6092 10600
rect 6144 10588 6150 10600
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 6144 10560 6469 10588
rect 6144 10548 6150 10560
rect 6457 10557 6469 10560
rect 6503 10557 6515 10591
rect 6457 10551 6515 10557
rect 3068 10452 3096 10506
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 3476 10492 3617 10520
rect 3476 10480 3482 10492
rect 3605 10489 3617 10492
rect 3651 10489 3663 10523
rect 4614 10520 4620 10532
rect 4575 10492 4620 10520
rect 3605 10483 3663 10489
rect 4614 10480 4620 10492
rect 4672 10480 4678 10532
rect 6365 10523 6423 10529
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 3068 10424 4077 10452
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 5828 10452 5856 10506
rect 6365 10489 6377 10523
rect 6411 10520 6423 10523
rect 16666 10520 16672 10532
rect 6411 10492 16672 10520
rect 6411 10489 6423 10492
rect 6365 10483 6423 10489
rect 16666 10480 16672 10492
rect 16724 10480 16730 10532
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 5828 10424 6653 10452
rect 4065 10415 4123 10421
rect 6641 10421 6653 10424
rect 6687 10421 6699 10455
rect 6641 10415 6699 10421
rect 920 10362 7084 10384
rect 920 10310 3598 10362
rect 3650 10310 3662 10362
rect 3714 10310 3726 10362
rect 3778 10310 3790 10362
rect 3842 10310 7084 10362
rect 920 10288 7084 10310
rect 1228 10220 5764 10248
rect 1228 10124 1256 10220
rect 3326 10180 3332 10192
rect 2714 10152 3332 10180
rect 3326 10140 3332 10152
rect 3384 10140 3390 10192
rect 4154 10140 4160 10192
rect 4212 10140 4218 10192
rect 5736 10180 5764 10220
rect 5994 10180 6000 10192
rect 5736 10152 6000 10180
rect 1210 10112 1216 10124
rect 1123 10084 1216 10112
rect 1210 10072 1216 10084
rect 1268 10072 1274 10124
rect 3418 10112 3424 10124
rect 2746 10084 3424 10112
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 2746 10044 2774 10084
rect 3418 10072 3424 10084
rect 3476 10112 3482 10124
rect 3697 10115 3755 10121
rect 3697 10112 3709 10115
rect 3476 10084 3709 10112
rect 3476 10072 3482 10084
rect 3697 10081 3709 10084
rect 3743 10081 3755 10115
rect 3697 10075 3755 10081
rect 3786 10072 3792 10124
rect 3844 10072 3850 10124
rect 4522 10072 4528 10124
rect 4580 10112 4586 10124
rect 5736 10121 5764 10152
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 5537 10115 5595 10121
rect 5537 10112 5549 10115
rect 4580 10084 5549 10112
rect 4580 10072 4586 10084
rect 5537 10081 5549 10084
rect 5583 10081 5595 10115
rect 5537 10075 5595 10081
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10081 5779 10115
rect 5721 10075 5779 10081
rect 1535 10016 2774 10044
rect 3237 10047 3295 10053
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 3237 10013 3249 10047
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 3804 10044 3832 10072
rect 3375 10016 3832 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 3252 9976 3280 10007
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5077 10047 5135 10053
rect 5077 10044 5089 10047
rect 5040 10016 5089 10044
rect 5040 10004 5046 10016
rect 5077 10013 5089 10016
rect 5123 10013 5135 10047
rect 5552 10044 5580 10075
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 5868 10084 6193 10112
rect 5868 10072 5874 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 5552 10016 6776 10044
rect 5077 10007 5135 10013
rect 3252 9948 3372 9976
rect 3344 9908 3372 9948
rect 4246 9908 4252 9920
rect 3344 9880 4252 9908
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5776 9880 5825 9908
rect 5776 9868 5782 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6748 9917 6776 10016
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 6144 9880 6377 9908
rect 6144 9868 6150 9880
rect 6365 9877 6377 9880
rect 6411 9877 6423 9911
rect 6365 9871 6423 9877
rect 6733 9911 6791 9917
rect 6733 9877 6745 9911
rect 6779 9908 6791 9911
rect 16574 9908 16580 9920
rect 6779 9880 16580 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 920 9818 7084 9840
rect 920 9766 2098 9818
rect 2150 9766 2162 9818
rect 2214 9766 2226 9818
rect 2278 9766 2290 9818
rect 2342 9766 5098 9818
rect 5150 9766 5162 9818
rect 5214 9766 5226 9818
rect 5278 9766 5290 9818
rect 5342 9766 7084 9818
rect 920 9744 7084 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3786 9704 3792 9716
rect 2924 9676 3792 9704
rect 2924 9664 2930 9676
rect 3786 9664 3792 9676
rect 3844 9704 3850 9716
rect 4338 9704 4344 9716
rect 3844 9676 4344 9704
rect 3844 9664 3850 9676
rect 4338 9664 4344 9676
rect 4396 9704 4402 9716
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 4396 9676 6285 9704
rect 4396 9664 4402 9676
rect 6273 9673 6285 9676
rect 6319 9673 6331 9707
rect 6273 9667 6331 9673
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9636 2099 9639
rect 3142 9636 3148 9648
rect 2087 9608 3148 9636
rect 2087 9605 2099 9608
rect 2041 9599 2099 9605
rect 3142 9596 3148 9608
rect 3200 9636 3206 9648
rect 3878 9636 3884 9648
rect 3200 9608 3884 9636
rect 3200 9596 3206 9608
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 6362 9636 6368 9648
rect 5184 9608 6368 9636
rect 1762 9528 1768 9580
rect 1820 9568 1826 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 1820 9540 3525 9568
rect 1820 9528 1826 9540
rect 3513 9537 3525 9540
rect 3559 9568 3571 9571
rect 5184 9568 5212 9608
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 3559 9540 5212 9568
rect 5905 9571 5963 9577
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 5951 9540 12434 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9469 1915 9503
rect 2682 9500 2688 9512
rect 2643 9472 2688 9500
rect 1857 9463 1915 9469
rect 1872 9364 1900 9463
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9469 3755 9503
rect 3697 9463 3755 9469
rect 2225 9435 2283 9441
rect 2225 9401 2237 9435
rect 2271 9432 2283 9435
rect 2406 9432 2412 9444
rect 2271 9404 2412 9432
rect 2271 9401 2283 9404
rect 2225 9395 2283 9401
rect 2406 9392 2412 9404
rect 2464 9392 2470 9444
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 3068 9432 3096 9463
rect 3712 9432 3740 9463
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3844 9472 3893 9500
rect 3844 9460 3850 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 5994 9500 6000 9512
rect 5955 9472 6000 9500
rect 3881 9463 3939 9469
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9469 6147 9503
rect 6089 9463 6147 9469
rect 4062 9432 4068 9444
rect 2648 9404 3648 9432
rect 3712 9404 4068 9432
rect 2648 9392 2654 9404
rect 3050 9364 3056 9376
rect 1872 9336 3056 9364
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3620 9364 3648 9404
rect 4062 9392 4068 9404
rect 4120 9392 4126 9444
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 4212 9404 4257 9432
rect 4212 9392 4218 9404
rect 4982 9364 4988 9376
rect 3620 9336 4988 9364
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5368 9364 5396 9418
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 6104 9432 6132 9463
rect 5500 9404 6132 9432
rect 12406 9432 12434 9540
rect 16574 9432 16580 9444
rect 12406 9404 16580 9432
rect 5500 9392 5506 9404
rect 16574 9392 16580 9404
rect 16632 9392 16638 9444
rect 6270 9364 6276 9376
rect 5368 9336 6276 9364
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 920 9274 7084 9296
rect 920 9222 3598 9274
rect 3650 9222 3662 9274
rect 3714 9222 3726 9274
rect 3778 9222 3790 9274
rect 3842 9222 7084 9274
rect 920 9200 7084 9222
rect 1210 9120 1216 9172
rect 1268 9160 1274 9172
rect 1397 9163 1455 9169
rect 1397 9160 1409 9163
rect 1268 9132 1409 9160
rect 1268 9120 1274 9132
rect 1397 9129 1409 9132
rect 1443 9129 1455 9163
rect 1762 9160 1768 9172
rect 1723 9132 1768 9160
rect 1397 9123 1455 9129
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 4062 9160 4068 9172
rect 2823 9132 4068 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 2590 9092 2596 9104
rect 1688 9064 2596 9092
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 1688 9033 1716 9064
rect 2590 9052 2596 9064
rect 2648 9052 2654 9104
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3418 9092 3424 9104
rect 3191 9064 3424 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 3878 9052 3884 9104
rect 3936 9052 3942 9104
rect 4985 9095 5043 9101
rect 4985 9061 4997 9095
rect 5031 9092 5043 9095
rect 10321 9095 10379 9101
rect 5031 9064 10272 9092
rect 5031 9061 5043 9064
rect 4985 9055 5043 9061
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1912 8996 1961 9024
rect 1912 8984 1918 8996
rect 1949 8993 1961 8996
rect 1995 9024 2007 9027
rect 2317 9027 2375 9033
rect 2317 9024 2329 9027
rect 1995 8996 2329 9024
rect 1995 8993 2007 8996
rect 1949 8987 2007 8993
rect 2317 8993 2329 8996
rect 2363 8993 2375 9027
rect 2317 8987 2375 8993
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 5132 8996 5457 9024
rect 5132 8984 5138 8996
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 8993 5779 9027
rect 5902 9024 5908 9036
rect 5863 8996 5908 9024
rect 5721 8987 5779 8993
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 4890 8956 4896 8968
rect 4851 8928 4896 8956
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 5736 8956 5764 8987
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6362 9024 6368 9036
rect 6323 8996 6368 9024
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6273 8959 6331 8965
rect 5736 8928 6224 8956
rect 6196 8832 6224 8928
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 10244 8956 10272 9064
rect 10321 9061 10333 9095
rect 10367 9092 10379 9095
rect 26326 9092 26332 9104
rect 10367 9064 26332 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 26326 9052 26332 9064
rect 26384 9052 26390 9104
rect 16574 8956 16580 8968
rect 10244 8928 16580 8956
rect 6273 8919 6331 8925
rect 6288 8888 6316 8919
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 6288 8860 7144 8888
rect 1946 8780 1952 8832
rect 2004 8820 2010 8832
rect 2133 8823 2191 8829
rect 2133 8820 2145 8823
rect 2004 8792 2145 8820
rect 2004 8780 2010 8792
rect 2133 8789 2145 8792
rect 2179 8789 2191 8823
rect 2498 8820 2504 8832
rect 2459 8792 2504 8820
rect 2133 8783 2191 8789
rect 2498 8780 2504 8792
rect 2556 8780 2562 8832
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 4430 8820 4436 8832
rect 3016 8792 4436 8820
rect 3016 8780 3022 8792
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 6236 8792 6653 8820
rect 6236 8780 6242 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 6641 8783 6699 8789
rect 920 8730 7084 8752
rect 920 8678 2098 8730
rect 2150 8678 2162 8730
rect 2214 8678 2226 8730
rect 2278 8678 2290 8730
rect 2342 8678 5098 8730
rect 5150 8678 5162 8730
rect 5214 8678 5226 8730
rect 5278 8678 5290 8730
rect 5342 8678 7084 8730
rect 920 8656 7084 8678
rect 1578 8576 1584 8628
rect 1636 8616 1642 8628
rect 1636 8588 2544 8616
rect 1636 8576 1642 8588
rect 2516 8548 2544 8588
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3384 8588 3525 8616
rect 3384 8576 3390 8588
rect 3513 8585 3525 8588
rect 3559 8585 3571 8619
rect 3513 8579 3571 8585
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4120 8588 5304 8616
rect 4120 8576 4126 8588
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 2516 8520 5181 8548
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5276 8548 5304 8588
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5592 8588 5917 8616
rect 5592 8576 5598 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 6270 8616 6276 8628
rect 6231 8588 6276 8616
rect 5905 8579 5963 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 7116 8616 7144 8860
rect 10321 8619 10379 8625
rect 10321 8616 10333 8619
rect 6779 8588 10333 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 10321 8585 10333 8588
rect 10367 8585 10379 8619
rect 10321 8579 10379 8585
rect 26510 8548 26516 8560
rect 5276 8520 26516 8548
rect 5169 8511 5227 8517
rect 26510 8508 26516 8520
rect 26568 8508 26574 8560
rect 1210 8480 1216 8492
rect 1171 8452 1216 8480
rect 1210 8440 1216 8452
rect 1268 8440 1274 8492
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8480 1547 8483
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 1535 8452 3464 8480
rect 1535 8449 1547 8452
rect 1489 8443 1547 8449
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3329 8415 3387 8421
rect 3329 8412 3341 8415
rect 3200 8384 3341 8412
rect 3200 8372 3206 8384
rect 3329 8381 3341 8384
rect 3375 8381 3387 8415
rect 3329 8375 3387 8381
rect 2498 8304 2504 8356
rect 2556 8304 2562 8356
rect 3234 8344 3240 8356
rect 3195 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 3436 8344 3464 8452
rect 3896 8452 6561 8480
rect 3896 8421 3924 8452
rect 6549 8449 6561 8452
rect 6595 8480 6607 8483
rect 26234 8480 26240 8492
rect 6595 8452 26240 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 26234 8440 26240 8452
rect 26292 8440 26298 8492
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 5534 8412 5540 8424
rect 4120 8384 5540 8412
rect 4120 8372 4126 8384
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5718 8412 5724 8424
rect 5679 8384 5724 8412
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 6086 8412 6092 8424
rect 5999 8384 6092 8412
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 4246 8344 4252 8356
rect 3436 8316 4252 8344
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 6104 8344 6132 8372
rect 5552 8316 6132 8344
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 3418 8276 3424 8288
rect 2464 8248 3424 8276
rect 2464 8236 2470 8248
rect 3418 8236 3424 8248
rect 3476 8236 3482 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 5552 8276 5580 8316
rect 16574 8276 16580 8288
rect 4028 8248 5580 8276
rect 12406 8248 16580 8276
rect 4028 8236 4034 8248
rect 920 8186 7084 8208
rect 920 8134 3598 8186
rect 3650 8134 3662 8186
rect 3714 8134 3726 8186
rect 3778 8134 3790 8186
rect 3842 8134 7084 8186
rect 920 8112 7084 8134
rect 3234 8072 3240 8084
rect 1504 8044 3240 8072
rect 1504 8013 1532 8044
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 3476 8044 5396 8072
rect 3476 8032 3482 8044
rect 1489 8007 1547 8013
rect 1489 7973 1501 8007
rect 1535 7973 1547 8007
rect 1489 7967 1547 7973
rect 1946 7964 1952 8016
rect 2004 7964 2010 8016
rect 5368 8004 5396 8044
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 5960 8044 6009 8072
rect 5960 8032 5966 8044
rect 5997 8041 6009 8044
rect 6043 8041 6055 8075
rect 5997 8035 6055 8041
rect 12406 8004 12434 8248
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 1210 7936 1216 7948
rect 1171 7908 1216 7936
rect 1210 7896 1216 7908
rect 1268 7896 1274 7948
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 3329 7939 3387 7945
rect 3329 7936 3341 7939
rect 3108 7908 3341 7936
rect 3108 7896 3114 7908
rect 3329 7905 3341 7908
rect 3375 7936 3387 7939
rect 4246 7936 4252 7948
rect 3375 7908 4108 7936
rect 4207 7908 4252 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 4080 7880 4108 7908
rect 4246 7896 4252 7908
rect 4304 7896 4310 7948
rect 5276 7936 5304 7990
rect 5368 7976 12434 8004
rect 5994 7936 6000 7948
rect 5276 7908 6000 7936
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7936 6147 7939
rect 6135 7908 6776 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 3234 7868 3240 7880
rect 3195 7840 3240 7868
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3881 7871 3939 7877
rect 3881 7837 3893 7871
rect 3927 7837 3939 7871
rect 3881 7831 3939 7837
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 3513 7735 3571 7741
rect 3513 7732 3525 7735
rect 1912 7704 3525 7732
rect 1912 7692 1918 7704
rect 3513 7701 3525 7704
rect 3559 7701 3571 7735
rect 3896 7732 3924 7831
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 6104 7868 6132 7899
rect 5684 7840 6132 7868
rect 5684 7828 5690 7840
rect 4246 7732 4252 7744
rect 3896 7704 4252 7732
rect 3513 7695 3571 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6748 7741 6776 7908
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 16666 7868 16672 7880
rect 6880 7840 16672 7868
rect 6880 7828 6886 7840
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 6273 7735 6331 7741
rect 6273 7732 6285 7735
rect 5960 7704 6285 7732
rect 5960 7692 5966 7704
rect 6273 7701 6285 7704
rect 6319 7701 6331 7735
rect 6273 7695 6331 7701
rect 6733 7735 6791 7741
rect 6733 7701 6745 7735
rect 6779 7732 6791 7735
rect 16574 7732 16580 7744
rect 6779 7704 16580 7732
rect 6779 7701 6791 7704
rect 6733 7695 6791 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 920 7642 7084 7664
rect 920 7590 2098 7642
rect 2150 7590 2162 7642
rect 2214 7590 2226 7642
rect 2278 7590 2290 7642
rect 2342 7590 5098 7642
rect 5150 7590 5162 7642
rect 5214 7590 5226 7642
rect 5278 7590 5290 7642
rect 5342 7590 7084 7642
rect 920 7568 7084 7590
rect 3605 7531 3663 7537
rect 3605 7497 3617 7531
rect 3651 7528 3663 7531
rect 3878 7528 3884 7540
rect 3651 7500 3884 7528
rect 3651 7497 3663 7500
rect 3605 7491 3663 7497
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6052 7500 6653 7528
rect 6052 7488 6058 7500
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 3234 7392 3240 7404
rect 1627 7364 3240 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 1305 7327 1363 7333
rect 1305 7293 1317 7327
rect 1351 7293 1363 7327
rect 1305 7287 1363 7293
rect 3421 7327 3479 7333
rect 3421 7293 3433 7327
rect 3467 7324 3479 7327
rect 3970 7324 3976 7336
rect 3467 7296 3976 7324
rect 3467 7293 3479 7296
rect 3421 7287 3479 7293
rect 1210 7148 1216 7200
rect 1268 7188 1274 7200
rect 1320 7188 1348 7287
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7293 4399 7327
rect 6454 7324 6460 7336
rect 6415 7296 6460 7324
rect 4341 7287 4399 7293
rect 2314 7216 2320 7268
rect 2372 7216 2378 7268
rect 3326 7256 3332 7268
rect 3287 7228 3332 7256
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 4356 7256 4384 7287
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 3528 7228 4384 7256
rect 4617 7259 4675 7265
rect 3528 7188 3556 7228
rect 4617 7225 4629 7259
rect 4663 7256 4675 7259
rect 4706 7256 4712 7268
rect 4663 7228 4712 7256
rect 4663 7225 4675 7228
rect 4617 7219 4675 7225
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 6365 7259 6423 7265
rect 5460 7200 5488 7242
rect 6365 7225 6377 7259
rect 6411 7256 6423 7259
rect 6730 7256 6736 7268
rect 6411 7228 6736 7256
rect 6411 7225 6423 7228
rect 6365 7219 6423 7225
rect 6730 7216 6736 7228
rect 6788 7256 6794 7268
rect 26418 7256 26424 7268
rect 6788 7228 26424 7256
rect 6788 7216 6794 7228
rect 26418 7216 26424 7228
rect 26476 7216 26482 7268
rect 4154 7188 4160 7200
rect 1268 7160 3556 7188
rect 4115 7160 4160 7188
rect 1268 7148 1274 7160
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 5442 7148 5448 7200
rect 5500 7148 5506 7200
rect 920 7098 7084 7120
rect 920 7046 3598 7098
rect 3650 7046 3662 7098
rect 3714 7046 3726 7098
rect 3778 7046 3790 7098
rect 3842 7046 7084 7098
rect 920 7024 7084 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 2372 6956 2421 6984
rect 2372 6944 2378 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 4154 6944 4160 6996
rect 4212 6944 4218 6996
rect 5810 6984 5816 6996
rect 5552 6956 5816 6984
rect 3234 6916 3240 6928
rect 3195 6888 3240 6916
rect 3234 6876 3240 6888
rect 3292 6876 3298 6928
rect 4172 6902 4200 6944
rect 5552 6916 5580 6956
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 5905 6919 5963 6925
rect 5905 6916 5917 6919
rect 5460 6888 5580 6916
rect 5644 6888 5917 6916
rect 1854 6848 1860 6860
rect 1815 6820 1860 6848
rect 1854 6808 1860 6820
rect 1912 6848 1918 6860
rect 5460 6857 5488 6888
rect 2225 6851 2283 6857
rect 2225 6848 2237 6851
rect 1912 6820 2237 6848
rect 1912 6808 1918 6820
rect 2225 6817 2237 6820
rect 2271 6817 2283 6851
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 2225 6811 2283 6817
rect 4448 6820 5089 6848
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2041 6647 2099 6653
rect 2041 6644 2053 6647
rect 2004 6616 2053 6644
rect 2004 6604 2010 6616
rect 2041 6613 2053 6616
rect 2087 6613 2099 6647
rect 2976 6644 3004 6743
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4448 6780 4476 6820
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6848 5595 6851
rect 5644 6848 5672 6888
rect 5905 6885 5917 6888
rect 5951 6885 5963 6919
rect 5905 6879 5963 6885
rect 5583 6820 5672 6848
rect 6733 6851 6791 6857
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 6733 6817 6745 6851
rect 6779 6848 6791 6851
rect 6822 6848 6828 6860
rect 6779 6820 6828 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 4028 6752 4476 6780
rect 4985 6783 5043 6789
rect 4028 6740 4034 6752
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5626 6780 5632 6792
rect 5031 6752 5632 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 5810 6780 5816 6792
rect 5771 6752 5816 6780
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 6086 6780 6092 6792
rect 6047 6752 6092 6780
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 4890 6672 4896 6724
rect 4948 6712 4954 6724
rect 16666 6712 16672 6724
rect 4948 6684 16672 6712
rect 4948 6672 4954 6684
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 4338 6644 4344 6656
rect 2976 6616 4344 6644
rect 2041 6607 2099 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5718 6644 5724 6656
rect 5307 6616 5724 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6822 6644 6828 6656
rect 5868 6616 6828 6644
rect 5868 6604 5874 6616
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 920 6554 7084 6576
rect 920 6502 2098 6554
rect 2150 6502 2162 6554
rect 2214 6502 2226 6554
rect 2278 6502 2290 6554
rect 2342 6502 5098 6554
rect 5150 6502 5162 6554
rect 5214 6502 5226 6554
rect 5278 6502 5290 6554
rect 5342 6502 7084 6554
rect 920 6480 7084 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 5810 6440 5816 6452
rect 2740 6412 5816 6440
rect 2740 6400 2746 6412
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 3326 6304 3332 6316
rect 1535 6276 3332 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 3326 6264 3332 6276
rect 3384 6304 3390 6316
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 3384 6276 4537 6304
rect 3384 6264 3390 6276
rect 4525 6273 4537 6276
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 1210 6236 1216 6248
rect 1171 6208 1216 6236
rect 1210 6196 1216 6208
rect 1268 6196 1274 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3344 6208 3433 6236
rect 3344 6180 3372 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6205 4307 6239
rect 5736 6236 5764 6264
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5736 6208 6377 6236
rect 4249 6199 4307 6205
rect 6365 6205 6377 6208
rect 6411 6236 6423 6239
rect 6454 6236 6460 6248
rect 6411 6208 6460 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 1946 6128 1952 6180
rect 2004 6128 2010 6180
rect 3237 6171 3295 6177
rect 3237 6137 3249 6171
rect 3283 6137 3295 6171
rect 3237 6131 3295 6137
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 3252 6100 3280 6131
rect 3326 6128 3332 6180
rect 3384 6128 3390 6180
rect 4264 6168 4292 6199
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 6273 6171 6331 6177
rect 4264 6140 4384 6168
rect 4356 6112 4384 6140
rect 1544 6072 3280 6100
rect 1544 6060 1550 6072
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3476 6072 3617 6100
rect 3476 6060 3482 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 3605 6063 3663 6069
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4522 6100 4528 6112
rect 4396 6072 4528 6100
rect 4396 6060 4402 6072
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 5736 6100 5764 6154
rect 6273 6137 6285 6171
rect 6319 6168 6331 6171
rect 16574 6168 16580 6180
rect 6319 6140 16580 6168
rect 6319 6137 6331 6140
rect 6273 6131 6331 6137
rect 16574 6128 16580 6140
rect 16632 6128 16638 6180
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 5736 6072 6561 6100
rect 6549 6069 6561 6072
rect 6595 6069 6607 6103
rect 6549 6063 6607 6069
rect 920 6010 7084 6032
rect 920 5958 3598 6010
rect 3650 5958 3662 6010
rect 3714 5958 3726 6010
rect 3778 5958 3790 6010
rect 3842 5958 7084 6010
rect 920 5936 7084 5958
rect 1854 5856 1860 5908
rect 1912 5896 1918 5908
rect 5169 5899 5227 5905
rect 1912 5868 2084 5896
rect 1912 5856 1918 5868
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1741 5763 1799 5769
rect 1741 5760 1753 5763
rect 1636 5732 1753 5760
rect 1636 5720 1642 5732
rect 1741 5729 1753 5732
rect 1787 5729 1799 5763
rect 1741 5723 1799 5729
rect 1882 5763 1940 5769
rect 1882 5729 1894 5763
rect 1928 5760 1940 5763
rect 2056 5760 2084 5868
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5442 5896 5448 5908
rect 5215 5868 5448 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6730 5896 6736 5908
rect 6691 5868 6736 5896
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 3142 5828 3148 5840
rect 2240 5800 3148 5828
rect 2240 5769 2268 5800
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 3418 5788 3424 5840
rect 3476 5788 3482 5840
rect 4614 5828 4620 5840
rect 4575 5800 4620 5828
rect 4614 5788 4620 5800
rect 4672 5788 4678 5840
rect 5902 5828 5908 5840
rect 5863 5800 5908 5828
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 1928 5732 2084 5760
rect 2225 5763 2283 5769
rect 1928 5729 1940 5732
rect 1882 5723 1940 5729
rect 2225 5729 2237 5763
rect 2271 5729 2283 5763
rect 2225 5723 2283 5729
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4985 5763 5043 5769
rect 4985 5760 4997 5763
rect 4212 5732 4997 5760
rect 4212 5720 4218 5732
rect 4985 5729 4997 5732
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 5353 5763 5411 5769
rect 5353 5729 5365 5763
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 2590 5692 2596 5704
rect 1596 5664 2596 5692
rect 1302 5584 1308 5636
rect 1360 5624 1366 5636
rect 1596 5633 1624 5664
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 4246 5692 4252 5704
rect 2915 5664 4252 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 5368 5692 5396 5723
rect 5813 5695 5871 5701
rect 5368 5664 5764 5692
rect 5736 5636 5764 5664
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 6086 5692 6092 5704
rect 5859 5664 6092 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 6638 5692 6644 5704
rect 6503 5664 6644 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 1581 5627 1639 5633
rect 1581 5624 1593 5627
rect 1360 5596 1593 5624
rect 1360 5584 1366 5596
rect 1581 5593 1593 5596
rect 1627 5593 1639 5627
rect 1581 5587 1639 5593
rect 5718 5584 5724 5636
rect 5776 5584 5782 5636
rect 1946 5516 1952 5568
rect 2004 5556 2010 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 2004 5528 2053 5556
rect 2004 5516 2010 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2406 5556 2412 5568
rect 2367 5528 2412 5556
rect 2041 5519 2099 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 4798 5556 4804 5568
rect 4759 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 920 5466 7084 5488
rect 920 5414 2098 5466
rect 2150 5414 2162 5466
rect 2214 5414 2226 5466
rect 2278 5414 2290 5466
rect 2342 5414 5098 5466
rect 5150 5414 5162 5466
rect 5214 5414 5226 5466
rect 5278 5414 5290 5466
rect 5342 5414 7084 5466
rect 920 5392 7084 5414
rect 4982 5312 4988 5364
rect 5040 5352 5046 5364
rect 6730 5352 6736 5364
rect 5040 5324 6736 5352
rect 5040 5312 5046 5324
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 1210 5216 1216 5228
rect 1171 5188 1216 5216
rect 1210 5176 1216 5188
rect 1268 5176 1274 5228
rect 1486 5216 1492 5228
rect 1447 5188 1492 5216
rect 1486 5176 1492 5188
rect 1544 5176 1550 5228
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 2740 5188 3249 5216
rect 2740 5176 2746 5188
rect 3237 5185 3249 5188
rect 3283 5185 3295 5219
rect 4062 5216 4068 5228
rect 3237 5179 3295 5185
rect 3344 5188 4068 5216
rect 3344 5157 3372 5188
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4798 5216 4804 5228
rect 4356 5188 4804 5216
rect 4356 5157 4384 5188
rect 4798 5176 4804 5188
rect 4856 5216 4862 5228
rect 4856 5188 6776 5216
rect 4856 5176 4862 5188
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3973 5151 4031 5157
rect 3973 5148 3985 5151
rect 3329 5111 3387 5117
rect 3528 5120 3985 5148
rect 1946 5040 1952 5092
rect 2004 5040 2010 5092
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3528 5021 3556 5120
rect 3973 5117 3985 5120
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 4580 5120 4629 5148
rect 4580 5108 4586 5120
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 4982 5148 4988 5160
rect 4943 5120 4988 5148
rect 4617 5111 4675 5117
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5534 5040 5540 5092
rect 5592 5040 5598 5092
rect 3513 5015 3571 5021
rect 3513 5012 3525 5015
rect 3384 4984 3525 5012
rect 3384 4972 3390 4984
rect 3513 4981 3525 4984
rect 3559 4981 3571 5015
rect 4154 5012 4160 5024
rect 4115 4984 4160 5012
rect 3513 4975 3571 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 5442 5012 5448 5024
rect 4479 4984 5448 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 6748 5021 6776 5188
rect 6733 5015 6791 5021
rect 6733 4981 6745 5015
rect 6779 5012 6791 5015
rect 16574 5012 16580 5024
rect 6779 4984 16580 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 920 4922 7084 4944
rect 920 4870 3598 4922
rect 3650 4870 3662 4922
rect 3714 4870 3726 4922
rect 3778 4870 3790 4922
rect 3842 4870 7084 4922
rect 920 4848 7084 4870
rect 2406 4768 2412 4820
rect 2464 4768 2470 4820
rect 2590 4768 2596 4820
rect 2648 4808 2654 4820
rect 4614 4808 4620 4820
rect 2648 4780 3464 4808
rect 2648 4768 2654 4780
rect 2424 4726 2452 4768
rect 3436 4684 3464 4780
rect 3712 4780 4620 4808
rect 3712 4749 3740 4780
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 3697 4743 3755 4749
rect 3697 4709 3709 4743
rect 3743 4709 3755 4743
rect 3697 4703 3755 4709
rect 4154 4700 4160 4752
rect 4212 4700 4218 4752
rect 1302 4672 1308 4684
rect 1263 4644 1308 4672
rect 1302 4632 1308 4644
rect 1360 4632 1366 4684
rect 3418 4672 3424 4684
rect 3331 4644 3424 4672
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 5994 4672 6000 4684
rect 5955 4644 6000 4672
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6454 4672 6460 4684
rect 6367 4644 6460 4672
rect 6454 4632 6460 4644
rect 6512 4672 6518 4684
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6512 4644 6745 4672
rect 6512 4632 6518 4644
rect 6733 4641 6745 4644
rect 6779 4672 6791 4675
rect 16574 4672 16580 4684
rect 6779 4644 16580 4672
rect 6779 4641 6791 4644
rect 6733 4635 6791 4641
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 1946 4604 1952 4616
rect 1627 4576 1952 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1946 4564 1952 4576
rect 2004 4604 2010 4616
rect 2590 4604 2596 4616
rect 2004 4576 2596 4604
rect 2004 4564 2010 4576
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 3344 4468 3372 4567
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 4212 4576 5457 4604
rect 4212 4564 4218 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 5810 4536 5816 4548
rect 5771 4508 5816 4536
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 4246 4468 4252 4480
rect 3344 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 5626 4468 5632 4480
rect 5587 4440 5632 4468
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 920 4378 7084 4400
rect 920 4326 2098 4378
rect 2150 4326 2162 4378
rect 2214 4326 2226 4378
rect 2278 4326 2290 4378
rect 2342 4326 5098 4378
rect 5150 4326 5162 4378
rect 5214 4326 5226 4378
rect 5278 4326 5290 4378
rect 5342 4326 7084 4378
rect 920 4304 7084 4326
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 6052 4236 6469 4264
rect 6052 4224 6058 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 16666 4264 16672 4276
rect 6457 4227 6515 4233
rect 12406 4236 16672 4264
rect 2590 4156 2596 4208
rect 2648 4196 2654 4208
rect 2648 4168 2820 4196
rect 2648 4156 2654 4168
rect 1210 4128 1216 4140
rect 1171 4100 1216 4128
rect 1210 4088 1216 4100
rect 1268 4088 1274 4140
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 2682 4128 2688 4140
rect 1535 4100 2688 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 2792 4128 2820 4168
rect 5626 4156 5632 4208
rect 5684 4196 5690 4208
rect 6546 4196 6552 4208
rect 5684 4168 6552 4196
rect 5684 4156 5690 4168
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 2792 4100 3249 4128
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3476 4100 3893 4128
rect 3476 4088 3482 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 4154 4128 4160 4140
rect 4115 4100 4160 4128
rect 3881 4091 3939 4097
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 4764 4100 5396 4128
rect 4764 4088 4770 4100
rect 3326 4060 3332 4072
rect 3239 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 5368 4060 5396 4100
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5500 4100 6224 4128
rect 5500 4088 5506 4100
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5368 4032 5917 4060
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 6086 4060 6092 4072
rect 6047 4032 6092 4060
rect 5905 4023 5963 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6196 4069 6224 4100
rect 6288 4069 6316 4168
rect 6546 4156 6552 4168
rect 6604 4196 6610 4208
rect 12406 4196 12434 4236
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 6604 4168 12434 4196
rect 6604 4156 6610 4168
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4029 6239 4063
rect 6181 4023 6239 4029
rect 6273 4063 6331 4069
rect 6273 4029 6285 4063
rect 6319 4029 6331 4063
rect 6273 4023 6331 4029
rect 3344 3992 3372 4020
rect 2700 3924 2728 3978
rect 3344 3964 4646 3992
rect 3513 3927 3571 3933
rect 3513 3924 3525 3927
rect 2700 3896 3525 3924
rect 3513 3893 3525 3896
rect 3559 3893 3571 3927
rect 3513 3887 3571 3893
rect 920 3834 7084 3856
rect 920 3782 3598 3834
rect 3650 3782 3662 3834
rect 3714 3782 3726 3834
rect 3778 3782 3790 3834
rect 3842 3782 7084 3834
rect 920 3760 7084 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3689 2191 3723
rect 2133 3683 2191 3689
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 2148 3652 2176 3683
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 16574 3720 16580 3732
rect 2372 3692 3924 3720
rect 2372 3680 2378 3692
rect 1728 3624 2084 3652
rect 2148 3624 3082 3652
rect 1728 3612 1734 3624
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3553 2007 3587
rect 2056 3584 2084 3624
rect 2314 3584 2320 3596
rect 2056 3556 2320 3584
rect 1949 3547 2007 3553
rect 1964 3380 1992 3547
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2682 3516 2688 3528
rect 2639 3488 2688 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 3896 3516 3924 3692
rect 4356 3692 16580 3720
rect 4356 3661 4384 3692
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 4341 3655 4399 3661
rect 4341 3621 4353 3655
rect 4387 3621 4399 3655
rect 4709 3655 4767 3661
rect 4709 3652 4721 3655
rect 4341 3615 4399 3621
rect 4448 3624 4721 3652
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4448 3584 4476 3624
rect 4709 3621 4721 3624
rect 4755 3621 4767 3655
rect 6454 3652 6460 3664
rect 6415 3624 6460 3652
rect 4709 3615 4767 3621
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 4212 3556 4476 3584
rect 4212 3544 4218 3556
rect 5810 3544 5816 3596
rect 5868 3544 5874 3596
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 3896 3488 4445 3516
rect 4433 3485 4445 3488
rect 4479 3516 4491 3519
rect 4479 3488 4568 3516
rect 4479 3485 4491 3488
rect 4433 3479 4491 3485
rect 4540 3392 4568 3488
rect 3050 3380 3056 3392
rect 1964 3352 3056 3380
rect 3050 3340 3056 3352
rect 3108 3380 3114 3392
rect 3326 3380 3332 3392
rect 3108 3352 3332 3380
rect 3108 3340 3114 3352
rect 3326 3340 3332 3352
rect 3384 3380 3390 3392
rect 4062 3380 4068 3392
rect 3384 3352 4068 3380
rect 3384 3340 3390 3352
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 6086 3340 6092 3392
rect 6144 3380 6150 3392
rect 6733 3383 6791 3389
rect 6733 3380 6745 3383
rect 6144 3352 6745 3380
rect 6144 3340 6150 3352
rect 6733 3349 6745 3352
rect 6779 3380 6791 3383
rect 16666 3380 16672 3392
rect 6779 3352 16672 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 920 3290 7084 3312
rect 920 3238 2098 3290
rect 2150 3238 2162 3290
rect 2214 3238 2226 3290
rect 2278 3238 2290 3290
rect 2342 3238 5098 3290
rect 5150 3238 5162 3290
rect 5214 3238 5226 3290
rect 5278 3238 5290 3290
rect 5342 3238 7084 3290
rect 920 3216 7084 3238
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 6546 3176 6552 3188
rect 3936 3148 5580 3176
rect 6507 3148 6552 3176
rect 3936 3136 3942 3148
rect 5552 3108 5580 3148
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 16574 3176 16580 3188
rect 12406 3148 16580 3176
rect 12406 3108 12434 3148
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 5552 3080 12434 3108
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1544 3012 1961 3040
rect 1544 3000 1550 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 16574 3040 16580 3052
rect 3743 3012 16580 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 1670 2972 1676 2984
rect 1631 2944 1676 2972
rect 1670 2932 1676 2944
rect 1728 2932 1734 2984
rect 3881 2975 3939 2981
rect 3082 2944 3832 2972
rect 3804 2904 3832 2944
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 4062 2972 4068 2984
rect 3927 2944 4068 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2972 4491 2975
rect 4522 2972 4528 2984
rect 4479 2944 4528 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 4764 2944 4813 2972
rect 4764 2932 4770 2944
rect 4801 2941 4813 2944
rect 4847 2941 4859 2975
rect 4801 2935 4859 2941
rect 3970 2904 3976 2916
rect 3804 2876 3976 2904
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 5534 2864 5540 2916
rect 5592 2864 5598 2916
rect 4062 2836 4068 2848
rect 4023 2808 4068 2836
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 6730 2836 6736 2848
rect 6691 2808 6736 2836
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 920 2746 7084 2768
rect 920 2694 3598 2746
rect 3650 2694 3662 2746
rect 3714 2694 3726 2746
rect 3778 2694 3790 2746
rect 3842 2694 7084 2746
rect 920 2672 7084 2694
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 5534 2632 5540 2644
rect 5491 2604 5540 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 1946 2564 1952 2576
rect 1907 2536 1952 2564
rect 1946 2524 1952 2536
rect 2004 2524 2010 2576
rect 4062 2564 4068 2576
rect 3174 2536 4068 2564
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 5994 2564 6000 2576
rect 5955 2536 6000 2564
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 3697 2499 3755 2505
rect 3697 2465 3709 2499
rect 3743 2496 3755 2499
rect 3786 2496 3792 2508
rect 3743 2468 3792 2496
rect 3743 2465 3755 2468
rect 3697 2459 3755 2465
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2465 3939 2499
rect 3881 2459 3939 2465
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 5626 2496 5632 2508
rect 5307 2468 5632 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3896 2428 3924 2459
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 6181 2499 6239 2505
rect 6181 2465 6193 2499
rect 6227 2496 6239 2499
rect 6730 2496 6736 2508
rect 6227 2468 6736 2496
rect 6227 2465 6239 2468
rect 6181 2459 6239 2465
rect 6730 2456 6736 2468
rect 6788 2496 6794 2508
rect 16574 2496 16580 2508
rect 6788 2468 16580 2496
rect 6788 2456 6794 2468
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 4982 2428 4988 2440
rect 3476 2400 3924 2428
rect 4943 2400 4988 2428
rect 3476 2388 3482 2400
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 4065 2363 4123 2369
rect 4065 2360 4077 2363
rect 4028 2332 4077 2360
rect 4028 2320 4034 2332
rect 4065 2329 4077 2332
rect 4111 2329 4123 2363
rect 4065 2323 4123 2329
rect 4430 2320 4436 2372
rect 4488 2360 4494 2372
rect 4488 2332 6316 2360
rect 4488 2320 4494 2332
rect 5169 2295 5227 2301
rect 5169 2261 5181 2295
rect 5215 2292 5227 2295
rect 5442 2292 5448 2304
rect 5215 2264 5448 2292
rect 5215 2261 5227 2264
rect 5169 2255 5227 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 6288 2301 6316 2332
rect 6273 2295 6331 2301
rect 6273 2261 6285 2295
rect 6319 2261 6331 2295
rect 6273 2255 6331 2261
rect 920 2202 7084 2224
rect 920 2150 2098 2202
rect 2150 2150 2162 2202
rect 2214 2150 2226 2202
rect 2278 2150 2290 2202
rect 2342 2150 5098 2202
rect 5150 2150 5162 2202
rect 5214 2150 5226 2202
rect 5278 2150 5290 2202
rect 5342 2150 7084 2202
rect 920 2128 7084 2150
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 16666 1340 16672 1352
rect 5040 1312 16672 1340
rect 5040 1300 5046 1312
rect 16666 1300 16672 1312
rect 16724 1300 16730 1352
rect 5442 1232 5448 1284
rect 5500 1272 5506 1284
rect 16758 1272 16764 1284
rect 5500 1244 16764 1272
rect 5500 1232 5506 1244
rect 16758 1232 16764 1244
rect 16816 1232 16822 1284
rect 6638 1164 6644 1216
rect 6696 1204 6702 1216
rect 16574 1204 16580 1216
rect 6696 1176 16580 1204
rect 6696 1164 6702 1176
rect 16574 1164 16580 1176
rect 16632 1164 16638 1216
<< via1 >>
rect 6460 12452 6512 12504
rect 16580 12452 16632 12504
rect 3598 11398 3650 11450
rect 3662 11398 3714 11450
rect 3726 11398 3778 11450
rect 3790 11398 3842 11450
rect 4528 11296 4580 11348
rect 4712 11296 4764 11348
rect 6828 11296 6880 11348
rect 3332 11271 3384 11280
rect 3332 11237 3341 11271
rect 3341 11237 3375 11271
rect 3375 11237 3384 11271
rect 3332 11228 3384 11237
rect 16580 11228 16632 11280
rect 3976 11203 4028 11212
rect 3976 11169 3985 11203
rect 3985 11169 4019 11203
rect 4019 11169 4028 11203
rect 3976 11160 4028 11169
rect 4528 11160 4580 11212
rect 4712 11203 4764 11212
rect 4712 11169 4721 11203
rect 4721 11169 4755 11203
rect 4755 11169 4764 11203
rect 4712 11160 4764 11169
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 4160 11067 4212 11076
rect 4160 11033 4169 11067
rect 4169 11033 4203 11067
rect 4203 11033 4212 11067
rect 4160 11024 4212 11033
rect 5448 11024 5500 11076
rect 4712 10956 4764 11008
rect 2098 10854 2150 10906
rect 2162 10854 2214 10906
rect 2226 10854 2278 10906
rect 2290 10854 2342 10906
rect 5098 10854 5150 10906
rect 5162 10854 5214 10906
rect 5226 10854 5278 10906
rect 5290 10854 5342 10906
rect 3332 10616 3384 10668
rect 1216 10548 1268 10600
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4344 10591 4396 10600
rect 4344 10557 4353 10591
rect 4353 10557 4387 10591
rect 4387 10557 4396 10591
rect 4344 10548 4396 10557
rect 6092 10548 6144 10600
rect 3424 10480 3476 10532
rect 4620 10523 4672 10532
rect 4620 10489 4629 10523
rect 4629 10489 4663 10523
rect 4663 10489 4672 10523
rect 4620 10480 4672 10489
rect 16672 10480 16724 10532
rect 3598 10310 3650 10362
rect 3662 10310 3714 10362
rect 3726 10310 3778 10362
rect 3790 10310 3842 10362
rect 3332 10140 3384 10192
rect 4160 10140 4212 10192
rect 1216 10115 1268 10124
rect 1216 10081 1225 10115
rect 1225 10081 1259 10115
rect 1259 10081 1268 10115
rect 1216 10072 1268 10081
rect 3424 10072 3476 10124
rect 3792 10072 3844 10124
rect 4528 10072 4580 10124
rect 6000 10140 6052 10192
rect 4988 10004 5040 10056
rect 5816 10072 5868 10124
rect 4252 9868 4304 9920
rect 5724 9868 5776 9920
rect 6092 9868 6144 9920
rect 16580 9868 16632 9920
rect 2098 9766 2150 9818
rect 2162 9766 2214 9818
rect 2226 9766 2278 9818
rect 2290 9766 2342 9818
rect 5098 9766 5150 9818
rect 5162 9766 5214 9818
rect 5226 9766 5278 9818
rect 5290 9766 5342 9818
rect 2872 9664 2924 9716
rect 3792 9664 3844 9716
rect 4344 9664 4396 9716
rect 3148 9596 3200 9648
rect 3884 9596 3936 9648
rect 1768 9528 1820 9580
rect 6368 9596 6420 9648
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 2412 9392 2464 9444
rect 2596 9392 2648 9444
rect 3792 9460 3844 9512
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 3056 9324 3108 9376
rect 4068 9392 4120 9444
rect 4160 9435 4212 9444
rect 4160 9401 4169 9435
rect 4169 9401 4203 9435
rect 4203 9401 4212 9435
rect 4160 9392 4212 9401
rect 4988 9324 5040 9376
rect 5448 9392 5500 9444
rect 16580 9392 16632 9444
rect 6276 9324 6328 9376
rect 3598 9222 3650 9274
rect 3662 9222 3714 9274
rect 3726 9222 3778 9274
rect 3790 9222 3842 9274
rect 1216 9120 1268 9172
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 4068 9120 4120 9172
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 2596 9052 2648 9104
rect 3424 9052 3476 9104
rect 3884 9052 3936 9104
rect 1860 8984 1912 9036
rect 5080 8984 5132 9036
rect 5908 9027 5960 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 26332 9052 26384 9104
rect 16580 8916 16632 8968
rect 1952 8780 2004 8832
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 2964 8780 3016 8832
rect 4436 8780 4488 8832
rect 6184 8780 6236 8832
rect 2098 8678 2150 8730
rect 2162 8678 2214 8730
rect 2226 8678 2278 8730
rect 2290 8678 2342 8730
rect 5098 8678 5150 8730
rect 5162 8678 5214 8730
rect 5226 8678 5278 8730
rect 5290 8678 5342 8730
rect 1584 8576 1636 8628
rect 3332 8576 3384 8628
rect 4068 8576 4120 8628
rect 5540 8576 5592 8628
rect 6276 8619 6328 8628
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 26516 8508 26568 8560
rect 1216 8483 1268 8492
rect 1216 8449 1225 8483
rect 1225 8449 1259 8483
rect 1259 8449 1268 8483
rect 1216 8440 1268 8449
rect 3148 8372 3200 8424
rect 2504 8304 2556 8356
rect 3240 8347 3292 8356
rect 3240 8313 3249 8347
rect 3249 8313 3283 8347
rect 3283 8313 3292 8347
rect 3240 8304 3292 8313
rect 26240 8440 26292 8492
rect 4068 8372 4120 8424
rect 5540 8372 5592 8424
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 4252 8304 4304 8356
rect 2412 8236 2464 8288
rect 3424 8236 3476 8288
rect 3976 8236 4028 8288
rect 3598 8134 3650 8186
rect 3662 8134 3714 8186
rect 3726 8134 3778 8186
rect 3790 8134 3842 8186
rect 3240 8032 3292 8084
rect 3424 8032 3476 8084
rect 1952 7964 2004 8016
rect 5908 8032 5960 8084
rect 16580 8236 16632 8288
rect 1216 7939 1268 7948
rect 1216 7905 1225 7939
rect 1225 7905 1259 7939
rect 1259 7905 1268 7939
rect 1216 7896 1268 7905
rect 3056 7896 3108 7948
rect 4252 7939 4304 7948
rect 4252 7905 4261 7939
rect 4261 7905 4295 7939
rect 4295 7905 4304 7939
rect 4252 7896 4304 7905
rect 6000 7896 6052 7948
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 1860 7692 1912 7744
rect 4068 7828 4120 7880
rect 5632 7828 5684 7880
rect 4252 7692 4304 7744
rect 5908 7692 5960 7744
rect 6828 7828 6880 7880
rect 16672 7828 16724 7880
rect 16580 7692 16632 7744
rect 2098 7590 2150 7642
rect 2162 7590 2214 7642
rect 2226 7590 2278 7642
rect 2290 7590 2342 7642
rect 5098 7590 5150 7642
rect 5162 7590 5214 7642
rect 5226 7590 5278 7642
rect 5290 7590 5342 7642
rect 3884 7488 3936 7540
rect 6000 7488 6052 7540
rect 3240 7352 3292 7404
rect 3976 7327 4028 7336
rect 1216 7148 1268 7200
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 6460 7327 6512 7336
rect 2320 7216 2372 7268
rect 3332 7259 3384 7268
rect 3332 7225 3341 7259
rect 3341 7225 3375 7259
rect 3375 7225 3384 7259
rect 3332 7216 3384 7225
rect 6460 7293 6469 7327
rect 6469 7293 6503 7327
rect 6503 7293 6512 7327
rect 6460 7284 6512 7293
rect 4712 7216 4764 7268
rect 6736 7216 6788 7268
rect 26424 7216 26476 7268
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 5448 7148 5500 7200
rect 3598 7046 3650 7098
rect 3662 7046 3714 7098
rect 3726 7046 3778 7098
rect 3790 7046 3842 7098
rect 2320 6944 2372 6996
rect 4160 6944 4212 6996
rect 3240 6919 3292 6928
rect 3240 6885 3249 6919
rect 3249 6885 3283 6919
rect 3283 6885 3292 6919
rect 3240 6876 3292 6885
rect 5816 6944 5868 6996
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 1952 6604 2004 6656
rect 3976 6740 4028 6792
rect 6828 6808 6880 6860
rect 5632 6740 5684 6792
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 4896 6672 4948 6724
rect 16672 6672 16724 6724
rect 4344 6604 4396 6656
rect 5724 6604 5776 6656
rect 5816 6604 5868 6656
rect 6828 6604 6880 6656
rect 2098 6502 2150 6554
rect 2162 6502 2214 6554
rect 2226 6502 2278 6554
rect 2290 6502 2342 6554
rect 5098 6502 5150 6554
rect 5162 6502 5214 6554
rect 5226 6502 5278 6554
rect 5290 6502 5342 6554
rect 2688 6400 2740 6452
rect 5816 6400 5868 6452
rect 3332 6264 3384 6316
rect 5724 6264 5776 6316
rect 1216 6239 1268 6248
rect 1216 6205 1225 6239
rect 1225 6205 1259 6239
rect 1259 6205 1268 6239
rect 1216 6196 1268 6205
rect 1952 6128 2004 6180
rect 1492 6060 1544 6112
rect 3332 6128 3384 6180
rect 6460 6196 6512 6248
rect 3424 6060 3476 6112
rect 4344 6060 4396 6112
rect 4528 6060 4580 6112
rect 16580 6128 16632 6180
rect 3598 5958 3650 6010
rect 3662 5958 3714 6010
rect 3726 5958 3778 6010
rect 3790 5958 3842 6010
rect 1860 5856 1912 5908
rect 1584 5720 1636 5772
rect 5448 5856 5500 5908
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 3148 5788 3200 5840
rect 3424 5788 3476 5840
rect 4620 5831 4672 5840
rect 4620 5797 4629 5831
rect 4629 5797 4663 5831
rect 4663 5797 4672 5831
rect 4620 5788 4672 5797
rect 5908 5831 5960 5840
rect 5908 5797 5917 5831
rect 5917 5797 5951 5831
rect 5951 5797 5960 5831
rect 5908 5788 5960 5797
rect 4160 5720 4212 5772
rect 2596 5695 2648 5704
rect 1308 5584 1360 5636
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 4252 5652 4304 5704
rect 6092 5652 6144 5704
rect 6644 5652 6696 5704
rect 5724 5584 5776 5636
rect 1952 5516 2004 5568
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 4804 5559 4856 5568
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 2098 5414 2150 5466
rect 2162 5414 2214 5466
rect 2226 5414 2278 5466
rect 2290 5414 2342 5466
rect 5098 5414 5150 5466
rect 5162 5414 5214 5466
rect 5226 5414 5278 5466
rect 5290 5414 5342 5466
rect 4988 5312 5040 5364
rect 6736 5312 6788 5364
rect 1216 5219 1268 5228
rect 1216 5185 1225 5219
rect 1225 5185 1259 5219
rect 1259 5185 1268 5219
rect 1216 5176 1268 5185
rect 1492 5219 1544 5228
rect 1492 5185 1501 5219
rect 1501 5185 1535 5219
rect 1535 5185 1544 5219
rect 1492 5176 1544 5185
rect 2688 5176 2740 5228
rect 4068 5176 4120 5228
rect 4804 5176 4856 5228
rect 1952 5040 2004 5092
rect 3332 4972 3384 5024
rect 4528 5108 4580 5160
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5540 5040 5592 5092
rect 4160 5015 4212 5024
rect 4160 4981 4169 5015
rect 4169 4981 4203 5015
rect 4203 4981 4212 5015
rect 4160 4972 4212 4981
rect 5448 4972 5500 5024
rect 16580 4972 16632 5024
rect 3598 4870 3650 4922
rect 3662 4870 3714 4922
rect 3726 4870 3778 4922
rect 3790 4870 3842 4922
rect 2412 4768 2464 4820
rect 2596 4768 2648 4820
rect 4620 4768 4672 4820
rect 4160 4700 4212 4752
rect 1308 4675 1360 4684
rect 1308 4641 1317 4675
rect 1317 4641 1351 4675
rect 1351 4641 1360 4675
rect 1308 4632 1360 4641
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 16580 4632 16632 4684
rect 1952 4564 2004 4616
rect 2596 4564 2648 4616
rect 4160 4564 4212 4616
rect 5816 4539 5868 4548
rect 5816 4505 5825 4539
rect 5825 4505 5859 4539
rect 5859 4505 5868 4539
rect 5816 4496 5868 4505
rect 4252 4428 4304 4480
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 2098 4326 2150 4378
rect 2162 4326 2214 4378
rect 2226 4326 2278 4378
rect 2290 4326 2342 4378
rect 5098 4326 5150 4378
rect 5162 4326 5214 4378
rect 5226 4326 5278 4378
rect 5290 4326 5342 4378
rect 6000 4224 6052 4276
rect 2596 4156 2648 4208
rect 1216 4131 1268 4140
rect 1216 4097 1225 4131
rect 1225 4097 1259 4131
rect 1259 4097 1268 4131
rect 1216 4088 1268 4097
rect 2688 4088 2740 4140
rect 5632 4156 5684 4208
rect 3424 4088 3476 4140
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4712 4088 4764 4140
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 5448 4088 5500 4140
rect 6092 4063 6144 4072
rect 6092 4029 6101 4063
rect 6101 4029 6135 4063
rect 6135 4029 6144 4063
rect 6092 4020 6144 4029
rect 6552 4156 6604 4208
rect 16672 4224 16724 4276
rect 3598 3782 3650 3834
rect 3662 3782 3714 3834
rect 3726 3782 3778 3834
rect 3790 3782 3842 3834
rect 1676 3612 1728 3664
rect 2320 3680 2372 3732
rect 2320 3587 2372 3596
rect 2320 3553 2329 3587
rect 2329 3553 2363 3587
rect 2363 3553 2372 3587
rect 2320 3544 2372 3553
rect 2688 3476 2740 3528
rect 16580 3680 16632 3732
rect 4160 3544 4212 3596
rect 6460 3655 6512 3664
rect 6460 3621 6469 3655
rect 6469 3621 6503 3655
rect 6503 3621 6512 3655
rect 6460 3612 6512 3621
rect 5816 3544 5868 3596
rect 3056 3340 3108 3392
rect 3332 3340 3384 3392
rect 4068 3340 4120 3392
rect 4528 3340 4580 3392
rect 6092 3340 6144 3392
rect 16672 3340 16724 3392
rect 2098 3238 2150 3290
rect 2162 3238 2214 3290
rect 2226 3238 2278 3290
rect 2290 3238 2342 3290
rect 5098 3238 5150 3290
rect 5162 3238 5214 3290
rect 5226 3238 5278 3290
rect 5290 3238 5342 3290
rect 3884 3136 3936 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 16580 3136 16632 3188
rect 1492 3000 1544 3052
rect 16580 3000 16632 3052
rect 1676 2975 1728 2984
rect 1676 2941 1685 2975
rect 1685 2941 1719 2975
rect 1719 2941 1728 2975
rect 1676 2932 1728 2941
rect 4068 2932 4120 2984
rect 4528 2932 4580 2984
rect 4712 2932 4764 2984
rect 3976 2864 4028 2916
rect 5540 2864 5592 2916
rect 4068 2839 4120 2848
rect 4068 2805 4077 2839
rect 4077 2805 4111 2839
rect 4111 2805 4120 2839
rect 4068 2796 4120 2805
rect 6736 2839 6788 2848
rect 6736 2805 6745 2839
rect 6745 2805 6779 2839
rect 6779 2805 6788 2839
rect 6736 2796 6788 2805
rect 3598 2694 3650 2746
rect 3662 2694 3714 2746
rect 3726 2694 3778 2746
rect 3790 2694 3842 2746
rect 5540 2592 5592 2644
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 1952 2567 2004 2576
rect 1952 2533 1961 2567
rect 1961 2533 1995 2567
rect 1995 2533 2004 2567
rect 1952 2524 2004 2533
rect 4068 2524 4120 2576
rect 6000 2567 6052 2576
rect 6000 2533 6009 2567
rect 6009 2533 6043 2567
rect 6043 2533 6052 2567
rect 6000 2524 6052 2533
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 3792 2456 3844 2508
rect 5632 2499 5684 2508
rect 3424 2388 3476 2440
rect 5632 2465 5641 2499
rect 5641 2465 5675 2499
rect 5675 2465 5684 2499
rect 5632 2456 5684 2465
rect 6736 2456 6788 2508
rect 16580 2456 16632 2508
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 3976 2320 4028 2372
rect 4436 2320 4488 2372
rect 5448 2252 5500 2304
rect 2098 2150 2150 2202
rect 2162 2150 2214 2202
rect 2226 2150 2278 2202
rect 2290 2150 2342 2202
rect 5098 2150 5150 2202
rect 5162 2150 5214 2202
rect 5226 2150 5278 2202
rect 5290 2150 5342 2202
rect 4988 1300 5040 1352
rect 16672 1300 16724 1352
rect 5448 1232 5500 1284
rect 16764 1232 16816 1284
rect 6644 1164 6696 1216
rect 16580 1164 16632 1216
<< metal2 >>
rect 26514 13696 26570 13705
rect 26514 13631 26570 13640
rect 26330 13152 26386 13161
rect 26330 13087 26386 13096
rect 16578 12608 16634 12617
rect 16578 12543 16634 12552
rect 16592 12510 16620 12543
rect 6460 12504 6512 12510
rect 6460 12446 6512 12452
rect 16580 12504 16632 12510
rect 16580 12446 16632 12452
rect 3572 11452 3868 11472
rect 3628 11450 3652 11452
rect 3708 11450 3732 11452
rect 3788 11450 3812 11452
rect 3650 11398 3652 11450
rect 3714 11398 3726 11450
rect 3788 11398 3790 11450
rect 3628 11396 3652 11398
rect 3708 11396 3732 11398
rect 3788 11396 3812 11398
rect 3572 11376 3868 11396
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 2072 10908 2368 10928
rect 2128 10906 2152 10908
rect 2208 10906 2232 10908
rect 2288 10906 2312 10908
rect 2150 10854 2152 10906
rect 2214 10854 2226 10906
rect 2288 10854 2290 10906
rect 2128 10852 2152 10854
rect 2208 10852 2232 10854
rect 2288 10852 2312 10854
rect 2072 10832 2368 10852
rect 3344 10674 3372 11222
rect 4540 11218 4568 11290
rect 4724 11218 4752 11290
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 1216 10600 1268 10606
rect 1216 10542 1268 10548
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 1228 10130 1256 10542
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 1216 10124 1268 10130
rect 1216 10066 1268 10072
rect 1228 9178 1256 10066
rect 2072 9820 2368 9840
rect 2128 9818 2152 9820
rect 2208 9818 2232 9820
rect 2288 9818 2312 9820
rect 2150 9766 2152 9818
rect 2214 9766 2226 9818
rect 2288 9766 2290 9818
rect 2128 9764 2152 9766
rect 2208 9764 2232 9766
rect 2288 9764 2312 9766
rect 2072 9744 2368 9764
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1780 9178 1808 9522
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 1216 9172 1268 9178
rect 1216 9114 1268 9120
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1228 8498 1256 9114
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1596 8634 1624 8978
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1216 8492 1268 8498
rect 1216 8434 1268 8440
rect 1228 7954 1256 8434
rect 1216 7948 1268 7954
rect 1216 7890 1268 7896
rect 1216 7200 1268 7206
rect 1216 7142 1268 7148
rect 1228 6254 1256 7142
rect 1216 6248 1268 6254
rect 1216 6190 1268 6196
rect 1228 5658 1256 6190
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1228 5642 1348 5658
rect 1228 5636 1360 5642
rect 1228 5630 1308 5636
rect 1308 5578 1360 5584
rect 1320 5250 1348 5578
rect 1228 5234 1348 5250
rect 1504 5234 1532 6054
rect 1596 5778 1624 8570
rect 1872 7750 1900 8978
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8022 1992 8774
rect 2072 8732 2368 8752
rect 2128 8730 2152 8732
rect 2208 8730 2232 8732
rect 2288 8730 2312 8732
rect 2150 8678 2152 8730
rect 2214 8678 2226 8730
rect 2288 8678 2290 8730
rect 2128 8676 2152 8678
rect 2208 8676 2232 8678
rect 2288 8676 2312 8678
rect 2072 8656 2368 8676
rect 2424 8294 2452 9386
rect 2608 9110 2636 9386
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 8362 2544 8774
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 6866 1900 7686
rect 2072 7644 2368 7664
rect 2128 7642 2152 7644
rect 2208 7642 2232 7644
rect 2288 7642 2312 7644
rect 2150 7590 2152 7642
rect 2214 7590 2226 7642
rect 2288 7590 2290 7642
rect 2128 7588 2152 7590
rect 2208 7588 2232 7590
rect 2288 7588 2312 7590
rect 2072 7568 2368 7588
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 7002 2360 7210
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1872 5914 1900 6802
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 6186 1992 6598
rect 2072 6556 2368 6576
rect 2128 6554 2152 6556
rect 2208 6554 2232 6556
rect 2288 6554 2312 6556
rect 2150 6502 2152 6554
rect 2214 6502 2226 6554
rect 2288 6502 2290 6554
rect 2128 6500 2152 6502
rect 2208 6500 2232 6502
rect 2288 6500 2312 6502
rect 2072 6480 2368 6500
rect 2700 6458 2728 9454
rect 2884 8974 2912 9658
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2976 8838 3004 9454
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 3068 7954 3096 9318
rect 3160 8430 3188 9590
rect 3344 8634 3372 10134
rect 3436 10130 3464 10474
rect 3572 10364 3868 10384
rect 3628 10362 3652 10364
rect 3708 10362 3732 10364
rect 3788 10362 3812 10364
rect 3650 10310 3652 10362
rect 3714 10310 3726 10362
rect 3788 10310 3790 10362
rect 3628 10308 3652 10310
rect 3708 10308 3732 10310
rect 3788 10308 3812 10310
rect 3572 10288 3868 10308
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3804 9722 3832 10066
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3804 9518 3832 9658
rect 3896 9654 3924 10542
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3572 9276 3868 9296
rect 3628 9274 3652 9276
rect 3708 9274 3732 9276
rect 3788 9274 3812 9276
rect 3650 9222 3652 9274
rect 3714 9222 3726 9274
rect 3788 9222 3790 9274
rect 3628 9220 3652 9222
rect 3708 9220 3732 9222
rect 3788 9220 3812 9222
rect 3572 9200 3868 9220
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3436 8514 3464 9046
rect 3252 8486 3464 8514
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 1952 6180 2004 6186
rect 1952 6122 2004 6128
rect 3160 5930 3188 8366
rect 3252 8362 3280 8486
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 8090 3280 8298
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 8090 3464 8230
rect 3572 8188 3868 8208
rect 3628 8186 3652 8188
rect 3708 8186 3732 8188
rect 3788 8186 3812 8188
rect 3650 8134 3652 8186
rect 3714 8134 3726 8186
rect 3788 8134 3790 8186
rect 3628 8132 3652 8134
rect 3708 8132 3732 8134
rect 3788 8132 3812 8134
rect 3572 8112 3868 8132
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7410 3280 7822
rect 3896 7546 3924 9046
rect 3988 8294 4016 11154
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10198 4200 11018
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4080 9178 4108 9386
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4080 8634 4108 9114
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3252 6934 3280 7346
rect 3988 7342 4016 8230
rect 4080 7886 4108 8366
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3344 6322 3372 7210
rect 3572 7100 3868 7120
rect 3628 7098 3652 7100
rect 3708 7098 3732 7100
rect 3788 7098 3812 7100
rect 3650 7046 3652 7098
rect 3714 7046 3726 7098
rect 3788 7046 3790 7098
rect 3628 7044 3652 7046
rect 3708 7044 3732 7046
rect 3788 7044 3812 7046
rect 3572 7024 3868 7044
rect 4080 6882 4108 7822
rect 4172 7290 4200 9386
rect 4264 8362 4292 9862
rect 4356 9722 4384 10542
rect 4540 10130 4568 11154
rect 4724 11014 4752 11154
rect 6472 11150 6500 12446
rect 16578 11520 16634 11529
rect 16578 11455 16634 11464
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 5072 10908 5368 10928
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5150 10854 5152 10906
rect 5214 10854 5226 10906
rect 5288 10854 5290 10906
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5072 10832 5368 10852
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 7954 4292 8298
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4252 7744 4304 7750
rect 4356 7732 4384 9658
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4304 7704 4384 7732
rect 4252 7686 4304 7692
rect 4172 7262 4292 7290
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 7002 4200 7142
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 3988 6854 4108 6882
rect 3988 6798 4016 6854
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 3068 5902 3188 5930
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 1216 5228 1348 5234
rect 1268 5222 1348 5228
rect 1216 5170 1268 5176
rect 1320 4690 1348 5222
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1320 4570 1348 4626
rect 1228 4542 1348 4570
rect 1228 4146 1256 4542
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 1504 3058 1532 5170
rect 1964 5098 1992 5510
rect 2072 5468 2368 5488
rect 2128 5466 2152 5468
rect 2208 5466 2232 5468
rect 2288 5466 2312 5468
rect 2150 5414 2152 5466
rect 2214 5414 2226 5466
rect 2288 5414 2290 5466
rect 2128 5412 2152 5414
rect 2208 5412 2232 5414
rect 2288 5412 2312 5414
rect 2072 5392 2368 5412
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 2424 4826 2452 5510
rect 2608 4826 2636 5646
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1688 2990 1716 3606
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 2514 1716 2926
rect 1964 2582 1992 4558
rect 2072 4380 2368 4400
rect 2128 4378 2152 4380
rect 2208 4378 2232 4380
rect 2288 4378 2312 4380
rect 2150 4326 2152 4378
rect 2214 4326 2226 4378
rect 2288 4326 2290 4378
rect 2128 4324 2152 4326
rect 2208 4324 2232 4326
rect 2288 4324 2312 4326
rect 2072 4304 2368 4324
rect 2608 4214 2636 4558
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 2700 4146 2728 5170
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2332 3602 2360 3674
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2700 3534 2728 4082
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 3068 3398 3096 5902
rect 3148 5840 3200 5846
rect 3344 5794 3372 6122
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5846 3464 6054
rect 3572 6012 3868 6032
rect 3628 6010 3652 6012
rect 3708 6010 3732 6012
rect 3788 6010 3812 6012
rect 3650 5958 3652 6010
rect 3714 5958 3726 6010
rect 3788 5958 3790 6010
rect 3628 5956 3652 5958
rect 3708 5956 3732 5958
rect 3788 5956 3812 5958
rect 3572 5936 3868 5956
rect 3200 5788 3372 5794
rect 3148 5782 3372 5788
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 4080 5794 4108 6854
rect 3160 5766 3372 5782
rect 3344 5030 3372 5766
rect 4080 5778 4200 5794
rect 4080 5772 4212 5778
rect 4080 5766 4160 5772
rect 4080 5234 4108 5766
rect 4160 5714 4212 5720
rect 4264 5710 4292 7262
rect 4356 6662 4384 7704
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6118 4384 6598
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3344 4078 3372 4966
rect 3572 4924 3868 4944
rect 3628 4922 3652 4924
rect 3708 4922 3732 4924
rect 3788 4922 3812 4924
rect 3650 4870 3652 4922
rect 3714 4870 3726 4922
rect 3788 4870 3790 4922
rect 3628 4868 3652 4870
rect 3708 4868 3732 4870
rect 3788 4868 3812 4870
rect 3572 4848 3868 4868
rect 4172 4758 4200 4966
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3436 4146 3464 4626
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4172 4146 4200 4558
rect 4264 4486 4292 5646
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3572 3836 3868 3856
rect 3628 3834 3652 3836
rect 3708 3834 3732 3836
rect 3788 3834 3812 3836
rect 3650 3782 3652 3834
rect 3714 3782 3726 3834
rect 3788 3782 3790 3834
rect 3628 3780 3652 3782
rect 3708 3780 3732 3782
rect 3788 3780 3812 3782
rect 3572 3760 3868 3780
rect 4172 3602 4200 4082
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 2072 3292 2368 3312
rect 2128 3290 2152 3292
rect 2208 3290 2232 3292
rect 2288 3290 2312 3292
rect 2150 3238 2152 3290
rect 2214 3238 2226 3290
rect 2288 3238 2290 3290
rect 2128 3236 2152 3238
rect 2208 3236 2232 3238
rect 2288 3236 2312 3238
rect 2072 3216 2368 3236
rect 3344 2774 3372 3334
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3344 2746 3464 2774
rect 1952 2576 2004 2582
rect 1952 2518 2004 2524
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 3436 2446 3464 2746
rect 3572 2748 3868 2768
rect 3628 2746 3652 2748
rect 3708 2746 3732 2748
rect 3788 2746 3812 2748
rect 3650 2694 3652 2746
rect 3714 2694 3726 2746
rect 3788 2694 3790 2746
rect 3628 2692 3652 2694
rect 3708 2692 3732 2694
rect 3788 2692 3812 2694
rect 3572 2672 3868 2692
rect 3896 2530 3924 3130
rect 4080 2990 4108 3334
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3804 2514 3924 2530
rect 3792 2508 3924 2514
rect 3844 2502 3924 2508
rect 3792 2450 3844 2456
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3988 2378 4016 2858
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4080 2582 4108 2790
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 4448 2378 4476 8774
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5166 4568 6054
rect 4632 5846 4660 10474
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9382 5028 9998
rect 5072 9820 5368 9840
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5150 9766 5152 9818
rect 5214 9766 5226 9818
rect 5288 9766 5290 9818
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5072 9744 5368 9764
rect 5460 9450 5488 11018
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5828 10010 5856 10066
rect 5736 9982 5856 10010
rect 5736 9926 5764 9982
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 9024 5028 9318
rect 5080 9036 5132 9042
rect 5000 8996 5080 9024
rect 5080 8978 5132 8984
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4540 3398 4568 5102
rect 4632 4826 4660 5782
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4724 4146 4752 7210
rect 4908 6730 4936 8910
rect 5072 8732 5368 8752
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5150 8678 5152 8730
rect 5214 8678 5226 8730
rect 5288 8678 5290 8730
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5072 8656 5368 8676
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5552 8430 5580 8570
rect 5736 8430 5764 9862
rect 6012 9518 6040 10134
rect 6104 9926 6132 10542
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5920 8090 5948 8978
rect 6104 8430 6132 9862
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5632 7880 5684 7886
rect 5920 7834 5948 8026
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5632 7822 5684 7828
rect 5072 7644 5368 7664
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5150 7590 5152 7642
rect 5214 7590 5226 7642
rect 5288 7590 5290 7642
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5072 7568 5368 7588
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 5072 6556 5368 6576
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5150 6502 5152 6554
rect 5214 6502 5226 6554
rect 5288 6502 5290 6554
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5072 6480 5368 6500
rect 5460 5914 5488 7142
rect 5644 6798 5672 7822
rect 5828 7806 5948 7834
rect 5828 7002 5856 7806
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5828 6662 5856 6734
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5736 6322 5764 6598
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5736 5642 5764 6258
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4816 5234 4844 5510
rect 5072 5468 5368 5488
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5150 5414 5152 5466
rect 5214 5414 5226 5466
rect 5288 5414 5290 5466
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5072 5392 5368 5412
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 5000 5166 5028 5306
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5552 5098 5580 5510
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5072 4380 5368 4400
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5150 4326 5152 4378
rect 5214 4326 5226 4378
rect 5288 4326 5290 4378
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5072 4304 5368 4324
rect 5460 4146 5488 4966
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 4214 5672 4422
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4540 2990 4568 3334
rect 4724 2990 4752 4082
rect 5072 3292 5368 3312
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5150 3238 5152 3290
rect 5214 3238 5226 3290
rect 5288 3238 5290 3290
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5072 3216 5368 3236
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5552 2650 5580 2858
rect 5736 2774 5764 5578
rect 5828 4554 5856 6394
rect 5920 5846 5948 7686
rect 6012 7546 6040 7890
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 6104 5710 6132 6734
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6196 5556 6224 8774
rect 6288 8634 6316 9318
rect 6380 9042 6408 9590
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6840 7886 6868 11290
rect 16592 11286 16620 11455
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 26238 10976 26294 10985
rect 26238 10911 26294 10920
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16578 10432 16634 10441
rect 16578 10367 16634 10376
rect 16592 9926 16620 10367
rect 16580 9920 16632 9926
rect 16684 9897 16712 10474
rect 16580 9862 16632 9868
rect 16670 9888 16726 9897
rect 16670 9823 16726 9832
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16592 9353 16620 9386
rect 16578 9344 16634 9353
rect 16578 9279 16634 9288
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16592 8809 16620 8910
rect 16578 8800 16634 8809
rect 16578 8735 16634 8744
rect 26252 8498 26280 10911
rect 26344 9110 26372 13087
rect 26422 12064 26478 12073
rect 26422 11999 26478 12008
rect 26332 9104 26384 9110
rect 26332 9046 26384 9052
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 16580 8288 16632 8294
rect 16578 8256 16580 8265
rect 16632 8256 16634 8265
rect 16578 8191 16634 8200
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6472 6254 6500 7278
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6748 5914 6776 7210
rect 6840 6866 6868 7822
rect 16580 7744 16632 7750
rect 16578 7712 16580 7721
rect 16632 7712 16634 7721
rect 16578 7647 16634 7656
rect 16684 7177 16712 7822
rect 26436 7274 26464 11999
rect 26528 8566 26556 13631
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26424 7268 26476 7274
rect 26424 7210 26476 7216
rect 16670 7168 16726 7177
rect 16670 7103 16726 7112
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6662 6868 6802
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16592 6186 16620 6559
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16684 6089 16712 6666
rect 16670 6080 16726 6089
rect 16670 6015 16726 6024
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6104 5528 6224 5556
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 6012 4282 6040 4626
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5644 2746 5764 2774
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5644 2514 5672 2746
rect 5828 2650 5856 3538
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6012 2582 6040 4218
rect 6104 4078 6132 5528
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6104 3398 6132 4014
rect 6472 3670 6500 4626
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6564 3194 6592 4150
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 2072 2204 2368 2224
rect 2128 2202 2152 2204
rect 2208 2202 2232 2204
rect 2288 2202 2312 2204
rect 2150 2150 2152 2202
rect 2214 2150 2226 2202
rect 2288 2150 2290 2202
rect 2128 2148 2152 2150
rect 2208 2148 2232 2150
rect 2288 2148 2312 2150
rect 2072 2128 2368 2148
rect 5000 1358 5028 2382
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5072 2204 5368 2224
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5150 2150 5152 2202
rect 5214 2150 5226 2202
rect 5288 2150 5290 2202
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5072 2128 5368 2148
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5460 1290 5488 2246
rect 5448 1284 5500 1290
rect 5448 1226 5500 1232
rect 6656 1222 6684 5646
rect 6748 5370 6776 5850
rect 16578 5536 16634 5545
rect 16578 5471 16634 5480
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 16592 5030 16620 5471
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16670 4992 16726 5001
rect 16670 4927 16726 4936
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16592 4457 16620 4626
rect 16578 4448 16634 4457
rect 16578 4383 16634 4392
rect 16684 4282 16712 4927
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16578 3904 16634 3913
rect 16578 3839 16634 3848
rect 16592 3738 16620 3839
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16672 3392 16724 3398
rect 16578 3360 16634 3369
rect 16672 3334 16724 3340
rect 16578 3295 16634 3304
rect 16592 3194 16620 3295
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 6736 2848 6788 2854
rect 16592 2825 16620 2994
rect 6736 2790 6788 2796
rect 16578 2816 16634 2825
rect 6748 2514 6776 2790
rect 16578 2751 16634 2760
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16592 2281 16620 2450
rect 16578 2272 16634 2281
rect 16578 2207 16634 2216
rect 16684 1737 16712 3334
rect 16670 1728 16726 1737
rect 16670 1663 16726 1672
rect 16672 1352 16724 1358
rect 16672 1294 16724 1300
rect 6644 1216 6696 1222
rect 16580 1216 16632 1222
rect 6644 1158 6696 1164
rect 16578 1184 16580 1193
rect 16632 1184 16634 1193
rect 16578 1119 16634 1128
rect 16684 649 16712 1294
rect 16764 1284 16816 1290
rect 16764 1226 16816 1232
rect 16670 640 16726 649
rect 16670 575 16726 584
rect 16776 241 16804 1226
rect 16762 232 16818 241
rect 16762 167 16818 176
<< via2 >>
rect 26514 13640 26570 13696
rect 26330 13096 26386 13152
rect 16578 12552 16634 12608
rect 3572 11450 3628 11452
rect 3652 11450 3708 11452
rect 3732 11450 3788 11452
rect 3812 11450 3868 11452
rect 3572 11398 3598 11450
rect 3598 11398 3628 11450
rect 3652 11398 3662 11450
rect 3662 11398 3708 11450
rect 3732 11398 3778 11450
rect 3778 11398 3788 11450
rect 3812 11398 3842 11450
rect 3842 11398 3868 11450
rect 3572 11396 3628 11398
rect 3652 11396 3708 11398
rect 3732 11396 3788 11398
rect 3812 11396 3868 11398
rect 2072 10906 2128 10908
rect 2152 10906 2208 10908
rect 2232 10906 2288 10908
rect 2312 10906 2368 10908
rect 2072 10854 2098 10906
rect 2098 10854 2128 10906
rect 2152 10854 2162 10906
rect 2162 10854 2208 10906
rect 2232 10854 2278 10906
rect 2278 10854 2288 10906
rect 2312 10854 2342 10906
rect 2342 10854 2368 10906
rect 2072 10852 2128 10854
rect 2152 10852 2208 10854
rect 2232 10852 2288 10854
rect 2312 10852 2368 10854
rect 2072 9818 2128 9820
rect 2152 9818 2208 9820
rect 2232 9818 2288 9820
rect 2312 9818 2368 9820
rect 2072 9766 2098 9818
rect 2098 9766 2128 9818
rect 2152 9766 2162 9818
rect 2162 9766 2208 9818
rect 2232 9766 2278 9818
rect 2278 9766 2288 9818
rect 2312 9766 2342 9818
rect 2342 9766 2368 9818
rect 2072 9764 2128 9766
rect 2152 9764 2208 9766
rect 2232 9764 2288 9766
rect 2312 9764 2368 9766
rect 2072 8730 2128 8732
rect 2152 8730 2208 8732
rect 2232 8730 2288 8732
rect 2312 8730 2368 8732
rect 2072 8678 2098 8730
rect 2098 8678 2128 8730
rect 2152 8678 2162 8730
rect 2162 8678 2208 8730
rect 2232 8678 2278 8730
rect 2278 8678 2288 8730
rect 2312 8678 2342 8730
rect 2342 8678 2368 8730
rect 2072 8676 2128 8678
rect 2152 8676 2208 8678
rect 2232 8676 2288 8678
rect 2312 8676 2368 8678
rect 2072 7642 2128 7644
rect 2152 7642 2208 7644
rect 2232 7642 2288 7644
rect 2312 7642 2368 7644
rect 2072 7590 2098 7642
rect 2098 7590 2128 7642
rect 2152 7590 2162 7642
rect 2162 7590 2208 7642
rect 2232 7590 2278 7642
rect 2278 7590 2288 7642
rect 2312 7590 2342 7642
rect 2342 7590 2368 7642
rect 2072 7588 2128 7590
rect 2152 7588 2208 7590
rect 2232 7588 2288 7590
rect 2312 7588 2368 7590
rect 2072 6554 2128 6556
rect 2152 6554 2208 6556
rect 2232 6554 2288 6556
rect 2312 6554 2368 6556
rect 2072 6502 2098 6554
rect 2098 6502 2128 6554
rect 2152 6502 2162 6554
rect 2162 6502 2208 6554
rect 2232 6502 2278 6554
rect 2278 6502 2288 6554
rect 2312 6502 2342 6554
rect 2342 6502 2368 6554
rect 2072 6500 2128 6502
rect 2152 6500 2208 6502
rect 2232 6500 2288 6502
rect 2312 6500 2368 6502
rect 3572 10362 3628 10364
rect 3652 10362 3708 10364
rect 3732 10362 3788 10364
rect 3812 10362 3868 10364
rect 3572 10310 3598 10362
rect 3598 10310 3628 10362
rect 3652 10310 3662 10362
rect 3662 10310 3708 10362
rect 3732 10310 3778 10362
rect 3778 10310 3788 10362
rect 3812 10310 3842 10362
rect 3842 10310 3868 10362
rect 3572 10308 3628 10310
rect 3652 10308 3708 10310
rect 3732 10308 3788 10310
rect 3812 10308 3868 10310
rect 3572 9274 3628 9276
rect 3652 9274 3708 9276
rect 3732 9274 3788 9276
rect 3812 9274 3868 9276
rect 3572 9222 3598 9274
rect 3598 9222 3628 9274
rect 3652 9222 3662 9274
rect 3662 9222 3708 9274
rect 3732 9222 3778 9274
rect 3778 9222 3788 9274
rect 3812 9222 3842 9274
rect 3842 9222 3868 9274
rect 3572 9220 3628 9222
rect 3652 9220 3708 9222
rect 3732 9220 3788 9222
rect 3812 9220 3868 9222
rect 3572 8186 3628 8188
rect 3652 8186 3708 8188
rect 3732 8186 3788 8188
rect 3812 8186 3868 8188
rect 3572 8134 3598 8186
rect 3598 8134 3628 8186
rect 3652 8134 3662 8186
rect 3662 8134 3708 8186
rect 3732 8134 3778 8186
rect 3778 8134 3788 8186
rect 3812 8134 3842 8186
rect 3842 8134 3868 8186
rect 3572 8132 3628 8134
rect 3652 8132 3708 8134
rect 3732 8132 3788 8134
rect 3812 8132 3868 8134
rect 3572 7098 3628 7100
rect 3652 7098 3708 7100
rect 3732 7098 3788 7100
rect 3812 7098 3868 7100
rect 3572 7046 3598 7098
rect 3598 7046 3628 7098
rect 3652 7046 3662 7098
rect 3662 7046 3708 7098
rect 3732 7046 3778 7098
rect 3778 7046 3788 7098
rect 3812 7046 3842 7098
rect 3842 7046 3868 7098
rect 3572 7044 3628 7046
rect 3652 7044 3708 7046
rect 3732 7044 3788 7046
rect 3812 7044 3868 7046
rect 16578 11464 16634 11520
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5098 10906
rect 5098 10854 5128 10906
rect 5152 10854 5162 10906
rect 5162 10854 5208 10906
rect 5232 10854 5278 10906
rect 5278 10854 5288 10906
rect 5312 10854 5342 10906
rect 5342 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 2072 5466 2128 5468
rect 2152 5466 2208 5468
rect 2232 5466 2288 5468
rect 2312 5466 2368 5468
rect 2072 5414 2098 5466
rect 2098 5414 2128 5466
rect 2152 5414 2162 5466
rect 2162 5414 2208 5466
rect 2232 5414 2278 5466
rect 2278 5414 2288 5466
rect 2312 5414 2342 5466
rect 2342 5414 2368 5466
rect 2072 5412 2128 5414
rect 2152 5412 2208 5414
rect 2232 5412 2288 5414
rect 2312 5412 2368 5414
rect 2072 4378 2128 4380
rect 2152 4378 2208 4380
rect 2232 4378 2288 4380
rect 2312 4378 2368 4380
rect 2072 4326 2098 4378
rect 2098 4326 2128 4378
rect 2152 4326 2162 4378
rect 2162 4326 2208 4378
rect 2232 4326 2278 4378
rect 2278 4326 2288 4378
rect 2312 4326 2342 4378
rect 2342 4326 2368 4378
rect 2072 4324 2128 4326
rect 2152 4324 2208 4326
rect 2232 4324 2288 4326
rect 2312 4324 2368 4326
rect 3572 6010 3628 6012
rect 3652 6010 3708 6012
rect 3732 6010 3788 6012
rect 3812 6010 3868 6012
rect 3572 5958 3598 6010
rect 3598 5958 3628 6010
rect 3652 5958 3662 6010
rect 3662 5958 3708 6010
rect 3732 5958 3778 6010
rect 3778 5958 3788 6010
rect 3812 5958 3842 6010
rect 3842 5958 3868 6010
rect 3572 5956 3628 5958
rect 3652 5956 3708 5958
rect 3732 5956 3788 5958
rect 3812 5956 3868 5958
rect 3572 4922 3628 4924
rect 3652 4922 3708 4924
rect 3732 4922 3788 4924
rect 3812 4922 3868 4924
rect 3572 4870 3598 4922
rect 3598 4870 3628 4922
rect 3652 4870 3662 4922
rect 3662 4870 3708 4922
rect 3732 4870 3778 4922
rect 3778 4870 3788 4922
rect 3812 4870 3842 4922
rect 3842 4870 3868 4922
rect 3572 4868 3628 4870
rect 3652 4868 3708 4870
rect 3732 4868 3788 4870
rect 3812 4868 3868 4870
rect 3572 3834 3628 3836
rect 3652 3834 3708 3836
rect 3732 3834 3788 3836
rect 3812 3834 3868 3836
rect 3572 3782 3598 3834
rect 3598 3782 3628 3834
rect 3652 3782 3662 3834
rect 3662 3782 3708 3834
rect 3732 3782 3778 3834
rect 3778 3782 3788 3834
rect 3812 3782 3842 3834
rect 3842 3782 3868 3834
rect 3572 3780 3628 3782
rect 3652 3780 3708 3782
rect 3732 3780 3788 3782
rect 3812 3780 3868 3782
rect 2072 3290 2128 3292
rect 2152 3290 2208 3292
rect 2232 3290 2288 3292
rect 2312 3290 2368 3292
rect 2072 3238 2098 3290
rect 2098 3238 2128 3290
rect 2152 3238 2162 3290
rect 2162 3238 2208 3290
rect 2232 3238 2278 3290
rect 2278 3238 2288 3290
rect 2312 3238 2342 3290
rect 2342 3238 2368 3290
rect 2072 3236 2128 3238
rect 2152 3236 2208 3238
rect 2232 3236 2288 3238
rect 2312 3236 2368 3238
rect 3572 2746 3628 2748
rect 3652 2746 3708 2748
rect 3732 2746 3788 2748
rect 3812 2746 3868 2748
rect 3572 2694 3598 2746
rect 3598 2694 3628 2746
rect 3652 2694 3662 2746
rect 3662 2694 3708 2746
rect 3732 2694 3778 2746
rect 3778 2694 3788 2746
rect 3812 2694 3842 2746
rect 3842 2694 3868 2746
rect 3572 2692 3628 2694
rect 3652 2692 3708 2694
rect 3732 2692 3788 2694
rect 3812 2692 3868 2694
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5098 9818
rect 5098 9766 5128 9818
rect 5152 9766 5162 9818
rect 5162 9766 5208 9818
rect 5232 9766 5278 9818
rect 5278 9766 5288 9818
rect 5312 9766 5342 9818
rect 5342 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5098 8730
rect 5098 8678 5128 8730
rect 5152 8678 5162 8730
rect 5162 8678 5208 8730
rect 5232 8678 5278 8730
rect 5278 8678 5288 8730
rect 5312 8678 5342 8730
rect 5342 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5098 7642
rect 5098 7590 5128 7642
rect 5152 7590 5162 7642
rect 5162 7590 5208 7642
rect 5232 7590 5278 7642
rect 5278 7590 5288 7642
rect 5312 7590 5342 7642
rect 5342 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5098 6554
rect 5098 6502 5128 6554
rect 5152 6502 5162 6554
rect 5162 6502 5208 6554
rect 5232 6502 5278 6554
rect 5278 6502 5288 6554
rect 5312 6502 5342 6554
rect 5342 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5098 5466
rect 5098 5414 5128 5466
rect 5152 5414 5162 5466
rect 5162 5414 5208 5466
rect 5232 5414 5278 5466
rect 5278 5414 5288 5466
rect 5312 5414 5342 5466
rect 5342 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5098 4378
rect 5098 4326 5128 4378
rect 5152 4326 5162 4378
rect 5162 4326 5208 4378
rect 5232 4326 5278 4378
rect 5278 4326 5288 4378
rect 5312 4326 5342 4378
rect 5342 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5098 3290
rect 5098 3238 5128 3290
rect 5152 3238 5162 3290
rect 5162 3238 5208 3290
rect 5232 3238 5278 3290
rect 5278 3238 5288 3290
rect 5312 3238 5342 3290
rect 5342 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 26238 10920 26294 10976
rect 16578 10376 16634 10432
rect 16670 9832 16726 9888
rect 16578 9288 16634 9344
rect 16578 8744 16634 8800
rect 26422 12008 26478 12064
rect 16578 8236 16580 8256
rect 16580 8236 16632 8256
rect 16632 8236 16634 8256
rect 16578 8200 16634 8236
rect 16578 7692 16580 7712
rect 16580 7692 16632 7712
rect 16632 7692 16634 7712
rect 16578 7656 16634 7692
rect 16670 7112 16726 7168
rect 16578 6568 16634 6624
rect 16670 6024 16726 6080
rect 2072 2202 2128 2204
rect 2152 2202 2208 2204
rect 2232 2202 2288 2204
rect 2312 2202 2368 2204
rect 2072 2150 2098 2202
rect 2098 2150 2128 2202
rect 2152 2150 2162 2202
rect 2162 2150 2208 2202
rect 2232 2150 2278 2202
rect 2278 2150 2288 2202
rect 2312 2150 2342 2202
rect 2342 2150 2368 2202
rect 2072 2148 2128 2150
rect 2152 2148 2208 2150
rect 2232 2148 2288 2150
rect 2312 2148 2368 2150
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5098 2202
rect 5098 2150 5128 2202
rect 5152 2150 5162 2202
rect 5162 2150 5208 2202
rect 5232 2150 5278 2202
rect 5278 2150 5288 2202
rect 5312 2150 5342 2202
rect 5342 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 16578 5480 16634 5536
rect 16670 4936 16726 4992
rect 16578 4392 16634 4448
rect 16578 3848 16634 3904
rect 16578 3304 16634 3360
rect 16578 2760 16634 2816
rect 16578 2216 16634 2272
rect 16670 1672 16726 1728
rect 16578 1164 16580 1184
rect 16580 1164 16632 1184
rect 16632 1164 16634 1184
rect 16578 1128 16634 1164
rect 16670 584 16726 640
rect 16762 176 16818 232
<< metal3 >>
rect 14000 13696 34000 13728
rect 14000 13640 26514 13696
rect 26570 13640 34000 13696
rect 14000 13608 34000 13640
rect 14000 13152 34000 13184
rect 14000 13096 26330 13152
rect 26386 13096 34000 13152
rect 14000 13064 34000 13096
rect 14000 12608 34000 12640
rect 14000 12552 16578 12608
rect 16634 12552 34000 12608
rect 14000 12520 34000 12552
rect 14000 12064 34000 12096
rect 14000 12008 26422 12064
rect 26478 12008 34000 12064
rect 14000 11976 34000 12008
rect 14000 11520 34000 11552
rect 14000 11464 16578 11520
rect 16634 11464 34000 11520
rect 3560 11456 3880 11457
rect 3560 11392 3568 11456
rect 3632 11392 3648 11456
rect 3712 11392 3728 11456
rect 3792 11392 3808 11456
rect 3872 11392 3880 11456
rect 14000 11432 34000 11464
rect 3560 11391 3880 11392
rect 14000 10976 34000 11008
rect 14000 10920 26238 10976
rect 26294 10920 34000 10976
rect 2060 10912 2380 10913
rect 2060 10848 2068 10912
rect 2132 10848 2148 10912
rect 2212 10848 2228 10912
rect 2292 10848 2308 10912
rect 2372 10848 2380 10912
rect 2060 10847 2380 10848
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 14000 10888 34000 10920
rect 5060 10847 5380 10848
rect 14000 10432 34000 10464
rect 14000 10376 16578 10432
rect 16634 10376 34000 10432
rect 3560 10368 3880 10369
rect 3560 10304 3568 10368
rect 3632 10304 3648 10368
rect 3712 10304 3728 10368
rect 3792 10304 3808 10368
rect 3872 10304 3880 10368
rect 14000 10344 34000 10376
rect 3560 10303 3880 10304
rect 14000 9888 34000 9920
rect 14000 9832 16670 9888
rect 16726 9832 34000 9888
rect 2060 9824 2380 9825
rect 2060 9760 2068 9824
rect 2132 9760 2148 9824
rect 2212 9760 2228 9824
rect 2292 9760 2308 9824
rect 2372 9760 2380 9824
rect 2060 9759 2380 9760
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9832
rect 5060 9759 5380 9760
rect 14000 9344 34000 9376
rect 14000 9288 16578 9344
rect 16634 9288 34000 9344
rect 3560 9280 3880 9281
rect 3560 9216 3568 9280
rect 3632 9216 3648 9280
rect 3712 9216 3728 9280
rect 3792 9216 3808 9280
rect 3872 9216 3880 9280
rect 14000 9256 34000 9288
rect 3560 9215 3880 9216
rect 14000 8800 34000 8832
rect 14000 8744 16578 8800
rect 16634 8744 34000 8800
rect 2060 8736 2380 8737
rect 2060 8672 2068 8736
rect 2132 8672 2148 8736
rect 2212 8672 2228 8736
rect 2292 8672 2308 8736
rect 2372 8672 2380 8736
rect 2060 8671 2380 8672
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 14000 8712 34000 8744
rect 5060 8671 5380 8672
rect 14000 8256 34000 8288
rect 14000 8200 16578 8256
rect 16634 8200 34000 8256
rect 3560 8192 3880 8193
rect 3560 8128 3568 8192
rect 3632 8128 3648 8192
rect 3712 8128 3728 8192
rect 3792 8128 3808 8192
rect 3872 8128 3880 8192
rect 14000 8168 34000 8200
rect 3560 8127 3880 8128
rect 14000 7712 34000 7744
rect 14000 7656 16578 7712
rect 16634 7656 34000 7712
rect 2060 7648 2380 7649
rect 2060 7584 2068 7648
rect 2132 7584 2148 7648
rect 2212 7584 2228 7648
rect 2292 7584 2308 7648
rect 2372 7584 2380 7648
rect 2060 7583 2380 7584
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 14000 7624 34000 7656
rect 5060 7583 5380 7584
rect 14000 7168 34000 7200
rect 14000 7112 16670 7168
rect 16726 7112 34000 7168
rect 3560 7104 3880 7105
rect 3560 7040 3568 7104
rect 3632 7040 3648 7104
rect 3712 7040 3728 7104
rect 3792 7040 3808 7104
rect 3872 7040 3880 7104
rect 14000 7080 34000 7112
rect 3560 7039 3880 7040
rect 14000 6624 34000 6656
rect 14000 6568 16578 6624
rect 16634 6568 34000 6624
rect 2060 6560 2380 6561
rect 2060 6496 2068 6560
rect 2132 6496 2148 6560
rect 2212 6496 2228 6560
rect 2292 6496 2308 6560
rect 2372 6496 2380 6560
rect 2060 6495 2380 6496
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6568
rect 5060 6495 5380 6496
rect 14000 6080 34000 6112
rect 14000 6024 16670 6080
rect 16726 6024 34000 6080
rect 3560 6016 3880 6017
rect 3560 5952 3568 6016
rect 3632 5952 3648 6016
rect 3712 5952 3728 6016
rect 3792 5952 3808 6016
rect 3872 5952 3880 6016
rect 14000 5992 34000 6024
rect 3560 5951 3880 5952
rect 14000 5536 34000 5568
rect 14000 5480 16578 5536
rect 16634 5480 34000 5536
rect 2060 5472 2380 5473
rect 2060 5408 2068 5472
rect 2132 5408 2148 5472
rect 2212 5408 2228 5472
rect 2292 5408 2308 5472
rect 2372 5408 2380 5472
rect 2060 5407 2380 5408
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 14000 5448 34000 5480
rect 5060 5407 5380 5408
rect 14000 4992 34000 5024
rect 14000 4936 16670 4992
rect 16726 4936 34000 4992
rect 3560 4928 3880 4929
rect 3560 4864 3568 4928
rect 3632 4864 3648 4928
rect 3712 4864 3728 4928
rect 3792 4864 3808 4928
rect 3872 4864 3880 4928
rect 14000 4904 34000 4936
rect 3560 4863 3880 4864
rect 14000 4448 34000 4480
rect 14000 4392 16578 4448
rect 16634 4392 34000 4448
rect 2060 4384 2380 4385
rect 2060 4320 2068 4384
rect 2132 4320 2148 4384
rect 2212 4320 2228 4384
rect 2292 4320 2308 4384
rect 2372 4320 2380 4384
rect 2060 4319 2380 4320
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 14000 4360 34000 4392
rect 5060 4319 5380 4320
rect 14000 3904 34000 3936
rect 14000 3848 16578 3904
rect 16634 3848 34000 3904
rect 3560 3840 3880 3841
rect 3560 3776 3568 3840
rect 3632 3776 3648 3840
rect 3712 3776 3728 3840
rect 3792 3776 3808 3840
rect 3872 3776 3880 3840
rect 14000 3816 34000 3848
rect 3560 3775 3880 3776
rect 14000 3360 34000 3392
rect 14000 3304 16578 3360
rect 16634 3304 34000 3360
rect 2060 3296 2380 3297
rect 2060 3232 2068 3296
rect 2132 3232 2148 3296
rect 2212 3232 2228 3296
rect 2292 3232 2308 3296
rect 2372 3232 2380 3296
rect 2060 3231 2380 3232
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 14000 3272 34000 3304
rect 5060 3231 5380 3232
rect 14000 2816 34000 2848
rect 14000 2760 16578 2816
rect 16634 2760 34000 2816
rect 3560 2752 3880 2753
rect 3560 2688 3568 2752
rect 3632 2688 3648 2752
rect 3712 2688 3728 2752
rect 3792 2688 3808 2752
rect 3872 2688 3880 2752
rect 14000 2728 34000 2760
rect 3560 2687 3880 2688
rect 14000 2272 34000 2304
rect 14000 2216 16578 2272
rect 16634 2216 34000 2272
rect 2060 2208 2380 2209
rect 2060 2144 2068 2208
rect 2132 2144 2148 2208
rect 2212 2144 2228 2208
rect 2292 2144 2308 2208
rect 2372 2144 2380 2208
rect 2060 2143 2380 2144
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 14000 2184 34000 2216
rect 5060 2143 5380 2144
rect 14000 1728 34000 1760
rect 14000 1672 16670 1728
rect 16726 1672 34000 1728
rect 14000 1640 34000 1672
rect 14000 1184 34000 1216
rect 14000 1128 16578 1184
rect 16634 1128 34000 1184
rect 14000 1096 34000 1128
rect 14000 640 34000 672
rect 14000 584 16670 640
rect 16726 584 34000 640
rect 14000 552 34000 584
rect 14000 232 34000 264
rect 14000 176 16762 232
rect 16818 176 34000 232
rect 14000 144 34000 176
<< via3 >>
rect 3568 11452 3632 11456
rect 3568 11396 3572 11452
rect 3572 11396 3628 11452
rect 3628 11396 3632 11452
rect 3568 11392 3632 11396
rect 3648 11452 3712 11456
rect 3648 11396 3652 11452
rect 3652 11396 3708 11452
rect 3708 11396 3712 11452
rect 3648 11392 3712 11396
rect 3728 11452 3792 11456
rect 3728 11396 3732 11452
rect 3732 11396 3788 11452
rect 3788 11396 3792 11452
rect 3728 11392 3792 11396
rect 3808 11452 3872 11456
rect 3808 11396 3812 11452
rect 3812 11396 3868 11452
rect 3868 11396 3872 11452
rect 3808 11392 3872 11396
rect 2068 10908 2132 10912
rect 2068 10852 2072 10908
rect 2072 10852 2128 10908
rect 2128 10852 2132 10908
rect 2068 10848 2132 10852
rect 2148 10908 2212 10912
rect 2148 10852 2152 10908
rect 2152 10852 2208 10908
rect 2208 10852 2212 10908
rect 2148 10848 2212 10852
rect 2228 10908 2292 10912
rect 2228 10852 2232 10908
rect 2232 10852 2288 10908
rect 2288 10852 2292 10908
rect 2228 10848 2292 10852
rect 2308 10908 2372 10912
rect 2308 10852 2312 10908
rect 2312 10852 2368 10908
rect 2368 10852 2372 10908
rect 2308 10848 2372 10852
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 3568 10364 3632 10368
rect 3568 10308 3572 10364
rect 3572 10308 3628 10364
rect 3628 10308 3632 10364
rect 3568 10304 3632 10308
rect 3648 10364 3712 10368
rect 3648 10308 3652 10364
rect 3652 10308 3708 10364
rect 3708 10308 3712 10364
rect 3648 10304 3712 10308
rect 3728 10364 3792 10368
rect 3728 10308 3732 10364
rect 3732 10308 3788 10364
rect 3788 10308 3792 10364
rect 3728 10304 3792 10308
rect 3808 10364 3872 10368
rect 3808 10308 3812 10364
rect 3812 10308 3868 10364
rect 3868 10308 3872 10364
rect 3808 10304 3872 10308
rect 2068 9820 2132 9824
rect 2068 9764 2072 9820
rect 2072 9764 2128 9820
rect 2128 9764 2132 9820
rect 2068 9760 2132 9764
rect 2148 9820 2212 9824
rect 2148 9764 2152 9820
rect 2152 9764 2208 9820
rect 2208 9764 2212 9820
rect 2148 9760 2212 9764
rect 2228 9820 2292 9824
rect 2228 9764 2232 9820
rect 2232 9764 2288 9820
rect 2288 9764 2292 9820
rect 2228 9760 2292 9764
rect 2308 9820 2372 9824
rect 2308 9764 2312 9820
rect 2312 9764 2368 9820
rect 2368 9764 2372 9820
rect 2308 9760 2372 9764
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 3568 9276 3632 9280
rect 3568 9220 3572 9276
rect 3572 9220 3628 9276
rect 3628 9220 3632 9276
rect 3568 9216 3632 9220
rect 3648 9276 3712 9280
rect 3648 9220 3652 9276
rect 3652 9220 3708 9276
rect 3708 9220 3712 9276
rect 3648 9216 3712 9220
rect 3728 9276 3792 9280
rect 3728 9220 3732 9276
rect 3732 9220 3788 9276
rect 3788 9220 3792 9276
rect 3728 9216 3792 9220
rect 3808 9276 3872 9280
rect 3808 9220 3812 9276
rect 3812 9220 3868 9276
rect 3868 9220 3872 9276
rect 3808 9216 3872 9220
rect 2068 8732 2132 8736
rect 2068 8676 2072 8732
rect 2072 8676 2128 8732
rect 2128 8676 2132 8732
rect 2068 8672 2132 8676
rect 2148 8732 2212 8736
rect 2148 8676 2152 8732
rect 2152 8676 2208 8732
rect 2208 8676 2212 8732
rect 2148 8672 2212 8676
rect 2228 8732 2292 8736
rect 2228 8676 2232 8732
rect 2232 8676 2288 8732
rect 2288 8676 2292 8732
rect 2228 8672 2292 8676
rect 2308 8732 2372 8736
rect 2308 8676 2312 8732
rect 2312 8676 2368 8732
rect 2368 8676 2372 8732
rect 2308 8672 2372 8676
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 3568 8188 3632 8192
rect 3568 8132 3572 8188
rect 3572 8132 3628 8188
rect 3628 8132 3632 8188
rect 3568 8128 3632 8132
rect 3648 8188 3712 8192
rect 3648 8132 3652 8188
rect 3652 8132 3708 8188
rect 3708 8132 3712 8188
rect 3648 8128 3712 8132
rect 3728 8188 3792 8192
rect 3728 8132 3732 8188
rect 3732 8132 3788 8188
rect 3788 8132 3792 8188
rect 3728 8128 3792 8132
rect 3808 8188 3872 8192
rect 3808 8132 3812 8188
rect 3812 8132 3868 8188
rect 3868 8132 3872 8188
rect 3808 8128 3872 8132
rect 2068 7644 2132 7648
rect 2068 7588 2072 7644
rect 2072 7588 2128 7644
rect 2128 7588 2132 7644
rect 2068 7584 2132 7588
rect 2148 7644 2212 7648
rect 2148 7588 2152 7644
rect 2152 7588 2208 7644
rect 2208 7588 2212 7644
rect 2148 7584 2212 7588
rect 2228 7644 2292 7648
rect 2228 7588 2232 7644
rect 2232 7588 2288 7644
rect 2288 7588 2292 7644
rect 2228 7584 2292 7588
rect 2308 7644 2372 7648
rect 2308 7588 2312 7644
rect 2312 7588 2368 7644
rect 2368 7588 2372 7644
rect 2308 7584 2372 7588
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 3568 7100 3632 7104
rect 3568 7044 3572 7100
rect 3572 7044 3628 7100
rect 3628 7044 3632 7100
rect 3568 7040 3632 7044
rect 3648 7100 3712 7104
rect 3648 7044 3652 7100
rect 3652 7044 3708 7100
rect 3708 7044 3712 7100
rect 3648 7040 3712 7044
rect 3728 7100 3792 7104
rect 3728 7044 3732 7100
rect 3732 7044 3788 7100
rect 3788 7044 3792 7100
rect 3728 7040 3792 7044
rect 3808 7100 3872 7104
rect 3808 7044 3812 7100
rect 3812 7044 3868 7100
rect 3868 7044 3872 7100
rect 3808 7040 3872 7044
rect 2068 6556 2132 6560
rect 2068 6500 2072 6556
rect 2072 6500 2128 6556
rect 2128 6500 2132 6556
rect 2068 6496 2132 6500
rect 2148 6556 2212 6560
rect 2148 6500 2152 6556
rect 2152 6500 2208 6556
rect 2208 6500 2212 6556
rect 2148 6496 2212 6500
rect 2228 6556 2292 6560
rect 2228 6500 2232 6556
rect 2232 6500 2288 6556
rect 2288 6500 2292 6556
rect 2228 6496 2292 6500
rect 2308 6556 2372 6560
rect 2308 6500 2312 6556
rect 2312 6500 2368 6556
rect 2368 6500 2372 6556
rect 2308 6496 2372 6500
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 3568 6012 3632 6016
rect 3568 5956 3572 6012
rect 3572 5956 3628 6012
rect 3628 5956 3632 6012
rect 3568 5952 3632 5956
rect 3648 6012 3712 6016
rect 3648 5956 3652 6012
rect 3652 5956 3708 6012
rect 3708 5956 3712 6012
rect 3648 5952 3712 5956
rect 3728 6012 3792 6016
rect 3728 5956 3732 6012
rect 3732 5956 3788 6012
rect 3788 5956 3792 6012
rect 3728 5952 3792 5956
rect 3808 6012 3872 6016
rect 3808 5956 3812 6012
rect 3812 5956 3868 6012
rect 3868 5956 3872 6012
rect 3808 5952 3872 5956
rect 2068 5468 2132 5472
rect 2068 5412 2072 5468
rect 2072 5412 2128 5468
rect 2128 5412 2132 5468
rect 2068 5408 2132 5412
rect 2148 5468 2212 5472
rect 2148 5412 2152 5468
rect 2152 5412 2208 5468
rect 2208 5412 2212 5468
rect 2148 5408 2212 5412
rect 2228 5468 2292 5472
rect 2228 5412 2232 5468
rect 2232 5412 2288 5468
rect 2288 5412 2292 5468
rect 2228 5408 2292 5412
rect 2308 5468 2372 5472
rect 2308 5412 2312 5468
rect 2312 5412 2368 5468
rect 2368 5412 2372 5468
rect 2308 5408 2372 5412
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 3568 4924 3632 4928
rect 3568 4868 3572 4924
rect 3572 4868 3628 4924
rect 3628 4868 3632 4924
rect 3568 4864 3632 4868
rect 3648 4924 3712 4928
rect 3648 4868 3652 4924
rect 3652 4868 3708 4924
rect 3708 4868 3712 4924
rect 3648 4864 3712 4868
rect 3728 4924 3792 4928
rect 3728 4868 3732 4924
rect 3732 4868 3788 4924
rect 3788 4868 3792 4924
rect 3728 4864 3792 4868
rect 3808 4924 3872 4928
rect 3808 4868 3812 4924
rect 3812 4868 3868 4924
rect 3868 4868 3872 4924
rect 3808 4864 3872 4868
rect 2068 4380 2132 4384
rect 2068 4324 2072 4380
rect 2072 4324 2128 4380
rect 2128 4324 2132 4380
rect 2068 4320 2132 4324
rect 2148 4380 2212 4384
rect 2148 4324 2152 4380
rect 2152 4324 2208 4380
rect 2208 4324 2212 4380
rect 2148 4320 2212 4324
rect 2228 4380 2292 4384
rect 2228 4324 2232 4380
rect 2232 4324 2288 4380
rect 2288 4324 2292 4380
rect 2228 4320 2292 4324
rect 2308 4380 2372 4384
rect 2308 4324 2312 4380
rect 2312 4324 2368 4380
rect 2368 4324 2372 4380
rect 2308 4320 2372 4324
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 3568 3836 3632 3840
rect 3568 3780 3572 3836
rect 3572 3780 3628 3836
rect 3628 3780 3632 3836
rect 3568 3776 3632 3780
rect 3648 3836 3712 3840
rect 3648 3780 3652 3836
rect 3652 3780 3708 3836
rect 3708 3780 3712 3836
rect 3648 3776 3712 3780
rect 3728 3836 3792 3840
rect 3728 3780 3732 3836
rect 3732 3780 3788 3836
rect 3788 3780 3792 3836
rect 3728 3776 3792 3780
rect 3808 3836 3872 3840
rect 3808 3780 3812 3836
rect 3812 3780 3868 3836
rect 3868 3780 3872 3836
rect 3808 3776 3872 3780
rect 2068 3292 2132 3296
rect 2068 3236 2072 3292
rect 2072 3236 2128 3292
rect 2128 3236 2132 3292
rect 2068 3232 2132 3236
rect 2148 3292 2212 3296
rect 2148 3236 2152 3292
rect 2152 3236 2208 3292
rect 2208 3236 2212 3292
rect 2148 3232 2212 3236
rect 2228 3292 2292 3296
rect 2228 3236 2232 3292
rect 2232 3236 2288 3292
rect 2288 3236 2292 3292
rect 2228 3232 2292 3236
rect 2308 3292 2372 3296
rect 2308 3236 2312 3292
rect 2312 3236 2368 3292
rect 2368 3236 2372 3292
rect 2308 3232 2372 3236
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 3568 2748 3632 2752
rect 3568 2692 3572 2748
rect 3572 2692 3628 2748
rect 3628 2692 3632 2748
rect 3568 2688 3632 2692
rect 3648 2748 3712 2752
rect 3648 2692 3652 2748
rect 3652 2692 3708 2748
rect 3708 2692 3712 2748
rect 3648 2688 3712 2692
rect 3728 2748 3792 2752
rect 3728 2692 3732 2748
rect 3732 2692 3788 2748
rect 3788 2692 3792 2748
rect 3728 2688 3792 2692
rect 3808 2748 3872 2752
rect 3808 2692 3812 2748
rect 3812 2692 3868 2748
rect 3868 2692 3872 2748
rect 3808 2688 3872 2692
rect 2068 2204 2132 2208
rect 2068 2148 2072 2204
rect 2072 2148 2128 2204
rect 2128 2148 2132 2204
rect 2068 2144 2132 2148
rect 2148 2204 2212 2208
rect 2148 2148 2152 2204
rect 2152 2148 2208 2204
rect 2208 2148 2212 2204
rect 2148 2144 2212 2148
rect 2228 2204 2292 2208
rect 2228 2148 2232 2204
rect 2232 2148 2288 2204
rect 2288 2148 2292 2204
rect 2228 2144 2292 2148
rect 2308 2204 2372 2208
rect 2308 2148 2312 2204
rect 2312 2148 2368 2204
rect 2368 2148 2372 2204
rect 2308 2144 2372 2148
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
<< metal4 >>
rect -1620 13922 -1300 13964
rect -1620 13686 -1578 13922
rect -1342 13686 -1300 13922
rect -1620 9694 -1300 13686
rect -1620 9458 -1578 9694
rect -1342 9458 -1300 9694
rect -1620 6494 -1300 9458
rect -1620 6258 -1578 6494
rect -1342 6258 -1300 6494
rect -1620 -86 -1300 6258
rect -960 13262 -640 13304
rect -960 13026 -918 13262
rect -682 13026 -640 13262
rect -960 8094 -640 13026
rect 2960 13262 3280 13964
rect 2960 13026 3002 13262
rect 3238 13026 3280 13262
rect -960 7858 -918 8094
rect -682 7858 -640 8094
rect -960 4894 -640 7858
rect -960 4658 -918 4894
rect -682 4658 -640 4894
rect -960 574 -640 4658
rect -300 12602 20 12644
rect -300 12366 -258 12602
rect -22 12366 20 12602
rect -300 8794 20 12366
rect -300 8558 -258 8794
rect -22 8558 20 8794
rect -300 5594 20 8558
rect -300 5358 -258 5594
rect -22 5358 20 5594
rect -300 1234 20 5358
rect 360 11942 680 11984
rect 360 11706 402 11942
rect 638 11706 680 11942
rect 360 10394 680 11706
rect 360 10158 402 10394
rect 638 10158 680 10394
rect 360 7194 680 10158
rect 360 6958 402 7194
rect 638 6958 680 7194
rect 360 3994 680 6958
rect 360 3758 402 3994
rect 638 3758 680 3994
rect 360 1894 680 3758
rect 360 1658 402 1894
rect 638 1658 680 1894
rect 360 1616 680 1658
rect 2060 11942 2380 12644
rect 2060 11706 2102 11942
rect 2338 11706 2380 11942
rect 2060 10912 2380 11706
rect 2060 10848 2068 10912
rect 2132 10848 2148 10912
rect 2212 10848 2228 10912
rect 2292 10848 2308 10912
rect 2372 10848 2380 10912
rect 2060 10394 2380 10848
rect 2060 10158 2102 10394
rect 2338 10158 2380 10394
rect 2060 9824 2380 10158
rect 2060 9760 2068 9824
rect 2132 9760 2148 9824
rect 2212 9760 2228 9824
rect 2292 9760 2308 9824
rect 2372 9760 2380 9824
rect 2060 8736 2380 9760
rect 2060 8672 2068 8736
rect 2132 8672 2148 8736
rect 2212 8672 2228 8736
rect 2292 8672 2308 8736
rect 2372 8672 2380 8736
rect 2060 7648 2380 8672
rect 2060 7584 2068 7648
rect 2132 7584 2148 7648
rect 2212 7584 2228 7648
rect 2292 7584 2308 7648
rect 2372 7584 2380 7648
rect 2060 7194 2380 7584
rect 2060 6958 2102 7194
rect 2338 6958 2380 7194
rect 2060 6560 2380 6958
rect 2060 6496 2068 6560
rect 2132 6496 2148 6560
rect 2212 6496 2228 6560
rect 2292 6496 2308 6560
rect 2372 6496 2380 6560
rect 2060 5472 2380 6496
rect 2060 5408 2068 5472
rect 2132 5408 2148 5472
rect 2212 5408 2228 5472
rect 2292 5408 2308 5472
rect 2372 5408 2380 5472
rect 2060 4384 2380 5408
rect 2060 4320 2068 4384
rect 2132 4320 2148 4384
rect 2212 4320 2228 4384
rect 2292 4320 2308 4384
rect 2372 4320 2380 4384
rect 2060 3994 2380 4320
rect 2060 3758 2102 3994
rect 2338 3758 2380 3994
rect 2060 3296 2380 3758
rect 2060 3232 2068 3296
rect 2132 3232 2148 3296
rect 2212 3232 2228 3296
rect 2292 3232 2308 3296
rect 2372 3232 2380 3296
rect 2060 2208 2380 3232
rect 2060 2144 2068 2208
rect 2132 2144 2148 2208
rect 2212 2144 2228 2208
rect 2292 2144 2308 2208
rect 2372 2144 2380 2208
rect 2060 1894 2380 2144
rect 2060 1658 2102 1894
rect 2338 1658 2380 1894
rect -300 998 -258 1234
rect -22 998 20 1234
rect -300 956 20 998
rect 2060 956 2380 1658
rect 2960 8094 3280 13026
rect 4460 13922 4780 13964
rect 4460 13686 4502 13922
rect 4738 13686 4780 13922
rect 2960 7858 3002 8094
rect 3238 7858 3280 8094
rect 2960 4894 3280 7858
rect 2960 4658 3002 4894
rect 3238 4658 3280 4894
rect -960 338 -918 574
rect -682 338 -640 574
rect -960 296 -640 338
rect 2960 574 3280 4658
rect 3560 12602 3880 12644
rect 3560 12366 3602 12602
rect 3838 12366 3880 12602
rect 3560 11456 3880 12366
rect 3560 11392 3568 11456
rect 3632 11392 3648 11456
rect 3712 11392 3728 11456
rect 3792 11392 3808 11456
rect 3872 11392 3880 11456
rect 3560 10368 3880 11392
rect 3560 10304 3568 10368
rect 3632 10304 3648 10368
rect 3712 10304 3728 10368
rect 3792 10304 3808 10368
rect 3872 10304 3880 10368
rect 3560 9280 3880 10304
rect 3560 9216 3568 9280
rect 3632 9216 3648 9280
rect 3712 9216 3728 9280
rect 3792 9216 3808 9280
rect 3872 9216 3880 9280
rect 3560 8794 3880 9216
rect 3560 8558 3602 8794
rect 3838 8558 3880 8794
rect 3560 8192 3880 8558
rect 3560 8128 3568 8192
rect 3632 8128 3648 8192
rect 3712 8128 3728 8192
rect 3792 8128 3808 8192
rect 3872 8128 3880 8192
rect 3560 7104 3880 8128
rect 3560 7040 3568 7104
rect 3632 7040 3648 7104
rect 3712 7040 3728 7104
rect 3792 7040 3808 7104
rect 3872 7040 3880 7104
rect 3560 6016 3880 7040
rect 3560 5952 3568 6016
rect 3632 5952 3648 6016
rect 3712 5952 3728 6016
rect 3792 5952 3808 6016
rect 3872 5952 3880 6016
rect 3560 5594 3880 5952
rect 3560 5358 3602 5594
rect 3838 5358 3880 5594
rect 3560 4928 3880 5358
rect 3560 4864 3568 4928
rect 3632 4864 3648 4928
rect 3712 4864 3728 4928
rect 3792 4864 3808 4928
rect 3872 4864 3880 4928
rect 3560 3840 3880 4864
rect 3560 3776 3568 3840
rect 3632 3776 3648 3840
rect 3712 3776 3728 3840
rect 3792 3776 3808 3840
rect 3872 3776 3880 3840
rect 3560 2752 3880 3776
rect 3560 2688 3568 2752
rect 3632 2688 3648 2752
rect 3712 2688 3728 2752
rect 3792 2688 3808 2752
rect 3872 2688 3880 2752
rect 3560 1234 3880 2688
rect 3560 998 3602 1234
rect 3838 998 3880 1234
rect 3560 956 3880 998
rect 4460 9694 4780 13686
rect 5960 13262 6280 13964
rect 9304 13922 9624 13964
rect 9304 13686 9346 13922
rect 9582 13686 9624 13922
rect 5960 13026 6002 13262
rect 6238 13026 6280 13262
rect 4460 9458 4502 9694
rect 4738 9458 4780 9694
rect 4460 6494 4780 9458
rect 4460 6258 4502 6494
rect 4738 6258 4780 6494
rect 2960 338 3002 574
rect 3238 338 3280 574
rect -1620 -322 -1578 -86
rect -1342 -322 -1300 -86
rect -1620 -364 -1300 -322
rect 2960 -364 3280 338
rect 4460 -86 4780 6258
rect 5060 11942 5380 12644
rect 5060 11706 5102 11942
rect 5338 11706 5380 11942
rect 5060 10912 5380 11706
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10394 5380 10848
rect 5060 10158 5102 10394
rect 5338 10158 5380 10394
rect 5060 9824 5380 10158
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 5060 8736 5380 9760
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7194 5380 7584
rect 5060 6958 5102 7194
rect 5338 6958 5380 7194
rect 5060 6560 5380 6958
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 5060 5472 5380 6496
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3994 5380 4320
rect 5060 3758 5102 3994
rect 5338 3758 5380 3994
rect 5060 3296 5380 3758
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 2208 5380 3232
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1894 5380 2144
rect 5060 1658 5102 1894
rect 5338 1658 5380 1894
rect 5060 956 5380 1658
rect 5960 8094 6280 13026
rect 8644 13262 8964 13304
rect 8644 13026 8686 13262
rect 8922 13026 8964 13262
rect 7984 12602 8304 12644
rect 7984 12366 8026 12602
rect 8262 12366 8304 12602
rect 5960 7858 6002 8094
rect 6238 7858 6280 8094
rect 5960 4894 6280 7858
rect 5960 4658 6002 4894
rect 6238 4658 6280 4894
rect 4460 -322 4502 -86
rect 4738 -322 4780 -86
rect 4460 -364 4780 -322
rect 5960 574 6280 4658
rect 7324 11942 7644 11984
rect 7324 11706 7366 11942
rect 7602 11706 7644 11942
rect 7324 10394 7644 11706
rect 7324 10158 7366 10394
rect 7602 10158 7644 10394
rect 7324 7194 7644 10158
rect 7324 6958 7366 7194
rect 7602 6958 7644 7194
rect 7324 3994 7644 6958
rect 7324 3758 7366 3994
rect 7602 3758 7644 3994
rect 7324 1894 7644 3758
rect 7324 1658 7366 1894
rect 7602 1658 7644 1894
rect 7324 1616 7644 1658
rect 7984 8794 8304 12366
rect 7984 8558 8026 8794
rect 8262 8558 8304 8794
rect 7984 5594 8304 8558
rect 7984 5358 8026 5594
rect 8262 5358 8304 5594
rect 7984 1234 8304 5358
rect 7984 998 8026 1234
rect 8262 998 8304 1234
rect 7984 956 8304 998
rect 8644 8094 8964 13026
rect 8644 7858 8686 8094
rect 8922 7858 8964 8094
rect 8644 4894 8964 7858
rect 8644 4658 8686 4894
rect 8922 4658 8964 4894
rect 5960 338 6002 574
rect 6238 338 6280 574
rect 5960 -364 6280 338
rect 8644 574 8964 4658
rect 8644 338 8686 574
rect 8922 338 8964 574
rect 8644 296 8964 338
rect 9304 9694 9624 13686
rect 9304 9458 9346 9694
rect 9582 9458 9624 9694
rect 9304 6494 9624 9458
rect 9304 6258 9346 6494
rect 9582 6258 9624 6494
rect 9304 -86 9624 6258
rect 9304 -322 9346 -86
rect 9582 -322 9624 -86
rect 9304 -364 9624 -322
<< via4 >>
rect -1578 13686 -1342 13922
rect -1578 9458 -1342 9694
rect -1578 6258 -1342 6494
rect -918 13026 -682 13262
rect 3002 13026 3238 13262
rect -918 7858 -682 8094
rect -918 4658 -682 4894
rect -258 12366 -22 12602
rect -258 8558 -22 8794
rect -258 5358 -22 5594
rect 402 11706 638 11942
rect 402 10158 638 10394
rect 402 6958 638 7194
rect 402 3758 638 3994
rect 402 1658 638 1894
rect 2102 11706 2338 11942
rect 2102 10158 2338 10394
rect 2102 6958 2338 7194
rect 2102 3758 2338 3994
rect 2102 1658 2338 1894
rect -258 998 -22 1234
rect 4502 13686 4738 13922
rect 3002 7858 3238 8094
rect 3002 4658 3238 4894
rect -918 338 -682 574
rect 3602 12366 3838 12602
rect 3602 8558 3838 8794
rect 3602 5358 3838 5594
rect 3602 998 3838 1234
rect 9346 13686 9582 13922
rect 6002 13026 6238 13262
rect 4502 9458 4738 9694
rect 4502 6258 4738 6494
rect 3002 338 3238 574
rect -1578 -322 -1342 -86
rect 5102 11706 5338 11942
rect 5102 10158 5338 10394
rect 5102 6958 5338 7194
rect 5102 3758 5338 3994
rect 5102 1658 5338 1894
rect 8686 13026 8922 13262
rect 8026 12366 8262 12602
rect 6002 7858 6238 8094
rect 6002 4658 6238 4894
rect 4502 -322 4738 -86
rect 7366 11706 7602 11942
rect 7366 10158 7602 10394
rect 7366 6958 7602 7194
rect 7366 3758 7602 3994
rect 7366 1658 7602 1894
rect 8026 8558 8262 8794
rect 8026 5358 8262 5594
rect 8026 998 8262 1234
rect 8686 7858 8922 8094
rect 8686 4658 8922 4894
rect 6002 338 6238 574
rect 8686 338 8922 574
rect 9346 9458 9582 9694
rect 9346 6258 9582 6494
rect 9346 -322 9582 -86
<< metal5 >>
rect -1620 13922 9624 13964
rect -1620 13686 -1578 13922
rect -1342 13686 4502 13922
rect 4738 13686 9346 13922
rect 9582 13686 9624 13922
rect -1620 13644 9624 13686
rect -960 13262 8964 13304
rect -960 13026 -918 13262
rect -682 13026 3002 13262
rect 3238 13026 6002 13262
rect 6238 13026 8686 13262
rect 8922 13026 8964 13262
rect -960 12984 8964 13026
rect -300 12602 8304 12644
rect -300 12366 -258 12602
rect -22 12366 3602 12602
rect 3838 12366 8026 12602
rect 8262 12366 8304 12602
rect -300 12324 8304 12366
rect 360 11942 7644 11984
rect 360 11706 402 11942
rect 638 11706 2102 11942
rect 2338 11706 5102 11942
rect 5338 11706 7366 11942
rect 7602 11706 7644 11942
rect 360 11664 7644 11706
rect -300 10394 8304 10436
rect -300 10158 402 10394
rect 638 10158 2102 10394
rect 2338 10158 5102 10394
rect 5338 10158 7366 10394
rect 7602 10158 8304 10394
rect -300 10116 8304 10158
rect -1620 9694 9624 9736
rect -1620 9458 -1578 9694
rect -1342 9458 4502 9694
rect 4738 9458 9346 9694
rect 9582 9458 9624 9694
rect -1620 9416 9624 9458
rect -300 8794 8304 8836
rect -300 8558 -258 8794
rect -22 8558 3602 8794
rect 3838 8558 8026 8794
rect 8262 8558 8304 8794
rect -300 8516 8304 8558
rect -1620 8094 9624 8136
rect -1620 7858 -918 8094
rect -682 7858 3002 8094
rect 3238 7858 6002 8094
rect 6238 7858 8686 8094
rect 8922 7858 9624 8094
rect -1620 7816 9624 7858
rect -300 7194 8304 7236
rect -300 6958 402 7194
rect 638 6958 2102 7194
rect 2338 6958 5102 7194
rect 5338 6958 7366 7194
rect 7602 6958 8304 7194
rect -300 6916 8304 6958
rect -1620 6494 9624 6536
rect -1620 6258 -1578 6494
rect -1342 6258 4502 6494
rect 4738 6258 9346 6494
rect 9582 6258 9624 6494
rect -1620 6216 9624 6258
rect -300 5594 8304 5636
rect -300 5358 -258 5594
rect -22 5358 3602 5594
rect 3838 5358 8026 5594
rect 8262 5358 8304 5594
rect -300 5316 8304 5358
rect -1620 4894 9624 4936
rect -1620 4658 -918 4894
rect -682 4658 3002 4894
rect 3238 4658 6002 4894
rect 6238 4658 8686 4894
rect 8922 4658 9624 4894
rect -1620 4616 9624 4658
rect -300 3994 8304 4036
rect -300 3758 402 3994
rect 638 3758 2102 3994
rect 2338 3758 5102 3994
rect 5338 3758 7366 3994
rect 7602 3758 8304 3994
rect -300 3716 8304 3758
rect 360 1894 7644 1936
rect 360 1658 402 1894
rect 638 1658 2102 1894
rect 2338 1658 5102 1894
rect 5338 1658 7366 1894
rect 7602 1658 7644 1894
rect 360 1616 7644 1658
rect -300 1234 8304 1276
rect -300 998 -258 1234
rect -22 998 3602 1234
rect 3838 998 8026 1234
rect 8262 998 8304 1234
rect -300 956 8304 998
rect -960 574 8964 616
rect -960 338 -918 574
rect -682 338 3002 574
rect 3238 338 6002 574
rect 6238 338 8686 574
rect 8922 338 8964 574
rect -960 296 8964 338
rect -1620 -86 9624 -44
rect -1620 -322 -1578 -86
rect -1342 -322 4502 -86
rect 4738 -322 9346 -86
rect 9582 -322 9624 -86
rect -1620 -364 9624 -322
use sky130_fd_sc_hd__dfrtp_4  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 1656 0 1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _100_
timestamp 1611237355
transform 1 0 1656 0 -1 2720
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 920 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1611237355
transform 1 0 920 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 1196 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 1564 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1611237355
transform 1 0 1196 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7
timestamp 1611237355
transform 1 0 1564 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1611237355
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1611237355
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 4416 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 4968 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1611237355
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 4232 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1611237355
transform 1 0 5612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 5980 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1611237355
transform -1 0 7084 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1611237355
transform -1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1611237355
transform 1 0 6624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 6624 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1611237355
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1611237355
transform 1 0 1932 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _099_
timestamp 1611237355
transform 1 0 2300 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1611237355
transform 1 0 920 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1611237355
transform 1 0 1196 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _095_
timestamp 1611237355
transform 1 0 4416 0 -1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1611237355
transform -1 0 7084 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1611237355
transform 1 0 6532 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A_0
timestamp 1611237355
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _108_
timestamp 1611237355
transform 1 0 1196 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1611237355
transform 1 0 920 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _048_
timestamp 1611237355
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _112_
timestamp 1611237355
transform 1 0 3864 0 1 3808
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1611237355
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1611237355
transform 1 0 3680 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 5980 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1611237355
transform -1 0 7084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _109_
timestamp 1611237355
transform 1 0 1288 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1611237355
transform 1 0 920 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1611237355
transform 1 0 1196 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _111_
timestamp 1611237355
transform 1 0 3404 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__nand2_4  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1611237355
transform -1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1611237355
transform 1 0 6532 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A_0
timestamp 1611237355
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__C_0
timestamp 1611237355
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _107_
timestamp 1611237355
transform 1 0 1196 0 1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1611237355
transform 1 0 920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _044_
timestamp 1611237355
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _045_
timestamp 1611237355
transform 1 0 3956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _097_
timestamp 1611237355
transform 1 0 4600 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1611237355
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_30
timestamp 1611237355
transform 1 0 3680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_32
timestamp 1611237355
transform 1 0 3864 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1611237355
transform -1 0 7084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _047_
timestamp 1611237355
transform 1 0 2208 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _050_
timestamp 1611237355
transform 1 0 1840 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _106_
timestamp 1611237355
transform 1 0 1196 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _110_
timestamp 1611237355
transform 1 0 2576 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1611237355
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1611237355
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 1564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1611237355
transform 1 0 1196 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _046_
timestamp 1611237355
transform 1 0 3404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1611237355
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1611237355
transform 1 0 4968 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _093_
timestamp 1611237355
transform 1 0 4232 0 1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1611237355
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A_0
timestamp 1611237355
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_43
timestamp 1611237355
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1611237355
transform 1 0 3312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_32
timestamp 1611237355
transform 1 0 3864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1611237355
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 5704 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1611237355
transform -1 0 7084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1611237355
transform -1 0 7084 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1611237355
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__D_0
timestamp 1611237355
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_63
timestamp 1611237355
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _051_
timestamp 1611237355
transform 1 0 1840 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _052_
timestamp 1611237355
transform 1 0 2208 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _092_
timestamp 1611237355
transform 1 0 2944 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1611237355
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 1196 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1611237355
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1611237355
transform 1 0 2576 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1611237355
transform 1 0 5060 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1611237355
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _086_
timestamp 1611237355
transform 1 0 5704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1611237355
transform -1 0 7084 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1611237355
transform 1 0 6532 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A_0
timestamp 1611237355
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _105_
timestamp 1611237355
transform 1 0 1288 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1611237355
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1611237355
transform 1 0 1196 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1611237355
transform 1 0 3956 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1611237355
transform 1 0 3404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _113_
timestamp 1611237355
transform 1 0 4324 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1611237355
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_32
timestamp 1611237355
transform 1 0 3864 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1611237355
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1611237355
transform -1 0 7084 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _104_
timestamp 1611237355
transform 1 0 1196 0 -1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1611237355
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _049_
timestamp 1611237355
transform 1 0 3312 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _094_
timestamp 1611237355
transform 1 0 3864 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_10_30
timestamp 1611237355
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1611237355
transform 1 0 6072 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1611237355
transform -1 0 7084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1611237355
transform 1 0 6532 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A_0
timestamp 1611237355
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_60
timestamp 1611237355
transform 1 0 6440 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _103_
timestamp 1611237355
transform 1 0 1196 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1611237355
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1611237355
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1611237355
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 3864 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1611237355
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _043_
timestamp 1611237355
transform 1 0 5704 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1611237355
transform 1 0 6072 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1611237355
transform -1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A_0
timestamp 1611237355
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B1_0
timestamp 1611237355
transform 1 0 6624 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _053_
timestamp 1611237355
transform 1 0 1932 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _054_
timestamp 1611237355
transform 1 0 2300 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1611237355
transform 1 0 1656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _089_
timestamp 1611237355
transform 1 0 2852 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1611237355
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_serial_clock
timestamp 1611237355
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B2_0
timestamp 1611237355
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1611237355
transform 1 0 1196 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 4968 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1611237355
transform -1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1611237355
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A2_0
timestamp 1611237355
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _055_
timestamp 1611237355
transform 1 0 1840 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_4  _081_
timestamp 1611237355
transform 1 0 2208 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_4  _102_
timestamp 1611237355
transform 1 0 1196 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1611237355
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1611237355
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1611237355
transform 1 0 1196 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1611237355
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _088_
timestamp 1611237355
transform 1 0 3312 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_4  _090_
timestamp 1611237355
transform 1 0 3864 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1611237355
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _042_
timestamp 1611237355
transform 1 0 5520 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1611237355
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 5980 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1611237355
transform -1 0 7084 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1611237355
transform -1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1611237355
transform 1 0 6532 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__042__B_0
timestamp 1611237355
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1611237355
transform 1 0 6624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _101_
timestamp 1611237355
transform 1 0 1564 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1611237355
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1611237355
transform 1 0 1196 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1611237355
transform 1 0 3864 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _091_
timestamp 1611237355
transform 1 0 4324 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1611237355
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_30
timestamp 1611237355
transform 1 0 3680 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_36
timestamp 1611237355
transform 1 0 4232 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1611237355
transform 1 0 6440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1611237355
transform -1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high
timestamp 1611237355
transform 1 0 1196 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1611237355
transform 1 0 920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 1472 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_18
timestamp 1611237355
transform 1 0 2576 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_24
timestamp 1611237355
transform 1 0 3128 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1611237355
transform 1 0 4324 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1611237355
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__D_0
timestamp 1611237355
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A_0
timestamp 1611237355
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A_0
timestamp 1611237355
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1611237355
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1611237355
transform 1 0 3956 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1611237355
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1611237355
transform 1 0 4692 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611237355
transform 1 0 4968 0 -1 11424
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1611237355
transform -1 0 7084 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1611237355
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_63
timestamp 1611237355
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
<< labels >>
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_in
port 0 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 1 nsew signal input
rlabel metal3 s 14000 2184 34000 2304 6 mgmt_gpio_out
port 2 nsew signal input
rlabel metal3 s 14000 552 34000 672 6 one
port 3 nsew signal tristate
rlabel metal3 s 14000 2728 34000 2848 6 pad_gpio_ana_en
port 4 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_pol
port 5 nsew signal tristate
rlabel metal3 s 14000 3816 34000 3936 6 pad_gpio_ana_sel
port 6 nsew signal tristate
rlabel metal3 s 14000 4360 34000 4480 6 pad_gpio_dm[0]
port 7 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_dm[1]
port 8 nsew signal tristate
rlabel metal3 s 14000 5448 34000 5568 6 pad_gpio_dm[2]
port 9 nsew signal tristate
rlabel metal3 s 14000 5992 34000 6112 6 pad_gpio_holdover
port 10 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ib_mode_sel
port 11 nsew signal tristate
rlabel metal3 s 14000 7080 34000 7200 6 pad_gpio_in
port 12 nsew signal input
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_inenb
port 13 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_out
port 14 nsew signal tristate
rlabel metal3 s 14000 8712 34000 8832 6 pad_gpio_outenb
port 15 nsew signal tristate
rlabel metal3 s 14000 9256 34000 9376 6 pad_gpio_slow_sel
port 16 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_vtrip_sel
port 17 nsew signal tristate
rlabel metal3 s 14000 10344 34000 10464 6 resetn
port 18 nsew signal input
rlabel metal3 s 14000 10888 34000 11008 6 serial_clock
port 19 nsew signal input
rlabel metal3 s 14000 11432 34000 11552 6 serial_data_in
port 20 nsew signal input
rlabel metal3 s 14000 11976 34000 12096 6 serial_data_out
port 21 nsew signal tristate
rlabel metal3 s 14000 12520 34000 12640 6 user_gpio_in
port 22 nsew signal tristate
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_oeb
port 23 nsew signal input
rlabel metal3 s 14000 13608 34000 13728 6 user_gpio_out
port 24 nsew signal input
rlabel metal3 s 14000 144 34000 264 6 zero
port 25 nsew signal tristate
rlabel metal4 s 5060 956 5380 12644 6 vccd
port 26 nsew power bidirectional
rlabel metal4 s 2060 956 2380 12644 6 vccd
port 27 nsew power bidirectional
rlabel metal4 s 7324 1616 7644 11984 6 vccd
port 28 nsew power bidirectional
rlabel metal4 s 360 1616 680 11984 6 vccd
port 29 nsew power bidirectional
rlabel metal5 s 360 11664 7644 11984 6 vccd
port 30 nsew power bidirectional
rlabel metal5 s -300 10116 8304 10436 6 vccd
port 31 nsew power bidirectional
rlabel metal5 s -300 6916 8304 7236 6 vccd
port 32 nsew power bidirectional
rlabel metal5 s -300 3716 8304 4036 6 vccd
port 33 nsew power bidirectional
rlabel metal5 s 360 1616 7644 1936 6 vccd
port 34 nsew power bidirectional
rlabel metal4 s 7984 956 8304 12644 6 vssd
port 35 nsew ground bidirectional
rlabel metal4 s 3560 956 3880 12644 6 vssd
port 36 nsew ground bidirectional
rlabel metal4 s -300 956 20 12644 4 vssd
port 37 nsew ground bidirectional
rlabel metal5 s -300 12324 8304 12644 6 vssd
port 38 nsew ground bidirectional
rlabel metal5 s -300 8516 8304 8836 6 vssd
port 39 nsew ground bidirectional
rlabel metal5 s -300 5316 8304 5636 6 vssd
port 40 nsew ground bidirectional
rlabel metal5 s -300 956 8304 1276 6 vssd
port 41 nsew ground bidirectional
rlabel metal4 s 5960 -364 6280 13964 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 2960 -364 3280 13964 6 vccd1
port 43 nsew power bidirectional
rlabel metal4 s 8644 296 8964 13304 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 45 nsew power bidirectional
rlabel metal5 s -960 12984 8964 13304 6 vccd1
port 46 nsew power bidirectional
rlabel metal5 s -1620 7816 9624 8136 6 vccd1
port 47 nsew power bidirectional
rlabel metal5 s -1620 4616 9624 4936 6 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -960 296 8964 616 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 9304 -364 9624 13964 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 4460 -364 4780 13964 6 vssd1
port 51 nsew ground bidirectional
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 52 nsew ground bidirectional
rlabel metal5 s -1620 13644 9624 13964 6 vssd1
port 53 nsew ground bidirectional
rlabel metal5 s -1620 9416 9624 9736 6 vssd1
port 54 nsew ground bidirectional
rlabel metal5 s -1620 6216 9624 6536 6 vssd1
port 55 nsew ground bidirectional
rlabel metal5 s -1620 -364 9624 -44 8 vssd1
port 56 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 34000 14000
<< end >>
